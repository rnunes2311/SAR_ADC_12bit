magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< pwell >>
rect -1031 -2382 1031 2382
<< psubdiff >>
rect -995 2312 -899 2346
rect 899 2312 995 2346
rect -995 2250 -961 2312
rect 961 2250 995 2312
rect -995 -2312 -961 -2250
rect 961 -2312 995 -2250
rect -995 -2346 -899 -2312
rect 899 -2346 995 -2312
<< psubdiffcont >>
rect -899 2312 899 2346
rect -995 -2250 -961 2250
rect 961 -2250 995 2250
rect -899 -2346 899 -2312
<< xpolycontact >>
rect -865 1784 -795 2216
rect -865 -2216 -795 -1784
rect -699 1784 -629 2216
rect -699 -2216 -629 -1784
rect -533 1784 -463 2216
rect -533 -2216 -463 -1784
rect -367 1784 -297 2216
rect -367 -2216 -297 -1784
rect -201 1784 -131 2216
rect -201 -2216 -131 -1784
rect -35 1784 35 2216
rect -35 -2216 35 -1784
rect 131 1784 201 2216
rect 131 -2216 201 -1784
rect 297 1784 367 2216
rect 297 -2216 367 -1784
rect 463 1784 533 2216
rect 463 -2216 533 -1784
rect 629 1784 699 2216
rect 629 -2216 699 -1784
rect 795 1784 865 2216
rect 795 -2216 865 -1784
<< ppolyres >>
rect -865 -1784 -795 1784
rect -699 -1784 -629 1784
rect -533 -1784 -463 1784
rect -367 -1784 -297 1784
rect -201 -1784 -131 1784
rect -35 -1784 35 1784
rect 131 -1784 201 1784
rect 297 -1784 367 1784
rect 463 -1784 533 1784
rect 629 -1784 699 1784
rect 795 -1784 865 1784
<< locali >>
rect -995 2312 -899 2346
rect 899 2312 995 2346
rect -995 2250 -961 2312
rect 961 2250 995 2312
rect -995 -2312 -961 -2250
rect 961 -2312 995 -2250
rect -995 -2346 -899 -2312
rect 899 -2346 995 -2312
<< viali >>
rect -849 1801 -811 2198
rect -683 1801 -645 2198
rect -517 1801 -479 2198
rect -351 1801 -313 2198
rect -185 1801 -147 2198
rect -19 1801 19 2198
rect 147 1801 185 2198
rect 313 1801 351 2198
rect 479 1801 517 2198
rect 645 1801 683 2198
rect 811 1801 849 2198
rect -849 -2198 -811 -1801
rect -683 -2198 -645 -1801
rect -517 -2198 -479 -1801
rect -351 -2198 -313 -1801
rect -185 -2198 -147 -1801
rect -19 -2198 19 -1801
rect 147 -2198 185 -1801
rect 313 -2198 351 -1801
rect 479 -2198 517 -1801
rect 645 -2198 683 -1801
rect 811 -2198 849 -1801
<< metal1 >>
rect -855 2198 -805 2210
rect -855 1801 -849 2198
rect -811 1801 -805 2198
rect -855 1789 -805 1801
rect -689 2198 -639 2210
rect -689 1801 -683 2198
rect -645 1801 -639 2198
rect -689 1789 -639 1801
rect -523 2198 -473 2210
rect -523 1801 -517 2198
rect -479 1801 -473 2198
rect -523 1789 -473 1801
rect -357 2198 -307 2210
rect -357 1801 -351 2198
rect -313 1801 -307 2198
rect -357 1789 -307 1801
rect -191 2198 -141 2210
rect -191 1801 -185 2198
rect -147 1801 -141 2198
rect -191 1789 -141 1801
rect -25 2198 25 2210
rect -25 1801 -19 2198
rect 19 1801 25 2198
rect -25 1789 25 1801
rect 141 2198 191 2210
rect 141 1801 147 2198
rect 185 1801 191 2198
rect 141 1789 191 1801
rect 307 2198 357 2210
rect 307 1801 313 2198
rect 351 1801 357 2198
rect 307 1789 357 1801
rect 473 2198 523 2210
rect 473 1801 479 2198
rect 517 1801 523 2198
rect 473 1789 523 1801
rect 639 2198 689 2210
rect 639 1801 645 2198
rect 683 1801 689 2198
rect 639 1789 689 1801
rect 805 2198 855 2210
rect 805 1801 811 2198
rect 849 1801 855 2198
rect 805 1789 855 1801
rect -855 -1801 -805 -1789
rect -855 -2198 -849 -1801
rect -811 -2198 -805 -1801
rect -855 -2210 -805 -2198
rect -689 -1801 -639 -1789
rect -689 -2198 -683 -1801
rect -645 -2198 -639 -1801
rect -689 -2210 -639 -2198
rect -523 -1801 -473 -1789
rect -523 -2198 -517 -1801
rect -479 -2198 -473 -1801
rect -523 -2210 -473 -2198
rect -357 -1801 -307 -1789
rect -357 -2198 -351 -1801
rect -313 -2198 -307 -1801
rect -357 -2210 -307 -2198
rect -191 -1801 -141 -1789
rect -191 -2198 -185 -1801
rect -147 -2198 -141 -1801
rect -191 -2210 -141 -2198
rect -25 -1801 25 -1789
rect -25 -2198 -19 -1801
rect 19 -2198 25 -1801
rect -25 -2210 25 -2198
rect 141 -1801 191 -1789
rect 141 -2198 147 -1801
rect 185 -2198 191 -1801
rect 141 -2210 191 -2198
rect 307 -1801 357 -1789
rect 307 -2198 313 -1801
rect 351 -2198 357 -1801
rect 307 -2210 357 -2198
rect 473 -1801 523 -1789
rect 473 -2198 479 -1801
rect 517 -2198 523 -1801
rect 473 -2210 523 -2198
rect 639 -1801 689 -1789
rect 639 -2198 645 -1801
rect 683 -2198 689 -1801
rect 639 -2210 689 -2198
rect 805 -1801 855 -1789
rect 805 -2198 811 -1801
rect 849 -2198 855 -1801
rect 805 -2210 855 -2198
<< properties >>
string FIXED_BBOX -978 -2329 978 2329
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 18.0 m 1 nx 11 wmin 0.350 lmin 0.50 rho 319.8 val 17.56k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
