magic
tech sky130A
timestamp 1710675123
<< pwell >>
rect -159 -329 159 329
<< mvnnmos >>
rect -45 -200 45 200
<< mvndiff >>
rect -74 194 -45 200
rect -74 -194 -68 194
rect -51 -194 -45 194
rect -74 -200 -45 -194
rect 45 194 74 200
rect 45 -194 51 194
rect 68 -194 74 194
rect 45 -200 74 -194
<< mvndiffc >>
rect -68 -194 -51 194
rect 51 -194 68 194
<< mvpsubdiff >>
rect -141 305 141 311
rect -141 288 -87 305
rect 87 288 141 305
rect -141 282 141 288
rect -141 257 -112 282
rect -141 -257 -135 257
rect -118 -257 -112 257
rect 112 257 141 282
rect -141 -282 -112 -257
rect 112 -257 118 257
rect 135 -257 141 257
rect 112 -282 141 -257
rect -141 -288 141 -282
rect -141 -305 -87 -288
rect 87 -305 141 -288
rect -141 -311 141 -305
<< mvpsubdiffcont >>
rect -87 288 87 305
rect -135 -257 -118 257
rect 118 -257 135 257
rect -87 -305 87 -288
<< poly >>
rect -45 236 45 244
rect -45 219 -37 236
rect 37 219 45 236
rect -45 200 45 219
rect -45 -219 45 -200
rect -45 -236 -37 -219
rect 37 -236 45 -219
rect -45 -244 45 -236
<< polycont >>
rect -37 219 37 236
rect -37 -236 37 -219
<< locali >>
rect -135 288 -87 305
rect 87 288 135 305
rect -135 257 -118 288
rect 118 257 135 288
rect -45 219 -37 236
rect 37 219 45 236
rect -68 194 -51 202
rect -68 -202 -51 -194
rect 51 194 68 202
rect 51 -202 68 -194
rect -45 -236 -37 -219
rect 37 -236 45 -219
rect -135 -288 -118 -257
rect 118 -288 135 -257
rect -135 -305 -87 -288
rect 87 -305 135 -288
<< viali >>
rect -37 219 37 236
rect -68 -194 -51 194
rect 51 -194 68 194
rect -37 -236 37 -219
<< metal1 >>
rect -43 236 43 239
rect -43 219 -37 236
rect 37 219 43 236
rect -43 216 43 219
rect -71 194 -48 200
rect -71 -194 -68 194
rect -51 -194 -48 194
rect -71 -200 -48 -194
rect 48 194 71 200
rect 48 -194 51 194
rect 68 -194 71 194
rect 48 -200 71 -194
rect -43 -219 43 -216
rect -43 -236 -37 -219
rect 37 -236 43 -219
rect -43 -239 43 -236
<< properties >>
string FIXED_BBOX -126 -296 126 296
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 4.0 l 0.9 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
