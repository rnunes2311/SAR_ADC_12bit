magic
tech sky130A
magscale 1 2
timestamp 1711883585
<< nwell >>
rect -926 -2855 926 2855
<< pmos >>
rect -730 1036 -630 2636
rect -458 1036 -358 2636
rect -186 1036 -86 2636
rect 86 1036 186 2636
rect 358 1036 458 2636
rect 630 1036 730 2636
rect -730 -800 -630 800
rect -458 -800 -358 800
rect -186 -800 -86 800
rect 86 -800 186 800
rect 358 -800 458 800
rect 630 -800 730 800
rect -730 -2636 -630 -1036
rect -458 -2636 -358 -1036
rect -186 -2636 -86 -1036
rect 86 -2636 186 -1036
rect 358 -2636 458 -1036
rect 630 -2636 730 -1036
<< pdiff >>
rect -788 2624 -730 2636
rect -788 1048 -776 2624
rect -742 1048 -730 2624
rect -788 1036 -730 1048
rect -630 2624 -572 2636
rect -630 1048 -618 2624
rect -584 1048 -572 2624
rect -630 1036 -572 1048
rect -516 2624 -458 2636
rect -516 1048 -504 2624
rect -470 1048 -458 2624
rect -516 1036 -458 1048
rect -358 2624 -300 2636
rect -358 1048 -346 2624
rect -312 1048 -300 2624
rect -358 1036 -300 1048
rect -244 2624 -186 2636
rect -244 1048 -232 2624
rect -198 1048 -186 2624
rect -244 1036 -186 1048
rect -86 2624 -28 2636
rect -86 1048 -74 2624
rect -40 1048 -28 2624
rect -86 1036 -28 1048
rect 28 2624 86 2636
rect 28 1048 40 2624
rect 74 1048 86 2624
rect 28 1036 86 1048
rect 186 2624 244 2636
rect 186 1048 198 2624
rect 232 1048 244 2624
rect 186 1036 244 1048
rect 300 2624 358 2636
rect 300 1048 312 2624
rect 346 1048 358 2624
rect 300 1036 358 1048
rect 458 2624 516 2636
rect 458 1048 470 2624
rect 504 1048 516 2624
rect 458 1036 516 1048
rect 572 2624 630 2636
rect 572 1048 584 2624
rect 618 1048 630 2624
rect 572 1036 630 1048
rect 730 2624 788 2636
rect 730 1048 742 2624
rect 776 1048 788 2624
rect 730 1036 788 1048
rect -788 788 -730 800
rect -788 -788 -776 788
rect -742 -788 -730 788
rect -788 -800 -730 -788
rect -630 788 -572 800
rect -630 -788 -618 788
rect -584 -788 -572 788
rect -630 -800 -572 -788
rect -516 788 -458 800
rect -516 -788 -504 788
rect -470 -788 -458 788
rect -516 -800 -458 -788
rect -358 788 -300 800
rect -358 -788 -346 788
rect -312 -788 -300 788
rect -358 -800 -300 -788
rect -244 788 -186 800
rect -244 -788 -232 788
rect -198 -788 -186 788
rect -244 -800 -186 -788
rect -86 788 -28 800
rect -86 -788 -74 788
rect -40 -788 -28 788
rect -86 -800 -28 -788
rect 28 788 86 800
rect 28 -788 40 788
rect 74 -788 86 788
rect 28 -800 86 -788
rect 186 788 244 800
rect 186 -788 198 788
rect 232 -788 244 788
rect 186 -800 244 -788
rect 300 788 358 800
rect 300 -788 312 788
rect 346 -788 358 788
rect 300 -800 358 -788
rect 458 788 516 800
rect 458 -788 470 788
rect 504 -788 516 788
rect 458 -800 516 -788
rect 572 788 630 800
rect 572 -788 584 788
rect 618 -788 630 788
rect 572 -800 630 -788
rect 730 788 788 800
rect 730 -788 742 788
rect 776 -788 788 788
rect 730 -800 788 -788
rect -788 -1048 -730 -1036
rect -788 -2624 -776 -1048
rect -742 -2624 -730 -1048
rect -788 -2636 -730 -2624
rect -630 -1048 -572 -1036
rect -630 -2624 -618 -1048
rect -584 -2624 -572 -1048
rect -630 -2636 -572 -2624
rect -516 -1048 -458 -1036
rect -516 -2624 -504 -1048
rect -470 -2624 -458 -1048
rect -516 -2636 -458 -2624
rect -358 -1048 -300 -1036
rect -358 -2624 -346 -1048
rect -312 -2624 -300 -1048
rect -358 -2636 -300 -2624
rect -244 -1048 -186 -1036
rect -244 -2624 -232 -1048
rect -198 -2624 -186 -1048
rect -244 -2636 -186 -2624
rect -86 -1048 -28 -1036
rect -86 -2624 -74 -1048
rect -40 -2624 -28 -1048
rect -86 -2636 -28 -2624
rect 28 -1048 86 -1036
rect 28 -2624 40 -1048
rect 74 -2624 86 -1048
rect 28 -2636 86 -2624
rect 186 -1048 244 -1036
rect 186 -2624 198 -1048
rect 232 -2624 244 -1048
rect 186 -2636 244 -2624
rect 300 -1048 358 -1036
rect 300 -2624 312 -1048
rect 346 -2624 358 -1048
rect 300 -2636 358 -2624
rect 458 -1048 516 -1036
rect 458 -2624 470 -1048
rect 504 -2624 516 -1048
rect 458 -2636 516 -2624
rect 572 -1048 630 -1036
rect 572 -2624 584 -1048
rect 618 -2624 630 -1048
rect 572 -2636 630 -2624
rect 730 -1048 788 -1036
rect 730 -2624 742 -1048
rect 776 -2624 788 -1048
rect 730 -2636 788 -2624
<< pdiffc >>
rect -776 1048 -742 2624
rect -618 1048 -584 2624
rect -504 1048 -470 2624
rect -346 1048 -312 2624
rect -232 1048 -198 2624
rect -74 1048 -40 2624
rect 40 1048 74 2624
rect 198 1048 232 2624
rect 312 1048 346 2624
rect 470 1048 504 2624
rect 584 1048 618 2624
rect 742 1048 776 2624
rect -776 -788 -742 788
rect -618 -788 -584 788
rect -504 -788 -470 788
rect -346 -788 -312 788
rect -232 -788 -198 788
rect -74 -788 -40 788
rect 40 -788 74 788
rect 198 -788 232 788
rect 312 -788 346 788
rect 470 -788 504 788
rect 584 -788 618 788
rect 742 -788 776 788
rect -776 -2624 -742 -1048
rect -618 -2624 -584 -1048
rect -504 -2624 -470 -1048
rect -346 -2624 -312 -1048
rect -232 -2624 -198 -1048
rect -74 -2624 -40 -1048
rect 40 -2624 74 -1048
rect 198 -2624 232 -1048
rect 312 -2624 346 -1048
rect 470 -2624 504 -1048
rect 584 -2624 618 -1048
rect 742 -2624 776 -1048
<< nsubdiff >>
rect -890 2785 -794 2819
rect 794 2785 890 2819
rect -890 2723 -856 2785
rect 856 2723 890 2785
rect -890 -2785 -856 -2723
rect 856 -2785 890 -2723
rect -890 -2819 -794 -2785
rect 794 -2819 890 -2785
<< nsubdiffcont >>
rect -794 2785 794 2819
rect -890 -2723 -856 2723
rect 856 -2723 890 2723
rect -794 -2819 794 -2785
<< poly >>
rect -730 2717 -630 2733
rect -730 2683 -714 2717
rect -646 2683 -630 2717
rect -730 2636 -630 2683
rect -458 2717 -358 2733
rect -458 2683 -442 2717
rect -374 2683 -358 2717
rect -458 2636 -358 2683
rect -186 2717 -86 2733
rect -186 2683 -170 2717
rect -102 2683 -86 2717
rect -186 2636 -86 2683
rect 86 2717 186 2733
rect 86 2683 102 2717
rect 170 2683 186 2717
rect 86 2636 186 2683
rect 358 2717 458 2733
rect 358 2683 374 2717
rect 442 2683 458 2717
rect 358 2636 458 2683
rect 630 2717 730 2733
rect 630 2683 646 2717
rect 714 2683 730 2717
rect 630 2636 730 2683
rect -730 989 -630 1036
rect -730 955 -714 989
rect -646 955 -630 989
rect -730 939 -630 955
rect -458 989 -358 1036
rect -458 955 -442 989
rect -374 955 -358 989
rect -458 939 -358 955
rect -186 989 -86 1036
rect -186 955 -170 989
rect -102 955 -86 989
rect -186 939 -86 955
rect 86 989 186 1036
rect 86 955 102 989
rect 170 955 186 989
rect 86 939 186 955
rect 358 989 458 1036
rect 358 955 374 989
rect 442 955 458 989
rect 358 939 458 955
rect 630 989 730 1036
rect 630 955 646 989
rect 714 955 730 989
rect 630 939 730 955
rect -730 881 -630 897
rect -730 847 -714 881
rect -646 847 -630 881
rect -730 800 -630 847
rect -458 881 -358 897
rect -458 847 -442 881
rect -374 847 -358 881
rect -458 800 -358 847
rect -186 881 -86 897
rect -186 847 -170 881
rect -102 847 -86 881
rect -186 800 -86 847
rect 86 881 186 897
rect 86 847 102 881
rect 170 847 186 881
rect 86 800 186 847
rect 358 881 458 897
rect 358 847 374 881
rect 442 847 458 881
rect 358 800 458 847
rect 630 881 730 897
rect 630 847 646 881
rect 714 847 730 881
rect 630 800 730 847
rect -730 -847 -630 -800
rect -730 -881 -714 -847
rect -646 -881 -630 -847
rect -730 -897 -630 -881
rect -458 -847 -358 -800
rect -458 -881 -442 -847
rect -374 -881 -358 -847
rect -458 -897 -358 -881
rect -186 -847 -86 -800
rect -186 -881 -170 -847
rect -102 -881 -86 -847
rect -186 -897 -86 -881
rect 86 -847 186 -800
rect 86 -881 102 -847
rect 170 -881 186 -847
rect 86 -897 186 -881
rect 358 -847 458 -800
rect 358 -881 374 -847
rect 442 -881 458 -847
rect 358 -897 458 -881
rect 630 -847 730 -800
rect 630 -881 646 -847
rect 714 -881 730 -847
rect 630 -897 730 -881
rect -730 -955 -630 -939
rect -730 -989 -714 -955
rect -646 -989 -630 -955
rect -730 -1036 -630 -989
rect -458 -955 -358 -939
rect -458 -989 -442 -955
rect -374 -989 -358 -955
rect -458 -1036 -358 -989
rect -186 -955 -86 -939
rect -186 -989 -170 -955
rect -102 -989 -86 -955
rect -186 -1036 -86 -989
rect 86 -955 186 -939
rect 86 -989 102 -955
rect 170 -989 186 -955
rect 86 -1036 186 -989
rect 358 -955 458 -939
rect 358 -989 374 -955
rect 442 -989 458 -955
rect 358 -1036 458 -989
rect 630 -955 730 -939
rect 630 -989 646 -955
rect 714 -989 730 -955
rect 630 -1036 730 -989
rect -730 -2683 -630 -2636
rect -730 -2717 -714 -2683
rect -646 -2717 -630 -2683
rect -730 -2733 -630 -2717
rect -458 -2683 -358 -2636
rect -458 -2717 -442 -2683
rect -374 -2717 -358 -2683
rect -458 -2733 -358 -2717
rect -186 -2683 -86 -2636
rect -186 -2717 -170 -2683
rect -102 -2717 -86 -2683
rect -186 -2733 -86 -2717
rect 86 -2683 186 -2636
rect 86 -2717 102 -2683
rect 170 -2717 186 -2683
rect 86 -2733 186 -2717
rect 358 -2683 458 -2636
rect 358 -2717 374 -2683
rect 442 -2717 458 -2683
rect 358 -2733 458 -2717
rect 630 -2683 730 -2636
rect 630 -2717 646 -2683
rect 714 -2717 730 -2683
rect 630 -2733 730 -2717
<< polycont >>
rect -714 2683 -646 2717
rect -442 2683 -374 2717
rect -170 2683 -102 2717
rect 102 2683 170 2717
rect 374 2683 442 2717
rect 646 2683 714 2717
rect -714 955 -646 989
rect -442 955 -374 989
rect -170 955 -102 989
rect 102 955 170 989
rect 374 955 442 989
rect 646 955 714 989
rect -714 847 -646 881
rect -442 847 -374 881
rect -170 847 -102 881
rect 102 847 170 881
rect 374 847 442 881
rect 646 847 714 881
rect -714 -881 -646 -847
rect -442 -881 -374 -847
rect -170 -881 -102 -847
rect 102 -881 170 -847
rect 374 -881 442 -847
rect 646 -881 714 -847
rect -714 -989 -646 -955
rect -442 -989 -374 -955
rect -170 -989 -102 -955
rect 102 -989 170 -955
rect 374 -989 442 -955
rect 646 -989 714 -955
rect -714 -2717 -646 -2683
rect -442 -2717 -374 -2683
rect -170 -2717 -102 -2683
rect 102 -2717 170 -2683
rect 374 -2717 442 -2683
rect 646 -2717 714 -2683
<< locali >>
rect -890 2785 -794 2819
rect 794 2785 890 2819
rect -890 2723 -856 2785
rect 856 2723 890 2785
rect -730 2683 -714 2717
rect -646 2683 -630 2717
rect -458 2683 -442 2717
rect -374 2683 -358 2717
rect -186 2683 -170 2717
rect -102 2683 -86 2717
rect 86 2683 102 2717
rect 170 2683 186 2717
rect 358 2683 374 2717
rect 442 2683 458 2717
rect 630 2683 646 2717
rect 714 2683 730 2717
rect -776 2624 -742 2640
rect -776 1032 -742 1048
rect -618 2624 -584 2640
rect -618 1032 -584 1048
rect -504 2624 -470 2640
rect -504 1032 -470 1048
rect -346 2624 -312 2640
rect -346 1032 -312 1048
rect -232 2624 -198 2640
rect -232 1032 -198 1048
rect -74 2624 -40 2640
rect -74 1032 -40 1048
rect 40 2624 74 2640
rect 40 1032 74 1048
rect 198 2624 232 2640
rect 198 1032 232 1048
rect 312 2624 346 2640
rect 312 1032 346 1048
rect 470 2624 504 2640
rect 470 1032 504 1048
rect 584 2624 618 2640
rect 584 1032 618 1048
rect 742 2624 776 2640
rect 742 1032 776 1048
rect -730 955 -714 989
rect -646 955 -630 989
rect -458 955 -442 989
rect -374 955 -358 989
rect -186 955 -170 989
rect -102 955 -86 989
rect 86 955 102 989
rect 170 955 186 989
rect 358 955 374 989
rect 442 955 458 989
rect 630 955 646 989
rect 714 955 730 989
rect -730 847 -714 881
rect -646 847 -630 881
rect -458 847 -442 881
rect -374 847 -358 881
rect -186 847 -170 881
rect -102 847 -86 881
rect 86 847 102 881
rect 170 847 186 881
rect 358 847 374 881
rect 442 847 458 881
rect 630 847 646 881
rect 714 847 730 881
rect -776 788 -742 804
rect -776 -804 -742 -788
rect -618 788 -584 804
rect -618 -804 -584 -788
rect -504 788 -470 804
rect -504 -804 -470 -788
rect -346 788 -312 804
rect -346 -804 -312 -788
rect -232 788 -198 804
rect -232 -804 -198 -788
rect -74 788 -40 804
rect -74 -804 -40 -788
rect 40 788 74 804
rect 40 -804 74 -788
rect 198 788 232 804
rect 198 -804 232 -788
rect 312 788 346 804
rect 312 -804 346 -788
rect 470 788 504 804
rect 470 -804 504 -788
rect 584 788 618 804
rect 584 -804 618 -788
rect 742 788 776 804
rect 742 -804 776 -788
rect -730 -881 -714 -847
rect -646 -881 -630 -847
rect -458 -881 -442 -847
rect -374 -881 -358 -847
rect -186 -881 -170 -847
rect -102 -881 -86 -847
rect 86 -881 102 -847
rect 170 -881 186 -847
rect 358 -881 374 -847
rect 442 -881 458 -847
rect 630 -881 646 -847
rect 714 -881 730 -847
rect -730 -989 -714 -955
rect -646 -989 -630 -955
rect -458 -989 -442 -955
rect -374 -989 -358 -955
rect -186 -989 -170 -955
rect -102 -989 -86 -955
rect 86 -989 102 -955
rect 170 -989 186 -955
rect 358 -989 374 -955
rect 442 -989 458 -955
rect 630 -989 646 -955
rect 714 -989 730 -955
rect -776 -1048 -742 -1032
rect -776 -2640 -742 -2624
rect -618 -1048 -584 -1032
rect -618 -2640 -584 -2624
rect -504 -1048 -470 -1032
rect -504 -2640 -470 -2624
rect -346 -1048 -312 -1032
rect -346 -2640 -312 -2624
rect -232 -1048 -198 -1032
rect -232 -2640 -198 -2624
rect -74 -1048 -40 -1032
rect -74 -2640 -40 -2624
rect 40 -1048 74 -1032
rect 40 -2640 74 -2624
rect 198 -1048 232 -1032
rect 198 -2640 232 -2624
rect 312 -1048 346 -1032
rect 312 -2640 346 -2624
rect 470 -1048 504 -1032
rect 470 -2640 504 -2624
rect 584 -1048 618 -1032
rect 584 -2640 618 -2624
rect 742 -1048 776 -1032
rect 742 -2640 776 -2624
rect -730 -2717 -714 -2683
rect -646 -2717 -630 -2683
rect -458 -2717 -442 -2683
rect -374 -2717 -358 -2683
rect -186 -2717 -170 -2683
rect -102 -2717 -86 -2683
rect 86 -2717 102 -2683
rect 170 -2717 186 -2683
rect 358 -2717 374 -2683
rect 442 -2717 458 -2683
rect 630 -2717 646 -2683
rect 714 -2717 730 -2683
rect -890 -2785 -856 -2723
rect 856 -2785 890 -2723
rect -890 -2819 -794 -2785
rect 794 -2819 890 -2785
<< viali >>
rect -714 2683 -646 2717
rect -442 2683 -374 2717
rect -170 2683 -102 2717
rect 102 2683 170 2717
rect 374 2683 442 2717
rect 646 2683 714 2717
rect -776 1048 -742 2624
rect -618 1048 -584 2624
rect -504 1048 -470 2624
rect -346 1048 -312 2624
rect -232 1048 -198 2624
rect -74 1048 -40 2624
rect 40 1048 74 2624
rect 198 1048 232 2624
rect 312 1048 346 2624
rect 470 1048 504 2624
rect 584 1048 618 2624
rect 742 1048 776 2624
rect -714 955 -646 989
rect -442 955 -374 989
rect -170 955 -102 989
rect 102 955 170 989
rect 374 955 442 989
rect 646 955 714 989
rect -714 847 -646 881
rect -442 847 -374 881
rect -170 847 -102 881
rect 102 847 170 881
rect 374 847 442 881
rect 646 847 714 881
rect -776 -788 -742 788
rect -618 -788 -584 788
rect -504 -788 -470 788
rect -346 -788 -312 788
rect -232 -788 -198 788
rect -74 -788 -40 788
rect 40 -788 74 788
rect 198 -788 232 788
rect 312 -788 346 788
rect 470 -788 504 788
rect 584 -788 618 788
rect 742 -788 776 788
rect -714 -881 -646 -847
rect -442 -881 -374 -847
rect -170 -881 -102 -847
rect 102 -881 170 -847
rect 374 -881 442 -847
rect 646 -881 714 -847
rect -714 -989 -646 -955
rect -442 -989 -374 -955
rect -170 -989 -102 -955
rect 102 -989 170 -955
rect 374 -989 442 -955
rect 646 -989 714 -955
rect -776 -2624 -742 -1048
rect -618 -2624 -584 -1048
rect -504 -2624 -470 -1048
rect -346 -2624 -312 -1048
rect -232 -2624 -198 -1048
rect -74 -2624 -40 -1048
rect 40 -2624 74 -1048
rect 198 -2624 232 -1048
rect 312 -2624 346 -1048
rect 470 -2624 504 -1048
rect 584 -2624 618 -1048
rect 742 -2624 776 -1048
rect -714 -2717 -646 -2683
rect -442 -2717 -374 -2683
rect -170 -2717 -102 -2683
rect 102 -2717 170 -2683
rect 374 -2717 442 -2683
rect 646 -2717 714 -2683
<< metal1 >>
rect -726 2717 -634 2723
rect -726 2683 -714 2717
rect -646 2683 -634 2717
rect -726 2677 -634 2683
rect -454 2717 -362 2723
rect -454 2683 -442 2717
rect -374 2683 -362 2717
rect -454 2677 -362 2683
rect -182 2717 -90 2723
rect -182 2683 -170 2717
rect -102 2683 -90 2717
rect -182 2677 -90 2683
rect 90 2717 182 2723
rect 90 2683 102 2717
rect 170 2683 182 2717
rect 90 2677 182 2683
rect 362 2717 454 2723
rect 362 2683 374 2717
rect 442 2683 454 2717
rect 362 2677 454 2683
rect 634 2717 726 2723
rect 634 2683 646 2717
rect 714 2683 726 2717
rect 634 2677 726 2683
rect -782 2624 -736 2636
rect -782 1048 -776 2624
rect -742 1048 -736 2624
rect -782 1036 -736 1048
rect -624 2624 -578 2636
rect -624 1048 -618 2624
rect -584 1048 -578 2624
rect -624 1036 -578 1048
rect -510 2624 -464 2636
rect -510 1048 -504 2624
rect -470 1048 -464 2624
rect -510 1036 -464 1048
rect -352 2624 -306 2636
rect -352 1048 -346 2624
rect -312 1048 -306 2624
rect -352 1036 -306 1048
rect -238 2624 -192 2636
rect -238 1048 -232 2624
rect -198 1048 -192 2624
rect -238 1036 -192 1048
rect -80 2624 -34 2636
rect -80 1048 -74 2624
rect -40 1048 -34 2624
rect -80 1036 -34 1048
rect 34 2624 80 2636
rect 34 1048 40 2624
rect 74 1048 80 2624
rect 34 1036 80 1048
rect 192 2624 238 2636
rect 192 1048 198 2624
rect 232 1048 238 2624
rect 192 1036 238 1048
rect 306 2624 352 2636
rect 306 1048 312 2624
rect 346 1048 352 2624
rect 306 1036 352 1048
rect 464 2624 510 2636
rect 464 1048 470 2624
rect 504 1048 510 2624
rect 464 1036 510 1048
rect 578 2624 624 2636
rect 578 1048 584 2624
rect 618 1048 624 2624
rect 578 1036 624 1048
rect 736 2624 782 2636
rect 736 1048 742 2624
rect 776 1048 782 2624
rect 736 1036 782 1048
rect -726 989 -634 995
rect -726 955 -714 989
rect -646 955 -634 989
rect -726 949 -634 955
rect -454 989 -362 995
rect -454 955 -442 989
rect -374 955 -362 989
rect -454 949 -362 955
rect -182 989 -90 995
rect -182 955 -170 989
rect -102 955 -90 989
rect -182 949 -90 955
rect 90 989 182 995
rect 90 955 102 989
rect 170 955 182 989
rect 90 949 182 955
rect 362 989 454 995
rect 362 955 374 989
rect 442 955 454 989
rect 362 949 454 955
rect 634 989 726 995
rect 634 955 646 989
rect 714 955 726 989
rect 634 949 726 955
rect -726 881 -634 887
rect -726 847 -714 881
rect -646 847 -634 881
rect -726 841 -634 847
rect -454 881 -362 887
rect -454 847 -442 881
rect -374 847 -362 881
rect -454 841 -362 847
rect -182 881 -90 887
rect -182 847 -170 881
rect -102 847 -90 881
rect -182 841 -90 847
rect 90 881 182 887
rect 90 847 102 881
rect 170 847 182 881
rect 90 841 182 847
rect 362 881 454 887
rect 362 847 374 881
rect 442 847 454 881
rect 362 841 454 847
rect 634 881 726 887
rect 634 847 646 881
rect 714 847 726 881
rect 634 841 726 847
rect -782 788 -736 800
rect -782 -788 -776 788
rect -742 -788 -736 788
rect -782 -800 -736 -788
rect -624 788 -578 800
rect -624 -788 -618 788
rect -584 -788 -578 788
rect -624 -800 -578 -788
rect -510 788 -464 800
rect -510 -788 -504 788
rect -470 -788 -464 788
rect -510 -800 -464 -788
rect -352 788 -306 800
rect -352 -788 -346 788
rect -312 -788 -306 788
rect -352 -800 -306 -788
rect -238 788 -192 800
rect -238 -788 -232 788
rect -198 -788 -192 788
rect -238 -800 -192 -788
rect -80 788 -34 800
rect -80 -788 -74 788
rect -40 -788 -34 788
rect -80 -800 -34 -788
rect 34 788 80 800
rect 34 -788 40 788
rect 74 -788 80 788
rect 34 -800 80 -788
rect 192 788 238 800
rect 192 -788 198 788
rect 232 -788 238 788
rect 192 -800 238 -788
rect 306 788 352 800
rect 306 -788 312 788
rect 346 -788 352 788
rect 306 -800 352 -788
rect 464 788 510 800
rect 464 -788 470 788
rect 504 -788 510 788
rect 464 -800 510 -788
rect 578 788 624 800
rect 578 -788 584 788
rect 618 -788 624 788
rect 578 -800 624 -788
rect 736 788 782 800
rect 736 -788 742 788
rect 776 -788 782 788
rect 736 -800 782 -788
rect -726 -847 -634 -841
rect -726 -881 -714 -847
rect -646 -881 -634 -847
rect -726 -887 -634 -881
rect -454 -847 -362 -841
rect -454 -881 -442 -847
rect -374 -881 -362 -847
rect -454 -887 -362 -881
rect -182 -847 -90 -841
rect -182 -881 -170 -847
rect -102 -881 -90 -847
rect -182 -887 -90 -881
rect 90 -847 182 -841
rect 90 -881 102 -847
rect 170 -881 182 -847
rect 90 -887 182 -881
rect 362 -847 454 -841
rect 362 -881 374 -847
rect 442 -881 454 -847
rect 362 -887 454 -881
rect 634 -847 726 -841
rect 634 -881 646 -847
rect 714 -881 726 -847
rect 634 -887 726 -881
rect -726 -955 -634 -949
rect -726 -989 -714 -955
rect -646 -989 -634 -955
rect -726 -995 -634 -989
rect -454 -955 -362 -949
rect -454 -989 -442 -955
rect -374 -989 -362 -955
rect -454 -995 -362 -989
rect -182 -955 -90 -949
rect -182 -989 -170 -955
rect -102 -989 -90 -955
rect -182 -995 -90 -989
rect 90 -955 182 -949
rect 90 -989 102 -955
rect 170 -989 182 -955
rect 90 -995 182 -989
rect 362 -955 454 -949
rect 362 -989 374 -955
rect 442 -989 454 -955
rect 362 -995 454 -989
rect 634 -955 726 -949
rect 634 -989 646 -955
rect 714 -989 726 -955
rect 634 -995 726 -989
rect -782 -1048 -736 -1036
rect -782 -2624 -776 -1048
rect -742 -2624 -736 -1048
rect -782 -2636 -736 -2624
rect -624 -1048 -578 -1036
rect -624 -2624 -618 -1048
rect -584 -2624 -578 -1048
rect -624 -2636 -578 -2624
rect -510 -1048 -464 -1036
rect -510 -2624 -504 -1048
rect -470 -2624 -464 -1048
rect -510 -2636 -464 -2624
rect -352 -1048 -306 -1036
rect -352 -2624 -346 -1048
rect -312 -2624 -306 -1048
rect -352 -2636 -306 -2624
rect -238 -1048 -192 -1036
rect -238 -2624 -232 -1048
rect -198 -2624 -192 -1048
rect -238 -2636 -192 -2624
rect -80 -1048 -34 -1036
rect -80 -2624 -74 -1048
rect -40 -2624 -34 -1048
rect -80 -2636 -34 -2624
rect 34 -1048 80 -1036
rect 34 -2624 40 -1048
rect 74 -2624 80 -1048
rect 34 -2636 80 -2624
rect 192 -1048 238 -1036
rect 192 -2624 198 -1048
rect 232 -2624 238 -1048
rect 192 -2636 238 -2624
rect 306 -1048 352 -1036
rect 306 -2624 312 -1048
rect 346 -2624 352 -1048
rect 306 -2636 352 -2624
rect 464 -1048 510 -1036
rect 464 -2624 470 -1048
rect 504 -2624 510 -1048
rect 464 -2636 510 -2624
rect 578 -1048 624 -1036
rect 578 -2624 584 -1048
rect 618 -2624 624 -1048
rect 578 -2636 624 -2624
rect 736 -1048 782 -1036
rect 736 -2624 742 -1048
rect 776 -2624 782 -1048
rect 736 -2636 782 -2624
rect -726 -2683 -634 -2677
rect -726 -2717 -714 -2683
rect -646 -2717 -634 -2683
rect -726 -2723 -634 -2717
rect -454 -2683 -362 -2677
rect -454 -2717 -442 -2683
rect -374 -2717 -362 -2683
rect -454 -2723 -362 -2717
rect -182 -2683 -90 -2677
rect -182 -2717 -170 -2683
rect -102 -2717 -90 -2683
rect -182 -2723 -90 -2717
rect 90 -2683 182 -2677
rect 90 -2717 102 -2683
rect 170 -2717 182 -2683
rect 90 -2723 182 -2717
rect 362 -2683 454 -2677
rect 362 -2717 374 -2683
rect 442 -2717 454 -2683
rect 362 -2723 454 -2717
rect 634 -2683 726 -2677
rect 634 -2717 646 -2683
rect 714 -2717 726 -2683
rect 634 -2723 726 -2717
<< properties >>
string FIXED_BBOX -873 -2802 873 2802
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 3 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
