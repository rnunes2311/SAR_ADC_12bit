magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect 721 878 779 884
rect -605 872 -547 878
rect -413 872 -355 878
rect -221 872 -163 878
rect -29 872 29 878
rect 163 872 221 878
rect 355 872 413 878
rect 547 872 605 878
rect -605 838 -593 872
rect -413 838 -401 872
rect -221 838 -209 872
rect -29 838 -17 872
rect 163 838 175 872
rect 355 838 367 872
rect 547 838 559 872
rect 721 844 733 878
rect 721 838 779 844
rect -605 832 -547 838
rect -413 832 -355 838
rect -221 832 -163 838
rect -29 832 29 838
rect 163 832 221 838
rect 355 832 413 838
rect 547 832 605 838
<< pwell >>
rect -887 -940 6957 1030
<< nmos >>
rect -687 -800 -657 800
rect -591 -800 -561 800
rect -495 -800 -465 800
rect -399 -800 -369 800
rect -303 -800 -273 800
rect -207 -800 -177 800
rect -111 -800 -81 800
rect -15 -800 15 800
rect 81 -800 111 800
rect 177 -800 207 800
rect 273 -800 303 800
rect 369 -800 399 800
rect 465 -800 495 800
rect 561 -800 591 800
rect 657 -800 687 800
<< ndiff >>
rect -749 788 -687 800
rect -749 -788 -737 788
rect -703 -788 -687 788
rect -749 -800 -687 -788
rect -657 788 -591 800
rect -657 -788 -641 788
rect -607 -788 -591 788
rect -657 -800 -591 -788
rect -561 788 -495 800
rect -561 -788 -545 788
rect -511 -788 -495 788
rect -561 -800 -495 -788
rect -465 788 -399 800
rect -465 -788 -449 788
rect -415 -788 -399 788
rect -465 -800 -399 -788
rect -369 788 -303 800
rect -369 -788 -353 788
rect -319 -788 -303 788
rect -369 -800 -303 -788
rect -273 788 -207 800
rect -273 -788 -257 788
rect -223 -788 -207 788
rect -273 -800 -207 -788
rect -177 788 -111 800
rect -177 -788 -161 788
rect -127 -788 -111 788
rect -177 -800 -111 -788
rect -81 788 -15 800
rect -81 -788 -65 788
rect -31 -788 -15 788
rect -81 -800 -15 -788
rect 15 788 81 800
rect 15 -788 31 788
rect 65 -788 81 788
rect 15 -800 81 -788
rect 111 788 177 800
rect 111 -788 127 788
rect 161 -788 177 788
rect 111 -800 177 -788
rect 207 788 273 800
rect 207 -788 223 788
rect 257 -788 273 788
rect 207 -800 273 -788
rect 303 788 369 800
rect 303 -788 319 788
rect 353 -788 369 788
rect 303 -800 369 -788
rect 399 788 465 800
rect 399 -788 415 788
rect 449 -788 465 788
rect 399 -800 465 -788
rect 495 788 561 800
rect 495 -788 511 788
rect 545 -788 561 788
rect 495 -800 561 -788
rect 591 788 657 800
rect 591 -788 607 788
rect 641 -788 657 788
rect 591 -800 657 -788
rect 687 788 749 800
rect 687 -788 703 788
rect 737 -788 749 788
rect 687 -800 749 -788
<< ndiffc >>
rect -737 -788 -703 788
rect -641 -788 -607 788
rect -545 -788 -511 788
rect -449 -788 -415 788
rect -353 -788 -319 788
rect -257 -788 -223 788
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
rect 223 -788 257 788
rect 319 -788 353 788
rect 415 -788 449 788
rect 511 -788 545 788
rect 607 -788 641 788
rect 703 -788 737 788
<< psubdiff >>
rect -851 960 -755 994
rect 6855 960 6921 994
rect -851 878 -817 960
rect 6887 878 6921 960
rect -851 -870 -817 -812
rect 6887 -870 6921 -812
rect -851 -904 -755 -870
rect 6855 -904 6921 -870
<< psubdiffcont >>
rect -755 960 6855 994
rect -851 -812 -817 878
rect 6887 -812 6921 878
rect -755 -904 6855 -870
<< poly >>
rect -609 878 -543 888
rect -417 878 -351 888
rect -225 878 -159 888
rect -33 878 33 888
rect 159 878 225 888
rect 351 878 417 888
rect 543 878 609 888
rect 717 878 783 894
rect -687 872 33 878
rect -687 838 -593 872
rect -559 838 -401 872
rect -367 838 -209 872
rect -175 838 -17 872
rect 17 838 33 872
rect -687 828 33 838
rect -687 800 -657 828
rect -609 822 -543 828
rect -591 800 -561 822
rect -495 800 -465 828
rect -417 822 -351 828
rect -399 800 -369 822
rect -303 800 -273 828
rect -225 822 -159 828
rect -207 800 -177 822
rect -111 800 -81 828
rect -33 822 33 828
rect 81 872 417 878
rect 81 838 175 872
rect 209 838 367 872
rect 401 838 417 872
rect 81 828 417 838
rect -15 800 15 822
rect 81 800 111 828
rect 159 822 225 828
rect 177 800 207 822
rect 273 800 303 828
rect 351 822 417 828
rect 465 872 609 878
rect 465 838 559 872
rect 593 838 609 872
rect 465 828 609 838
rect 369 800 399 822
rect 465 800 495 828
rect 543 822 609 828
rect 657 844 733 878
rect 767 844 783 878
rect 657 828 783 844
rect 561 800 591 822
rect 657 800 687 828
rect -687 -826 -657 -800
rect -591 -826 -561 -800
rect -495 -826 -465 -800
rect -399 -826 -369 -800
rect -303 -826 -273 -800
rect -207 -826 -177 -800
rect -111 -826 -81 -800
rect -15 -826 15 -800
rect 81 -826 111 -800
rect 177 -826 207 -800
rect 273 -826 303 -800
rect 369 -826 399 -800
rect 465 -826 495 -800
rect 561 -826 591 -800
rect 657 -826 687 -800
<< polycont >>
rect -593 838 -559 872
rect -401 838 -367 872
rect -209 838 -175 872
rect -17 838 17 872
rect 175 838 209 872
rect 367 838 401 872
rect 559 838 593 872
rect 733 844 767 878
<< locali >>
rect -851 960 -755 994
rect 6855 960 6921 994
rect -851 878 -817 960
rect 6887 878 6921 960
rect -609 838 -593 872
rect -559 838 -543 872
rect -417 838 -401 872
rect -367 838 -351 872
rect -225 838 -209 872
rect -175 838 -159 872
rect -33 838 -17 872
rect 17 838 33 872
rect 159 838 175 872
rect 209 838 225 872
rect 351 838 367 872
rect 401 838 417 872
rect 543 838 559 872
rect 593 838 609 872
rect 717 844 733 878
rect 767 844 783 878
rect -737 788 -703 804
rect -737 -804 -703 -788
rect -641 788 -607 804
rect -641 -804 -607 -788
rect -545 788 -511 804
rect -545 -804 -511 -788
rect -449 788 -415 804
rect -449 -804 -415 -788
rect -353 788 -319 804
rect -353 -804 -319 -788
rect -257 788 -223 804
rect -257 -804 -223 -788
rect -161 788 -127 804
rect -161 -804 -127 -788
rect -65 788 -31 804
rect -65 -804 -31 -788
rect 31 788 65 804
rect 31 -804 65 -788
rect 127 788 161 804
rect 127 -804 161 -788
rect 223 788 257 804
rect 223 -804 257 -788
rect 319 788 353 804
rect 319 -804 353 -788
rect 415 788 449 804
rect 415 -804 449 -788
rect 511 788 545 804
rect 511 -804 545 -788
rect 607 788 641 804
rect 607 -804 641 -788
rect 703 788 737 804
rect 703 -804 737 -788
rect -851 -870 -817 -812
rect 6887 -870 6921 -812
rect -851 -904 -755 -870
rect 6855 -904 6921 -870
<< viali >>
rect -593 838 -559 872
rect -401 838 -367 872
rect -209 838 -175 872
rect -17 838 17 872
rect 175 838 209 872
rect 367 838 401 872
rect 559 838 593 872
rect 733 844 767 878
rect -737 -788 -703 788
rect -641 -788 -607 788
rect -545 -788 -511 788
rect -449 -788 -415 788
rect -353 -788 -319 788
rect -257 -788 -223 788
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
rect 223 -788 257 788
rect 319 -788 353 788
rect 415 -788 449 788
rect 511 -788 545 788
rect 607 -788 641 788
rect 703 -788 737 788
<< metal1 >>
rect 721 878 779 884
rect -605 872 -547 878
rect -605 838 -593 872
rect -559 838 -547 872
rect -605 832 -547 838
rect -413 872 -355 878
rect -413 838 -401 872
rect -367 838 -355 872
rect -413 832 -355 838
rect -221 872 -163 878
rect -221 838 -209 872
rect -175 838 -163 872
rect -221 832 -163 838
rect -29 872 29 878
rect -29 838 -17 872
rect 17 838 29 872
rect -29 832 29 838
rect 163 872 221 878
rect 163 838 175 872
rect 209 838 221 872
rect 163 832 221 838
rect 355 872 413 878
rect 355 838 367 872
rect 401 838 413 872
rect 355 832 413 838
rect 547 872 605 878
rect 547 838 559 872
rect 593 838 605 872
rect 721 844 733 878
rect 767 844 779 878
rect 721 838 779 844
rect 547 832 605 838
rect -743 788 -697 800
rect -743 -788 -737 788
rect -703 -788 -697 788
rect -743 -800 -697 -788
rect -647 788 -601 800
rect -647 -788 -641 788
rect -607 -788 -601 788
rect -647 -800 -601 -788
rect -551 788 -505 800
rect -551 -788 -545 788
rect -511 -788 -505 788
rect -551 -800 -505 -788
rect -455 788 -409 800
rect -455 -788 -449 788
rect -415 -788 -409 788
rect -455 -800 -409 -788
rect -359 788 -313 800
rect -359 -788 -353 788
rect -319 -788 -313 788
rect -359 -800 -313 -788
rect -263 788 -217 800
rect -263 -788 -257 788
rect -223 -788 -217 788
rect -263 -800 -217 -788
rect -167 788 -121 800
rect -167 -788 -161 788
rect -127 -788 -121 788
rect -167 -800 -121 -788
rect -71 788 -25 800
rect -71 -788 -65 788
rect -31 -788 -25 788
rect -71 -800 -25 -788
rect 25 788 71 800
rect 25 -788 31 788
rect 65 -788 71 788
rect 25 -800 71 -788
rect 121 788 167 800
rect 121 -788 127 788
rect 161 -788 167 788
rect 121 -800 167 -788
rect 217 788 263 800
rect 217 -788 223 788
rect 257 -788 263 788
rect 217 -800 263 -788
rect 313 788 359 800
rect 313 -788 319 788
rect 353 -788 359 788
rect 313 -800 359 -788
rect 409 788 455 800
rect 409 -788 415 788
rect 449 -788 455 788
rect 409 -800 455 -788
rect 505 788 551 800
rect 505 -788 511 788
rect 545 -788 551 788
rect 505 -800 551 -788
rect 601 788 647 800
rect 601 -788 607 788
rect 641 -788 647 788
rect 601 -800 647 -788
rect 697 788 743 800
rect 697 -788 703 788
rect 737 -788 743 788
rect 697 -800 743 -788
<< properties >>
string FIXED_BBOX -834 -957 834 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.150 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
