magic
tech sky130A
magscale 1 2
timestamp 1714331631
<< metal1 >>
rect 13740 48110 13750 48170
rect 13810 48158 13820 48170
rect 13810 48130 24074 48158
rect 13810 48110 13820 48130
rect -3925 48060 -3865 48070
rect -3925 47990 -3865 48000
rect -4005 47800 -3945 47810
rect -4005 47730 -3945 47740
rect -4075 47530 -4015 47540
rect -4075 47460 -4015 47470
rect -4135 47250 -4075 47260
rect -4135 47180 -4075 47190
rect -4195 46980 -4135 46990
rect -4195 46910 -4135 46920
rect -4255 46700 -4195 46710
rect -4255 46630 -4195 46640
rect -4315 46440 -4255 46450
rect -4315 46370 -4255 46380
rect -4375 46170 -4315 46180
rect -4375 46100 -4315 46110
rect -4435 45890 -4375 45900
rect -4435 45820 -4375 45830
rect -4495 45620 -4435 45630
rect -4495 45550 -4435 45560
rect -4555 45360 -4495 45370
rect -4555 45290 -4495 45300
rect -4615 45080 -4555 45090
rect -4615 45010 -4555 45020
rect -4675 44810 -4615 44820
rect -4675 44740 -4615 44750
rect -4735 44530 -4675 44540
rect -4735 44460 -4675 44470
rect -4795 44270 -4735 44280
rect -4795 44200 -4735 44210
rect -4855 44000 -4795 44010
rect -4855 43930 -4795 43940
rect -4915 43730 -4855 43740
rect -4915 43660 -4855 43670
rect -4975 43440 -4915 43450
rect -4975 43370 -4915 43380
rect -5035 43170 -4975 43180
rect -5035 43100 -4975 43110
rect -5095 42910 -5035 42920
rect -5095 42840 -5035 42850
rect -5155 42620 -5095 42630
rect -5155 42550 -5095 42560
rect -5215 42350 -5155 42360
rect -5215 42280 -5155 42290
rect -5275 42070 -5215 42080
rect -5275 42000 -5215 42010
rect -5245 41408 -5215 42000
rect -5185 41408 -5155 42280
rect -5125 41408 -5095 42550
rect -5065 41408 -5035 42840
rect -5005 41408 -4975 43100
rect -4945 41408 -4915 43370
rect -4885 41408 -4855 43660
rect -4825 41408 -4795 43930
rect -4765 41408 -4735 44200
rect -4705 41408 -4675 44460
rect -4645 41408 -4615 44740
rect -4585 41408 -4555 45010
rect -4525 41408 -4495 45290
rect -4465 41408 -4435 45550
rect -4405 41408 -4375 45820
rect -4345 41408 -4315 46100
rect -4285 41408 -4255 46370
rect -4225 41408 -4195 46630
rect -4165 41408 -4135 46910
rect -4105 41408 -4075 47180
rect -4045 41408 -4015 47460
rect -3985 41408 -3955 47730
rect -3895 41435 -3865 47990
rect 16130 41675 16140 41700
rect -1350 41590 -1340 41650
rect -1280 41625 -1270 41650
rect 15440 41645 16140 41675
rect -1280 41595 -560 41625
rect -1280 41590 -1270 41595
rect -3190 41530 -3180 41590
rect -3120 41530 -3110 41590
rect -2270 41530 -2260 41590
rect -2200 41555 -2190 41590
rect -2200 41530 -622 41555
rect -3160 41495 -3130 41530
rect -2245 41525 -622 41530
rect -3160 41465 -695 41495
rect -3895 41405 -755 41435
rect -785 36645 -755 41405
rect -3775 36615 -755 36645
rect -5245 35961 -5215 36092
rect -5185 35914 -5155 36117
rect -5125 35944 -5095 36112
rect -5065 35933 -5035 36114
rect -5005 35955 -4975 36110
rect -4945 35945 -4915 36111
rect -4885 35956 -4855 36133
rect -4825 35959 -4795 36110
rect -4765 35939 -4735 36135
rect -4705 35929 -4675 36109
rect -4645 35935 -4615 36104
rect -4585 35946 -4555 36106
rect -4525 35926 -4495 36106
rect -4465 35926 -4435 36108
rect -4405 35943 -4375 36100
rect -4345 35939 -4315 36098
rect -4285 35948 -4255 36108
rect -4225 35934 -4195 36129
rect -4165 35938 -4135 36112
rect -4105 35940 -4075 36109
rect -4045 35940 -4015 36114
rect -3985 35949 -3955 36089
rect -3775 36075 -3745 36615
rect -725 36585 -695 41465
rect -652 38746 -622 41525
rect -590 39830 -560 41595
rect 15210 41410 15220 41470
rect 15280 41435 15290 41470
rect 15280 41410 15410 41435
rect 15235 41405 15410 41410
rect 13360 41330 13370 41390
rect 13430 41375 13440 41390
rect 13430 41345 15350 41375
rect 13430 41330 13440 41345
rect 490 41240 500 41300
rect 560 41285 570 41300
rect 560 41255 15290 41285
rect 560 41240 570 41255
rect 2320 41150 2330 41210
rect 2390 41195 2400 41210
rect 2390 41165 15230 41195
rect 2390 41150 2400 41165
rect 10610 41105 10620 41120
rect 185 41075 10620 41105
rect -590 39770 -580 39830
rect -520 39770 -510 39830
rect -667 38736 -607 38746
rect -667 38676 -662 38736
rect -667 38666 -607 38676
rect -3895 36045 -3745 36075
rect -3715 36555 95 36585
rect -3895 35935 -3865 36045
rect -3715 36015 -3685 36555
rect 65 36265 95 36555
rect 185 36490 215 41075
rect 10610 41060 10620 41075
rect 10680 41060 10690 41120
rect 15080 41040 15090 41100
rect 15150 41040 15160 41100
rect 8770 41015 8780 41030
rect 245 40985 8780 41015
rect 245 36550 275 40985
rect 8770 40970 8780 40985
rect 8840 40970 8850 41030
rect 6930 40925 6940 40940
rect 305 40895 6940 40925
rect 305 36610 335 40895
rect 6930 40880 6940 40895
rect 7000 40880 7010 40940
rect 14990 40835 15000 40850
rect 365 40805 15000 40835
rect 365 36670 395 40805
rect 14990 40790 15000 40805
rect 15060 40790 15070 40850
rect 5080 40745 5090 40750
rect 425 40715 5090 40745
rect 425 36730 455 40715
rect 5080 40690 5090 40715
rect 5150 40690 5160 40750
rect 14700 40745 14710 40760
rect 9125 40715 14710 40745
rect 4170 40655 4180 40660
rect 485 40625 4180 40655
rect 485 36790 515 40625
rect 4170 40600 4180 40625
rect 4240 40600 4250 40660
rect 9125 40565 9155 40715
rect 14700 40700 14710 40715
rect 14770 40700 14780 40760
rect 2545 40535 9155 40565
rect 2545 40485 2575 40535
rect 690 40455 2575 40485
rect 545 39760 555 39820
rect 615 39760 625 39820
rect 550 36915 580 39760
rect 690 38740 720 40455
rect 9250 40340 9260 40680
rect 9630 40340 9640 40680
rect 1530 40170 1540 40270
rect 1910 40170 1920 40270
rect 670 38680 680 38740
rect 740 38680 750 38740
rect 3400 38020 3410 38080
rect 3470 38020 3480 38080
rect 14830 38020 14860 38030
rect 3420 37670 3460 38020
rect 14800 37960 14810 38020
rect 14870 38005 14880 38020
rect 15120 38005 15150 41040
rect 14870 37975 15150 38005
rect 14870 37960 14880 37975
rect 3400 37610 3410 37670
rect 3470 37610 3480 37670
rect 1960 37330 2300 37510
rect 1950 36990 1960 37330
rect 2300 36990 2310 37330
rect 7400 36990 7410 37330
rect 7750 36990 7760 37330
rect 15070 36915 15080 36940
rect 550 36885 15080 36915
rect 15070 36880 15080 36885
rect 15140 36880 15150 36940
rect 15200 36850 15230 41165
rect 10095 36840 15230 36850
rect 485 36780 10035 36790
rect 485 36760 9975 36780
rect 425 36720 9945 36730
rect 425 36700 9885 36720
rect 365 36660 9855 36670
rect 365 36640 9795 36660
rect 305 36600 9765 36610
rect 305 36580 9705 36600
rect 245 36540 9675 36550
rect 245 36520 9615 36540
rect 185 36480 9585 36490
rect 185 36460 9525 36480
rect 10155 36820 15230 36840
rect 15260 36790 15290 41255
rect 10095 36770 10155 36780
rect 10185 36780 15290 36790
rect 9975 36710 10035 36720
rect 10245 36760 15290 36780
rect 15320 36730 15350 41345
rect 10185 36710 10245 36720
rect 10275 36720 15350 36730
rect 9885 36650 9945 36660
rect 10335 36700 15350 36720
rect 15380 36670 15410 41405
rect 10275 36650 10335 36660
rect 10365 36660 15410 36670
rect 9795 36590 9855 36600
rect 10425 36640 15410 36660
rect 15440 36610 15470 41645
rect 16130 41640 16140 41645
rect 16200 41640 16210 41700
rect 17970 41605 17980 41630
rect 10365 36590 10425 36600
rect 10455 36600 15470 36610
rect 9705 36530 9765 36540
rect 10515 36580 15470 36600
rect 15500 41575 17980 41605
rect 15500 36550 15530 41575
rect 17970 41570 17980 41575
rect 18040 41570 18050 41630
rect 20730 41535 20740 41560
rect 10455 36530 10515 36540
rect 10545 36540 15530 36550
rect 9615 36470 9675 36480
rect 10605 36520 15530 36540
rect 15560 41505 20740 41535
rect 15560 36490 15590 41505
rect 20730 41500 20740 41505
rect 20800 41500 20810 41560
rect 19810 41445 19820 41470
rect 15620 41415 19820 41445
rect 15620 40860 15650 41415
rect 19810 41410 19820 41415
rect 19880 41410 19890 41470
rect 22570 41410 22580 41470
rect 22640 41460 22650 41470
rect 23190 41460 23200 41470
rect 22640 41430 23200 41460
rect 22640 41410 22650 41430
rect 23190 41410 23200 41430
rect 23260 41410 23270 41470
rect 23630 41380 23640 41410
rect 15715 41350 23640 41380
rect 23700 41350 23710 41410
rect 15620 40850 15680 40860
rect 15620 40780 15680 40790
rect 15715 40770 15745 41350
rect 24046 41315 24074 48130
rect 24152 48070 24212 48080
rect 24152 48000 24212 48010
rect 15790 41285 24075 41315
rect 15790 41110 15820 41285
rect 17070 41150 17080 41240
rect 17450 41150 17460 41240
rect 15780 41100 15840 41110
rect 22470 41080 22480 41230
rect 23040 41080 23050 41230
rect 23180 41040 23190 41100
rect 23250 41040 23260 41100
rect 23510 41040 23520 41100
rect 23580 41085 23590 41100
rect 23580 41040 23591 41085
rect 23630 41040 23640 41100
rect 23700 41040 23710 41100
rect 15780 41030 15840 41040
rect 23210 40900 23240 41040
rect 15710 40760 15770 40770
rect 15710 40690 15770 40700
rect 23561 39255 23591 41040
rect 23650 40390 23680 41040
rect 24065 41020 24095 41025
rect 24040 40960 24050 41020
rect 24110 40960 24120 41020
rect 23620 40330 23630 40390
rect 23690 40330 23700 40390
rect 15760 38894 15770 38954
rect 15830 38894 15840 38954
rect 15670 38004 15680 38064
rect 15740 38004 15750 38064
rect 15700 37880 15730 38004
rect 15670 37820 15680 37880
rect 15740 37820 15750 37880
rect 15790 37750 15820 38894
rect 15740 37690 15750 37750
rect 15810 37690 15820 37750
rect 10545 36470 10605 36480
rect 10635 36480 15590 36490
rect 9525 36410 9585 36420
rect 10695 36460 15590 36480
rect 10635 36410 10695 36420
rect 15070 36330 15080 36390
rect 15140 36380 15150 36390
rect 24075 36380 24105 40960
rect 15140 36350 24105 36380
rect 15140 36330 15150 36350
rect 65 36235 22455 36265
rect -3805 35985 -3685 36015
rect -3805 35295 -3775 35985
rect 22425 35295 22455 36235
rect 24152 35942 24182 48000
rect 24232 47810 24292 47820
rect 24232 47740 24292 47750
rect 24242 35935 24272 47740
rect 24302 47540 24362 47550
rect 24302 47470 24362 47480
rect 24302 35925 24332 47470
rect 24362 47260 24422 47270
rect 24362 47190 24422 47200
rect 24362 35925 24392 47190
rect 24422 46990 24482 47000
rect 24422 46920 24482 46930
rect 24422 35945 24452 46920
rect 24482 46710 24542 46720
rect 24482 46640 24542 46650
rect 24482 35915 24512 46640
rect 24542 46450 24602 46460
rect 24542 46380 24602 46390
rect 24542 35945 24572 46380
rect 24602 46180 24662 46190
rect 24602 46110 24662 46120
rect 24602 35935 24632 46110
rect 24662 45900 24722 45910
rect 24662 45830 24722 45840
rect 24662 35925 24692 45830
rect 24722 45630 24782 45640
rect 24722 45560 24782 45570
rect 24722 35945 24752 45560
rect 24782 45370 24842 45380
rect 24782 45300 24842 45310
rect 24782 35915 24812 45300
rect 24842 45090 24902 45100
rect 24842 45020 24902 45030
rect 24842 35915 24872 45020
rect 24902 44820 24962 44830
rect 24902 44750 24962 44760
rect 24902 35925 24932 44750
rect 24962 44540 25022 44550
rect 24962 44470 25022 44480
rect 24962 35925 24992 44470
rect 25022 44280 25082 44290
rect 25022 44210 25082 44220
rect 25022 35945 25052 44210
rect 25082 44010 25142 44020
rect 25082 43940 25142 43950
rect 25082 35945 25112 43940
rect 25142 43740 25202 43750
rect 25142 43670 25202 43680
rect 25142 35915 25172 43670
rect 25202 43450 25262 43460
rect 25202 43380 25262 43390
rect 25202 35935 25232 43380
rect 25262 43180 25322 43190
rect 25262 43110 25322 43120
rect 25262 35962 25292 43110
rect 25322 42920 25382 42930
rect 25322 42850 25382 42860
rect 25322 35945 25352 42850
rect 25382 42630 25442 42640
rect 25382 42560 25442 42570
rect 25382 35945 25412 42560
rect 25442 42360 25502 42370
rect 25442 42290 25502 42300
rect 25442 35905 25472 42290
rect 25502 42080 25562 42090
rect 25502 42010 25562 42020
rect 25502 35915 25532 42010
rect -3805 35265 -1965 35295
rect 22265 35265 22455 35295
rect 10610 33890 10620 33950
rect 10680 33890 10690 33950
rect 10520 33800 10530 33860
rect 10590 33800 10600 33860
rect 10430 33710 10440 33770
rect 10500 33710 10510 33770
rect 10340 33620 10350 33680
rect 10410 33620 10420 33680
rect 10250 33530 10260 33590
rect 10320 33530 10330 33590
rect 10160 33440 10170 33500
rect 10230 33440 10240 33500
rect 10070 33350 10080 33410
rect 10140 33350 10150 33410
rect 9980 33260 9990 33320
rect 10050 33260 10060 33320
rect 9890 33170 9900 33230
rect 9960 33170 9970 33230
rect 9800 33080 9810 33140
rect 9870 33080 9880 33140
rect 9710 32990 9720 33050
rect 9780 32990 9790 33050
rect 9620 32900 9630 32960
rect 9690 32900 9700 32960
rect 9530 32810 9540 32870
rect 9600 32810 9610 32870
<< via1 >>
rect 13750 48110 13810 48170
rect -3925 48000 -3865 48060
rect -4005 47740 -3945 47800
rect -4075 47470 -4015 47530
rect -4135 47190 -4075 47250
rect -4195 46920 -4135 46980
rect -4255 46640 -4195 46700
rect -4315 46380 -4255 46440
rect -4375 46110 -4315 46170
rect -4435 45830 -4375 45890
rect -4495 45560 -4435 45620
rect -4555 45300 -4495 45360
rect -4615 45020 -4555 45080
rect -4675 44750 -4615 44810
rect -4735 44470 -4675 44530
rect -4795 44210 -4735 44270
rect -4855 43940 -4795 44000
rect -4915 43670 -4855 43730
rect -4975 43380 -4915 43440
rect -5035 43110 -4975 43170
rect -5095 42850 -5035 42910
rect -5155 42560 -5095 42620
rect -5215 42290 -5155 42350
rect -5275 42010 -5215 42070
rect -1340 41590 -1280 41650
rect -3180 41530 -3120 41590
rect -2260 41530 -2200 41590
rect 15220 41410 15280 41470
rect 13370 41330 13430 41390
rect 500 41240 560 41300
rect 2330 41150 2390 41210
rect -580 39770 -520 39830
rect -662 38676 -607 38736
rect 10620 41060 10680 41120
rect 15090 41040 15150 41100
rect 8780 40970 8840 41030
rect 6940 40880 7000 40940
rect 15000 40790 15060 40850
rect 5090 40690 5150 40750
rect 4180 40600 4240 40660
rect 14710 40700 14770 40760
rect 555 39760 615 39820
rect 9260 40340 9630 40680
rect 1540 40170 1910 40270
rect 680 38680 740 38740
rect 3410 38020 3470 38080
rect 14810 37960 14870 38020
rect 3410 37610 3470 37670
rect 1960 36990 2300 37330
rect 7410 36990 7750 37330
rect 15080 36880 15140 36940
rect 9525 36420 9585 36480
rect 9615 36480 9675 36540
rect 9705 36540 9765 36600
rect 9795 36600 9855 36660
rect 9885 36660 9945 36720
rect 9975 36720 10035 36780
rect 10095 36780 10155 36840
rect 10185 36720 10245 36780
rect 10275 36660 10335 36720
rect 10365 36600 10425 36660
rect 16140 41640 16200 41700
rect 10455 36540 10515 36600
rect 17980 41570 18040 41630
rect 10545 36480 10605 36540
rect 20740 41500 20800 41560
rect 19820 41410 19880 41470
rect 22580 41410 22640 41470
rect 23200 41410 23260 41470
rect 23640 41350 23700 41410
rect 15620 40790 15680 40850
rect 24152 48010 24212 48070
rect 17080 41150 17450 41240
rect 15780 41040 15840 41100
rect 22480 41080 23040 41230
rect 23190 41040 23250 41100
rect 23520 41040 23580 41100
rect 23640 41040 23700 41100
rect 15710 40700 15770 40760
rect 24050 40960 24110 41020
rect 23630 40330 23690 40390
rect 15770 38894 15830 38954
rect 15680 38004 15740 38064
rect 15680 37820 15740 37880
rect 15750 37690 15810 37750
rect 10635 36420 10695 36480
rect 15080 36330 15140 36390
rect 24232 47750 24292 47810
rect 24302 47480 24362 47540
rect 24362 47200 24422 47260
rect 24422 46930 24482 46990
rect 24482 46650 24542 46710
rect 24542 46390 24602 46450
rect 24602 46120 24662 46180
rect 24662 45840 24722 45900
rect 24722 45570 24782 45630
rect 24782 45310 24842 45370
rect 24842 45030 24902 45090
rect 24902 44760 24962 44820
rect 24962 44480 25022 44540
rect 25022 44220 25082 44280
rect 25082 43950 25142 44010
rect 25142 43680 25202 43740
rect 25202 43390 25262 43450
rect 25262 43120 25322 43180
rect 25322 42860 25382 42920
rect 25382 42570 25442 42630
rect 25442 42300 25502 42360
rect 25502 42020 25562 42080
rect 10620 33890 10680 33950
rect 10530 33800 10590 33860
rect 10440 33710 10500 33770
rect 10350 33620 10410 33680
rect 10260 33530 10320 33590
rect 10170 33440 10230 33500
rect 10080 33350 10140 33410
rect 9990 33260 10050 33320
rect 9900 33170 9960 33230
rect 9810 33080 9870 33140
rect 9720 32990 9780 33050
rect 9630 32900 9690 32960
rect 9540 32810 9600 32870
<< metal2 >>
rect -3540 48070 -3480 48080
rect -3925 48060 -3865 48070
rect -3865 48010 -3540 48040
rect -2990 48010 -2940 48190
rect -600 48010 -550 48190
rect 1790 48010 1840 48190
rect 4190 48010 4240 48190
rect 6580 48010 6630 48190
rect 8970 48010 9020 48190
rect 11360 48010 11410 48190
rect 13750 48170 13810 48180
rect 13750 48100 13810 48110
rect -3540 48000 -3480 48010
rect -3925 47990 -3865 48000
rect 13750 47880 13806 48100
rect 16140 48010 16190 48190
rect 18540 48010 18590 48190
rect 20930 48010 20980 48190
rect 23320 48010 23370 48190
rect 24152 48070 24212 48080
rect 23950 48060 24010 48070
rect 24010 48020 24152 48050
rect 24152 48000 24212 48010
rect 23950 47990 24010 48000
rect 24232 47810 24292 47820
rect -4005 47800 -3945 47810
rect -3540 47790 -3480 47800
rect -3945 47750 -3540 47780
rect -4005 47730 -3945 47740
rect -3540 47720 -3480 47730
rect 23950 47790 24010 47800
rect 24010 47760 24232 47790
rect 24232 47740 24292 47750
rect 23950 47720 24010 47730
rect 24302 47540 24362 47550
rect -4075 47530 -4015 47540
rect -3540 47530 -3480 47540
rect -4015 47480 -3540 47510
rect -4075 47460 -4015 47470
rect -3540 47460 -3480 47470
rect 23950 47520 24010 47530
rect 24010 47490 24302 47520
rect 24302 47470 24362 47480
rect 23950 47450 24010 47460
rect 24362 47260 24422 47270
rect -4135 47250 -4075 47260
rect -3540 47250 -3480 47260
rect -4075 47200 -3540 47230
rect -4135 47180 -4075 47190
rect -3540 47180 -3480 47190
rect 23950 47250 24010 47260
rect 24010 47210 24362 47240
rect 24362 47190 24422 47200
rect 23950 47180 24010 47190
rect 24422 46990 24482 47000
rect -4195 46980 -4135 46990
rect -3550 46980 -3490 46990
rect -4135 46930 -3550 46960
rect -4195 46910 -4135 46920
rect -3550 46910 -3490 46920
rect 23950 46970 24010 46980
rect 24010 46940 24422 46970
rect 24422 46920 24482 46930
rect 23950 46900 24010 46910
rect -3550 46710 -3490 46720
rect -4255 46700 -4195 46710
rect -4195 46650 -3550 46680
rect 24482 46710 24542 46720
rect -3550 46640 -3490 46650
rect 23950 46690 24010 46700
rect -4255 46630 -4195 46640
rect 24010 46660 24482 46690
rect 24482 46640 24542 46650
rect 23950 46620 24010 46630
rect 24542 46450 24602 46460
rect -4315 46440 -4255 46450
rect -3540 46440 -3480 46450
rect -4255 46390 -3540 46420
rect -4315 46370 -4255 46380
rect -3540 46370 -3480 46380
rect 23950 46430 24010 46440
rect 24010 46400 24542 46430
rect 24542 46380 24602 46390
rect 23950 46360 24010 46370
rect 24602 46180 24662 46190
rect -4375 46170 -4315 46180
rect -3550 46170 -3490 46180
rect -4315 46120 -3550 46150
rect -4375 46100 -4315 46110
rect -3550 46100 -3490 46110
rect 23950 46160 24010 46170
rect 24010 46130 24602 46160
rect 24602 46110 24662 46120
rect 23950 46090 24010 46100
rect -3540 45900 -3480 45910
rect 24662 45900 24722 45910
rect -4435 45890 -4375 45900
rect -4375 45840 -3540 45870
rect -3540 45830 -3480 45840
rect 23950 45890 24010 45900
rect 24010 45850 24662 45880
rect 24662 45830 24722 45840
rect -4435 45820 -4375 45830
rect 23950 45820 24010 45830
rect -3540 45630 -3480 45640
rect -4495 45620 -4435 45630
rect -4435 45570 -3540 45600
rect 24722 45630 24782 45640
rect -3540 45560 -3480 45570
rect 23950 45610 24010 45620
rect -4495 45550 -4435 45560
rect 24010 45580 24722 45610
rect 24722 45560 24782 45570
rect 23950 45540 24010 45550
rect 24782 45370 24842 45380
rect -4555 45360 -4495 45370
rect -3540 45350 -3480 45360
rect -4495 45310 -3540 45340
rect -4555 45290 -4495 45300
rect -3540 45280 -3480 45290
rect 23950 45350 24010 45360
rect 24010 45320 24782 45350
rect 24782 45300 24842 45310
rect 23950 45280 24010 45290
rect 24842 45090 24902 45100
rect -4615 45080 -4555 45090
rect -3540 45080 -3480 45090
rect -4555 45030 -3540 45060
rect -4615 45010 -4555 45020
rect -3540 45010 -3480 45020
rect 23950 45080 24010 45090
rect 24010 45040 24842 45070
rect 24842 45020 24902 45030
rect 23950 45010 24010 45020
rect 24902 44820 24962 44830
rect -4675 44810 -4615 44820
rect 23950 44810 24010 44820
rect -3540 44800 -3480 44810
rect -4615 44760 -3540 44790
rect -4675 44740 -4615 44750
rect 24010 44770 24902 44800
rect 24902 44750 24962 44760
rect 23950 44740 24010 44750
rect -3540 44730 -3480 44740
rect 24962 44540 25022 44550
rect -4735 44530 -4675 44540
rect -3540 44530 -3480 44540
rect -4675 44480 -3540 44510
rect -4735 44460 -4675 44470
rect -3540 44460 -3480 44470
rect 23950 44530 24010 44540
rect 24010 44490 24962 44520
rect 24962 44470 25022 44480
rect 23950 44460 24010 44470
rect 25022 44280 25082 44290
rect -4795 44270 -4735 44280
rect 23950 44270 24010 44280
rect -3540 44260 -3480 44270
rect -4735 44220 -3540 44250
rect -4795 44200 -4735 44210
rect 24010 44230 25022 44260
rect 25022 44210 25082 44220
rect 23950 44200 24010 44210
rect -3540 44190 -3480 44200
rect 25082 44010 25142 44020
rect -4855 44000 -4795 44010
rect -3540 43990 -3480 44000
rect -4795 43950 -3540 43980
rect -4855 43930 -4795 43940
rect -3540 43920 -3480 43930
rect 23950 43990 24010 44000
rect 24010 43960 25082 43990
rect 25082 43940 25142 43950
rect 23950 43920 24010 43930
rect 25142 43740 25202 43750
rect -4915 43730 -4855 43740
rect -3540 43720 -3480 43730
rect -4855 43680 -3540 43710
rect -4915 43660 -4855 43670
rect -3540 43650 -3480 43660
rect 23950 43720 24010 43730
rect 24010 43690 25142 43720
rect 25142 43670 25202 43680
rect 23950 43650 24010 43660
rect -3540 43450 -3480 43460
rect 25202 43450 25262 43460
rect -4975 43440 -4915 43450
rect -4915 43390 -3540 43420
rect -3540 43380 -3480 43390
rect 23950 43440 24010 43450
rect 24010 43400 25202 43430
rect 25202 43380 25262 43390
rect -4975 43370 -4915 43380
rect 23950 43370 24010 43380
rect -3540 43180 -3480 43190
rect 25262 43180 25322 43190
rect -5035 43170 -4975 43180
rect -4975 43120 -3540 43150
rect 23960 43170 24020 43180
rect 23957 43130 23960 43160
rect -3540 43110 -3480 43120
rect 24020 43130 25262 43160
rect 25262 43110 25322 43120
rect -5035 43100 -4975 43110
rect 23960 43100 24020 43110
rect 25322 42920 25382 42930
rect -5095 42910 -5035 42920
rect -3540 42910 -3480 42920
rect -5035 42860 -3540 42890
rect -5095 42840 -5035 42850
rect -3540 42840 -3480 42850
rect 23950 42910 24010 42920
rect 24010 42870 25322 42900
rect 25322 42850 25382 42860
rect 23950 42840 24010 42850
rect -3540 42640 -3480 42650
rect -5155 42620 -5095 42630
rect -5095 42580 -3540 42600
rect 25382 42630 25442 42640
rect -5095 42570 -3480 42580
rect 23950 42620 24010 42630
rect -5155 42550 -5095 42560
rect 24010 42580 25382 42610
rect 25382 42560 25442 42570
rect 23950 42550 24010 42560
rect -3540 42370 -3480 42380
rect -5215 42350 -5155 42360
rect -5155 42310 -3540 42330
rect -5155 42300 -3480 42310
rect 23950 42360 24010 42370
rect 25442 42360 25502 42370
rect 24010 42310 25442 42340
rect 23950 42290 24010 42300
rect 25442 42290 25502 42300
rect -5215 42280 -5155 42290
rect 8796 42126 9734 42154
rect 10636 42096 11564 42124
rect 23940 42080 24000 42090
rect -5275 42070 -5215 42080
rect -3540 42060 -3480 42070
rect -5215 42020 -3540 42050
rect -5275 42000 -5215 42010
rect 1436 42046 2384 42074
rect 6956 42036 7884 42064
rect 14316 42016 15254 42044
rect 25502 42080 25562 42090
rect 24000 42030 25502 42060
rect 23940 42010 24000 42020
rect 25502 42010 25562 42020
rect -3540 41990 -3480 42000
rect 3276 41906 4214 41934
rect 20756 41906 21684 41934
rect 16156 41876 17094 41904
rect 17996 41846 18924 41874
rect -404 41736 534 41764
rect 16140 41700 16200 41710
rect -1340 41650 -1280 41660
rect -3180 41590 -3120 41600
rect -3180 41520 -3120 41530
rect -2260 41590 -2200 41600
rect 5116 41616 6030 41644
rect 16140 41630 16200 41640
rect 17980 41630 18040 41640
rect -1340 41580 -1280 41590
rect 12510 41546 13424 41574
rect -2260 41520 -2200 41530
rect 510 41310 540 41530
rect 500 41300 560 41310
rect 500 41230 560 41240
rect 2350 41220 2380 41530
rect 2330 41210 2390 41220
rect 2330 41140 2390 41150
rect -2670 40680 -2500 40690
rect -2670 40330 -2500 40340
rect 1540 40680 1910 40690
rect 4190 40670 4220 41530
rect 5110 40760 5140 41530
rect 6950 40950 6980 41530
rect 8790 41040 8820 41530
rect 10630 41130 10660 41530
rect 15222 41480 15278 41588
rect 17980 41560 18040 41570
rect 19830 41480 19870 41610
rect 20740 41560 20800 41570
rect 20740 41490 20800 41500
rect 22590 41480 22630 41610
rect 15220 41470 15280 41480
rect 13390 41400 13420 41440
rect 15220 41400 15280 41410
rect 19820 41470 19880 41480
rect 19820 41400 19880 41410
rect 22580 41470 22640 41480
rect 22580 41400 22640 41410
rect 23200 41470 23260 41480
rect 23200 41400 23260 41410
rect 13370 41390 13430 41400
rect 13370 41320 13430 41330
rect 17080 41240 17450 41250
rect 10620 41120 10680 41130
rect 10620 41050 10680 41060
rect 15090 41100 15150 41110
rect 15780 41100 15840 41110
rect 15150 41050 15780 41080
rect 8780 41030 8840 41040
rect 15090 41030 15150 41040
rect 15780 41030 15840 41040
rect 8780 40960 8840 40970
rect 6940 40940 7000 40950
rect 6940 40870 7000 40880
rect 15000 40850 15060 40860
rect 15620 40850 15680 40860
rect 15060 40800 15620 40830
rect 15000 40780 15060 40790
rect 15620 40780 15680 40790
rect 14710 40760 14770 40770
rect 5090 40750 5150 40760
rect 15710 40760 15770 40770
rect 14770 40710 15710 40740
rect 14710 40690 14770 40700
rect 15710 40690 15770 40700
rect 5090 40680 5150 40690
rect 9260 40680 9630 40690
rect 4180 40660 4240 40670
rect 4180 40590 4240 40600
rect 1540 40270 1910 40340
rect 9260 40330 9630 40340
rect 17080 40680 17450 41150
rect 22480 41230 23040 41240
rect 23210 41110 23240 41400
rect 23520 41110 23550 41565
rect 23640 41410 23700 41420
rect 23640 41340 23700 41350
rect 23660 41110 23690 41340
rect 22480 41070 23040 41080
rect 23190 41100 23250 41110
rect 23190 41030 23250 41040
rect 23520 41100 23580 41110
rect 23520 41030 23580 41040
rect 23640 41100 23700 41110
rect 23640 41030 23700 41040
rect 24050 41020 24110 41030
rect 23875 40970 24050 41000
rect 24050 40950 24110 40960
rect 17080 40330 17450 40340
rect 23630 40390 23690 40400
rect 23630 40320 23690 40330
rect 1540 40160 1910 40170
rect -580 39830 -520 39840
rect 555 39820 615 39830
rect -520 39780 555 39820
rect -580 39760 -520 39770
rect 615 39780 1050 39820
rect 555 39750 615 39760
rect 10360 39670 10420 39680
rect 10360 39600 10420 39610
rect 15770 38954 15830 38964
rect 9980 38910 10040 38920
rect 15770 38884 15830 38894
rect 9980 38840 10040 38850
rect 14530 38750 15060 38850
rect -667 38736 -607 38746
rect -667 38676 -662 38736
rect 680 38740 740 38750
rect -607 38690 680 38730
rect -667 38666 -607 38676
rect 740 38690 1067 38730
rect 680 38670 740 38680
rect 3410 38080 3470 38090
rect 3290 38040 3410 38080
rect 3410 38010 3470 38020
rect 14810 38020 14870 38030
rect 14750 37970 14810 38000
rect 14810 37950 14870 37960
rect 15010 37920 15060 38750
rect 15680 38064 15740 38074
rect 15740 38015 15880 38055
rect 15680 37994 15740 38004
rect 14695 37890 14905 37918
rect 14695 37888 14920 37890
rect 14860 37880 14920 37888
rect 14695 37798 14805 37828
rect 14860 37810 14920 37820
rect 3345 37750 3486 37768
rect 3250 37738 3486 37750
rect 3250 37710 3390 37738
rect 14775 37735 14805 37798
rect 14860 37750 14920 37760
rect 14775 37705 14860 37735
rect 14860 37680 14920 37690
rect 3410 37670 3470 37680
rect 15010 37640 15630 37920
rect 15680 37880 15740 37890
rect 15680 37810 15740 37820
rect 15750 37750 15810 37760
rect 15750 37680 15810 37690
rect 3410 37600 3470 37610
rect 1960 37330 2300 37340
rect 1960 36980 2300 36990
rect 7410 37330 7750 37340
rect 7410 36980 7750 36990
rect 15080 36940 15140 36950
rect 15080 36870 15140 36880
rect 10095 36840 10155 36850
rect 9975 36780 10035 36790
rect 9885 36720 9945 36730
rect 9795 36660 9855 36670
rect 9705 36600 9765 36610
rect 9615 36540 9675 36550
rect 9525 36480 9585 36490
rect 9975 36710 10035 36720
rect 9885 36650 9945 36660
rect 9795 36590 9855 36600
rect 9705 36530 9765 36540
rect 9615 36470 9675 36480
rect 9525 36410 9585 36420
rect 560 36190 900 36200
rect 560 36090 900 36100
rect -100 35040 240 35050
rect -100 34690 240 34700
rect 9555 32880 9585 36410
rect 9645 32970 9675 36470
rect 9735 33060 9765 36530
rect 9825 33150 9855 36590
rect 9915 33240 9945 36650
rect 10005 33330 10035 36710
rect 10095 36770 10155 36780
rect 10185 36780 10245 36790
rect 10095 33420 10125 36770
rect 10185 36710 10245 36720
rect 10275 36720 10335 36730
rect 10185 33510 10215 36710
rect 10275 36650 10335 36660
rect 10365 36660 10425 36670
rect 10275 33600 10305 36650
rect 10365 36590 10425 36600
rect 10455 36600 10515 36610
rect 10365 33690 10395 36590
rect 10455 36530 10515 36540
rect 10545 36540 10605 36550
rect 10455 33780 10485 36530
rect 10545 36470 10605 36480
rect 10635 36480 10695 36490
rect 10545 33870 10575 36470
rect 10635 36410 10695 36420
rect 10635 33960 10665 36410
rect 15100 36400 15130 36870
rect 15080 36390 15140 36400
rect 15080 36320 15140 36330
rect 19810 36190 20150 36200
rect 19810 36090 20150 36100
rect 19540 35040 19910 35050
rect 19540 34660 19910 34670
rect 10620 33950 10680 33960
rect 10620 33880 10680 33890
rect 10530 33860 10590 33870
rect 10530 33790 10590 33800
rect 10440 33770 10500 33780
rect 10440 33700 10500 33710
rect 10350 33680 10410 33690
rect 10350 33610 10410 33620
rect 10260 33590 10320 33600
rect 10260 33520 10320 33530
rect 10170 33500 10230 33510
rect 10170 33430 10230 33440
rect 10080 33410 10140 33420
rect 10080 33340 10140 33350
rect 9990 33320 10050 33330
rect 9990 33250 10050 33260
rect 9900 33230 9960 33240
rect 9900 33160 9960 33170
rect 9810 33140 9870 33150
rect 9810 33070 9870 33080
rect 9720 33050 9780 33060
rect 9720 32980 9780 32990
rect 9630 32960 9690 32970
rect 9630 32890 9690 32900
rect 9540 32870 9600 32880
rect 9540 32800 9600 32810
rect 18840 32160 19200 32170
rect 1090 32140 1430 32150
rect 1090 31790 1430 31800
rect 18840 31790 19200 31800
<< via2 >>
rect -3540 48010 -3480 48070
rect 23950 48000 24010 48060
rect -3540 47730 -3480 47790
rect 23950 47730 24010 47790
rect -3540 47470 -3480 47530
rect 23950 47460 24010 47520
rect -3540 47190 -3480 47250
rect 23950 47190 24010 47250
rect -3550 46920 -3490 46980
rect 23950 46910 24010 46970
rect -3550 46650 -3490 46710
rect 23950 46630 24010 46690
rect -3540 46380 -3480 46440
rect 23950 46370 24010 46430
rect -3550 46110 -3490 46170
rect 23950 46100 24010 46160
rect -3540 45840 -3480 45900
rect 23950 45830 24010 45890
rect -3540 45570 -3480 45630
rect 23950 45550 24010 45610
rect -3540 45290 -3480 45350
rect 23950 45290 24010 45350
rect -3540 45020 -3480 45080
rect 23950 45020 24010 45080
rect -3540 44740 -3480 44800
rect 23950 44750 24010 44810
rect -3540 44470 -3480 44530
rect 23950 44470 24010 44530
rect -3540 44200 -3480 44260
rect 23950 44210 24010 44270
rect -3540 43930 -3480 43990
rect 23950 43930 24010 43990
rect -3540 43660 -3480 43720
rect 23950 43660 24010 43720
rect -3540 43390 -3480 43450
rect 23950 43380 24010 43440
rect -3540 43120 -3480 43180
rect 23960 43110 24020 43170
rect -3540 42850 -3480 42910
rect 23950 42850 24010 42910
rect -3540 42580 -3480 42640
rect 23950 42560 24010 42620
rect -3540 42310 -3480 42370
rect 23950 42300 24010 42360
rect -3540 42000 -3480 42060
rect 23940 42020 24000 42080
rect -2670 40340 -2500 40680
rect 1540 40340 1910 40680
rect 9260 40340 9630 40680
rect 22480 41080 23040 41230
rect 17080 40340 17450 40680
rect 10360 39610 10420 39670
rect 9980 38850 10040 38910
rect 14860 37820 14920 37880
rect 14860 37690 14920 37750
rect 15680 37820 15740 37880
rect 15750 37690 15810 37750
rect 1960 36990 2300 37330
rect 7410 36990 7750 37330
rect 560 36100 900 36190
rect -100 34700 240 35040
rect 19810 36100 20150 36190
rect 19540 34670 19910 35040
rect 1090 31800 1430 32140
rect 18840 31800 19200 32160
<< metal3 >>
rect -3550 48070 -3470 48075
rect -3550 48010 -3540 48070
rect -3480 48010 -3470 48070
rect -3550 48005 -3470 48010
rect 23940 48060 24020 48065
rect 23940 48000 23950 48060
rect 24010 48000 24020 48060
rect 23940 47995 24020 48000
rect -3550 47790 -3470 47795
rect -3550 47730 -3540 47790
rect -3480 47730 -3470 47790
rect -3550 47725 -3470 47730
rect 23940 47790 24020 47795
rect 23940 47730 23950 47790
rect 24010 47730 24020 47790
rect 23940 47725 24020 47730
rect -3550 47530 -3470 47535
rect -3550 47470 -3540 47530
rect -3480 47470 -3470 47530
rect -3550 47465 -3470 47470
rect 23940 47520 24020 47525
rect 23940 47460 23950 47520
rect 24010 47460 24020 47520
rect 23940 47455 24020 47460
rect -3550 47250 -3470 47255
rect -3550 47190 -3540 47250
rect -3480 47190 -3470 47250
rect -3550 47185 -3470 47190
rect 23940 47250 24020 47255
rect 23940 47190 23950 47250
rect 24010 47190 24020 47250
rect 23940 47185 24020 47190
rect -3560 46980 -3480 46985
rect -3560 46920 -3550 46980
rect -3490 46920 -3480 46980
rect -3560 46915 -3480 46920
rect 23940 46970 24020 46975
rect 23940 46910 23950 46970
rect 24010 46910 24020 46970
rect 23940 46905 24020 46910
rect -3560 46710 -3480 46715
rect -3560 46650 -3550 46710
rect -3490 46650 -3480 46710
rect -3560 46645 -3480 46650
rect 23940 46690 24020 46695
rect 23940 46630 23950 46690
rect 24010 46630 24020 46690
rect 23940 46625 24020 46630
rect -3550 46440 -3470 46445
rect -3550 46380 -3540 46440
rect -3480 46380 -3470 46440
rect -3550 46375 -3470 46380
rect 23940 46430 24020 46435
rect 23940 46370 23950 46430
rect 24010 46370 24020 46430
rect 23940 46365 24020 46370
rect -3560 46170 -3480 46175
rect -3560 46110 -3550 46170
rect -3490 46110 -3480 46170
rect -3560 46105 -3480 46110
rect 23940 46160 24020 46165
rect 23940 46100 23950 46160
rect 24010 46100 24020 46160
rect 23940 46095 24020 46100
rect -3550 45900 -3470 45905
rect -3550 45840 -3540 45900
rect -3480 45840 -3470 45900
rect -3550 45835 -3470 45840
rect 23940 45890 24020 45895
rect 23940 45830 23950 45890
rect 24010 45830 24020 45890
rect 23940 45825 24020 45830
rect -3550 45630 -3470 45635
rect -3550 45570 -3540 45630
rect -3480 45570 -3470 45630
rect -3550 45565 -3470 45570
rect 23940 45610 24020 45615
rect 23940 45550 23950 45610
rect 24010 45550 24020 45610
rect 23940 45545 24020 45550
rect -3550 45350 -3470 45355
rect -3550 45290 -3540 45350
rect -3480 45290 -3470 45350
rect -3550 45285 -3470 45290
rect 23940 45350 24020 45355
rect 23940 45290 23950 45350
rect 24010 45290 24020 45350
rect 23940 45285 24020 45290
rect -3550 45080 -3470 45085
rect -3550 45020 -3540 45080
rect -3480 45020 -3470 45080
rect -3550 45015 -3470 45020
rect 23940 45080 24020 45085
rect 23940 45020 23950 45080
rect 24010 45020 24020 45080
rect 23940 45015 24020 45020
rect 23940 44810 24020 44815
rect -3550 44800 -3470 44805
rect -3550 44740 -3540 44800
rect -3480 44740 -3470 44800
rect 23940 44750 23950 44810
rect 24010 44750 24020 44810
rect 23940 44745 24020 44750
rect -3550 44735 -3470 44740
rect -3550 44530 -3470 44535
rect -3550 44470 -3540 44530
rect -3480 44470 -3470 44530
rect -3550 44465 -3470 44470
rect 23940 44530 24020 44535
rect 23940 44470 23950 44530
rect 24010 44470 24020 44530
rect 23940 44465 24020 44470
rect 23940 44270 24020 44275
rect -3550 44260 -3470 44265
rect -3550 44200 -3540 44260
rect -3480 44200 -3470 44260
rect 23940 44210 23950 44270
rect 24010 44210 24020 44270
rect 23940 44205 24020 44210
rect -3550 44195 -3470 44200
rect -3550 43990 -3470 43995
rect -3550 43930 -3540 43990
rect -3480 43930 -3470 43990
rect -3550 43925 -3470 43930
rect 23940 43990 24020 43995
rect 23940 43930 23950 43990
rect 24010 43930 24020 43990
rect 23940 43925 24020 43930
rect -3550 43720 -3470 43725
rect -3550 43660 -3540 43720
rect -3480 43660 -3470 43720
rect -3550 43655 -3470 43660
rect 23940 43720 24020 43725
rect 23940 43660 23950 43720
rect 24010 43660 24020 43720
rect 23940 43655 24020 43660
rect -3550 43450 -3470 43455
rect -3550 43390 -3540 43450
rect -3480 43390 -3470 43450
rect -3550 43385 -3470 43390
rect 23940 43440 24020 43445
rect 23940 43380 23950 43440
rect 24010 43380 24020 43440
rect 23940 43375 24020 43380
rect -3550 43180 -3470 43185
rect -3550 43120 -3540 43180
rect -3480 43120 -3470 43180
rect -3550 43115 -3470 43120
rect 23950 43170 24030 43175
rect 23950 43110 23960 43170
rect 24020 43110 24030 43170
rect 23950 43105 24030 43110
rect -3550 42910 -3470 42915
rect -3550 42850 -3540 42910
rect -3480 42850 -3470 42910
rect -3550 42845 -3470 42850
rect 23940 42910 24020 42915
rect 23940 42850 23950 42910
rect 24010 42850 24020 42910
rect 23940 42845 24020 42850
rect -3550 42640 -3470 42645
rect -3550 42580 -3540 42640
rect -3480 42580 -3470 42640
rect -3550 42575 -3470 42580
rect 23940 42620 24020 42625
rect 23940 42560 23950 42620
rect 24010 42560 24020 42620
rect 23940 42555 24020 42560
rect -3550 42370 -3470 42375
rect -3550 42310 -3540 42370
rect -3480 42310 -3470 42370
rect -3550 42305 -3470 42310
rect 23940 42360 24020 42365
rect 23940 42300 23950 42360
rect 24010 42300 24020 42360
rect 23940 42295 24020 42300
rect 23930 42080 24010 42085
rect -3550 42060 -3470 42065
rect -3550 42000 -3540 42060
rect -3480 42000 -3470 42060
rect 23930 42020 23940 42080
rect 24000 42020 24010 42080
rect 23930 42015 24010 42020
rect -3550 41995 -3470 42000
rect 22470 41230 23050 41235
rect -3040 40850 560 41190
rect 900 40850 910 41190
rect 22470 41080 22480 41230
rect 23040 41080 23050 41230
rect 22470 41075 23050 41080
rect -3040 40315 -2870 40850
rect -2680 40680 -2490 40685
rect -110 40680 250 40685
rect 1530 40680 1920 40685
rect 9250 40680 9640 40685
rect 17070 40680 17460 40685
rect -2680 40340 -2670 40680
rect -2500 40340 -100 40680
rect 240 40340 1540 40680
rect 1910 40340 9260 40680
rect 9630 40340 17080 40680
rect 17450 40340 19170 40680
rect 19540 40340 22390 40680
rect -2680 40335 -2490 40340
rect -110 40335 250 40340
rect 1530 40335 1920 40340
rect 9250 40335 9640 40340
rect 17070 40335 17460 40340
rect 9670 39810 10690 40020
rect 9670 39460 10240 39810
rect 10340 39680 10440 39690
rect 10340 39610 10360 39680
rect 10430 39610 10440 39680
rect 10340 39590 10440 39610
rect 10570 39460 10690 39810
rect 9670 39060 10690 39460
rect 9670 38710 9840 39060
rect 9950 38920 10060 38930
rect 9950 38850 9970 38920
rect 10040 38850 10060 38920
rect 9950 38830 10060 38850
rect 10170 38710 10690 39060
rect 1950 37330 2310 37335
rect 7400 37330 7760 37335
rect 9670 37330 10690 38710
rect 14850 37880 14930 37885
rect 15670 37880 15750 37885
rect 14850 37820 14860 37880
rect 14920 37820 15680 37880
rect 15740 37820 15750 37880
rect 14850 37815 14930 37820
rect 15670 37815 15750 37820
rect 14850 37750 14930 37755
rect 15740 37750 15820 37755
rect 14850 37690 14860 37750
rect 14920 37690 15750 37750
rect 15810 37690 15820 37750
rect 14850 37685 14930 37690
rect 15740 37685 15820 37690
rect 550 36990 560 37330
rect 900 36990 1960 37330
rect 2300 36990 7410 37330
rect 7750 36990 22480 37330
rect 23040 36990 23050 37330
rect 1950 36985 2310 36990
rect 7400 36985 7760 36990
rect 550 36190 910 36195
rect 550 36100 560 36190
rect 900 36100 910 36190
rect 550 36095 910 36100
rect -110 35040 250 35045
rect -110 34700 -100 35040
rect 240 34700 250 35040
rect -110 34695 250 34700
rect -5310 4780 -5250 31560
rect -5180 4840 -5120 31410
rect -5050 4960 -4990 31820
rect -4790 31720 -4730 32440
rect 3370 32350 4190 32630
rect -4920 31660 -4730 31720
rect 1080 32140 1440 32150
rect 1080 31800 1090 32140
rect 1430 31800 1440 32140
rect -4920 5080 -4860 31660
rect 1080 30870 1440 31800
rect 3370 32100 3670 32350
rect 3890 32100 4190 32350
rect 3370 30870 4190 32100
rect 1080 30850 4190 30870
rect 9670 30860 10690 36990
rect 19810 36195 20150 36990
rect 19800 36190 20160 36195
rect 19800 36100 19810 36190
rect 20150 36100 20160 36190
rect 19800 36095 20160 36100
rect 19530 35040 19920 35045
rect 19530 34670 19540 35040
rect 19910 34670 19920 35040
rect 19530 34665 19920 34670
rect 16110 32350 16930 32630
rect 16110 32100 16390 32350
rect 16620 32100 16930 32350
rect 16110 30870 16930 32100
rect 18830 32160 19210 32165
rect 18830 31800 18840 32160
rect 19200 31800 19210 32160
rect 18830 31795 19210 31800
rect 18850 30870 19210 31795
rect 25017 31720 25077 32440
rect 25017 31660 25207 31720
rect 16110 30860 19210 30870
rect 9670 30850 19210 30860
rect 1080 30510 19210 30850
rect 3370 30140 16930 30510
rect 3370 30130 12210 30140
rect 8080 29840 12210 30130
rect 8080 29470 12010 29840
rect 25147 5080 25207 31660
rect -4920 5020 25207 5080
rect 25277 4960 25337 31820
rect -5050 4900 25337 4960
rect 25407 4840 25467 31410
rect -5180 4780 25467 4840
rect 25537 4780 25597 31560
<< via3 >>
rect 560 40850 900 41190
rect 22480 41080 23040 41230
rect -100 40340 240 40680
rect 19170 40340 19540 40680
rect 10360 39670 10430 39680
rect 10360 39610 10420 39670
rect 10420 39610 10430 39670
rect 9970 38910 10040 38920
rect 9970 38850 9980 38910
rect 9980 38850 10040 38910
rect 560 36990 900 37330
rect 22480 36990 23040 37330
rect 560 36100 900 36190
rect -100 34700 240 35040
rect 1090 31800 1430 32140
rect 19540 34670 19910 35040
<< metal4 >>
rect -92 47401 228 47630
rect 568 47438 888 47620
rect -101 41089 241 47401
rect 560 41191 900 47438
rect 22480 41231 23040 41270
rect 22479 41230 23041 41231
rect 559 41190 901 41191
rect -100 40681 240 41089
rect 559 40850 560 41190
rect 900 40850 901 41190
rect 22479 41080 22480 41230
rect 23040 41080 23041 41230
rect 22479 41079 23041 41080
rect 559 40849 901 40850
rect -101 40680 241 40681
rect -101 40340 -100 40680
rect 240 40340 241 40680
rect -101 40339 241 40340
rect -100 35041 240 40339
rect 560 37331 900 40849
rect 19169 40680 19541 40681
rect 19169 40340 19170 40680
rect 19540 40340 19541 40680
rect 19169 40339 19541 40340
rect 10359 39680 10431 39681
rect 10359 39610 10360 39680
rect 10430 39610 10431 39680
rect 10359 39609 10431 39610
rect 9969 38920 10041 38921
rect 9969 38850 9970 38920
rect 10040 38890 10041 38920
rect 10040 38850 10050 38890
rect 9969 38849 10050 38850
rect 559 37330 901 37331
rect 559 36990 560 37330
rect 900 36990 901 37330
rect 559 36989 901 36990
rect 560 36191 900 36989
rect 559 36190 901 36191
rect 559 36100 560 36190
rect 900 36100 901 36190
rect 559 36099 901 36100
rect -101 35040 241 35041
rect -101 34700 -100 35040
rect 240 34700 241 35040
rect -101 34699 241 34700
rect -100 34670 240 34699
rect 560 33351 900 36099
rect 559 32141 901 33351
rect 3739 32199 3821 32281
rect 559 32140 1431 32141
rect 559 31800 1090 32140
rect 1430 31800 1431 32140
rect 559 31799 1431 31800
rect 3750 30530 3810 32199
rect 9990 30530 10050 38849
rect 3750 30470 10050 30530
rect 9990 29740 10050 30470
rect 8370 29680 10050 29740
rect 10370 30530 10430 39609
rect 19170 35041 19540 40339
rect 22480 37331 23040 41079
rect 22479 37330 23041 37331
rect 22479 36990 22480 37330
rect 23040 36990 23041 37330
rect 22479 36989 23041 36990
rect 19170 35040 19911 35041
rect 19170 34670 19540 35040
rect 19910 34670 19911 35040
rect 19539 34669 19911 34670
rect 16480 32271 16540 32285
rect 16469 32189 16551 32271
rect 16480 30530 16540 32189
rect 10370 30470 16540 30530
rect 10370 29740 10430 30470
rect 10370 29680 11917 29740
rect 8370 29460 8430 29680
rect 11857 29470 11917 29680
use break_before_make  break_before_make_0 ~/Desktop/SAR_ADC_12bit/break_before_make/layout
timestamp 1714246951
transform 1 0 -7060 0 1 30160
box 1800 5890 6245 11260
use DAC_and_SW  DAC_and_SW_0
timestamp 1714329720
transform -1 0 24887 0 1 5100
box -720 0 15040 31096
use DAC_and_SW  DAC_and_SW_2
timestamp 1714329720
transform 1 0 -4600 0 1 5100
box -720 0 15040 31096
use latched_comparator  latched_comparator_0 ~/Desktop/SAR_ADC_12bit/layout/../latched_comparator/layout
timestamp 1712061640
transform -1 0 8780 0 1 39170
box 5450 -1740 7860 1100
use offset_calibration  offset_calibration_0 ~/Desktop/SAR_ADC_12bit/layout/../offset_calibration/layout
timestamp 1712002773
transform 1 0 12181 0 1 38345
box 3610 -1900 11750 2900
use preamplifier  preamplifier_0 ~/Desktop/SAR_ADC_12bit/layout/../preamplifier/layout
timestamp 1711972782
transform -1 0 11136 0 1 30538
box -3630 6580 7680 9930
use state_machine  state_machine_0 ~/Desktop/SAR_ADC_12bit/layout/../state_machine/layout
timestamp 1714331631
transform 1 0 -4300 0 1 40085
box 560 1200 28420 8110
<< labels >>
rlabel metal2 3350 38050 3380 38070 1 VDAC_Pi
rlabel metal2 3340 37720 3370 37740 1 VDAC_Ni
rlabel metal2 910 39790 940 39810 1 COMP_P
rlabel metal3 15640 37700 15660 37730 1 CAL_N
rlabel metal3 15640 37830 15660 37860 1 CAL_P
rlabel metal4 11870 29490 11910 29510 1 VDAC_N
rlabel metal4 8380 29490 8420 29510 1 VDAC_P
rlabel metal2 -3744 48018 -3716 48034 1 SMPL_ON_P
rlabel metal2 24104 48026 24132 48042 1 SMPL_ON_N
rlabel metal2 -2990 48010 -2940 48190 1 CLK_DATA
port 1 n
rlabel metal2 -600 48010 -550 48190 1 DATA[0]
port 2 n
rlabel metal4 -80 47340 200 47600 1 VDD
port 20 n
rlabel metal2 1790 48010 1840 48190 1 DATA[1]
port 3 n
rlabel metal2 4190 48010 4240 48190 1 DATA[2]
port 4 n
rlabel metal2 6580 48010 6630 48190 1 DATA[3]
port 5 n
rlabel metal2 8970 48010 9020 48190 1 DATA[4]
port 6 n
rlabel metal2 11360 48010 11410 48190 1 DATA[5]
port 7 n
rlabel metal2 13750 47890 13800 48070 1 RST_Z
port 9 n
rlabel metal2 16140 48010 16190 48190 1 CLK
port 22 n
rlabel metal2 18540 48010 18590 48190 1 START
port 10 n
rlabel metal2 23320 48010 23370 48190 1 EN_OFFSET_CAL
port 11 n
rlabel metal2 20930 48010 20980 48190 1 SINGLE_ENDED
port 23 n
rlabel metal2 9050 9490 9070 9560 1 C10_P_btm
rlabel metal2 9140 11680 9160 11780 1 C9_P_btm
rlabel metal2 9230 13490 9250 13580 1 C8_P_btm
rlabel metal2 9320 14600 9340 14720 1 C7_P_btm
rlabel metal2 9410 15330 9430 15410 1 C6_P_btm
rlabel metal2 9500 15720 9520 15800 1 C5_P_btm
rlabel metal2 9590 16430 9610 16510 1 C4_P_btm
rlabel metal2 9670 16900 9690 16960 1 C2_P_btm
rlabel metal2 9770 17190 9790 17260 1 C0_dummy_P_btm
rlabel metal2 9860 17560 9880 17620 1 C0_P_btm
rlabel metal2 9950 17920 9970 17980 1 C1_P_btm
rlabel metal2 10040 18290 10060 18350 1 C3_P_btm
rlabel metal2 11220 9470 11240 9540 1 C10_N_btm
rlabel metal2 11130 11690 11150 11790 1 C9_N_btm
rlabel metal2 11030 13500 11050 13590 1 C8_N_btm
rlabel metal2 10950 14630 10970 14750 1 C7_N_btm
rlabel metal2 10860 15340 10880 15420 1 C6_N_btm
rlabel metal2 10770 15700 10790 15780 1 C5_N_btm
rlabel metal2 10670 16430 10690 16510 1 C4_N_btm
rlabel metal2 10590 16830 10610 16890 1 C2_N_btm
rlabel metal2 10500 17190 10520 17260 1 C0_dummy_N_btm
rlabel metal2 10410 17570 10430 17630 1 C0_N_btm
rlabel metal2 10320 17930 10340 17990 1 C1_N_btm
rlabel metal2 10230 18300 10250 18360 1 C3_N_btm
rlabel metal3 -5310 4780 -5250 4840 1 VIN_P
port 24 n
rlabel metal3 25537 4780 25597 4840 1 VIN_N
port 25 n
rlabel metal3 10230 5020 10300 5080 1 VCM
port 26 n
rlabel metal3 10230 4900 10300 4960 1 VREF
port 27 n
rlabel metal3 10230 4780 10300 4840 1 VREF_GND
port 28 n
rlabel metal2 1366 34636 1394 34652 1 EN_VIN_BSTR_P
rlabel metal2 18890 34628 18920 34660 1 EN_VIN_BSTR_N
rlabel metal4 582 47342 868 47606 1 VSS
port 29 n
<< end >>
