magic
tech sky130A
magscale 1 2
timestamp 1711994487
<< nwell >>
rect -1196 -3455 1196 3455
<< pmoslvt >>
rect -1000 1236 1000 3236
rect -1000 -1000 1000 1000
rect -1000 -3236 1000 -1236
<< pdiff >>
rect -1058 3224 -1000 3236
rect -1058 1248 -1046 3224
rect -1012 1248 -1000 3224
rect -1058 1236 -1000 1248
rect 1000 3224 1058 3236
rect 1000 1248 1012 3224
rect 1046 1248 1058 3224
rect 1000 1236 1058 1248
rect -1058 988 -1000 1000
rect -1058 -988 -1046 988
rect -1012 -988 -1000 988
rect -1058 -1000 -1000 -988
rect 1000 988 1058 1000
rect 1000 -988 1012 988
rect 1046 -988 1058 988
rect 1000 -1000 1058 -988
rect -1058 -1248 -1000 -1236
rect -1058 -3224 -1046 -1248
rect -1012 -3224 -1000 -1248
rect -1058 -3236 -1000 -3224
rect 1000 -1248 1058 -1236
rect 1000 -3224 1012 -1248
rect 1046 -3224 1058 -1248
rect 1000 -3236 1058 -3224
<< pdiffc >>
rect -1046 1248 -1012 3224
rect 1012 1248 1046 3224
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect -1046 -3224 -1012 -1248
rect 1012 -3224 1046 -1248
<< nsubdiff >>
rect -1160 3385 -1064 3419
rect 1064 3385 1160 3419
rect -1160 3323 -1126 3385
rect 1126 3323 1160 3385
rect -1160 -3385 -1126 -3323
rect 1126 -3385 1160 -3323
rect -1160 -3419 -1064 -3385
rect 1064 -3419 1160 -3385
<< nsubdiffcont >>
rect -1064 3385 1064 3419
rect -1160 -3323 -1126 3323
rect 1126 -3323 1160 3323
rect -1064 -3419 1064 -3385
<< poly >>
rect -1000 3317 1000 3333
rect -1000 3283 -984 3317
rect 984 3283 1000 3317
rect -1000 3236 1000 3283
rect -1000 1189 1000 1236
rect -1000 1155 -984 1189
rect 984 1155 1000 1189
rect -1000 1139 1000 1155
rect -1000 1081 1000 1097
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1000 1000 1000 1047
rect -1000 -1047 1000 -1000
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1000 -1097 1000 -1081
rect -1000 -1155 1000 -1139
rect -1000 -1189 -984 -1155
rect 984 -1189 1000 -1155
rect -1000 -1236 1000 -1189
rect -1000 -3283 1000 -3236
rect -1000 -3317 -984 -3283
rect 984 -3317 1000 -3283
rect -1000 -3333 1000 -3317
<< polycont >>
rect -984 3283 984 3317
rect -984 1155 984 1189
rect -984 1047 984 1081
rect -984 -1081 984 -1047
rect -984 -1189 984 -1155
rect -984 -3317 984 -3283
<< locali >>
rect -1160 3385 -1064 3419
rect 1064 3385 1160 3419
rect -1160 3323 -1126 3385
rect 1126 3323 1160 3385
rect -1000 3283 -984 3317
rect 984 3283 1000 3317
rect -1046 3224 -1012 3240
rect -1046 1232 -1012 1248
rect 1012 3224 1046 3240
rect 1012 1232 1046 1248
rect -1000 1155 -984 1189
rect 984 1155 1000 1189
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1046 988 -1012 1004
rect -1046 -1004 -1012 -988
rect 1012 988 1046 1004
rect 1012 -1004 1046 -988
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1000 -1189 -984 -1155
rect 984 -1189 1000 -1155
rect -1046 -1248 -1012 -1232
rect -1046 -3240 -1012 -3224
rect 1012 -1248 1046 -1232
rect 1012 -3240 1046 -3224
rect -1000 -3317 -984 -3283
rect 984 -3317 1000 -3283
rect -1160 -3385 -1126 -3323
rect 1126 -3385 1160 -3323
rect -1160 -3419 -1064 -3385
rect 1064 -3419 1160 -3385
<< viali >>
rect -984 3283 984 3317
rect -1046 1248 -1012 3224
rect 1012 1248 1046 3224
rect -984 1155 984 1189
rect -984 1047 984 1081
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect -984 -1081 984 -1047
rect -984 -1189 984 -1155
rect -1046 -3224 -1012 -1248
rect 1012 -3224 1046 -1248
rect -984 -3317 984 -3283
<< metal1 >>
rect -996 3317 996 3323
rect -996 3283 -984 3317
rect 984 3283 996 3317
rect -996 3277 996 3283
rect -1052 3224 -1006 3236
rect -1052 1248 -1046 3224
rect -1012 1248 -1006 3224
rect -1052 1236 -1006 1248
rect 1006 3224 1052 3236
rect 1006 1248 1012 3224
rect 1046 1248 1052 3224
rect 1006 1236 1052 1248
rect -996 1189 996 1195
rect -996 1155 -984 1189
rect 984 1155 996 1189
rect -996 1149 996 1155
rect -996 1081 996 1087
rect -996 1047 -984 1081
rect 984 1047 996 1081
rect -996 1041 996 1047
rect -1052 988 -1006 1000
rect -1052 -988 -1046 988
rect -1012 -988 -1006 988
rect -1052 -1000 -1006 -988
rect 1006 988 1052 1000
rect 1006 -988 1012 988
rect 1046 -988 1052 988
rect 1006 -1000 1052 -988
rect -996 -1047 996 -1041
rect -996 -1081 -984 -1047
rect 984 -1081 996 -1047
rect -996 -1087 996 -1081
rect -996 -1155 996 -1149
rect -996 -1189 -984 -1155
rect 984 -1189 996 -1155
rect -996 -1195 996 -1189
rect -1052 -1248 -1006 -1236
rect -1052 -3224 -1046 -1248
rect -1012 -3224 -1006 -1248
rect -1052 -3236 -1006 -3224
rect 1006 -1248 1052 -1236
rect 1006 -3224 1012 -1248
rect 1046 -3224 1052 -1248
rect 1006 -3236 1052 -3224
rect -996 -3283 996 -3277
rect -996 -3317 -984 -3283
rect 984 -3317 996 -3283
rect -996 -3323 996 -3317
<< properties >>
string FIXED_BBOX -1143 -3402 1143 3402
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 10.0 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
