* NGSPICE file created from bootstrap.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_7FRQHJ a_n3087_118# a_n3029_21# a_29_n965# a_n3087_n868#
+ a_n29_n868# a_29_21# a_3029_n868# a_3029_118# w_n3225_n1087# a_n3029_n965# a_n29_118#
X0 a_n29_118# a_n3029_21# a_n3087_118# w_n3225_n1087# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=1.0875 ps=8.08 w=3.75 l=15
X1 a_3029_118# a_29_21# a_n29_118# w_n3225_n1087# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0.54375 ps=4.04 w=3.75 l=15
X2 a_n29_n868# a_n3029_n965# a_n3087_n868# w_n3225_n1087# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=1.0875 ps=8.08 w=3.75 l=15
X3 a_3029_n868# a_29_n965# a_n29_n868# w_n3225_n1087# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0.54375 ps=4.04 w=3.75 l=15
.ends

.subckt sky130_fd_pr__pfet_01v8_XG6TDL a_n159_n426# a_111_431# a_33_n426# a_n221_n400#
+ a_n129_n400# a_63_n400# a_n81_431# w_n359_n619# a_n33_n400# a_159_n400#
X0 a_n129_n400# a_n159_n426# a_n221_n400# w_n359_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1 a_n33_n400# a_n81_431# a_n129_n400# w_n359_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2 a_159_n400# a_111_431# a_63_n400# w_n359_n619# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3 a_63_n400# a_33_n426# a_n33_n400# w_n359_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_F93ZEE a_209_n400# a_n29_n400# a_n209_n488# a_n401_n622#
+ a_n267_n400# a_29_n488#
X0 a_n29_n400# a_n209_n488# a_n267_n400# a_n401_n622# sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X1 a_209_n400# a_29_n488# a_n29_n400# a_n401_n622# sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
.ends

.subckt sky130_fd_pr__nfet_01v8_6EHS5V a_n227_n574# a_n125_n400# a_63_n400# a_n63_n426#
+ a_n33_n400#
X0 a_63_n400# a_n63_n426# a_n33_n400# a_n227_n574# sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1 a_n33_n400# a_n63_n426# a_n125_n400# a_n227_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_JFFQEL a_n90_n488# a_90_n400# a_n282_n622# a_n148_n400#
X0 a_90_n400# a_n90_n488# a_n148_n400# a_n282_n622# sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
.ends

.subckt bootstrap VDD VSS VIN SW_ON EN VGATE
Xx1 EN VSS VSS VDD VDD EN_Z sky130_fd_sc_hd__inv_4
Xx3 x3/A VSS VSS VDD VDD SW_ON sky130_fd_sc_hd__inv_4
Xx2 VGATE_1V8 VSS VSS VDD VDD x3/A sky130_fd_sc_hd__inv_2
Xsky130_fd_pr__pfet_01v8_7FRQHJ_0 Vtop Vbottom Vbottom Vtop Vtop Vbottom Vtop Vtop
+ Vtop Vbottom Vtop sky130_fd_pr__pfet_01v8_7FRQHJ
Xsky130_fd_pr__pfet_01v8_XG6TDL_0 EN_Z EN_Z EN_Z Vtop VGATE VGATE EN_Z Vtop Vtop Vtop
+ sky130_fd_pr__pfet_01v8_XG6TDL
XXM1 Vtop VDD Vtop VGATE sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 VGATE Vd VDD VSS VGATE VDD sky130_fd_pr__nfet_05v0_nvt_F93ZEE
XXM4 VSS VSS VSS EN_Z Vd sky130_fd_pr__nfet_01v8_6EHS5V
XXM5 VSS VSS VSS EN_Z Vbottom sky130_fd_pr__nfet_01v8_6EHS5V
XXM7 VDD VGATE_1V8 VSS VGATE sky130_fd_pr__nfet_05v0_nvt_JFFQEL
XXM8 VSS VIN VIN VGATE Vbottom sky130_fd_pr__nfet_01v8_6EHS5V
.ends

