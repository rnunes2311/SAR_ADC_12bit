magic
tech sky130A
magscale 1 2
timestamp 1711994487
<< nwell >>
rect -3254 -1219 3254 1219
<< pmoslvt >>
rect -3058 -1000 -1058 1000
rect -1000 -1000 1000 1000
rect 1058 -1000 3058 1000
<< pdiff >>
rect -3116 988 -3058 1000
rect -3116 -988 -3104 988
rect -3070 -988 -3058 988
rect -3116 -1000 -3058 -988
rect -1058 988 -1000 1000
rect -1058 -988 -1046 988
rect -1012 -988 -1000 988
rect -1058 -1000 -1000 -988
rect 1000 988 1058 1000
rect 1000 -988 1012 988
rect 1046 -988 1058 988
rect 1000 -1000 1058 -988
rect 3058 988 3116 1000
rect 3058 -988 3070 988
rect 3104 -988 3116 988
rect 3058 -1000 3116 -988
<< pdiffc >>
rect -3104 -988 -3070 988
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect 3070 -988 3104 988
<< nsubdiff >>
rect -3218 1149 -3122 1183
rect 3122 1149 3218 1183
rect -3218 1087 -3184 1149
rect 3184 1087 3218 1149
rect -3218 -1149 -3184 -1087
rect 3184 -1149 3218 -1087
rect -3218 -1183 -3122 -1149
rect 3122 -1183 3218 -1149
<< nsubdiffcont >>
rect -3122 1149 3122 1183
rect -3218 -1087 -3184 1087
rect 3184 -1087 3218 1087
rect -3122 -1183 3122 -1149
<< poly >>
rect -3058 1081 -1058 1097
rect -3058 1047 -3042 1081
rect -1074 1047 -1058 1081
rect -3058 1000 -1058 1047
rect -1000 1081 1000 1097
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1000 1000 1000 1047
rect 1058 1081 3058 1097
rect 1058 1047 1074 1081
rect 3042 1047 3058 1081
rect 1058 1000 3058 1047
rect -3058 -1047 -1058 -1000
rect -3058 -1081 -3042 -1047
rect -1074 -1081 -1058 -1047
rect -3058 -1097 -1058 -1081
rect -1000 -1047 1000 -1000
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1000 -1097 1000 -1081
rect 1058 -1047 3058 -1000
rect 1058 -1081 1074 -1047
rect 3042 -1081 3058 -1047
rect 1058 -1097 3058 -1081
<< polycont >>
rect -3042 1047 -1074 1081
rect -984 1047 984 1081
rect 1074 1047 3042 1081
rect -3042 -1081 -1074 -1047
rect -984 -1081 984 -1047
rect 1074 -1081 3042 -1047
<< locali >>
rect -3218 1149 -3122 1183
rect 3122 1149 3218 1183
rect -3218 1087 -3184 1149
rect 3184 1087 3218 1149
rect -3058 1047 -3042 1081
rect -1074 1047 -1058 1081
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect 1058 1047 1074 1081
rect 3042 1047 3058 1081
rect -3104 988 -3070 1004
rect -3104 -1004 -3070 -988
rect -1046 988 -1012 1004
rect -1046 -1004 -1012 -988
rect 1012 988 1046 1004
rect 1012 -1004 1046 -988
rect 3070 988 3104 1004
rect 3070 -1004 3104 -988
rect -3058 -1081 -3042 -1047
rect -1074 -1081 -1058 -1047
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect 1058 -1081 1074 -1047
rect 3042 -1081 3058 -1047
rect -3218 -1149 -3184 -1087
rect 3184 -1149 3218 -1087
rect -3218 -1183 -3122 -1149
rect 3122 -1183 3218 -1149
<< viali >>
rect -3042 1047 -1074 1081
rect -984 1047 984 1081
rect 1074 1047 3042 1081
rect -3104 -988 -3070 988
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect 3070 -988 3104 988
rect -3042 -1081 -1074 -1047
rect -984 -1081 984 -1047
rect 1074 -1081 3042 -1047
<< metal1 >>
rect -3054 1081 -1062 1087
rect -3054 1047 -3042 1081
rect -1074 1047 -1062 1081
rect -3054 1041 -1062 1047
rect -996 1081 996 1087
rect -996 1047 -984 1081
rect 984 1047 996 1081
rect -996 1041 996 1047
rect 1062 1081 3054 1087
rect 1062 1047 1074 1081
rect 3042 1047 3054 1081
rect 1062 1041 3054 1047
rect -3110 988 -3064 1000
rect -3110 -988 -3104 988
rect -3070 -988 -3064 988
rect -3110 -1000 -3064 -988
rect -1052 988 -1006 1000
rect -1052 -988 -1046 988
rect -1012 -988 -1006 988
rect -1052 -1000 -1006 -988
rect 1006 988 1052 1000
rect 1006 -988 1012 988
rect 1046 -988 1052 988
rect 1006 -1000 1052 -988
rect 3064 988 3110 1000
rect 3064 -988 3070 988
rect 3104 -988 3110 988
rect 3064 -1000 3110 -988
rect -3054 -1047 -1062 -1041
rect -3054 -1081 -3042 -1047
rect -1074 -1081 -1062 -1047
rect -3054 -1087 -1062 -1081
rect -996 -1047 996 -1041
rect -996 -1081 -984 -1047
rect 984 -1081 996 -1047
rect -996 -1087 996 -1081
rect 1062 -1047 3054 -1041
rect 1062 -1081 1074 -1047
rect 3042 -1081 3054 -1047
rect 1062 -1087 3054 -1081
<< properties >>
string FIXED_BBOX -3201 -1166 3201 1166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 10.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
