magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< error_p >>
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect -29 1159 29 1165
rect -29 689 29 695
rect -29 655 -17 689
rect -29 649 29 655
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect -29 -695 29 -689
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect -29 -1205 29 -1199
<< pwell >>
rect -211 -1337 211 1337
<< nmos >>
rect -15 727 15 1127
rect -15 109 15 509
rect -15 -509 15 -109
rect -15 -1127 15 -727
<< ndiff >>
rect -73 1115 -15 1127
rect -73 739 -61 1115
rect -27 739 -15 1115
rect -73 727 -15 739
rect 15 1115 73 1127
rect 15 739 27 1115
rect 61 739 73 1115
rect 15 727 73 739
rect -73 497 -15 509
rect -73 121 -61 497
rect -27 121 -15 497
rect -73 109 -15 121
rect 15 497 73 509
rect 15 121 27 497
rect 61 121 73 497
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -497 -61 -121
rect -27 -497 -15 -121
rect -73 -509 -15 -497
rect 15 -121 73 -109
rect 15 -497 27 -121
rect 61 -497 73 -121
rect 15 -509 73 -497
rect -73 -739 -15 -727
rect -73 -1115 -61 -739
rect -27 -1115 -15 -739
rect -73 -1127 -15 -1115
rect 15 -739 73 -727
rect 15 -1115 27 -739
rect 61 -1115 73 -739
rect 15 -1127 73 -1115
<< ndiffc >>
rect -61 739 -27 1115
rect 27 739 61 1115
rect -61 121 -27 497
rect 27 121 61 497
rect -61 -497 -27 -121
rect 27 -497 61 -121
rect -61 -1115 -27 -739
rect 27 -1115 61 -739
<< psubdiff >>
rect -175 1267 -79 1301
rect 79 1267 175 1301
rect -175 1205 -141 1267
rect 141 1205 175 1267
rect -175 -1267 -141 -1205
rect 141 -1267 175 -1205
rect -175 -1301 -79 -1267
rect 79 -1301 175 -1267
<< psubdiffcont >>
rect -79 1267 79 1301
rect -175 -1205 -141 1205
rect 141 -1205 175 1205
rect -79 -1301 79 -1267
<< poly >>
rect -33 1199 33 1215
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -33 1149 33 1165
rect -15 1127 15 1149
rect -15 705 15 727
rect -33 689 33 705
rect -33 655 -17 689
rect 17 655 33 689
rect -33 639 33 655
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -15 509 15 531
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -531 15 -509
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect -33 -655 33 -639
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -33 -705 33 -689
rect -15 -727 15 -705
rect -15 -1149 15 -1127
rect -33 -1165 33 -1149
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -33 -1215 33 -1199
<< polycont >>
rect -17 1165 17 1199
rect -17 655 17 689
rect -17 547 17 581
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -17 -1199 17 -1165
<< locali >>
rect -175 1267 -79 1301
rect 79 1267 175 1301
rect -175 1205 -141 1267
rect 141 1205 175 1267
rect -33 1165 -17 1199
rect 17 1165 33 1199
rect -61 1115 -27 1131
rect -61 723 -27 739
rect 27 1115 61 1131
rect 27 723 61 739
rect -33 655 -17 689
rect 17 655 33 689
rect -33 547 -17 581
rect 17 547 33 581
rect -61 497 -27 513
rect -61 105 -27 121
rect 27 497 61 513
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -513 -27 -497
rect 27 -121 61 -105
rect 27 -513 61 -497
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -61 -739 -27 -723
rect -61 -1131 -27 -1115
rect 27 -739 61 -723
rect 27 -1131 61 -1115
rect -33 -1199 -17 -1165
rect 17 -1199 33 -1165
rect -175 -1267 -141 -1205
rect 141 -1267 175 -1205
rect -175 -1301 -79 -1267
rect 79 -1301 175 -1267
<< viali >>
rect -17 1165 17 1199
rect -61 739 -27 1115
rect 27 739 61 1115
rect -17 655 17 689
rect -17 547 17 581
rect -61 121 -27 497
rect 27 121 61 497
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -497 -27 -121
rect 27 -497 61 -121
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -61 -1115 -27 -739
rect 27 -1115 61 -739
rect -17 -1199 17 -1165
<< metal1 >>
rect -29 1199 29 1205
rect -29 1165 -17 1199
rect 17 1165 29 1199
rect -29 1159 29 1165
rect -67 1115 -21 1127
rect -67 739 -61 1115
rect -27 739 -21 1115
rect -67 727 -21 739
rect 21 1115 67 1127
rect 21 739 27 1115
rect 61 739 67 1115
rect 21 727 67 739
rect -29 689 29 695
rect -29 655 -17 689
rect 17 655 29 689
rect -29 649 29 655
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -67 497 -21 509
rect -67 121 -61 497
rect -27 121 -21 497
rect -67 109 -21 121
rect 21 497 67 509
rect 21 121 27 497
rect 61 121 67 497
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -497 -61 -121
rect -27 -497 -21 -121
rect -67 -509 -21 -497
rect 21 -121 67 -109
rect 21 -497 27 -121
rect 61 -497 67 -121
rect 21 -509 67 -497
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect 17 -689 29 -655
rect -29 -695 29 -689
rect -67 -739 -21 -727
rect -67 -1115 -61 -739
rect -27 -1115 -21 -739
rect -67 -1127 -21 -1115
rect 21 -739 67 -727
rect 21 -1115 27 -739
rect 61 -1115 67 -739
rect 21 -1127 67 -1115
rect -29 -1165 29 -1159
rect -29 -1199 -17 -1165
rect 17 -1199 29 -1165
rect -29 -1205 29 -1199
<< properties >>
string FIXED_BBOX -158 -1284 158 1284
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
