magic
tech sky130A
magscale 1 2
timestamp 1711965631
<< pwell >>
rect -357 -308 357 308
<< nnmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< mvndiff >>
rect -187 38 -129 50
rect -187 -38 -175 38
rect -141 -38 -129 38
rect -187 -50 -129 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 129 38 187 50
rect 129 -38 141 38
rect 175 -38 187 38
rect 129 -50 187 -38
<< mvndiffc >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< mvpsubdiff >>
rect -321 260 321 272
rect -321 226 -213 260
rect 213 226 321 260
rect -321 214 321 226
rect -321 164 -263 214
rect -321 -164 -309 164
rect -275 -164 -263 164
rect 263 164 321 214
rect -321 -214 -263 -164
rect 263 -164 275 164
rect 309 -164 321 164
rect 263 -214 321 -164
rect -321 -226 321 -214
rect -321 -260 -213 -226
rect 213 -260 321 -226
rect -321 -272 321 -260
<< mvpsubdiffcont >>
rect -213 226 213 260
rect -309 -164 -275 164
rect 275 -164 309 164
rect -213 -260 213 -226
<< poly >>
rect -129 122 -29 138
rect -129 88 -113 122
rect -45 88 -29 122
rect -129 50 -29 88
rect 29 122 129 138
rect 29 88 45 122
rect 113 88 129 122
rect 29 50 129 88
rect -129 -88 -29 -50
rect -129 -122 -113 -88
rect -45 -122 -29 -88
rect -129 -138 -29 -122
rect 29 -88 129 -50
rect 29 -122 45 -88
rect 113 -122 129 -88
rect 29 -138 129 -122
<< polycont >>
rect -113 88 -45 122
rect 45 88 113 122
rect -113 -122 -45 -88
rect 45 -122 113 -88
<< locali >>
rect -309 226 -213 260
rect 213 226 309 260
rect -309 164 -275 226
rect 275 164 309 226
rect -129 88 -113 122
rect -45 88 -29 122
rect 29 88 45 122
rect 113 88 129 122
rect -175 38 -141 54
rect -175 -54 -141 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 141 38 175 54
rect 141 -54 175 -38
rect -129 -122 -113 -88
rect -45 -122 -29 -88
rect 29 -122 45 -88
rect 113 -122 129 -88
rect -309 -226 -275 -164
rect 275 -226 309 -164
rect -309 -260 -213 -226
rect 213 -260 309 -226
<< viali >>
rect -113 88 -45 122
rect 45 88 113 122
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
rect -113 -122 -45 -88
rect 45 -122 113 -88
<< metal1 >>
rect -125 122 -33 128
rect -125 88 -113 122
rect -45 88 -33 122
rect -125 82 -33 88
rect 33 122 125 128
rect 33 88 45 122
rect 113 88 125 122
rect 33 82 125 88
rect -181 38 -135 50
rect -181 -38 -175 38
rect -141 -38 -135 38
rect -181 -50 -135 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 135 38 181 50
rect 135 -38 141 38
rect 175 -38 181 38
rect 135 -50 181 -38
rect -125 -88 -33 -82
rect -125 -122 -113 -88
rect -45 -122 -33 -88
rect -125 -128 -33 -122
rect 33 -88 125 -82
rect 33 -122 45 -88
rect 113 -122 125 -88
rect 33 -128 125 -122
<< properties >>
string FIXED_BBOX -292 -243 292 243
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
