magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -372 1399 -314 1405
rect -176 1399 -118 1405
rect 20 1399 78 1405
rect 216 1399 274 1405
rect -372 1365 -360 1399
rect -176 1365 -164 1399
rect 20 1365 32 1399
rect 216 1365 228 1399
rect -372 1359 -314 1365
rect -176 1359 -118 1365
rect 20 1359 78 1365
rect 216 1359 274 1365
rect -274 71 -216 77
rect -78 71 -20 77
rect 118 71 176 77
rect 314 71 372 77
rect -274 37 -262 71
rect -78 37 -66 71
rect 118 37 130 71
rect 314 37 326 71
rect -274 31 -216 37
rect -78 31 -20 37
rect 118 31 176 37
rect 314 31 372 37
rect -274 -37 -216 -31
rect -78 -37 -20 -31
rect 118 -37 176 -31
rect 314 -37 372 -31
rect -274 -71 -262 -37
rect -78 -71 -66 -37
rect 118 -71 130 -37
rect 314 -71 326 -37
rect -274 -77 -216 -71
rect -78 -77 -20 -71
rect 118 -77 176 -71
rect 314 -77 372 -71
rect -372 -1365 -314 -1359
rect -176 -1365 -118 -1359
rect 20 -1365 78 -1359
rect 216 -1365 274 -1359
rect -372 -1399 -360 -1365
rect -176 -1399 -164 -1365
rect 20 -1399 32 -1365
rect 216 -1399 228 -1365
rect -372 -1405 -314 -1399
rect -176 -1405 -118 -1399
rect 20 -1405 78 -1399
rect 216 -1405 274 -1399
<< nwell >>
rect -559 -1537 559 1537
<< pmos >>
rect -363 118 -323 1318
rect -265 118 -225 1318
rect -167 118 -127 1318
rect -69 118 -29 1318
rect 29 118 69 1318
rect 127 118 167 1318
rect 225 118 265 1318
rect 323 118 363 1318
rect -363 -1318 -323 -118
rect -265 -1318 -225 -118
rect -167 -1318 -127 -118
rect -69 -1318 -29 -118
rect 29 -1318 69 -118
rect 127 -1318 167 -118
rect 225 -1318 265 -118
rect 323 -1318 363 -118
<< pdiff >>
rect -421 1306 -363 1318
rect -421 130 -409 1306
rect -375 130 -363 1306
rect -421 118 -363 130
rect -323 1306 -265 1318
rect -323 130 -311 1306
rect -277 130 -265 1306
rect -323 118 -265 130
rect -225 1306 -167 1318
rect -225 130 -213 1306
rect -179 130 -167 1306
rect -225 118 -167 130
rect -127 1306 -69 1318
rect -127 130 -115 1306
rect -81 130 -69 1306
rect -127 118 -69 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 69 1306 127 1318
rect 69 130 81 1306
rect 115 130 127 1306
rect 69 118 127 130
rect 167 1306 225 1318
rect 167 130 179 1306
rect 213 130 225 1306
rect 167 118 225 130
rect 265 1306 323 1318
rect 265 130 277 1306
rect 311 130 323 1306
rect 265 118 323 130
rect 363 1306 421 1318
rect 363 130 375 1306
rect 409 130 421 1306
rect 363 118 421 130
rect -421 -130 -363 -118
rect -421 -1306 -409 -130
rect -375 -1306 -363 -130
rect -421 -1318 -363 -1306
rect -323 -130 -265 -118
rect -323 -1306 -311 -130
rect -277 -1306 -265 -130
rect -323 -1318 -265 -1306
rect -225 -130 -167 -118
rect -225 -1306 -213 -130
rect -179 -1306 -167 -130
rect -225 -1318 -167 -1306
rect -127 -130 -69 -118
rect -127 -1306 -115 -130
rect -81 -1306 -69 -130
rect -127 -1318 -69 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 69 -130 127 -118
rect 69 -1306 81 -130
rect 115 -1306 127 -130
rect 69 -1318 127 -1306
rect 167 -130 225 -118
rect 167 -1306 179 -130
rect 213 -1306 225 -130
rect 167 -1318 225 -1306
rect 265 -130 323 -118
rect 265 -1306 277 -130
rect 311 -1306 323 -130
rect 265 -1318 323 -1306
rect 363 -130 421 -118
rect 363 -1306 375 -130
rect 409 -1306 421 -130
rect 363 -1318 421 -1306
<< pdiffc >>
rect -409 130 -375 1306
rect -311 130 -277 1306
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect 277 130 311 1306
rect 375 130 409 1306
rect -409 -1306 -375 -130
rect -311 -1306 -277 -130
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect 277 -1306 311 -130
rect 375 -1306 409 -130
<< nsubdiff >>
rect -523 1467 -427 1501
rect 427 1467 523 1501
rect -523 -1467 -489 1467
rect 489 1405 523 1467
rect 489 -1467 523 -1405
rect -523 -1501 -427 -1467
rect 427 -1501 523 -1467
<< nsubdiffcont >>
rect -427 1467 427 1501
rect 489 -1405 523 1405
rect -427 -1501 427 -1467
<< poly >>
rect -376 1399 -310 1415
rect -376 1365 -360 1399
rect -326 1365 -310 1399
rect -376 1349 -310 1365
rect -180 1399 -114 1415
rect -180 1365 -164 1399
rect -130 1365 -114 1399
rect -180 1349 -114 1365
rect 16 1399 82 1415
rect 16 1365 32 1399
rect 66 1365 82 1399
rect 16 1349 82 1365
rect 212 1399 278 1415
rect 212 1365 228 1399
rect 262 1365 278 1399
rect 212 1349 278 1365
rect -363 1318 -323 1349
rect -265 1318 -225 1344
rect -167 1318 -127 1349
rect -69 1318 -29 1344
rect 29 1318 69 1349
rect 127 1318 167 1344
rect 225 1318 265 1349
rect 323 1318 363 1344
rect -363 92 -323 118
rect -265 87 -225 118
rect -167 92 -127 118
rect -69 87 -29 118
rect 29 92 69 118
rect 127 87 167 118
rect 225 92 265 118
rect 323 87 363 118
rect -278 71 -212 87
rect -278 37 -262 71
rect -228 37 -212 71
rect -278 21 -212 37
rect -82 71 -16 87
rect -82 37 -66 71
rect -32 37 -16 71
rect -82 21 -16 37
rect 114 71 180 87
rect 114 37 130 71
rect 164 37 180 71
rect 114 21 180 37
rect 310 71 376 87
rect 310 37 326 71
rect 360 37 376 71
rect 310 21 376 37
rect -278 -37 -212 -21
rect -278 -71 -262 -37
rect -228 -71 -212 -37
rect -278 -87 -212 -71
rect -82 -37 -16 -21
rect -82 -71 -66 -37
rect -32 -71 -16 -37
rect -82 -87 -16 -71
rect 114 -37 180 -21
rect 114 -71 130 -37
rect 164 -71 180 -37
rect 114 -87 180 -71
rect 310 -37 376 -21
rect 310 -71 326 -37
rect 360 -71 376 -37
rect 310 -87 376 -71
rect -363 -118 -323 -92
rect -265 -118 -225 -87
rect -167 -118 -127 -92
rect -69 -118 -29 -87
rect 29 -118 69 -92
rect 127 -118 167 -87
rect 225 -118 265 -92
rect 323 -118 363 -87
rect -363 -1349 -323 -1318
rect -265 -1344 -225 -1318
rect -167 -1349 -127 -1318
rect -69 -1344 -29 -1318
rect 29 -1349 69 -1318
rect 127 -1344 167 -1318
rect 225 -1349 265 -1318
rect 323 -1344 363 -1318
rect -376 -1365 -310 -1349
rect -376 -1399 -360 -1365
rect -326 -1399 -310 -1365
rect -376 -1415 -310 -1399
rect -180 -1365 -114 -1349
rect -180 -1399 -164 -1365
rect -130 -1399 -114 -1365
rect -180 -1415 -114 -1399
rect 16 -1365 82 -1349
rect 16 -1399 32 -1365
rect 66 -1399 82 -1365
rect 16 -1415 82 -1399
rect 212 -1365 278 -1349
rect 212 -1399 228 -1365
rect 262 -1399 278 -1365
rect 212 -1415 278 -1399
<< polycont >>
rect -360 1365 -326 1399
rect -164 1365 -130 1399
rect 32 1365 66 1399
rect 228 1365 262 1399
rect -262 37 -228 71
rect -66 37 -32 71
rect 130 37 164 71
rect 326 37 360 71
rect -262 -71 -228 -37
rect -66 -71 -32 -37
rect 130 -71 164 -37
rect 326 -71 360 -37
rect -360 -1399 -326 -1365
rect -164 -1399 -130 -1365
rect 32 -1399 66 -1365
rect 228 -1399 262 -1365
<< locali >>
rect -523 1467 -427 1501
rect 427 1467 523 1501
rect -523 -1467 -489 1467
rect 489 1405 523 1467
rect -376 1365 -360 1399
rect -326 1365 -310 1399
rect -180 1365 -164 1399
rect -130 1365 -114 1399
rect 16 1365 32 1399
rect 66 1365 82 1399
rect 212 1365 228 1399
rect 262 1365 278 1399
rect -409 1306 -375 1322
rect -409 114 -375 130
rect -311 1306 -277 1322
rect -311 114 -277 130
rect -213 1306 -179 1322
rect -213 114 -179 130
rect -115 1306 -81 1322
rect -115 114 -81 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 81 1306 115 1322
rect 81 114 115 130
rect 179 1306 213 1322
rect 179 114 213 130
rect 277 1306 311 1322
rect 277 114 311 130
rect 375 1306 409 1322
rect 375 114 409 130
rect -278 37 -262 71
rect -228 37 -212 71
rect -82 37 -66 71
rect -32 37 -16 71
rect 114 37 130 71
rect 164 37 180 71
rect 310 37 326 71
rect 360 37 376 71
rect -278 -71 -262 -37
rect -228 -71 -212 -37
rect -82 -71 -66 -37
rect -32 -71 -16 -37
rect 114 -71 130 -37
rect 164 -71 180 -37
rect 310 -71 326 -37
rect 360 -71 376 -37
rect -409 -130 -375 -114
rect -409 -1322 -375 -1306
rect -311 -130 -277 -114
rect -311 -1322 -277 -1306
rect -213 -130 -179 -114
rect -213 -1322 -179 -1306
rect -115 -130 -81 -114
rect -115 -1322 -81 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 81 -130 115 -114
rect 81 -1322 115 -1306
rect 179 -130 213 -114
rect 179 -1322 213 -1306
rect 277 -130 311 -114
rect 277 -1322 311 -1306
rect 375 -130 409 -114
rect 375 -1322 409 -1306
rect -376 -1399 -360 -1365
rect -326 -1399 -310 -1365
rect -180 -1399 -164 -1365
rect -130 -1399 -114 -1365
rect 16 -1399 32 -1365
rect 66 -1399 82 -1365
rect 212 -1399 228 -1365
rect 262 -1399 278 -1365
rect 489 -1467 523 -1405
rect -523 -1501 -427 -1467
rect 427 -1501 523 -1467
<< viali >>
rect -360 1365 -326 1399
rect -164 1365 -130 1399
rect 32 1365 66 1399
rect 228 1365 262 1399
rect -409 130 -375 1306
rect -311 130 -277 1306
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect 277 130 311 1306
rect 375 130 409 1306
rect -262 37 -228 71
rect -66 37 -32 71
rect 130 37 164 71
rect 326 37 360 71
rect -262 -71 -228 -37
rect -66 -71 -32 -37
rect 130 -71 164 -37
rect 326 -71 360 -37
rect -409 -1306 -375 -130
rect -311 -1306 -277 -130
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect 277 -1306 311 -130
rect 375 -1306 409 -130
rect -360 -1399 -326 -1365
rect -164 -1399 -130 -1365
rect 32 -1399 66 -1365
rect 228 -1399 262 -1365
<< metal1 >>
rect -372 1399 -314 1405
rect -372 1365 -360 1399
rect -326 1365 -314 1399
rect -372 1359 -314 1365
rect -176 1399 -118 1405
rect -176 1365 -164 1399
rect -130 1365 -118 1399
rect -176 1359 -118 1365
rect 20 1399 78 1405
rect 20 1365 32 1399
rect 66 1365 78 1399
rect 20 1359 78 1365
rect 216 1399 274 1405
rect 216 1365 228 1399
rect 262 1365 274 1399
rect 216 1359 274 1365
rect -415 1306 -369 1318
rect -415 130 -409 1306
rect -375 130 -369 1306
rect -415 118 -369 130
rect -317 1306 -271 1318
rect -317 130 -311 1306
rect -277 130 -271 1306
rect -317 118 -271 130
rect -219 1306 -173 1318
rect -219 130 -213 1306
rect -179 130 -173 1306
rect -219 118 -173 130
rect -121 1306 -75 1318
rect -121 130 -115 1306
rect -81 130 -75 1306
rect -121 118 -75 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 75 1306 121 1318
rect 75 130 81 1306
rect 115 130 121 1306
rect 75 118 121 130
rect 173 1306 219 1318
rect 173 130 179 1306
rect 213 130 219 1306
rect 173 118 219 130
rect 271 1306 317 1318
rect 271 130 277 1306
rect 311 130 317 1306
rect 271 118 317 130
rect 369 1306 415 1318
rect 369 130 375 1306
rect 409 130 415 1306
rect 369 118 415 130
rect -274 71 -216 77
rect -274 37 -262 71
rect -228 37 -216 71
rect -274 31 -216 37
rect -78 71 -20 77
rect -78 37 -66 71
rect -32 37 -20 71
rect -78 31 -20 37
rect 118 71 176 77
rect 118 37 130 71
rect 164 37 176 71
rect 118 31 176 37
rect 314 71 372 77
rect 314 37 326 71
rect 360 37 372 71
rect 314 31 372 37
rect -274 -37 -216 -31
rect -274 -71 -262 -37
rect -228 -71 -216 -37
rect -274 -77 -216 -71
rect -78 -37 -20 -31
rect -78 -71 -66 -37
rect -32 -71 -20 -37
rect -78 -77 -20 -71
rect 118 -37 176 -31
rect 118 -71 130 -37
rect 164 -71 176 -37
rect 118 -77 176 -71
rect 314 -37 372 -31
rect 314 -71 326 -37
rect 360 -71 372 -37
rect 314 -77 372 -71
rect -415 -130 -369 -118
rect -415 -1306 -409 -130
rect -375 -1306 -369 -130
rect -415 -1318 -369 -1306
rect -317 -130 -271 -118
rect -317 -1306 -311 -130
rect -277 -1306 -271 -130
rect -317 -1318 -271 -1306
rect -219 -130 -173 -118
rect -219 -1306 -213 -130
rect -179 -1306 -173 -130
rect -219 -1318 -173 -1306
rect -121 -130 -75 -118
rect -121 -1306 -115 -130
rect -81 -1306 -75 -130
rect -121 -1318 -75 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 75 -130 121 -118
rect 75 -1306 81 -130
rect 115 -1306 121 -130
rect 75 -1318 121 -1306
rect 173 -130 219 -118
rect 173 -1306 179 -130
rect 213 -1306 219 -130
rect 173 -1318 219 -1306
rect 271 -130 317 -118
rect 271 -1306 277 -130
rect 311 -1306 317 -130
rect 271 -1318 317 -1306
rect 369 -130 415 -118
rect 369 -1306 375 -130
rect 409 -1306 415 -130
rect 369 -1318 415 -1306
rect -372 -1365 -314 -1359
rect -372 -1399 -360 -1365
rect -326 -1399 -314 -1365
rect -372 -1405 -314 -1399
rect -176 -1365 -118 -1359
rect -176 -1399 -164 -1365
rect -130 -1399 -118 -1365
rect -176 -1405 -118 -1399
rect 20 -1365 78 -1359
rect 20 -1399 32 -1365
rect 66 -1399 78 -1365
rect 20 -1405 78 -1399
rect 216 -1365 274 -1359
rect 216 -1399 228 -1365
rect 262 -1399 274 -1365
rect 216 -1405 274 -1399
<< properties >>
string FIXED_BBOX -506 -1484 506 1484
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.2 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
