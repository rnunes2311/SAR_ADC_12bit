magic
tech sky130A
magscale 1 2
timestamp 1711308867
<< pwell >>
rect -201 -1832 201 1832
<< psubdiff >>
rect -165 1762 -69 1796
rect 69 1762 165 1796
rect -165 1700 -131 1762
rect -165 -1762 -131 -1700
rect 131 -1762 165 1762
rect -165 -1796 -69 -1762
rect 69 -1796 165 -1762
<< psubdiffcont >>
rect -69 1762 69 1796
rect -165 -1700 -131 1700
rect -69 -1796 69 -1762
<< xpolycontact >>
rect -35 1234 35 1666
rect -35 -1666 35 -1234
<< ppolyres >>
rect -35 -1234 35 1234
<< locali >>
rect -85 1762 -69 1796
rect 69 1762 85 1796
rect -165 1700 -131 1716
rect -165 -1716 -131 -1700
rect -85 -1796 -69 -1762
rect 69 -1796 85 -1762
<< viali >>
rect -19 1251 19 1648
rect -19 -1648 19 -1251
<< metal1 >>
rect -25 1648 25 1660
rect -25 1251 -19 1648
rect 19 1251 25 1648
rect -25 1239 25 1251
rect -25 -1251 25 -1239
rect -25 -1648 -19 -1251
rect 19 -1648 25 -1251
rect -25 -1660 25 -1648
<< properties >>
string FIXED_BBOX -148 -1779 148 1779
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 12.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 12.534k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 0 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
