magic
tech sky130A
timestamp 1711813427
<< error_p >>
rect -172 136 -143 139
rect 38 136 67 139
rect 248 136 277 139
rect -172 119 -166 136
rect 38 119 44 136
rect 248 119 254 136
rect -172 116 -143 119
rect 38 116 67 119
rect 248 116 277 119
rect -277 -119 -248 -116
rect -67 -119 -38 -116
rect 143 -119 172 -116
rect -277 -136 -271 -119
rect -67 -136 -61 -119
rect 143 -136 149 -119
rect -277 -139 -248 -136
rect -67 -139 -38 -136
rect 143 -139 172 -136
<< nmos >>
rect -270 -100 -255 100
rect -165 -100 -150 100
rect -60 -100 -45 100
rect 45 -100 60 100
rect 150 -100 165 100
rect 255 -100 270 100
<< ndiff >>
rect -301 94 -270 100
rect -301 -94 -295 94
rect -278 -94 -270 94
rect -301 -100 -270 -94
rect -255 94 -224 100
rect -255 -94 -247 94
rect -230 -94 -224 94
rect -255 -100 -224 -94
rect -196 94 -165 100
rect -196 -94 -190 94
rect -173 -94 -165 94
rect -196 -100 -165 -94
rect -150 94 -119 100
rect -150 -94 -142 94
rect -125 -94 -119 94
rect -150 -100 -119 -94
rect -91 94 -60 100
rect -91 -94 -85 94
rect -68 -94 -60 94
rect -91 -100 -60 -94
rect -45 94 -14 100
rect -45 -94 -37 94
rect -20 -94 -14 94
rect -45 -100 -14 -94
rect 14 94 45 100
rect 14 -94 20 94
rect 37 -94 45 94
rect 14 -100 45 -94
rect 60 94 91 100
rect 60 -94 68 94
rect 85 -94 91 94
rect 60 -100 91 -94
rect 119 94 150 100
rect 119 -94 125 94
rect 142 -94 150 94
rect 119 -100 150 -94
rect 165 94 196 100
rect 165 -94 173 94
rect 190 -94 196 94
rect 165 -100 196 -94
rect 224 94 255 100
rect 224 -94 230 94
rect 247 -94 255 94
rect 224 -100 255 -94
rect 270 94 301 100
rect 270 -94 278 94
rect 295 -94 301 94
rect 270 -100 301 -94
<< ndiffc >>
rect -295 -94 -278 94
rect -247 -94 -230 94
rect -190 -94 -173 94
rect -142 -94 -125 94
rect -85 -94 -68 94
rect -37 -94 -20 94
rect 20 -94 37 94
rect 68 -94 85 94
rect 125 -94 142 94
rect 173 -94 190 94
rect 230 -94 247 94
rect 278 -94 295 94
<< poly >>
rect -174 136 -141 144
rect -174 119 -166 136
rect -149 119 -141 136
rect -270 100 -255 113
rect -174 111 -141 119
rect 36 136 69 144
rect 36 119 44 136
rect 61 119 69 136
rect -165 100 -150 111
rect -60 100 -45 113
rect 36 111 69 119
rect 246 136 279 144
rect 246 119 254 136
rect 271 119 279 136
rect 45 100 60 111
rect 150 100 165 113
rect 246 111 279 119
rect 255 100 270 111
rect -270 -111 -255 -100
rect -279 -119 -246 -111
rect -165 -113 -150 -100
rect -60 -111 -45 -100
rect -279 -136 -271 -119
rect -254 -136 -246 -119
rect -279 -144 -246 -136
rect -69 -119 -36 -111
rect 45 -113 60 -100
rect 150 -111 165 -100
rect -69 -136 -61 -119
rect -44 -136 -36 -119
rect -69 -144 -36 -136
rect 141 -119 174 -111
rect 255 -113 270 -100
rect 141 -136 149 -119
rect 166 -136 174 -119
rect 141 -144 174 -136
<< polycont >>
rect -166 119 -149 136
rect 44 119 61 136
rect 254 119 271 136
rect -271 -136 -254 -119
rect -61 -136 -44 -119
rect 149 -136 166 -119
<< locali >>
rect -174 119 -166 136
rect -149 119 -141 136
rect 36 119 44 136
rect 61 119 69 136
rect 246 119 254 136
rect 271 119 279 136
rect -295 94 -278 102
rect -295 -102 -278 -94
rect -247 94 -230 102
rect -247 -102 -230 -94
rect -190 94 -173 102
rect -190 -102 -173 -94
rect -142 94 -125 102
rect -142 -102 -125 -94
rect -85 94 -68 102
rect -85 -102 -68 -94
rect -37 94 -20 102
rect -37 -102 -20 -94
rect 20 94 37 102
rect 20 -102 37 -94
rect 68 94 85 102
rect 68 -102 85 -94
rect 125 94 142 102
rect 125 -102 142 -94
rect 173 94 190 102
rect 173 -102 190 -94
rect 230 94 247 102
rect 230 -102 247 -94
rect 278 94 295 102
rect 278 -102 295 -94
rect -279 -136 -271 -119
rect -254 -136 -246 -119
rect -69 -136 -61 -119
rect -44 -136 -36 -119
rect 141 -136 149 -119
rect 166 -136 174 -119
<< viali >>
rect -166 119 -149 136
rect 44 119 61 136
rect 254 119 271 136
rect -295 -94 -278 94
rect -247 -94 -230 94
rect -190 -94 -173 94
rect -142 -94 -125 94
rect -85 -94 -68 94
rect -37 -94 -20 94
rect 20 -94 37 94
rect 68 -94 85 94
rect 125 -94 142 94
rect 173 -94 190 94
rect 230 -94 247 94
rect 278 -94 295 94
rect -271 -136 -254 -119
rect -61 -136 -44 -119
rect 149 -136 166 -119
<< metal1 >>
rect -172 136 -143 139
rect -172 119 -166 136
rect -149 119 -143 136
rect -172 116 -143 119
rect 38 136 67 139
rect 38 119 44 136
rect 61 119 67 136
rect 38 116 67 119
rect 248 136 277 139
rect 248 119 254 136
rect 271 119 277 136
rect 248 116 277 119
rect -298 94 -275 100
rect -298 -94 -295 94
rect -278 -94 -275 94
rect -298 -100 -275 -94
rect -250 94 -227 100
rect -250 -94 -247 94
rect -230 -94 -227 94
rect -250 -100 -227 -94
rect -193 94 -170 100
rect -193 -94 -190 94
rect -173 -94 -170 94
rect -193 -100 -170 -94
rect -145 94 -122 100
rect -145 -94 -142 94
rect -125 -94 -122 94
rect -145 -100 -122 -94
rect -88 94 -65 100
rect -88 -94 -85 94
rect -68 -94 -65 94
rect -88 -100 -65 -94
rect -40 94 -17 100
rect -40 -94 -37 94
rect -20 -94 -17 94
rect -40 -100 -17 -94
rect 17 94 40 100
rect 17 -94 20 94
rect 37 -94 40 94
rect 17 -100 40 -94
rect 65 94 88 100
rect 65 -94 68 94
rect 85 -94 88 94
rect 65 -100 88 -94
rect 122 94 145 100
rect 122 -94 125 94
rect 142 -94 145 94
rect 122 -100 145 -94
rect 170 94 193 100
rect 170 -94 173 94
rect 190 -94 193 94
rect 170 -100 193 -94
rect 227 94 250 100
rect 227 -94 230 94
rect 247 -94 250 94
rect 227 -100 250 -94
rect 275 94 298 100
rect 275 -94 278 94
rect 295 -94 298 94
rect 275 -100 298 -94
rect -277 -119 -248 -116
rect -277 -136 -271 -119
rect -254 -136 -248 -119
rect -277 -139 -248 -136
rect -67 -119 -38 -116
rect -67 -136 -61 -119
rect -44 -136 -38 -119
rect -67 -139 -38 -136
rect 143 -119 172 -116
rect 143 -136 149 -119
rect 166 -136 172 -119
rect 143 -139 172 -136
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
