magic
tech sky130A
magscale 1 2
timestamp 1711969435
<< pwell >>
rect -357 -277 357 277
<< nnmos >>
rect -129 -19 -29 81
rect 29 -19 129 81
<< mvndiff >>
rect -187 69 -129 81
rect -187 -7 -175 69
rect -141 -7 -129 69
rect -187 -19 -129 -7
rect -29 69 29 81
rect -29 -7 -17 69
rect 17 -7 29 69
rect -29 -19 29 -7
rect 129 69 187 81
rect 129 -7 141 69
rect 175 -7 187 69
rect 129 -19 187 -7
<< mvndiffc >>
rect -175 -7 -141 69
rect -17 -7 17 69
rect 141 -7 175 69
<< mvpsubdiff >>
rect -321 229 321 241
rect -321 195 -213 229
rect 213 195 321 229
rect -321 183 321 195
rect -321 133 -263 183
rect -321 -133 -309 133
rect -275 -133 -263 133
rect 263 133 321 183
rect -321 -183 -263 -133
rect 263 -133 275 133
rect 309 -133 321 133
rect 263 -183 321 -133
rect -321 -195 321 -183
rect -321 -229 -213 -195
rect 213 -229 321 -195
rect -321 -241 321 -229
<< mvpsubdiffcont >>
rect -213 195 213 229
rect -309 -133 -275 133
rect 275 -133 309 133
rect -213 -229 213 -195
<< poly >>
rect -129 81 -29 107
rect 29 81 129 107
rect -129 -57 -29 -19
rect -129 -91 -113 -57
rect -45 -91 -29 -57
rect -129 -107 -29 -91
rect 29 -57 129 -19
rect 29 -91 45 -57
rect 113 -91 129 -57
rect 29 -107 129 -91
<< polycont >>
rect -113 -91 -45 -57
rect 45 -91 113 -57
<< locali >>
rect -309 195 -213 229
rect 213 195 309 229
rect -309 133 -275 195
rect 275 133 309 195
rect -175 69 -141 85
rect -175 -23 -141 -7
rect -17 69 17 85
rect -17 -23 17 -7
rect 141 69 175 85
rect 141 -23 175 -7
rect -129 -91 -113 -57
rect -45 -91 -29 -57
rect 29 -91 45 -57
rect 113 -91 129 -57
rect -309 -195 -275 -133
rect 275 -195 309 -133
rect -309 -229 -213 -195
rect 213 -229 309 -195
<< viali >>
rect -175 -7 -141 69
rect -17 -7 17 69
rect 141 -7 175 69
rect -113 -91 -45 -57
rect 45 -91 113 -57
<< metal1 >>
rect -181 69 -135 81
rect -181 -7 -175 69
rect -141 -7 -135 69
rect -181 -19 -135 -7
rect -23 69 23 81
rect -23 -7 -17 69
rect 17 -7 23 69
rect -23 -19 23 -7
rect 135 69 181 81
rect 135 -7 141 69
rect 175 -7 181 69
rect 135 -19 181 -7
rect -125 -57 -33 -51
rect -125 -91 -113 -57
rect -45 -91 -33 -57
rect -125 -97 -33 -91
rect 33 -57 125 -51
rect 33 -91 45 -57
rect 113 -91 125 -57
rect 33 -97 125 -91
<< properties >>
string FIXED_BBOX -292 -212 292 212
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
