magic
tech sky130A
magscale 1 2
timestamp 1711964565
<< nwell >>
rect -1878 -1019 1878 1019
<< pmos >>
rect -1682 -800 -1582 800
rect -1410 -800 -1310 800
rect -1138 -800 -1038 800
rect -866 -800 -766 800
rect -594 -800 -494 800
rect -322 -800 -222 800
rect -50 -800 50 800
rect 222 -800 322 800
rect 494 -800 594 800
rect 766 -800 866 800
rect 1038 -800 1138 800
rect 1310 -800 1410 800
rect 1582 -800 1682 800
<< pdiff >>
rect -1740 788 -1682 800
rect -1740 -788 -1728 788
rect -1694 -788 -1682 788
rect -1740 -800 -1682 -788
rect -1582 788 -1524 800
rect -1582 -788 -1570 788
rect -1536 -788 -1524 788
rect -1582 -800 -1524 -788
rect -1468 788 -1410 800
rect -1468 -788 -1456 788
rect -1422 -788 -1410 788
rect -1468 -800 -1410 -788
rect -1310 788 -1252 800
rect -1310 -788 -1298 788
rect -1264 -788 -1252 788
rect -1310 -800 -1252 -788
rect -1196 788 -1138 800
rect -1196 -788 -1184 788
rect -1150 -788 -1138 788
rect -1196 -800 -1138 -788
rect -1038 788 -980 800
rect -1038 -788 -1026 788
rect -992 -788 -980 788
rect -1038 -800 -980 -788
rect -924 788 -866 800
rect -924 -788 -912 788
rect -878 -788 -866 788
rect -924 -800 -866 -788
rect -766 788 -708 800
rect -766 -788 -754 788
rect -720 -788 -708 788
rect -766 -800 -708 -788
rect -652 788 -594 800
rect -652 -788 -640 788
rect -606 -788 -594 788
rect -652 -800 -594 -788
rect -494 788 -436 800
rect -494 -788 -482 788
rect -448 -788 -436 788
rect -494 -800 -436 -788
rect -380 788 -322 800
rect -380 -788 -368 788
rect -334 -788 -322 788
rect -380 -800 -322 -788
rect -222 788 -164 800
rect -222 -788 -210 788
rect -176 -788 -164 788
rect -222 -800 -164 -788
rect -108 788 -50 800
rect -108 -788 -96 788
rect -62 -788 -50 788
rect -108 -800 -50 -788
rect 50 788 108 800
rect 50 -788 62 788
rect 96 -788 108 788
rect 50 -800 108 -788
rect 164 788 222 800
rect 164 -788 176 788
rect 210 -788 222 788
rect 164 -800 222 -788
rect 322 788 380 800
rect 322 -788 334 788
rect 368 -788 380 788
rect 322 -800 380 -788
rect 436 788 494 800
rect 436 -788 448 788
rect 482 -788 494 788
rect 436 -800 494 -788
rect 594 788 652 800
rect 594 -788 606 788
rect 640 -788 652 788
rect 594 -800 652 -788
rect 708 788 766 800
rect 708 -788 720 788
rect 754 -788 766 788
rect 708 -800 766 -788
rect 866 788 924 800
rect 866 -788 878 788
rect 912 -788 924 788
rect 866 -800 924 -788
rect 980 788 1038 800
rect 980 -788 992 788
rect 1026 -788 1038 788
rect 980 -800 1038 -788
rect 1138 788 1196 800
rect 1138 -788 1150 788
rect 1184 -788 1196 788
rect 1138 -800 1196 -788
rect 1252 788 1310 800
rect 1252 -788 1264 788
rect 1298 -788 1310 788
rect 1252 -800 1310 -788
rect 1410 788 1468 800
rect 1410 -788 1422 788
rect 1456 -788 1468 788
rect 1410 -800 1468 -788
rect 1524 788 1582 800
rect 1524 -788 1536 788
rect 1570 -788 1582 788
rect 1524 -800 1582 -788
rect 1682 788 1740 800
rect 1682 -788 1694 788
rect 1728 -788 1740 788
rect 1682 -800 1740 -788
<< pdiffc >>
rect -1728 -788 -1694 788
rect -1570 -788 -1536 788
rect -1456 -788 -1422 788
rect -1298 -788 -1264 788
rect -1184 -788 -1150 788
rect -1026 -788 -992 788
rect -912 -788 -878 788
rect -754 -788 -720 788
rect -640 -788 -606 788
rect -482 -788 -448 788
rect -368 -788 -334 788
rect -210 -788 -176 788
rect -96 -788 -62 788
rect 62 -788 96 788
rect 176 -788 210 788
rect 334 -788 368 788
rect 448 -788 482 788
rect 606 -788 640 788
rect 720 -788 754 788
rect 878 -788 912 788
rect 992 -788 1026 788
rect 1150 -788 1184 788
rect 1264 -788 1298 788
rect 1422 -788 1456 788
rect 1536 -788 1570 788
rect 1694 -788 1728 788
<< nsubdiff >>
rect -1842 949 -1746 983
rect 1746 949 1842 983
rect -1842 887 -1808 949
rect 1808 887 1842 949
rect -1842 -949 -1808 -887
rect 1808 -949 1842 -887
rect -1842 -983 -1746 -949
rect 1746 -983 1842 -949
<< nsubdiffcont >>
rect -1746 949 1746 983
rect -1842 -887 -1808 887
rect 1808 -887 1842 887
rect -1746 -983 1746 -949
<< poly >>
rect -1682 881 -1582 897
rect -1682 847 -1666 881
rect -1598 847 -1582 881
rect -1682 800 -1582 847
rect -1410 881 -1310 897
rect -1410 847 -1394 881
rect -1326 847 -1310 881
rect -1410 800 -1310 847
rect -1138 881 -1038 897
rect -1138 847 -1122 881
rect -1054 847 -1038 881
rect -1138 800 -1038 847
rect -866 881 -766 897
rect -866 847 -850 881
rect -782 847 -766 881
rect -866 800 -766 847
rect -594 881 -494 897
rect -594 847 -578 881
rect -510 847 -494 881
rect -594 800 -494 847
rect -322 881 -222 897
rect -322 847 -306 881
rect -238 847 -222 881
rect -322 800 -222 847
rect -50 881 50 897
rect -50 847 -34 881
rect 34 847 50 881
rect -50 800 50 847
rect 222 881 322 897
rect 222 847 238 881
rect 306 847 322 881
rect 222 800 322 847
rect 494 881 594 897
rect 494 847 510 881
rect 578 847 594 881
rect 494 800 594 847
rect 766 881 866 897
rect 766 847 782 881
rect 850 847 866 881
rect 766 800 866 847
rect 1038 881 1138 897
rect 1038 847 1054 881
rect 1122 847 1138 881
rect 1038 800 1138 847
rect 1310 881 1410 897
rect 1310 847 1326 881
rect 1394 847 1410 881
rect 1310 800 1410 847
rect 1582 881 1682 897
rect 1582 847 1598 881
rect 1666 847 1682 881
rect 1582 800 1682 847
rect -1682 -847 -1582 -800
rect -1682 -881 -1666 -847
rect -1598 -881 -1582 -847
rect -1682 -897 -1582 -881
rect -1410 -847 -1310 -800
rect -1410 -881 -1394 -847
rect -1326 -881 -1310 -847
rect -1410 -897 -1310 -881
rect -1138 -847 -1038 -800
rect -1138 -881 -1122 -847
rect -1054 -881 -1038 -847
rect -1138 -897 -1038 -881
rect -866 -847 -766 -800
rect -866 -881 -850 -847
rect -782 -881 -766 -847
rect -866 -897 -766 -881
rect -594 -847 -494 -800
rect -594 -881 -578 -847
rect -510 -881 -494 -847
rect -594 -897 -494 -881
rect -322 -847 -222 -800
rect -322 -881 -306 -847
rect -238 -881 -222 -847
rect -322 -897 -222 -881
rect -50 -847 50 -800
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect -50 -897 50 -881
rect 222 -847 322 -800
rect 222 -881 238 -847
rect 306 -881 322 -847
rect 222 -897 322 -881
rect 494 -847 594 -800
rect 494 -881 510 -847
rect 578 -881 594 -847
rect 494 -897 594 -881
rect 766 -847 866 -800
rect 766 -881 782 -847
rect 850 -881 866 -847
rect 766 -897 866 -881
rect 1038 -847 1138 -800
rect 1038 -881 1054 -847
rect 1122 -881 1138 -847
rect 1038 -897 1138 -881
rect 1310 -847 1410 -800
rect 1310 -881 1326 -847
rect 1394 -881 1410 -847
rect 1310 -897 1410 -881
rect 1582 -847 1682 -800
rect 1582 -881 1598 -847
rect 1666 -881 1682 -847
rect 1582 -897 1682 -881
<< polycont >>
rect -1666 847 -1598 881
rect -1394 847 -1326 881
rect -1122 847 -1054 881
rect -850 847 -782 881
rect -578 847 -510 881
rect -306 847 -238 881
rect -34 847 34 881
rect 238 847 306 881
rect 510 847 578 881
rect 782 847 850 881
rect 1054 847 1122 881
rect 1326 847 1394 881
rect 1598 847 1666 881
rect -1666 -881 -1598 -847
rect -1394 -881 -1326 -847
rect -1122 -881 -1054 -847
rect -850 -881 -782 -847
rect -578 -881 -510 -847
rect -306 -881 -238 -847
rect -34 -881 34 -847
rect 238 -881 306 -847
rect 510 -881 578 -847
rect 782 -881 850 -847
rect 1054 -881 1122 -847
rect 1326 -881 1394 -847
rect 1598 -881 1666 -847
<< locali >>
rect -1842 949 -1746 983
rect 1746 949 1842 983
rect -1842 887 -1808 949
rect 1808 887 1842 949
rect -1682 847 -1666 881
rect -1598 847 -1582 881
rect -1410 847 -1394 881
rect -1326 847 -1310 881
rect -1138 847 -1122 881
rect -1054 847 -1038 881
rect -866 847 -850 881
rect -782 847 -766 881
rect -594 847 -578 881
rect -510 847 -494 881
rect -322 847 -306 881
rect -238 847 -222 881
rect -50 847 -34 881
rect 34 847 50 881
rect 222 847 238 881
rect 306 847 322 881
rect 494 847 510 881
rect 578 847 594 881
rect 766 847 782 881
rect 850 847 866 881
rect 1038 847 1054 881
rect 1122 847 1138 881
rect 1310 847 1326 881
rect 1394 847 1410 881
rect 1582 847 1598 881
rect 1666 847 1682 881
rect -1728 788 -1694 804
rect -1728 -804 -1694 -788
rect -1570 788 -1536 804
rect -1570 -804 -1536 -788
rect -1456 788 -1422 804
rect -1456 -804 -1422 -788
rect -1298 788 -1264 804
rect -1298 -804 -1264 -788
rect -1184 788 -1150 804
rect -1184 -804 -1150 -788
rect -1026 788 -992 804
rect -1026 -804 -992 -788
rect -912 788 -878 804
rect -912 -804 -878 -788
rect -754 788 -720 804
rect -754 -804 -720 -788
rect -640 788 -606 804
rect -640 -804 -606 -788
rect -482 788 -448 804
rect -482 -804 -448 -788
rect -368 788 -334 804
rect -368 -804 -334 -788
rect -210 788 -176 804
rect -210 -804 -176 -788
rect -96 788 -62 804
rect -96 -804 -62 -788
rect 62 788 96 804
rect 62 -804 96 -788
rect 176 788 210 804
rect 176 -804 210 -788
rect 334 788 368 804
rect 334 -804 368 -788
rect 448 788 482 804
rect 448 -804 482 -788
rect 606 788 640 804
rect 606 -804 640 -788
rect 720 788 754 804
rect 720 -804 754 -788
rect 878 788 912 804
rect 878 -804 912 -788
rect 992 788 1026 804
rect 992 -804 1026 -788
rect 1150 788 1184 804
rect 1150 -804 1184 -788
rect 1264 788 1298 804
rect 1264 -804 1298 -788
rect 1422 788 1456 804
rect 1422 -804 1456 -788
rect 1536 788 1570 804
rect 1536 -804 1570 -788
rect 1694 788 1728 804
rect 1694 -804 1728 -788
rect -1682 -881 -1666 -847
rect -1598 -881 -1582 -847
rect -1410 -881 -1394 -847
rect -1326 -881 -1310 -847
rect -1138 -881 -1122 -847
rect -1054 -881 -1038 -847
rect -866 -881 -850 -847
rect -782 -881 -766 -847
rect -594 -881 -578 -847
rect -510 -881 -494 -847
rect -322 -881 -306 -847
rect -238 -881 -222 -847
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect 222 -881 238 -847
rect 306 -881 322 -847
rect 494 -881 510 -847
rect 578 -881 594 -847
rect 766 -881 782 -847
rect 850 -881 866 -847
rect 1038 -881 1054 -847
rect 1122 -881 1138 -847
rect 1310 -881 1326 -847
rect 1394 -881 1410 -847
rect 1582 -881 1598 -847
rect 1666 -881 1682 -847
rect -1842 -949 -1808 -887
rect 1808 -949 1842 -887
rect -1842 -983 -1746 -949
rect 1746 -983 1842 -949
<< viali >>
rect -1666 847 -1598 881
rect -1394 847 -1326 881
rect -1122 847 -1054 881
rect -850 847 -782 881
rect -578 847 -510 881
rect -306 847 -238 881
rect -34 847 34 881
rect 238 847 306 881
rect 510 847 578 881
rect 782 847 850 881
rect 1054 847 1122 881
rect 1326 847 1394 881
rect 1598 847 1666 881
rect -1728 -788 -1694 788
rect -1570 -788 -1536 788
rect -1456 -788 -1422 788
rect -1298 -788 -1264 788
rect -1184 -788 -1150 788
rect -1026 -788 -992 788
rect -912 -788 -878 788
rect -754 -788 -720 788
rect -640 -788 -606 788
rect -482 -788 -448 788
rect -368 -788 -334 788
rect -210 -788 -176 788
rect -96 -788 -62 788
rect 62 -788 96 788
rect 176 -788 210 788
rect 334 -788 368 788
rect 448 -788 482 788
rect 606 -788 640 788
rect 720 -788 754 788
rect 878 -788 912 788
rect 992 -788 1026 788
rect 1150 -788 1184 788
rect 1264 -788 1298 788
rect 1422 -788 1456 788
rect 1536 -788 1570 788
rect 1694 -788 1728 788
rect -1666 -881 -1598 -847
rect -1394 -881 -1326 -847
rect -1122 -881 -1054 -847
rect -850 -881 -782 -847
rect -578 -881 -510 -847
rect -306 -881 -238 -847
rect -34 -881 34 -847
rect 238 -881 306 -847
rect 510 -881 578 -847
rect 782 -881 850 -847
rect 1054 -881 1122 -847
rect 1326 -881 1394 -847
rect 1598 -881 1666 -847
<< metal1 >>
rect -1678 881 -1586 887
rect -1678 847 -1666 881
rect -1598 847 -1586 881
rect -1678 841 -1586 847
rect -1406 881 -1314 887
rect -1406 847 -1394 881
rect -1326 847 -1314 881
rect -1406 841 -1314 847
rect -1134 881 -1042 887
rect -1134 847 -1122 881
rect -1054 847 -1042 881
rect -1134 841 -1042 847
rect -862 881 -770 887
rect -862 847 -850 881
rect -782 847 -770 881
rect -862 841 -770 847
rect -590 881 -498 887
rect -590 847 -578 881
rect -510 847 -498 881
rect -590 841 -498 847
rect -318 881 -226 887
rect -318 847 -306 881
rect -238 847 -226 881
rect -318 841 -226 847
rect -46 881 46 887
rect -46 847 -34 881
rect 34 847 46 881
rect -46 841 46 847
rect 226 881 318 887
rect 226 847 238 881
rect 306 847 318 881
rect 226 841 318 847
rect 498 881 590 887
rect 498 847 510 881
rect 578 847 590 881
rect 498 841 590 847
rect 770 881 862 887
rect 770 847 782 881
rect 850 847 862 881
rect 770 841 862 847
rect 1042 881 1134 887
rect 1042 847 1054 881
rect 1122 847 1134 881
rect 1042 841 1134 847
rect 1314 881 1406 887
rect 1314 847 1326 881
rect 1394 847 1406 881
rect 1314 841 1406 847
rect 1586 881 1678 887
rect 1586 847 1598 881
rect 1666 847 1678 881
rect 1586 841 1678 847
rect -1734 788 -1688 800
rect -1734 -788 -1728 788
rect -1694 -788 -1688 788
rect -1734 -800 -1688 -788
rect -1576 788 -1530 800
rect -1576 -788 -1570 788
rect -1536 -788 -1530 788
rect -1576 -800 -1530 -788
rect -1462 788 -1416 800
rect -1462 -788 -1456 788
rect -1422 -788 -1416 788
rect -1462 -800 -1416 -788
rect -1304 788 -1258 800
rect -1304 -788 -1298 788
rect -1264 -788 -1258 788
rect -1304 -800 -1258 -788
rect -1190 788 -1144 800
rect -1190 -788 -1184 788
rect -1150 -788 -1144 788
rect -1190 -800 -1144 -788
rect -1032 788 -986 800
rect -1032 -788 -1026 788
rect -992 -788 -986 788
rect -1032 -800 -986 -788
rect -918 788 -872 800
rect -918 -788 -912 788
rect -878 -788 -872 788
rect -918 -800 -872 -788
rect -760 788 -714 800
rect -760 -788 -754 788
rect -720 -788 -714 788
rect -760 -800 -714 -788
rect -646 788 -600 800
rect -646 -788 -640 788
rect -606 -788 -600 788
rect -646 -800 -600 -788
rect -488 788 -442 800
rect -488 -788 -482 788
rect -448 -788 -442 788
rect -488 -800 -442 -788
rect -374 788 -328 800
rect -374 -788 -368 788
rect -334 -788 -328 788
rect -374 -800 -328 -788
rect -216 788 -170 800
rect -216 -788 -210 788
rect -176 -788 -170 788
rect -216 -800 -170 -788
rect -102 788 -56 800
rect -102 -788 -96 788
rect -62 -788 -56 788
rect -102 -800 -56 -788
rect 56 788 102 800
rect 56 -788 62 788
rect 96 -788 102 788
rect 56 -800 102 -788
rect 170 788 216 800
rect 170 -788 176 788
rect 210 -788 216 788
rect 170 -800 216 -788
rect 328 788 374 800
rect 328 -788 334 788
rect 368 -788 374 788
rect 328 -800 374 -788
rect 442 788 488 800
rect 442 -788 448 788
rect 482 -788 488 788
rect 442 -800 488 -788
rect 600 788 646 800
rect 600 -788 606 788
rect 640 -788 646 788
rect 600 -800 646 -788
rect 714 788 760 800
rect 714 -788 720 788
rect 754 -788 760 788
rect 714 -800 760 -788
rect 872 788 918 800
rect 872 -788 878 788
rect 912 -788 918 788
rect 872 -800 918 -788
rect 986 788 1032 800
rect 986 -788 992 788
rect 1026 -788 1032 788
rect 986 -800 1032 -788
rect 1144 788 1190 800
rect 1144 -788 1150 788
rect 1184 -788 1190 788
rect 1144 -800 1190 -788
rect 1258 788 1304 800
rect 1258 -788 1264 788
rect 1298 -788 1304 788
rect 1258 -800 1304 -788
rect 1416 788 1462 800
rect 1416 -788 1422 788
rect 1456 -788 1462 788
rect 1416 -800 1462 -788
rect 1530 788 1576 800
rect 1530 -788 1536 788
rect 1570 -788 1576 788
rect 1530 -800 1576 -788
rect 1688 788 1734 800
rect 1688 -788 1694 788
rect 1728 -788 1734 788
rect 1688 -800 1734 -788
rect -1678 -847 -1586 -841
rect -1678 -881 -1666 -847
rect -1598 -881 -1586 -847
rect -1678 -887 -1586 -881
rect -1406 -847 -1314 -841
rect -1406 -881 -1394 -847
rect -1326 -881 -1314 -847
rect -1406 -887 -1314 -881
rect -1134 -847 -1042 -841
rect -1134 -881 -1122 -847
rect -1054 -881 -1042 -847
rect -1134 -887 -1042 -881
rect -862 -847 -770 -841
rect -862 -881 -850 -847
rect -782 -881 -770 -847
rect -862 -887 -770 -881
rect -590 -847 -498 -841
rect -590 -881 -578 -847
rect -510 -881 -498 -847
rect -590 -887 -498 -881
rect -318 -847 -226 -841
rect -318 -881 -306 -847
rect -238 -881 -226 -847
rect -318 -887 -226 -881
rect -46 -847 46 -841
rect -46 -881 -34 -847
rect 34 -881 46 -847
rect -46 -887 46 -881
rect 226 -847 318 -841
rect 226 -881 238 -847
rect 306 -881 318 -847
rect 226 -887 318 -881
rect 498 -847 590 -841
rect 498 -881 510 -847
rect 578 -881 590 -847
rect 498 -887 590 -881
rect 770 -847 862 -841
rect 770 -881 782 -847
rect 850 -881 862 -847
rect 770 -887 862 -881
rect 1042 -847 1134 -841
rect 1042 -881 1054 -847
rect 1122 -881 1134 -847
rect 1042 -887 1134 -881
rect 1314 -847 1406 -841
rect 1314 -881 1326 -847
rect 1394 -881 1406 -847
rect 1314 -887 1406 -881
rect 1586 -847 1678 -841
rect 1586 -881 1598 -847
rect 1666 -881 1678 -847
rect 1586 -887 1678 -881
<< properties >>
string FIXED_BBOX -1825 -966 1825 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
