magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect 145 878 203 884
rect -29 872 29 878
rect -29 838 -17 872
rect 145 844 157 878
rect 145 838 203 844
rect -29 832 29 838
rect -173 -800 -111 800
rect -81 -800 -15 800
rect 15 -800 81 800
rect 111 -800 173 800
<< pwell >>
rect 68 816 215 901
<< nmos >>
rect -111 -800 -81 800
rect -15 -800 15 800
rect 81 -800 111 800
<< ndiff >>
rect -173 788 -111 800
rect -173 -788 -161 788
rect -127 -788 -111 788
rect -173 -800 -111 -788
rect -81 788 -15 800
rect -81 -788 -65 788
rect -31 -788 -15 788
rect -81 -800 -15 -788
rect 15 788 81 800
rect 15 -788 31 788
rect 65 -788 81 788
rect 15 -800 81 -788
rect 111 788 173 800
rect 111 -788 127 788
rect 161 -788 173 788
rect 111 -800 173 -788
<< ndiffc >>
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
<< poly >>
rect -33 878 33 888
rect 141 878 207 894
rect -111 872 33 878
rect -111 838 -17 872
rect 17 838 33 872
rect -111 828 33 838
rect -111 800 -81 828
rect -33 822 33 828
rect 81 844 157 878
rect 191 844 207 878
rect 81 828 207 844
rect -15 800 15 822
rect 81 800 111 828
rect -111 -826 -81 -800
rect -15 -826 15 -800
rect 81 -826 111 -800
<< polycont >>
rect -17 838 17 872
rect 157 844 191 878
<< locali >>
rect -33 838 -17 872
rect 17 838 33 872
rect 141 844 157 878
rect 191 844 207 878
rect -161 788 -127 804
rect -161 -804 -127 -788
rect -65 788 -31 804
rect -65 -804 -31 -788
rect 31 788 65 804
rect 31 -804 65 -788
rect 127 788 161 804
rect 127 -804 161 -788
<< viali >>
rect -17 838 17 872
rect 157 844 191 878
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
<< metal1 >>
rect 145 878 203 884
rect -29 872 29 878
rect -29 838 -17 872
rect 17 838 29 872
rect 145 844 157 878
rect 191 844 203 878
rect 145 838 203 844
rect -29 832 29 838
rect -167 788 -121 800
rect -167 -788 -161 788
rect -127 -788 -121 788
rect -167 -800 -121 -788
rect -71 788 -25 800
rect -71 -788 -65 788
rect -31 -788 -25 788
rect -71 -800 -25 -788
rect 25 788 71 800
rect 25 -788 31 788
rect 65 -788 71 788
rect 25 -800 71 -788
rect 121 788 167 800
rect 121 -788 127 788
rect 161 -788 167 788
rect 121 -800 167 -788
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
