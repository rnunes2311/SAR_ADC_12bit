magic
tech sky130A
magscale 1 2
timestamp 1711314126
<< nwell >>
rect -311 -619 311 619
<< pmos >>
rect -111 -400 -81 400
rect -15 -400 15 400
rect 81 -400 111 400
<< pdiff >>
rect -173 388 -111 400
rect -173 -388 -161 388
rect -127 -388 -111 388
rect -173 -400 -111 -388
rect -81 388 -15 400
rect -81 -388 -65 388
rect -31 -388 -15 388
rect -81 -400 -15 -388
rect 15 388 81 400
rect 15 -388 31 388
rect 65 -388 81 388
rect 15 -400 81 -388
rect 111 388 173 400
rect 111 -388 127 388
rect 161 -388 173 388
rect 111 -400 173 -388
<< pdiffc >>
rect -161 -388 -127 388
rect -65 -388 -31 388
rect 31 -388 65 388
rect 127 -388 161 388
<< nsubdiff >>
rect -275 549 -179 583
rect 179 549 275 583
rect -275 487 -241 549
rect 241 487 275 549
rect -275 -549 -241 -487
rect 241 -549 275 -487
rect -275 -583 -179 -549
rect 179 -583 275 -549
<< nsubdiffcont >>
rect -179 549 179 583
rect -275 -487 -241 487
rect 241 -487 275 487
rect -179 -583 179 -549
<< poly >>
rect -129 481 129 497
rect -129 447 -113 481
rect -79 447 -17 481
rect 17 447 79 481
rect 113 447 129 481
rect -129 431 129 447
rect -111 400 -81 431
rect -15 400 15 431
rect 81 400 111 431
rect -111 -426 -81 -400
rect -15 -426 15 -400
rect 81 -426 111 -400
<< polycont >>
rect -113 447 -79 481
rect -17 447 17 481
rect 79 447 113 481
<< locali >>
rect -275 549 -179 583
rect 179 549 275 583
rect -275 487 -241 549
rect 241 487 275 549
rect -129 447 -113 481
rect -79 447 -17 481
rect 17 447 79 481
rect 113 447 129 481
rect -161 388 -127 404
rect -161 -404 -127 -388
rect -65 388 -31 404
rect -65 -404 -31 -388
rect 31 388 65 404
rect 31 -404 65 -388
rect 127 388 161 404
rect 127 -404 161 -388
rect -275 -549 -241 -487
rect 241 -549 275 -487
rect -275 -583 -179 -549
rect 179 -583 275 -549
<< viali >>
rect -113 447 -79 481
rect -17 447 17 481
rect 79 447 113 481
rect -161 -388 -127 388
rect -65 -388 -31 388
rect 31 -388 65 388
rect 127 -388 161 388
<< metal1 >>
rect -132 481 134 490
rect -132 447 -113 481
rect -79 447 -17 481
rect 17 447 79 481
rect 113 447 134 481
rect -132 438 134 447
rect -167 388 -121 400
rect -167 -388 -161 388
rect -127 -388 -121 388
rect -167 -400 -121 -388
rect -71 388 -25 400
rect -71 -388 -65 388
rect -31 -388 -25 388
rect -71 -400 -25 -388
rect 25 388 71 400
rect 25 -388 31 388
rect 65 -388 71 388
rect 25 -400 71 -388
rect 121 388 167 400
rect 121 -388 127 388
rect 161 -388 167 388
rect 121 -400 167 -388
<< properties >>
string FIXED_BBOX -258 -566 258 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
