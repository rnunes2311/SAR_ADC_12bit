* SPICE3 file created from CDAC_mim_12bit.ext - technology: sky130A

.subckt CDAC_12bit C0_dummy C0 C1 C2 C3 C4 C5 C6 C7 C8 C9 C10 Ctop VSS
X0 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X9 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X10 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X11 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X12 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X13 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X14 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X15 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X16 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X17 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X18 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X19 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X20 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X21 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X22 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X23 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X24 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X25 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X26 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X27 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X28 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X29 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X30 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X31 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X32 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X33 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X34 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X35 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X36 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X37 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X38 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X39 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X40 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X41 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X42 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X43 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X44 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X45 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X46 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X47 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X48 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X49 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X50 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X51 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X52 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X53 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X54 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X55 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X56 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X57 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X58 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X59 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X60 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X61 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X62 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X63 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X64 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X65 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X66 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X67 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X68 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X69 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X70 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X71 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X72 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X73 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X74 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X75 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X76 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X77 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X78 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X79 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X80 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X81 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X82 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X83 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X84 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X85 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X86 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X87 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X88 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X89 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X90 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X91 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X92 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X93 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X94 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X95 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X96 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X97 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X98 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X99 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X100 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X101 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X102 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X103 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X104 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X105 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X106 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X107 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X108 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X109 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X110 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X111 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X112 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X113 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X114 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X115 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X116 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X117 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X118 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X119 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X120 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X121 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X122 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X123 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X124 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X125 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X126 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X127 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X128 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X129 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X130 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X131 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X132 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X133 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X134 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X135 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X136 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X137 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X138 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X139 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X140 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X141 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X142 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X143 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X144 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X145 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X146 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X147 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X148 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X149 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X150 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X151 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X152 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X153 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X154 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X155 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X156 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X157 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X158 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X159 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X160 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X161 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X162 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X163 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X164 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X165 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X166 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X167 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X168 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X169 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X170 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X171 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X172 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X173 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X174 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X175 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X176 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X177 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X178 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X179 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X180 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X181 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X182 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X183 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X184 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X185 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X186 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X187 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X188 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X189 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X190 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X191 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X192 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X193 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X194 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X195 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X196 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X197 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X198 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X199 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X200 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X201 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X202 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X203 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X204 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X205 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X206 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X207 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X208 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X209 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X210 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X211 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X212 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X213 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X214 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X215 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X216 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X217 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X218 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X219 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X220 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X221 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X222 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X223 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X224 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X225 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X226 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X227 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X228 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X229 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X230 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X231 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X232 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X233 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X234 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X235 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X236 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X237 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X238 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X239 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X240 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X241 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X242 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X243 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X244 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X245 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X246 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X247 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X248 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X249 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X250 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X251 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X252 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X253 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X254 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X255 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X256 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X257 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X258 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X259 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X260 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X261 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X262 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X263 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X264 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X265 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X266 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X267 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X268 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X269 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X270 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X271 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X272 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X273 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X274 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X275 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X276 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X277 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X278 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X279 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X280 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X281 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X282 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X283 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X284 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X285 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X286 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X287 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X288 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X289 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X290 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X291 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X292 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X293 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X294 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X295 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X296 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X297 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X298 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X299 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X300 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X301 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X302 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X303 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X304 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X305 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X306 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X307 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X308 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X309 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X310 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X311 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X312 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X313 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X314 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X315 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X316 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X317 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X318 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X319 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X320 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X321 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X322 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X323 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X324 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X325 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X326 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X327 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X328 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X329 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X330 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X331 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X332 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X333 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X334 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X335 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X336 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X337 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X338 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X339 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X340 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X341 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X342 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X343 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X344 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X345 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X346 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X347 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X348 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X349 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X350 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X351 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X352 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X353 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X354 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X355 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X356 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X357 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X358 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X359 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X360 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X361 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X362 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X363 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X364 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X365 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X366 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X367 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X368 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X369 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X370 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X371 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X372 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X373 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X374 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X375 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X376 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X377 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X378 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X379 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X380 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X381 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X382 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X383 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X384 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X385 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X386 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X387 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X388 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X389 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X390 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X391 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X392 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X393 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X394 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X395 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X396 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X397 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X398 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X399 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X400 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X401 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X402 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X403 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X404 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X405 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X406 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X407 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X408 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X409 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X410 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X411 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X412 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X413 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X414 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X415 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X416 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X417 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X418 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X419 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X420 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X421 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X422 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X423 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X424 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X425 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X426 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X427 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X428 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X429 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X430 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X431 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X432 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X433 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X434 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X435 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X436 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X437 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X438 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X439 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X440 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X441 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X442 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X443 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X444 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X445 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X446 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X447 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X448 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X449 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X450 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X451 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X452 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X453 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X454 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X455 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X456 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X457 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X458 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X459 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X460 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X461 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X462 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X463 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X464 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X465 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X466 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X467 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X468 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X469 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X470 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X471 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X472 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X473 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X474 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X475 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X476 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X477 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X478 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X479 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X480 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X481 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X482 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X483 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X484 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X485 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X486 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X487 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X488 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X489 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X490 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X491 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X492 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X493 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X494 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X495 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X496 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X497 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X498 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X499 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X500 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X501 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X502 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X503 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X504 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X505 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X506 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X507 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X508 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X509 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X510 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X511 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X512 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X513 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X514 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X515 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X516 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X517 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X518 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X519 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X520 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X521 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X522 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X523 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X524 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X525 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X526 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X527 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X528 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X529 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X530 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X531 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X532 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X533 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X534 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X535 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X536 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X537 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X538 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X539 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X540 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X541 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X542 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X543 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X544 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X545 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X546 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X547 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X548 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X549 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X550 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X551 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X552 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X553 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X554 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X555 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X556 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X557 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X558 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X559 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X560 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X561 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X562 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X563 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X564 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X565 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X566 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X567 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X568 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X569 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X570 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X571 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X572 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X573 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X574 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X575 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X576 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X577 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X578 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X579 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X580 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X581 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X582 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X583 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X584 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X585 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X586 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X587 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X588 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X589 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X590 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X591 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X592 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X593 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X594 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X595 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X596 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X597 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X598 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X599 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X600 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X601 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X602 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X603 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X604 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X605 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X606 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X607 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X608 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X609 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X610 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X611 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X612 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X613 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X614 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X615 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X616 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X617 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X618 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X619 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X620 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X621 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X622 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X623 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X624 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X625 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X626 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X627 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X628 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X629 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X630 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X631 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X632 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X633 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X634 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X635 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X636 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X637 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X638 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X639 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X640 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X641 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X642 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X643 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X644 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X645 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X646 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X647 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X648 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X649 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X650 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X651 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X652 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X653 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X654 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X655 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X656 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X657 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X658 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X659 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X660 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X661 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X662 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X663 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X664 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X665 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X666 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X667 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X668 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X669 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X670 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X671 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X672 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X673 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X674 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X675 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X676 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X677 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X678 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X679 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X680 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X681 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X682 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X683 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X684 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X685 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X686 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X687 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X688 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X689 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X690 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X691 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X692 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X693 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X694 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X695 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X696 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X697 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X698 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X699 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X700 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X701 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X702 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X703 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X704 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X705 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X706 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X707 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X708 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X709 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X710 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X711 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X712 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X713 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X714 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X715 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X716 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X717 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X718 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X719 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X720 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X721 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X722 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X723 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X724 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X725 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X726 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X727 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X728 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X729 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X730 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X731 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X732 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X733 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X734 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X735 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X736 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X737 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X738 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X739 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X740 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X741 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X742 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X743 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X744 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X745 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X746 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X747 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X748 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X749 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X750 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X751 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X752 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X753 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X754 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X755 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X756 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X757 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X758 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X759 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X760 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X761 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X762 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X763 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X764 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X765 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X766 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X767 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X768 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X769 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X770 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X771 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X772 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X773 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X774 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X775 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X776 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X777 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X778 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X779 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X780 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X781 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X782 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X783 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X784 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X785 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X786 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X787 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X788 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X789 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X790 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X791 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X792 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X793 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X794 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X795 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X796 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X797 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X798 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X799 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X800 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X801 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X802 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X803 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X804 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X805 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X806 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X807 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X808 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X809 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X810 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X811 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X812 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X813 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X814 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X815 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X816 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X817 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X818 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X819 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X820 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X821 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X822 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X823 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X824 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X825 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X826 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X827 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X828 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X829 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X830 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X831 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X832 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X833 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X834 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X835 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X836 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X837 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X838 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X839 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X840 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X841 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X842 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X843 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X844 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X845 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X846 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X847 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X848 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X849 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X850 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X851 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X852 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X853 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X854 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X855 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X856 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X857 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X858 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X859 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X860 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X861 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X862 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X863 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X864 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X865 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X866 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X867 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X868 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X869 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X870 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X871 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X872 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X873 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X874 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X875 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X876 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X877 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X878 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X879 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X880 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X881 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X882 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X883 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X884 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X885 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X886 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X887 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X888 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X889 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X890 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X891 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X892 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X893 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X894 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X895 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X896 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X897 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X898 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X899 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X900 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X901 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X902 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X903 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X904 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X905 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X906 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X907 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X908 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X909 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X910 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X911 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X912 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X913 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X914 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X915 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X916 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X917 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X918 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X919 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X920 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X921 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X922 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X923 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X924 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X925 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X926 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X927 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X928 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X929 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X930 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X931 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X932 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X933 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X934 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X935 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X936 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X937 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X938 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X939 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X940 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X941 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X942 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X943 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X944 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X945 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X946 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X947 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X948 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X949 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X950 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X951 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X952 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X953 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X954 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X955 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X956 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X957 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X958 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X959 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X960 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X961 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X962 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X963 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X964 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X965 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X966 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X967 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X968 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X969 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X970 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X971 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X972 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X973 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X974 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X975 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X976 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X977 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X978 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X979 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X980 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X981 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X982 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X983 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X984 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X985 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X986 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X987 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X988 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X989 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X990 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X991 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X992 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X993 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X994 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X995 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X996 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X997 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X998 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X999 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1000 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1001 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1002 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1003 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1004 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1005 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1006 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1007 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1008 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1009 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1010 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1011 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1012 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1013 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1014 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1015 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1016 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1017 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1018 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1019 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1020 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1021 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1022 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1023 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1024 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1025 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1026 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1027 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1028 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1029 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1030 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1031 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1032 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1033 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1034 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1035 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1036 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1037 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1038 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1039 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1040 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1041 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1042 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1043 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1044 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1045 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1046 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1047 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1048 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1049 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1050 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1051 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1052 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1053 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1054 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1055 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1056 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1057 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1058 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1059 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1060 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1061 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1062 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1063 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1064 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1065 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1066 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1067 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1068 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1069 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1070 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1071 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1072 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1073 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1074 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1075 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1076 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1077 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1078 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1079 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1080 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1081 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1082 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1083 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1084 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1085 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1086 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1087 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1088 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1089 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1090 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1091 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1092 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1093 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1094 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1095 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1096 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1097 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1098 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1099 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1100 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1101 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1102 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1103 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1104 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1105 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1106 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1107 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1108 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1109 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1110 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1111 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1112 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1113 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1114 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1115 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1116 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1117 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1118 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1119 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1120 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1121 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1122 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1123 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1124 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1125 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1126 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1127 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1128 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1129 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1130 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1131 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1132 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1133 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1134 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1135 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1136 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1137 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1138 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1139 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1140 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1141 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1142 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1143 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1144 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1145 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1146 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1147 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1148 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1149 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1150 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1151 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1152 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1153 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1154 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1155 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1156 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1157 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1158 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1159 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1160 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1161 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1162 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1163 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1164 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1165 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1166 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1167 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1168 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1169 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1170 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1171 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1172 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1173 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1174 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1175 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1176 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1177 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1178 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1179 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1180 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1181 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1182 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1183 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1184 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1185 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1186 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1187 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1188 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1189 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1190 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1191 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1192 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1193 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1194 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1195 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1196 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1197 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1198 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1199 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1200 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1201 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1202 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1203 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1204 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1205 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1206 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1207 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1208 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1209 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1210 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1211 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1212 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1213 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1214 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1215 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1216 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1217 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1218 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1219 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1220 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1221 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1222 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1223 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1224 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1225 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1226 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1227 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1228 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1229 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1230 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1231 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1232 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1233 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1234 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1235 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1236 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1237 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1238 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1239 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1240 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1241 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1242 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1243 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1244 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1245 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1246 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1247 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1248 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1249 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1250 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1251 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1252 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1253 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1254 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1255 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1256 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1257 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1258 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1259 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1260 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1261 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1262 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1263 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1264 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1265 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1266 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1267 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1268 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1269 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1270 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1271 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1272 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1273 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1274 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1275 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1276 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1277 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1278 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1279 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1280 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1281 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1282 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1283 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1284 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1285 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1286 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1287 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1288 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1289 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1290 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1291 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1292 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1293 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1294 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1295 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1296 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1297 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1298 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1299 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1300 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1301 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1302 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1303 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1304 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1305 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1306 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1307 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1308 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1309 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1310 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1311 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1312 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1313 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1314 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1315 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1316 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1317 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1318 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1319 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1320 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1321 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1322 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1323 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1324 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1325 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1326 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1327 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1328 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1329 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1330 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1331 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1332 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1333 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1334 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1335 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1336 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1337 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1338 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1339 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1340 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1341 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1342 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1343 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1344 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1345 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1346 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1347 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1348 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1349 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1350 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1351 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1352 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1353 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1354 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1355 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1356 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1357 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1358 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1359 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1360 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1361 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1362 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1363 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1364 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1365 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1366 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1367 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1368 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1369 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1370 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1371 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1372 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1373 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1374 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1375 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1376 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1377 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1378 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1379 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1380 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1381 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1382 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1383 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1384 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1385 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1386 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1387 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1388 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1389 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1390 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1391 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1392 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1393 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1394 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1395 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1396 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1397 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1398 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1399 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1400 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1401 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1402 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1403 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1404 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1405 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1406 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1407 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1408 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1409 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1410 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1411 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1412 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1413 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1414 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1415 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1416 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1417 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1418 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1419 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1420 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1421 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1422 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1423 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1424 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1425 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1426 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1427 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1428 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1429 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1430 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1431 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1432 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1433 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1434 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1435 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1436 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1437 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1438 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1439 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1440 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1441 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1442 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1443 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1444 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1445 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1446 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1447 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1448 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1449 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1450 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1451 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1452 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1453 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1454 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1455 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1456 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1457 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1458 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1459 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1460 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1461 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1462 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1463 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1464 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1465 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1466 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1467 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1468 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1469 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1470 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1471 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1472 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1473 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1474 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1475 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1476 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1477 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1478 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1479 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1480 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1481 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1482 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1483 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1484 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1485 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1486 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1487 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1488 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1489 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1490 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1491 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1492 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1493 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1494 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1495 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1496 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1497 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1498 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1499 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1500 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1501 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1502 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1503 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1504 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1505 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1506 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1507 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1508 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1509 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1510 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1511 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1512 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1513 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1514 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1515 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1516 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1517 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1518 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1519 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1520 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1521 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1522 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1523 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1524 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1525 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1526 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1527 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1528 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1529 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1530 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1531 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1532 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1533 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1534 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1535 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1536 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1537 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1538 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1539 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1540 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1541 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1542 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1543 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1544 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1545 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1546 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1547 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1548 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1549 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1550 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1551 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1552 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1553 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1554 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1555 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1556 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1557 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1558 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1559 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1560 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1561 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1562 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1563 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1564 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1565 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1566 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1567 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1568 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1569 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1570 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1571 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1572 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1573 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1574 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1575 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1576 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1577 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1578 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1579 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1580 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1581 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1582 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1583 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1584 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1585 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1586 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1587 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1588 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1589 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1590 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1591 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1592 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1593 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1594 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1595 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1596 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1597 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1598 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1599 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1600 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1601 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1602 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1603 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1604 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1605 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1606 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1607 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1608 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1609 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1610 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1611 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1612 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1613 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1614 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1615 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1616 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1617 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1618 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1619 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1620 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1621 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1622 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1623 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1624 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1625 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1626 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1627 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1628 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1629 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1630 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1631 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1632 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1633 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1634 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1635 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1636 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1637 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1638 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1639 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1640 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1641 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1642 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1643 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1644 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1645 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1646 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1647 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1648 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1649 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1650 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1651 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1652 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1653 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1654 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1655 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1656 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1657 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1658 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1659 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1660 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1661 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1662 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1663 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1664 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1665 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1666 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1667 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1668 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1669 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1670 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1671 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1672 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1673 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1674 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1675 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1676 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1677 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1678 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1679 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1680 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1681 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1682 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1683 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1684 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1685 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1686 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1687 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1688 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1689 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1690 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1691 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1692 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1693 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1694 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1695 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1696 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1697 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1698 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1699 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1700 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1701 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1702 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1703 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1704 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1705 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1706 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1707 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1708 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1709 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1710 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1711 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1712 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1713 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1714 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1715 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1716 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1717 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1718 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1719 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1720 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1721 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1722 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1723 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1724 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1725 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1726 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1727 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1728 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1729 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1730 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1731 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1732 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1733 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1734 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1735 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1736 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1737 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1738 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1739 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1740 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1741 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1742 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1743 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1744 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1745 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1746 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1747 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1748 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1749 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1750 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1751 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1752 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1753 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1754 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1755 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1756 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1757 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1758 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1759 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1760 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1761 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1762 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1763 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1764 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1765 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1766 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1767 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1768 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1769 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1770 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1771 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1772 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1773 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1774 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1775 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1776 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1777 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1778 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1779 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1780 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1781 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1782 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1783 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1784 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1785 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1786 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1787 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1788 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1789 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1790 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1791 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1792 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1793 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1794 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1795 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1796 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1797 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1798 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1799 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1800 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1801 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1802 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1803 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1804 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1805 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1806 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1807 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1808 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1809 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1810 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1811 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1812 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1813 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1814 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1815 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1816 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1817 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1818 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1819 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1820 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1821 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1822 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1823 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1824 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1825 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1826 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1827 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1828 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1829 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1830 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1831 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1832 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1833 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1834 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1835 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1836 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1837 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1838 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1839 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1840 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1841 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1842 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1843 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1844 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1845 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1846 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1847 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1848 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1849 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1850 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1851 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1852 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1853 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1854 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1855 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1856 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1857 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1858 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1859 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1860 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1861 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1862 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1863 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1864 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1865 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1866 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1867 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1868 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1869 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1870 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1871 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1872 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1873 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1874 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1875 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1876 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1877 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1878 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1879 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1880 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1881 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1882 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1883 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1884 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1885 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1886 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1887 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1888 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1889 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1890 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1891 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1892 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1893 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1894 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1895 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1896 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1897 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1898 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1899 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1900 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1901 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1902 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1903 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1904 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1905 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1906 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1907 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1908 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1909 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1910 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1911 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1912 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1913 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1914 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1915 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1916 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1917 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1918 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1919 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1920 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1921 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1922 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1923 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1924 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1925 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1926 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1927 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1928 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1929 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1930 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1931 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1932 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1933 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1934 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1935 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1936 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1937 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1938 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1939 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1940 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1941 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1942 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1943 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1944 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1945 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1946 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1947 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1948 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1949 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1950 Ctop C2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1951 Ctop C2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1952 Ctop C2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1953 Ctop C1 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1954 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1955 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1956 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1957 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1958 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1959 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1960 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1961 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1962 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1963 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1964 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1965 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1966 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1967 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1968 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1969 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1970 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1971 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1972 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1973 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1974 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1975 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1976 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1977 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1978 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1979 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1980 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1981 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1982 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1983 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1984 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1985 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1986 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1987 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1988 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1989 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1990 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1991 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1992 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1993 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1994 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1995 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1996 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1997 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1998 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1999 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2000 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2001 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2002 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2003 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2004 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2005 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2006 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2007 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2008 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2009 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2010 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2011 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2012 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2013 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2014 Ctop C2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2015 Ctop C0_dummy sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2016 Ctop C0 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2017 Ctop C1 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2018 Ctop C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2019 Ctop C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2020 Ctop C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2021 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2022 Ctop C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2023 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2024 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2025 Ctop C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2026 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2027 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2028 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2029 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2030 Ctop C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2031 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2032 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2033 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2034 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2035 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2036 Ctop C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2037 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2038 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2039 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2040 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2041 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2042 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2043 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2044 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2045 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2046 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2047 Ctop C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2048 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2049 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2050 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2051 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2052 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2053 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2054 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2055 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2056 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2057 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2058 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2059 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2060 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2061 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2062 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2063 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2064 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2065 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2066 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2067 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2068 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2069 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2070 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2071 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2072 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2073 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2074 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2075 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2076 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2077 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2078 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2079 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2080 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2081 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2082 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2083 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2084 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2085 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2086 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2087 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2088 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2089 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2090 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2091 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2092 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2093 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2094 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2095 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2096 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2097 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2098 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2099 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2100 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2101 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2102 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2103 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2104 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2105 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2106 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2107 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2108 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2109 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2110 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2111 Ctop VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2112 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2113 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2114 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2115 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2116 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2117 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2118 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2119 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2120 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2121 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2122 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2123 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2124 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2125 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2126 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2127 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2128 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2129 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2130 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2131 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2132 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2133 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2134 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2135 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2136 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2137 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2138 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2139 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2140 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2141 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2142 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2143 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2144 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2145 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2146 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2147 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2148 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2149 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2150 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2151 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2152 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2153 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2154 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2155 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2156 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2157 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2158 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2159 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2160 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2161 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2162 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2163 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2164 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2165 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2166 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2167 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2168 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2169 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2170 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2171 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2172 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2173 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2174 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2175 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2176 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2177 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2178 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2179 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2180 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2181 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2182 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2183 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2184 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2185 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2186 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2187 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2188 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2189 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2190 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2191 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2192 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2193 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2194 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2195 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2196 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2197 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2198 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2199 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2200 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2201 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2202 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2203 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2204 VSS C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2205 VSS C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2206 VSS C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2207 VSS C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2208 VSS C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2209 VSS C2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2210 VSS C0_dummy sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2211 VSS C0 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2212 VSS C1 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2213 VSS C3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2214 VSS C4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2215 VSS C5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2216 VSS C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2217 VSS C6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2218 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2219 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2220 VSS C7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2221 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2222 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2223 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2224 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2225 VSS C8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2226 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2227 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2228 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2229 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2230 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2231 VSS C9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2232 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2233 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2234 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2235 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2236 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2237 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2238 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2239 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2240 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2241 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2242 VSS C10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2243 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
C0 C0 C1 0.455366f
C1 C6 C2 0.170878f
C2 C0_dummy Ctop 0.233088f
C3 C0_dummy C1 0.146899f
C4 C0 C2 0.148128f
C5 Ctop C9 0.110161p
C6 C4 Ctop 3.483357f
C7 C0_dummy C2 0.457823f
C8 C4 C1 0.360409f
C9 Ctop C10 0.220974p
C10 C4 C2 1.211851f
C11 C7 C5 1.52167f
C12 C8 C7 18.72166f
C13 Ctop C3 1.731604f
C14 C3 C1 0.680234f
C15 C3 C2 0.244636f
C16 C6 C5 6.655549f
C17 C0 C5 0.093587f
C18 Ctop C1 0.446552f
C19 C6 C8 1.240844f
C20 C0_dummy C5 0.093587f
C21 Ctop C2 0.875194f
C22 C2 C1 0.422971f
C23 C4 C5 2.87264f
C24 C9 C8 26.831766f
C25 C6 C7 11.960523f
C26 C5 C3 0.548642f
C27 C4 C7 0.54418f
C28 C0 C6 0.030497f
C29 Ctop C5 6.894931f
C30 C0_dummy C6 0.030497f
C31 C5 C1 0.132512f
C32 C0_dummy C0 0.454741f
C33 C4 C6 1.677797f
C34 Ctop C8 55.147877f
C35 C5 C2 0.2261f
C36 C7 C3 0.076242f
C37 C0 C4 0.239773f
C38 C0_dummy C4 0.298117f
C39 Ctop C7 27.562223f
C40 C10 C9 37.167885f
C41 C6 C3 0.502664f
C42 C0 C3 0.14726f
C43 C0_dummy C3 0.088341f
C44 C6 Ctop 13.80047f
C45 C4 C3 1.551874f
C46 C6 C1 0.140381f
C47 C0 Ctop 0.233088f
C48 C6 VSS 51.84848f
C49 C4 VSS 14.24818f
C50 C0 VSS 1.482448f
C51 C0_dummy VSS 1.482448f
C52 C1 VSS 2.2231f
C53 C2 VSS 3.778132f
C54 C3 VSS 6.839335f
C55 C5 VSS 25.819008f
C56 C7 VSS 0.102345p
C57 C8 VSS 0.204738p
C58 C9 VSS 0.404615p
C59 C10 VSS 0.824602p
C60 Ctop VSS 0.317192p
.ends
