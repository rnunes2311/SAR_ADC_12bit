magic
tech sky130A
magscale 1 2
timestamp 1711831820
<< nwell >>
rect 15679 1323 15712 2253
rect 15638 1203 16023 1323
rect 15679 1140 15909 1203
rect 15679 714 15930 1140
rect 19900 964 20165 1107
rect 15690 610 15930 714
rect 19860 870 20165 964
rect 19860 696 20164 870
rect 15900 560 15930 610
<< pwell >>
rect 19345 1204 19839 1304
rect 19345 1022 19832 1204
rect 19334 135 19682 340
rect 19334 84 20115 135
rect 19367 83 20115 84
<< psubdiff >>
rect 19381 1234 19405 1268
rect 19811 1234 19835 1268
rect 19390 96 19419 130
rect 20005 96 20034 130
<< nsubdiff >>
rect 19940 910 20030 940
rect 19940 690 20030 781
<< psubdiffcont >>
rect 19405 1234 19811 1268
rect 19419 96 20005 130
<< nsubdiffcont >>
rect 19940 781 20030 910
<< poly >>
rect 16106 1129 16442 1200
<< locali >>
rect 19389 1234 19405 1268
rect 19811 1234 19827 1268
rect 19426 964 19460 1002
rect 19735 967 19773 1001
rect 19920 910 20049 931
rect 19920 781 19940 910
rect 20030 781 20049 910
rect 19920 698 20049 781
rect 19459 685 20049 698
rect 19459 664 20015 685
rect 19402 358 19440 392
rect 19554 352 19728 402
rect 20056 352 20090 390
rect 16700 120 16770 160
rect 17860 120 18070 160
rect 19270 154 19310 160
rect 19270 153 19405 154
rect 19270 130 19433 153
rect 19270 127 19419 130
rect 19270 122 19394 127
rect 19270 120 19419 122
rect 19367 119 19419 120
rect 19373 96 19419 119
rect 20005 96 20073 122
<< viali >>
rect 12499 2183 15466 2217
rect 16100 1272 16500 1306
rect 19426 1002 19460 1038
rect 9281 301 9315 980
rect 15626 315 15660 994
rect 16553 307 16587 986
rect 19699 967 19735 1001
rect 19773 967 19809 1001
rect 19426 928 19460 964
rect 19366 358 19402 392
rect 19440 358 19476 392
rect 20056 390 20090 426
rect 20056 316 20090 352
rect 12508 120 15475 154
rect 16110 120 16510 154
rect 16770 120 17860 160
rect 18070 120 19270 160
<< metal1 >>
rect 9245 2217 15690 2254
rect 9245 2183 12499 2217
rect 15466 2183 15690 2217
rect 9245 2157 15690 2183
rect 9245 1868 9342 2157
rect 9980 2050 9990 2120
rect 10050 2050 10080 2120
rect 10140 2050 10150 2120
rect 11770 2050 11780 2120
rect 11840 2050 11870 2120
rect 11930 2050 11940 2120
rect 12950 2050 12960 2120
rect 13020 2050 13050 2120
rect 13110 2050 13120 2120
rect 15220 2060 15230 2120
rect 15290 2060 15330 2120
rect 15390 2060 15400 2120
rect 15591 1868 15690 2157
rect 9245 1439 15690 1868
rect 9245 980 9342 1439
rect 15591 1322 15690 1439
rect 15591 1306 16624 1322
rect 15591 1272 16100 1306
rect 16500 1272 16624 1306
rect 15591 1266 16624 1272
rect 9464 1140 12425 1226
rect 12533 1140 15494 1229
rect 15591 1225 16157 1266
rect 16470 1225 16624 1266
rect 15591 1140 16003 1225
rect 16230 1193 16291 1203
rect 16189 1144 16230 1190
rect 9445 1130 15496 1140
rect 9445 1094 9995 1130
rect 10056 1094 10089 1130
rect 9995 1068 10056 1078
rect 10150 1094 11775 1130
rect 10089 1068 10150 1078
rect 11836 1094 11869 1130
rect 11775 1068 11836 1078
rect 11930 1094 12955 1130
rect 11869 1068 11930 1078
rect 13016 1094 13049 1130
rect 12955 1068 13016 1078
rect 13110 1094 15225 1130
rect 13049 1068 13110 1078
rect 15286 1094 15319 1130
rect 15225 1068 15286 1078
rect 15380 1094 15496 1130
rect 15319 1068 15380 1078
rect 9245 301 9281 980
rect 9315 864 9342 980
rect 15591 994 15690 1140
rect 15829 1038 15839 1099
rect 15891 1038 15901 1099
rect 15840 1005 15890 1038
rect 15591 864 15626 994
rect 9315 435 15626 864
rect 9315 301 9342 435
rect 9245 185 9342 301
rect 15591 315 15626 435
rect 15660 652 15690 994
rect 15829 944 15839 1005
rect 15891 944 15901 1005
rect 15660 474 15688 652
rect 15660 326 15748 474
rect 15840 350 15890 944
rect 15930 560 16003 1140
rect 16324 1193 16385 1203
rect 16291 1144 16324 1190
rect 16230 1131 16291 1141
rect 16385 1144 16428 1190
rect 16324 1131 16385 1141
rect 16527 986 16624 1225
rect 16141 696 16151 757
rect 16203 696 16213 757
rect 16333 696 16343 757
rect 16395 696 16405 757
rect 16141 602 16151 663
rect 16203 602 16213 663
rect 16333 602 16343 663
rect 16395 602 16405 663
rect 15932 552 16003 560
rect 15932 551 16104 552
rect 15932 490 16047 551
rect 16099 490 16109 551
rect 16229 490 16239 551
rect 16291 490 16301 551
rect 16421 490 16431 551
rect 16483 490 16493 551
rect 15932 457 16104 490
rect 15932 396 16047 457
rect 16099 396 16109 457
rect 16229 396 16239 457
rect 16291 396 16301 457
rect 16421 396 16431 457
rect 16483 396 16493 457
rect 15660 315 15688 326
rect 9993 278 10054 288
rect 9445 226 9993 262
rect 10087 278 10148 288
rect 10054 226 10087 262
rect 11765 278 11826 288
rect 10148 226 11765 262
rect 11859 278 11920 288
rect 11826 226 11859 262
rect 12945 278 13006 288
rect 11920 226 12945 262
rect 13039 278 13100 288
rect 13006 226 13039 262
rect 15221 276 15282 286
rect 13100 226 15221 262
rect 9445 224 15221 226
rect 15315 276 15376 286
rect 15282 224 15315 262
rect 15376 224 15496 262
rect 9445 216 15496 224
rect 15221 214 15282 216
rect 15315 214 15376 216
rect 15591 185 15688 315
rect 15723 265 15784 275
rect 15723 203 15784 213
rect 15817 265 15878 275
rect 15817 203 15878 213
rect 9245 167 15688 185
rect 15932 185 16003 396
rect 16527 307 16553 986
rect 16587 307 16624 986
rect 16527 185 16624 307
rect 15932 167 16624 185
rect 9245 154 16624 167
rect 9245 120 12508 154
rect 15475 120 16110 154
rect 16510 120 16624 154
rect 9245 88 16624 120
rect 16660 1306 19850 1388
rect 16660 185 16738 1306
rect 16856 1243 17266 1264
rect 16856 1191 16986 1243
rect 17047 1191 17080 1243
rect 17141 1191 17266 1243
rect 16856 1168 17266 1191
rect 17025 992 17035 1053
rect 17087 992 17097 1053
rect 17025 898 17035 959
rect 17087 898 17097 959
rect 16787 664 16797 725
rect 16849 664 16859 725
rect 17263 664 17273 725
rect 17325 664 17335 725
rect 16787 570 16797 631
rect 16849 570 16859 631
rect 17263 570 17273 631
rect 17325 570 17335 631
rect 17392 185 17480 1306
rect 17521 1243 17840 1264
rect 17521 1191 17651 1243
rect 17712 1191 17745 1243
rect 17806 1191 17840 1243
rect 17521 1162 17840 1191
rect 17906 1234 19850 1306
rect 17906 1050 18064 1234
rect 18178 1184 18333 1194
rect 18239 1132 18272 1184
rect 18178 1122 18333 1132
rect 17531 666 17541 727
rect 17593 666 17603 727
rect 17531 572 17541 633
rect 17593 572 17603 633
rect 17769 468 17779 529
rect 17831 468 17841 529
rect 17769 374 17779 435
rect 17831 374 17841 435
rect 17906 366 18144 1050
rect 18209 992 18219 1053
rect 18271 992 18281 1053
rect 18424 1050 18488 1234
rect 18209 898 18219 959
rect 18271 898 18281 959
rect 17906 185 18064 366
rect 18342 364 18488 1050
rect 18847 1004 18909 1234
rect 19015 1184 19170 1194
rect 19076 1132 19109 1184
rect 19015 1122 19170 1132
rect 19236 1004 19325 1234
rect 19402 1024 19412 1085
rect 19464 1024 19474 1085
rect 18639 828 18649 889
rect 18701 828 18711 889
rect 18639 734 18649 795
rect 18701 734 18711 795
rect 18535 575 18545 636
rect 18597 575 18607 636
rect 18733 575 18743 636
rect 18795 575 18805 636
rect 18535 481 18545 542
rect 18597 481 18607 542
rect 18733 481 18743 542
rect 18795 481 18805 542
rect 18424 185 18488 364
rect 18847 357 18991 1004
rect 19049 818 19059 879
rect 19111 818 19121 879
rect 19049 724 19059 785
rect 19111 724 19121 785
rect 18593 256 18654 266
rect 18593 194 18654 204
rect 18687 256 18748 266
rect 18687 194 18748 204
rect 16660 166 18488 185
rect 18847 185 18909 357
rect 19187 351 19325 1004
rect 19420 1002 19426 1024
rect 19460 1002 19466 1024
rect 19696 1012 19757 1022
rect 19420 991 19466 1002
rect 19402 930 19412 991
rect 19464 930 19474 991
rect 19687 961 19696 1007
rect 19790 1012 19851 1022
rect 19757 1001 19790 1007
rect 19757 967 19773 1001
rect 19757 961 19790 967
rect 19696 950 19757 960
rect 19790 950 19851 960
rect 19420 928 19426 930
rect 19460 928 19466 930
rect 19420 916 19466 928
rect 19439 644 19449 718
rect 20024 644 20034 718
rect 20051 438 20061 459
rect 20050 426 20061 438
rect 19363 404 19424 414
rect 19354 352 19363 398
rect 19457 404 19518 414
rect 19424 392 19457 398
rect 19424 358 19440 392
rect 19424 352 19457 358
rect 19236 185 19325 351
rect 19363 342 19424 352
rect 19457 342 19518 352
rect 20050 390 20056 426
rect 20113 398 20123 459
rect 20090 390 20096 398
rect 20050 365 20096 390
rect 20050 352 20061 365
rect 20050 316 20056 352
rect 20050 304 20061 316
rect 20113 304 20123 365
rect 18847 166 19417 185
rect 16660 160 19417 166
rect 16660 159 16770 160
rect 17860 159 18070 160
rect 19270 159 19417 160
rect 16660 99 16703 159
rect 19290 120 19417 159
rect 19434 120 19444 158
rect 19290 99 19444 120
rect 16660 96 19444 99
rect 20040 96 20050 158
rect 16660 89 19464 96
<< via1 >>
rect 9990 2050 10050 2120
rect 10080 2050 10140 2120
rect 11780 2050 11840 2120
rect 11870 2050 11930 2120
rect 12960 2050 13020 2120
rect 13050 2050 13110 2120
rect 15230 2060 15290 2120
rect 15330 2060 15390 2120
rect 9995 1078 10056 1130
rect 10089 1078 10150 1130
rect 11775 1078 11836 1130
rect 11869 1078 11930 1130
rect 12955 1078 13016 1130
rect 13049 1078 13110 1130
rect 15225 1078 15286 1130
rect 15319 1078 15380 1130
rect 15839 1038 15891 1099
rect 15839 944 15891 1005
rect 16230 1141 16291 1193
rect 16324 1141 16385 1193
rect 16151 696 16203 757
rect 16343 696 16395 757
rect 16151 602 16203 663
rect 16343 602 16395 663
rect 16047 490 16099 551
rect 16239 490 16291 551
rect 16431 490 16483 551
rect 16047 396 16099 457
rect 16239 396 16291 457
rect 16431 396 16483 457
rect 9993 226 10054 278
rect 10087 226 10148 278
rect 11765 226 11826 278
rect 11859 226 11920 278
rect 12945 226 13006 278
rect 13039 226 13100 278
rect 15221 224 15282 276
rect 15315 224 15376 276
rect 15723 213 15784 265
rect 15817 213 15878 265
rect 16986 1191 17047 1243
rect 17080 1191 17141 1243
rect 17035 992 17087 1053
rect 17035 898 17087 959
rect 16797 664 16849 725
rect 17273 664 17325 725
rect 16797 570 16849 631
rect 17273 570 17325 631
rect 17651 1191 17712 1243
rect 17745 1191 17806 1243
rect 18178 1132 18239 1184
rect 18272 1132 18333 1184
rect 17541 666 17593 727
rect 17541 572 17593 633
rect 17779 468 17831 529
rect 17779 374 17831 435
rect 18219 992 18271 1053
rect 18219 898 18271 959
rect 19015 1132 19076 1184
rect 19109 1132 19170 1184
rect 19412 1038 19464 1085
rect 19412 1024 19426 1038
rect 19426 1024 19460 1038
rect 19460 1024 19464 1038
rect 18649 828 18701 889
rect 18649 734 18701 795
rect 18545 575 18597 636
rect 18743 575 18795 636
rect 18545 481 18597 542
rect 18743 481 18795 542
rect 19059 818 19111 879
rect 19059 724 19111 785
rect 18593 204 18654 256
rect 18687 204 18748 256
rect 19412 964 19464 991
rect 19412 930 19426 964
rect 19426 930 19460 964
rect 19460 930 19464 964
rect 19696 1001 19757 1012
rect 19790 1001 19851 1012
rect 19696 967 19699 1001
rect 19699 967 19735 1001
rect 19735 967 19757 1001
rect 19790 967 19809 1001
rect 19809 967 19851 1001
rect 19696 960 19757 967
rect 19790 960 19851 967
rect 19449 644 20024 718
rect 20061 426 20113 459
rect 19363 392 19424 404
rect 19457 392 19518 404
rect 19363 358 19366 392
rect 19366 358 19402 392
rect 19402 358 19424 392
rect 19457 358 19476 392
rect 19476 358 19518 392
rect 19363 352 19424 358
rect 19457 352 19518 358
rect 20061 398 20090 426
rect 20090 398 20113 426
rect 20061 352 20113 365
rect 20061 316 20090 352
rect 20090 316 20113 352
rect 20061 304 20113 316
rect 16703 120 16770 159
rect 16770 120 17860 159
rect 17860 120 18070 159
rect 18070 120 19270 159
rect 19270 120 19290 159
rect 16703 99 19290 120
rect 19444 96 20040 158
<< metal2 >>
rect 9990 2120 10050 2130
rect 10080 2120 10140 2130
rect 10050 2050 10080 2090
rect 9990 2040 10140 2050
rect 11780 2120 11840 2130
rect 11870 2120 11930 2130
rect 11840 2050 11870 2090
rect 11780 2040 11930 2050
rect 12960 2120 13020 2130
rect 13050 2120 13110 2130
rect 13020 2050 13050 2100
rect 15230 2120 15390 2130
rect 15290 2060 15330 2120
rect 15230 2050 15390 2060
rect 12960 2040 13110 2050
rect 10020 1130 10120 2040
rect 11780 1130 11880 2040
rect 12970 1130 13070 2040
rect 15240 1130 15340 2050
rect 15618 1265 20034 1388
rect 15618 1212 16157 1265
rect 16470 1243 20034 1265
rect 16470 1212 16986 1243
rect 9985 1078 9995 1130
rect 10056 1078 10089 1130
rect 10150 1078 10160 1130
rect 11765 1078 11775 1130
rect 11836 1078 11869 1130
rect 11930 1078 11940 1130
rect 12945 1078 12955 1130
rect 13016 1078 13049 1130
rect 13110 1078 13120 1130
rect 15215 1078 15225 1130
rect 15286 1078 15319 1130
rect 15380 1078 15390 1130
rect 15850 1109 15880 1212
rect 16194 1141 16230 1193
rect 16291 1141 16324 1193
rect 16385 1170 16395 1193
rect 16976 1191 16986 1212
rect 17047 1191 17080 1243
rect 17141 1212 17651 1243
rect 17141 1191 17151 1212
rect 17641 1191 17651 1212
rect 17712 1191 17745 1243
rect 17806 1212 20034 1243
rect 17806 1191 17816 1212
rect 19634 1187 19834 1212
rect 16385 1141 16816 1170
rect 16194 1133 16816 1141
rect 18130 1133 18178 1184
rect 16194 1132 18178 1133
rect 18239 1132 18272 1184
rect 18333 1170 18343 1184
rect 19005 1170 19015 1184
rect 18333 1132 19015 1170
rect 19076 1132 19109 1184
rect 19170 1170 19180 1184
rect 19170 1132 19450 1170
rect 16194 1130 19450 1132
rect 15839 1099 15891 1109
rect 10020 278 10120 1078
rect 11780 278 11880 1078
rect 12970 278 13070 1078
rect 15240 850 15340 1078
rect 16767 1093 18178 1130
rect 19420 1095 19450 1130
rect 19412 1085 19464 1095
rect 15839 1005 15891 1038
rect 15839 934 15891 944
rect 17035 1053 17087 1063
rect 18219 1053 18271 1063
rect 17087 992 18219 1004
rect 17035 959 18271 992
rect 17087 956 18219 959
rect 17035 888 17087 898
rect 19412 991 19464 1024
rect 19412 920 19464 930
rect 19685 1012 19885 1078
rect 19685 960 19696 1012
rect 19757 960 19790 1012
rect 19851 960 19885 1012
rect 18219 888 18271 898
rect 18649 889 18701 899
rect 15240 828 18649 850
rect 19059 879 19111 889
rect 18701 828 19059 850
rect 15240 818 19059 828
rect 19685 878 19885 960
rect 15240 800 19111 818
rect 9983 226 9993 278
rect 10054 226 10087 278
rect 10148 226 10158 278
rect 11755 226 11765 278
rect 11826 226 11859 278
rect 11920 226 11930 278
rect 12935 226 12945 278
rect 13006 226 13039 278
rect 13100 226 13110 278
rect 15240 276 15340 800
rect 18649 795 18701 800
rect 16151 757 16203 767
rect 16343 757 16395 767
rect 16203 696 16343 700
rect 16710 725 16910 740
rect 16710 700 16797 725
rect 16395 696 16797 700
rect 16151 686 16797 696
rect 15936 664 16797 686
rect 16849 700 16910 725
rect 17273 725 17325 735
rect 16849 664 17273 700
rect 17541 727 17593 737
rect 17325 666 17541 700
rect 18649 724 18701 734
rect 19059 785 19111 800
rect 19942 728 20033 1212
rect 19059 714 19111 724
rect 19449 718 20033 728
rect 17325 664 17593 666
rect 15936 663 17593 664
rect 15936 654 16151 663
rect 15211 224 15221 276
rect 15282 224 15315 276
rect 15376 224 15386 276
rect 15713 213 15723 265
rect 15784 213 15817 265
rect 15878 257 15888 265
rect 15936 257 15968 654
rect 16203 648 16343 663
rect 16151 592 16203 602
rect 16395 648 17593 663
rect 16343 592 16395 602
rect 16710 631 16910 648
rect 16710 570 16797 631
rect 16849 570 16910 631
rect 16047 551 16099 561
rect 16239 551 16291 561
rect 16099 490 16239 494
rect 16431 551 16483 561
rect 16291 490 16431 494
rect 16710 540 16910 570
rect 17273 631 17325 648
rect 17273 560 17325 570
rect 17541 633 17593 648
rect 18574 646 18774 660
rect 17541 562 17593 572
rect 18545 636 18795 646
rect 18597 575 18743 636
rect 20024 644 20033 718
rect 19449 634 20033 644
rect 18545 542 18795 575
rect 16047 457 16483 490
rect 16099 442 16239 457
rect 16047 386 16099 396
rect 16291 442 16431 457
rect 16239 386 16291 396
rect 16431 386 16483 396
rect 17779 529 17831 539
rect 18597 481 18743 542
rect 18545 471 18795 481
rect 17779 435 17831 468
rect 18574 460 18774 471
rect 19979 459 20179 479
rect 17831 374 19363 404
rect 17779 364 19363 374
rect 17780 352 19363 364
rect 19424 352 19457 404
rect 19518 352 19528 404
rect 19979 398 20061 459
rect 20113 398 20179 459
rect 19979 365 20179 398
rect 15878 256 18583 257
rect 15878 225 18593 256
rect 15878 213 15888 225
rect 18583 204 18593 225
rect 18654 204 18687 256
rect 18748 204 18758 256
rect 19667 170 19867 347
rect 19979 304 20061 365
rect 20113 304 20179 365
rect 19979 279 20179 304
rect 16657 159 20126 170
rect 16657 99 16703 159
rect 19290 158 20126 159
rect 19290 99 19444 158
rect 16657 96 19444 99
rect 20040 96 20126 158
rect 16657 77 20126 96
use sky130_fd_pr__pfet_01v8_7FRQHJ  sky130_fd_pr__pfet_01v8_7FRQHJ_0
timestamp 1711831168
transform 1 0 12471 0 1 1171
box -3225 -1087 3225 1087
use sky130_fd_pr__pfet_01v8_XG6TDL  sky130_fd_pr__pfet_01v8_XG6TDL_0
timestamp 1710675123
transform 1 0 16265 0 1 703
box -359 -619 359 619
use sky130_fd_sc_hd__inv_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 19850 0 -1 1225
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19390 0 1 137
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x3
timestamp 1710522493
transform 1 0 19666 0 1 137
box -38 -48 498 592
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1710675955
transform 1 0 15801 0 1 403
box -211 -319 211 319
use sky130_fd_pr__nfet_05v0_nvt_F93ZEE  XM3
timestamp 1710675123
transform 1 0 17061 0 1 730
box -437 -658 437 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM4
timestamp 1710677421
transform 1 0 18249 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_01v8_6EHS5V  XM5
timestamp 1710677421
transform 1 0 19089 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_05v0_nvt_JFFQEL  XM7
timestamp 1710675123
transform 1 0 17686 0 1 730
box -318 -658 318 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM8
timestamp 1710677421
transform 1 0 18669 0 -1 694
box -263 -610 263 610
<< labels >>
flabel metal2 15707 1286 15763 1337 0 FreeSans 800 0 0 0 VDD
flabel metal1 11070 600 11130 660 0 FreeSans 800 0 0 0 Vtop
flabel metal2 16238 666 16278 688 0 FreeSans 800 0 0 0 Vgate
flabel metal2 17672 968 17696 982 0 FreeSans 800 0 0 0 Vd
flabel metal2 18486 360 18516 390 0 FreeSans 800 0 0 0 VGATE_1V8
flabel metal2 18844 810 18876 829 0 FreeSans 800 0 0 0 Vbottom
flabel metal2 18937 1141 18963 1157 0 FreeSans 800 0 0 0 EN_Z
flabel metal2 16710 540 16910 740 0 FreeSans 256 0 0 0 VGATE
port 5 nsew
flabel metal2 19685 878 19885 1078 0 FreeSans 256 0 0 0 EN
port 4 nsew
flabel metal2 19979 279 20179 479 0 FreeSans 256 0 0 0 SW_ON
port 3 nsew
flabel metal2 18574 460 18774 660 0 FreeSans 256 0 0 0 VIN
port 2 nsew
flabel metal2 19667 147 19867 347 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal2 19634 1187 19834 1387 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 11069 1604 11129 1664 0 FreeSans 800 0 0 0 Vtop
<< end >>
