magic
tech sky130A
magscale 1 2
timestamp 1714236875
<< metal1 >>
rect 1815 7597 1845 11260
rect 1875 9985 1905 11260
rect 1935 10045 1965 11260
rect 1995 10105 2025 11260
rect 2055 10165 2085 11260
rect 2115 10225 2145 11260
rect 2175 10285 2205 11260
rect 2235 10344 2265 11260
rect 2295 10405 2325 11260
rect 2355 10465 2385 11260
rect 2415 10525 2445 11260
rect 2475 10610 2505 11260
rect 2535 10670 2565 11260
rect 2595 10730 2625 11260
rect 2655 10790 2685 11260
rect 2715 10850 2745 11260
rect 2775 10910 2805 11260
rect 2835 10970 2865 11260
rect 2895 11030 2925 11260
rect 2955 11090 2985 11260
rect 3015 11150 3045 11260
rect 3075 11210 3105 11260
rect 3075 11180 6230 11210
rect 3015 11120 6155 11150
rect 2955 11060 6080 11090
rect 2895 11000 6004 11030
rect 2835 10940 5930 10970
rect 2775 10880 5855 10910
rect 2715 10820 5780 10850
rect 2655 10760 5704 10790
rect 2595 10700 5630 10730
rect 2535 10640 5555 10670
rect 2475 10580 5480 10610
rect 2415 10495 2595 10525
rect 2355 10435 2520 10465
rect 2295 10375 2445 10405
rect 2235 10315 2370 10344
rect 2175 10255 2295 10285
rect 2115 10195 2220 10225
rect 2055 10135 2145 10165
rect 1995 10075 2070 10105
rect 1935 10015 1995 10045
rect 1875 9945 1920 9985
rect 1890 7718 1920 9945
rect 1965 8053 1995 10015
rect 2040 8284 2070 10075
rect 2115 8685 2145 10135
rect 2190 8806 2220 10195
rect 2265 9141 2295 10255
rect 2341 9311 2370 10315
rect 2415 9773 2445 10375
rect 2490 9933 2520 10435
rect 2565 10399 2595 10495
rect 2550 10389 2610 10399
rect 2605 10329 2610 10389
rect 2550 10319 2610 10329
rect 2550 10149 2610 10159
rect 2605 10089 2610 10149
rect 2550 10079 2610 10089
rect 2475 9923 2535 9933
rect 2530 9863 2535 9923
rect 2475 9853 2535 9863
rect 2400 9763 2460 9773
rect 2455 9703 2460 9763
rect 2400 9693 2460 9703
rect 2475 9633 2535 9643
rect 2530 9573 2535 9633
rect 2475 9563 2535 9573
rect 2400 9513 2460 9523
rect 2455 9453 2460 9513
rect 2400 9443 2460 9453
rect 2326 9301 2386 9311
rect 2381 9241 2386 9301
rect 2326 9231 2386 9241
rect 2250 9131 2310 9141
rect 2305 9071 2310 9131
rect 2250 9061 2310 9071
rect 2326 9028 2386 9038
rect 2381 8968 2386 9028
rect 2326 8958 2386 8968
rect 2250 8924 2310 8934
rect 2305 8864 2310 8924
rect 2250 8854 2310 8864
rect 2176 8796 2236 8806
rect 2231 8736 2236 8796
rect 2176 8726 2236 8736
rect 2100 8675 2160 8685
rect 2155 8615 2160 8675
rect 2100 8605 2160 8615
rect 2176 8545 2236 8555
rect 2231 8485 2236 8545
rect 2176 8475 2236 8485
rect 2100 8425 2160 8435
rect 2155 8365 2160 8425
rect 2100 8355 2160 8365
rect 2041 8223 2070 8284
rect 2026 8213 2086 8223
rect 2081 8153 2086 8213
rect 2026 8143 2086 8153
rect 1950 8043 2010 8053
rect 2005 7983 2010 8043
rect 1950 7973 2010 7983
rect 2026 7940 2086 7950
rect 2081 7880 2086 7940
rect 2026 7870 2086 7880
rect 1950 7836 2010 7846
rect 2005 7776 2010 7836
rect 1950 7766 2010 7776
rect 1876 7708 1936 7718
rect 1931 7648 1936 7708
rect 1876 7638 1936 7648
rect 1800 7587 1860 7597
rect 1855 7527 1860 7587
rect 1800 7517 1860 7527
rect 1876 7457 1936 7467
rect 1931 7397 1936 7457
rect 1876 7387 1936 7397
rect 1800 7337 1860 7347
rect 1855 7277 1860 7337
rect 1800 7267 1860 7277
rect 1815 5890 1845 7267
rect 1890 7195 1920 7387
rect 1875 7145 1920 7195
rect 1875 5890 1905 7145
rect 1965 7115 1995 7766
rect 1935 7085 1995 7115
rect 1935 5890 1965 7085
rect 2040 7055 2070 7870
rect 1995 7025 2070 7055
rect 1995 5890 2025 7025
rect 2115 6995 2145 8355
rect 2055 6965 2145 6995
rect 2055 5890 2085 6965
rect 2190 6935 2220 8475
rect 2115 6905 2220 6935
rect 2115 5890 2145 6905
rect 2265 6875 2295 8854
rect 2175 6845 2295 6875
rect 2175 5890 2205 6845
rect 2341 6815 2370 8958
rect 2235 6786 2370 6815
rect 2235 6785 2365 6786
rect 2235 5890 2265 6785
rect 2415 6755 2445 9443
rect 2295 6725 2445 6755
rect 2295 5890 2325 6725
rect 2490 6695 2520 9563
rect 2355 6665 2520 6695
rect 2355 5890 2385 6665
rect 2565 6635 2595 10079
rect 5450 7632 5480 10580
rect 5525 7741 5555 10640
rect 5600 8182 5630 10700
rect 5675 8304 5704 10760
rect 5750 8720 5780 10820
rect 5825 8829 5855 10880
rect 5900 9270 5930 10940
rect 5975 9392 6004 11000
rect 6050 9808 6080 11060
rect 6125 9917 6155 11120
rect 6200 10433 6230 11180
rect 6185 10423 6245 10433
rect 6185 10363 6190 10423
rect 6185 10353 6245 10363
rect 6185 10213 6245 10223
rect 6185 10153 6190 10213
rect 6185 10143 6245 10153
rect 6110 9907 6170 9917
rect 6110 9847 6115 9907
rect 6110 9837 6170 9847
rect 6035 9798 6095 9808
rect 6035 9738 6040 9798
rect 6035 9728 6095 9738
rect 6110 9667 6170 9677
rect 6110 9607 6115 9667
rect 6110 9597 6170 9607
rect 6035 9517 6095 9527
rect 6035 9457 6040 9517
rect 6035 9447 6095 9457
rect 5975 9385 6005 9392
rect 5960 9375 6020 9385
rect 5960 9315 5965 9375
rect 5960 9305 6020 9315
rect 5885 9260 5945 9270
rect 5885 9200 5890 9260
rect 5885 9190 5945 9200
rect 5960 9125 6020 9135
rect 5960 9065 5965 9125
rect 5960 9055 6020 9065
rect 5975 9052 6005 9055
rect 5885 8995 5945 9005
rect 5885 8935 5890 8995
rect 5885 8925 5945 8935
rect 5810 8819 5870 8829
rect 5810 8759 5815 8819
rect 5810 8749 5870 8759
rect 5735 8710 5795 8720
rect 5735 8650 5740 8710
rect 5735 8640 5795 8650
rect 5810 8579 5870 8589
rect 5810 8519 5815 8579
rect 5810 8509 5870 8519
rect 5735 8429 5795 8439
rect 5735 8369 5740 8429
rect 5735 8359 5795 8369
rect 5675 8297 5705 8304
rect 5660 8287 5720 8297
rect 5660 8227 5665 8287
rect 5660 8217 5720 8227
rect 5585 8172 5645 8182
rect 5585 8112 5590 8172
rect 5585 8102 5645 8112
rect 5660 8037 5720 8047
rect 5660 7977 5665 8037
rect 5660 7967 5720 7977
rect 5675 7964 5705 7967
rect 5585 7907 5645 7917
rect 5585 7847 5590 7907
rect 5585 7837 5645 7847
rect 5510 7731 5570 7741
rect 5510 7671 5515 7731
rect 5510 7661 5570 7671
rect 5435 7622 5495 7632
rect 5435 7562 5440 7622
rect 5435 7552 5495 7562
rect 5510 7491 5570 7501
rect 5510 7431 5515 7491
rect 5510 7421 5570 7431
rect 5435 7341 5495 7351
rect 5435 7281 5440 7341
rect 5435 7271 5495 7281
rect 5450 7148 5480 7271
rect 2415 6605 2595 6635
rect 2625 7118 5480 7148
rect 2415 5890 2445 6605
rect 2625 6575 2655 7118
rect 5525 7088 5555 7421
rect 2475 6545 2655 6575
rect 2685 7058 5555 7088
rect 2475 5890 2505 6545
rect 2685 6515 2715 7058
rect 5600 7028 5630 7837
rect 2535 6485 2715 6515
rect 2745 7003 5630 7028
rect 5675 7241 5704 7964
rect 2745 6998 5626 7003
rect 2535 5890 2565 6485
rect 2745 6455 2775 6998
rect 5675 6968 5705 7241
rect 2595 6425 2775 6455
rect 2805 6938 5705 6968
rect 2595 5890 2625 6425
rect 2805 6395 2835 6938
rect 5750 6908 5780 8359
rect 2655 6365 2835 6395
rect 2865 6878 5780 6908
rect 2655 5890 2685 6365
rect 2865 6335 2895 6878
rect 5825 6848 5855 8509
rect 2715 6305 2895 6335
rect 2925 6818 5855 6848
rect 2715 5890 2745 6305
rect 2925 6275 2955 6818
rect 5900 6788 5930 8925
rect 2775 6245 2955 6275
rect 2985 6758 5930 6788
rect 5975 7241 6004 9052
rect 2775 5890 2805 6245
rect 2985 6215 3015 6758
rect 5975 6728 6005 7241
rect 2835 6185 3015 6215
rect 3045 6698 6005 6728
rect 2835 5890 2865 6185
rect 3045 6155 3075 6698
rect 6050 6668 6080 9447
rect 2895 6125 3075 6155
rect 3105 6638 6080 6668
rect 2895 5890 2925 6125
rect 3105 6095 3135 6638
rect 6125 6608 6155 9597
rect 2955 6065 3135 6095
rect 3165 6578 6155 6608
rect 2955 5890 2985 6065
rect 3165 6035 3195 6578
rect 6200 6548 6230 10143
rect 3226 6545 6230 6548
rect 3015 6005 3195 6035
rect 3225 6520 6230 6545
rect 3015 5890 3045 6005
rect 3225 5975 3255 6520
rect 3075 5945 3255 5975
rect 3075 5890 3105 5945
<< via1 >>
rect 2550 10329 2605 10389
rect 2550 10089 2605 10149
rect 2475 9863 2530 9923
rect 2400 9703 2455 9763
rect 2475 9573 2530 9633
rect 2400 9453 2455 9513
rect 2326 9241 2381 9301
rect 2250 9071 2305 9131
rect 2326 8968 2381 9028
rect 2250 8864 2305 8924
rect 2176 8736 2231 8796
rect 2100 8615 2155 8675
rect 2176 8485 2231 8545
rect 2100 8365 2155 8425
rect 2026 8153 2081 8213
rect 1950 7983 2005 8043
rect 2026 7880 2081 7940
rect 1950 7776 2005 7836
rect 1876 7648 1931 7708
rect 1800 7527 1855 7587
rect 1876 7397 1931 7457
rect 1800 7277 1855 7337
rect 6190 10363 6245 10423
rect 6190 10153 6245 10213
rect 6115 9847 6170 9907
rect 6040 9738 6095 9798
rect 6115 9607 6170 9667
rect 6040 9457 6095 9517
rect 5965 9315 6020 9375
rect 5890 9200 5945 9260
rect 5965 9065 6020 9125
rect 5890 8935 5945 8995
rect 5815 8759 5870 8819
rect 5740 8650 5795 8710
rect 5815 8519 5870 8579
rect 5740 8369 5795 8429
rect 5665 8227 5720 8287
rect 5590 8112 5645 8172
rect 5665 7977 5720 8037
rect 5590 7847 5645 7907
rect 5515 7671 5570 7731
rect 5440 7562 5495 7622
rect 5515 7431 5570 7491
rect 5440 7281 5495 7341
<< metal2 >>
rect 6185 10423 6245 10433
rect 6185 10411 6190 10423
rect 2550 10389 2610 10399
rect 2605 10371 2610 10389
rect 5410 10381 6190 10411
rect 2605 10341 2686 10371
rect 6185 10363 6190 10381
rect 6185 10353 6245 10363
rect 2605 10329 2610 10341
rect 2550 10319 2610 10329
rect 6185 10213 6245 10223
rect 6185 10211 6190 10213
rect 5410 10181 6190 10211
rect 2550 10149 2610 10159
rect 2605 10131 2610 10149
rect 6185 10153 6190 10181
rect 6185 10143 6245 10153
rect 2605 10101 2665 10131
rect 2605 10089 2610 10101
rect 2550 10079 2610 10089
rect 2475 9923 2535 9933
rect 2530 9905 2535 9923
rect 6110 9907 6170 9917
rect 2530 9875 2670 9905
rect 6110 9895 6115 9907
rect 2530 9863 2535 9875
rect 5392 9865 6115 9895
rect 2475 9853 2535 9863
rect 6110 9847 6115 9865
rect 6110 9837 6170 9847
rect 6035 9798 6095 9808
rect 6035 9786 6040 9798
rect 2400 9763 2460 9773
rect 2455 9745 2460 9763
rect 5395 9756 6040 9786
rect 2455 9715 2665 9745
rect 6035 9738 6040 9756
rect 6035 9728 6095 9738
rect 2455 9703 2460 9715
rect 2400 9693 2460 9703
rect 6110 9667 6170 9677
rect 6110 9665 6115 9667
rect 2475 9633 2535 9643
rect 5395 9635 6115 9665
rect 2530 9615 2535 9633
rect 2530 9585 2677 9615
rect 6110 9607 6115 9635
rect 6110 9597 6170 9607
rect 2530 9573 2535 9585
rect 2475 9563 2535 9573
rect 2400 9513 2460 9523
rect 6035 9517 6095 9527
rect 6035 9515 6040 9517
rect 2455 9495 2460 9513
rect 2455 9465 2683 9495
rect 5395 9485 6040 9515
rect 2455 9453 2460 9465
rect 2400 9443 2460 9453
rect 6035 9457 6040 9485
rect 6035 9447 6095 9457
rect 5960 9375 6020 9385
rect 5960 9363 5965 9375
rect 5390 9333 5965 9363
rect 5960 9315 5965 9333
rect 2326 9301 2386 9311
rect 5960 9305 6020 9315
rect 2381 9283 2386 9301
rect 2381 9253 2692 9283
rect 5885 9260 5945 9270
rect 2381 9241 2386 9253
rect 5885 9248 5890 9260
rect 2326 9231 2386 9241
rect 5395 9218 5890 9248
rect 5885 9200 5890 9218
rect 5885 9190 5945 9200
rect 2250 9131 2310 9141
rect 2305 9113 2310 9131
rect 5960 9125 6020 9135
rect 5960 9123 5965 9125
rect 2305 9083 2685 9113
rect 5395 9093 5965 9123
rect 2305 9071 2310 9083
rect 2250 9061 2310 9071
rect 5960 9065 5965 9093
rect 5960 9055 6020 9065
rect 2326 9028 2386 9038
rect 2381 9010 2386 9028
rect 2381 8980 2665 9010
rect 5885 8995 5945 9005
rect 5885 8993 5890 8995
rect 2381 8968 2386 8980
rect 2326 8958 2386 8968
rect 5395 8963 5890 8993
rect 5885 8935 5890 8963
rect 2250 8924 2310 8934
rect 5885 8925 5945 8935
rect 2305 8906 2310 8924
rect 2305 8876 2665 8906
rect 2305 8864 2310 8876
rect 2250 8854 2310 8864
rect 5810 8819 5870 8829
rect 5810 8807 5815 8819
rect 2176 8796 2236 8806
rect 2231 8778 2236 8796
rect 2231 8748 2665 8778
rect 5395 8777 5815 8807
rect 5810 8759 5815 8777
rect 5810 8749 5870 8759
rect 2231 8736 2236 8748
rect 2176 8726 2236 8736
rect 5735 8710 5795 8720
rect 5735 8698 5740 8710
rect 2100 8675 2160 8685
rect 2155 8657 2160 8675
rect 5395 8668 5740 8698
rect 2155 8627 2665 8657
rect 5735 8650 5740 8668
rect 5735 8640 5795 8650
rect 2155 8615 2160 8627
rect 2100 8605 2160 8615
rect 5810 8579 5870 8589
rect 5810 8577 5815 8579
rect 2176 8545 2236 8555
rect 5395 8547 5815 8577
rect 2231 8527 2236 8545
rect 2231 8497 2682 8527
rect 5810 8519 5815 8547
rect 5810 8509 5870 8519
rect 2231 8485 2236 8497
rect 2176 8475 2236 8485
rect 2100 8425 2160 8435
rect 5735 8429 5795 8439
rect 5735 8427 5740 8429
rect 2155 8407 2160 8425
rect 2155 8377 2665 8407
rect 5389 8397 5740 8427
rect 2155 8365 2160 8377
rect 2100 8355 2160 8365
rect 5735 8369 5740 8397
rect 5735 8359 5795 8369
rect 5660 8287 5720 8297
rect 5660 8275 5665 8287
rect 5411 8245 5665 8275
rect 5660 8227 5665 8245
rect 2026 8213 2086 8223
rect 5660 8217 5720 8227
rect 2081 8195 2086 8213
rect 2081 8165 2685 8195
rect 5585 8172 5645 8182
rect 2081 8153 2086 8165
rect 5585 8160 5590 8172
rect 2026 8143 2086 8153
rect 5411 8130 5590 8160
rect 5585 8112 5590 8130
rect 5585 8102 5645 8112
rect 1950 8043 2010 8053
rect 2005 8025 2010 8043
rect 5660 8037 5720 8047
rect 5660 8035 5665 8037
rect 2005 7995 2665 8025
rect 5411 8005 5665 8035
rect 2005 7983 2010 7995
rect 1950 7973 2010 7983
rect 5660 7977 5665 8005
rect 5660 7967 5720 7977
rect 2026 7940 2086 7950
rect 2081 7922 2086 7940
rect 2081 7892 2668 7922
rect 5585 7907 5645 7917
rect 5585 7905 5590 7907
rect 2081 7880 2086 7892
rect 2026 7870 2086 7880
rect 5411 7875 5590 7905
rect 5585 7847 5590 7875
rect 1950 7836 2010 7846
rect 5585 7837 5645 7847
rect 2005 7818 2010 7836
rect 2005 7788 2666 7818
rect 2005 7776 2010 7788
rect 1950 7766 2010 7776
rect 5510 7731 5570 7741
rect 5510 7719 5515 7731
rect 1876 7708 1936 7718
rect 1931 7690 1936 7708
rect 1931 7660 2665 7690
rect 5411 7689 5515 7719
rect 5510 7671 5515 7689
rect 5510 7661 5570 7671
rect 1931 7648 1936 7660
rect 1876 7638 1936 7648
rect 5435 7622 5495 7632
rect 5435 7610 5440 7622
rect 1800 7587 1860 7597
rect 1855 7569 1860 7587
rect 5411 7580 5440 7610
rect 1855 7539 2665 7569
rect 5435 7562 5440 7580
rect 5435 7552 5495 7562
rect 1855 7527 1860 7539
rect 1800 7517 1860 7527
rect 5510 7491 5570 7501
rect 5510 7489 5515 7491
rect 1876 7457 1936 7467
rect 5411 7459 5515 7489
rect 1931 7439 1936 7457
rect 1931 7409 2678 7439
rect 5510 7431 5515 7459
rect 5510 7421 5570 7431
rect 1931 7397 1936 7409
rect 1876 7387 1936 7397
rect 1800 7337 1860 7347
rect 5435 7341 5495 7351
rect 5435 7339 5440 7341
rect 1855 7319 1860 7337
rect 1855 7289 2666 7319
rect 5411 7309 5440 7339
rect 1855 7277 1860 7289
rect 1800 7267 1860 7277
rect 5435 7281 5440 7309
rect 5435 7271 5495 7281
use bbm_unit_x3  bbm_unit_x3_0
timestamp 1714230552
transform 1 0 4135 0 1 9381
box -1500 -20 1290 1164
use bbm_unit_x4  bbm_unit_x4_0
timestamp 1714234260
transform 1 0 4135 0 1 8293
box -1500 -20 1290 1164
use bbm_unit_x4  bbm_unit_x4_1
timestamp 1714234260
transform 1 0 4135 0 1 7205
box -1500 -20 1290 1164
<< end >>
