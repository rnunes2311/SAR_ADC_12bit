magic
tech sky130A
magscale 1 2
timestamp 1712002773
<< locali >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2830 10170 2870
rect 3700 2810 10170 2830
rect 3700 2770 3800 2810
rect 3700 -1770 3710 2770
rect 3780 -1770 3800 2770
rect 10310 -830 10340 -770
rect 3700 -1830 3800 -1770
rect 3700 -1840 10140 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1890 10140 -1840
rect 3700 -1900 10140 -1890
<< viali >>
rect 3830 2830 10100 2870
rect 3710 -1770 3780 2770
rect 10130 -540 10170 2740
rect 10360 2514 10426 2562
rect 10511 2512 10577 2562
rect 10680 2512 10747 2566
rect 10280 2410 10330 2470
rect 10600 2350 10650 2410
rect 10280 2077 10330 2127
rect 10362 1904 10423 1953
rect 10511 1904 10578 1954
rect 10680 1900 10747 1954
rect 10519 1789 10580 1838
rect 10280 1520 10340 1580
rect 10629 1570 10663 1604
rect 10360 1426 10426 1474
rect 10507 1424 10570 1490
rect 10620 1430 10680 1490
rect 10800 1430 10860 1500
rect 10360 961 10425 1009
rect 10634 977 10699 1025
rect 10278 816 10343 864
rect 10554 816 10619 864
rect 10250 -830 10310 -770
rect 3820 -1890 10100 -1840
<< metal1 >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2830 10170 2870
rect 3700 2810 10170 2830
rect 10210 2810 11700 2900
rect 3700 2770 3800 2810
rect 3700 -1770 3710 2770
rect 3780 1840 3800 2770
rect 10130 2752 10170 2810
rect 6880 2740 6890 2750
rect 3900 2690 6890 2740
rect 6950 2740 6960 2750
rect 10124 2740 10176 2752
rect 6950 2690 10020 2740
rect 10124 1840 10130 2740
rect 3780 1500 10130 1840
rect 3780 -600 3800 1500
rect 6880 610 6890 620
rect 3890 560 6890 610
rect 6950 610 6960 620
rect 6950 560 10010 610
rect 6880 410 6890 420
rect 3890 360 6890 410
rect 6950 410 6960 420
rect 6950 360 10010 410
rect 9730 70 9740 130
rect 9800 70 9810 130
rect 9750 -460 9790 70
rect 10124 -70 10130 1500
rect 10170 2280 10176 2740
rect 10670 2572 10680 2580
rect 10510 2568 10520 2570
rect 10348 2562 10438 2568
rect 10348 2514 10360 2562
rect 10426 2514 10438 2562
rect 10348 2508 10438 2514
rect 10499 2562 10520 2568
rect 10499 2512 10511 2562
rect 10499 2510 10520 2512
rect 10580 2510 10590 2570
rect 10668 2510 10680 2572
rect 10750 2510 10760 2580
rect 11000 2520 11010 2580
rect 11070 2520 11080 2580
rect 10274 2470 10336 2482
rect 10250 2410 10260 2470
rect 10330 2410 10336 2470
rect 10274 2398 10336 2410
rect 10378 2392 10410 2508
rect 10499 2506 10589 2510
rect 10668 2506 10759 2510
rect 10594 2410 10656 2422
rect 10594 2400 10600 2410
rect 10650 2400 10656 2410
rect 10580 2392 10590 2400
rect 10378 2347 10590 2392
rect 10580 2340 10590 2347
rect 10650 2340 10660 2400
rect 10594 2338 10656 2340
rect 10170 2190 10270 2280
rect 10170 1190 10176 2190
rect 10270 2133 10280 2137
rect 10268 2077 10280 2133
rect 10340 2077 10350 2137
rect 10268 2071 10342 2077
rect 11030 1960 11060 2520
rect 11100 2430 11110 2490
rect 11170 2430 11180 2490
rect 10350 1953 10435 1959
rect 10350 1904 10362 1953
rect 10423 1904 10435 1953
rect 10350 1898 10435 1904
rect 10499 1900 10510 1960
rect 10570 1954 10590 1960
rect 10578 1904 10590 1954
rect 10570 1900 10590 1904
rect 10499 1898 10590 1900
rect 10390 1830 10420 1898
rect 10668 1894 10680 1960
rect 10670 1890 10680 1894
rect 10750 1890 10760 1960
rect 11000 1900 11010 1960
rect 11070 1900 11080 1960
rect 10510 1844 10520 1850
rect 10507 1838 10520 1844
rect 10580 1844 10590 1850
rect 10507 1830 10519 1838
rect 10390 1800 10519 1830
rect 10507 1789 10519 1800
rect 10580 1789 10592 1844
rect 10920 1790 10930 1850
rect 10990 1790 11000 1850
rect 10507 1783 10592 1789
rect 10750 1650 10760 1720
rect 10830 1650 10840 1720
rect 10597 1604 10679 1611
rect 10597 1600 10629 1604
rect 10663 1600 10679 1604
rect 10597 1590 10620 1600
rect 10268 1580 10352 1586
rect 10268 1520 10280 1580
rect 10340 1520 10352 1580
rect 10268 1514 10352 1520
rect 10400 1560 10620 1590
rect 10400 1480 10430 1560
rect 10610 1540 10620 1560
rect 10680 1540 10690 1600
rect 10501 1500 10576 1502
rect 10794 1500 10880 1512
rect 10490 1490 10580 1500
rect 10348 1474 10438 1480
rect 10348 1426 10360 1474
rect 10426 1426 10438 1474
rect 10348 1420 10438 1426
rect 10490 1424 10507 1490
rect 10570 1424 10580 1490
rect 10608 1490 10692 1496
rect 10794 1490 10800 1500
rect 10608 1430 10620 1490
rect 10680 1430 10692 1490
rect 10790 1430 10800 1490
rect 10860 1430 10880 1500
rect 10608 1424 10692 1430
rect 10490 1406 10580 1424
rect 10490 1340 10500 1406
rect 10563 1340 10580 1406
rect 10640 1290 10670 1424
rect 10794 1418 10880 1430
rect 10810 1417 10880 1418
rect 10810 1300 10850 1417
rect 10540 1230 10550 1290
rect 10610 1240 10670 1290
rect 10790 1240 10800 1300
rect 10860 1240 10870 1300
rect 10610 1230 10620 1240
rect 10170 1100 10260 1190
rect 10170 150 10176 1100
rect 10622 1030 10711 1031
rect 10350 1015 10360 1020
rect 10348 960 10360 1015
rect 10420 1015 10430 1020
rect 10420 1009 10437 1015
rect 10425 961 10437 1009
rect 10620 970 10630 1030
rect 10700 971 10711 1030
rect 10700 970 10710 971
rect 10420 960 10437 961
rect 10348 955 10437 960
rect 10266 864 10355 870
rect 10266 860 10278 864
rect 10260 816 10278 860
rect 10343 816 10355 864
rect 10260 810 10355 816
rect 10540 810 10550 870
rect 10610 864 10631 870
rect 10619 816 10631 864
rect 10610 810 10631 816
rect 10260 740 10350 810
rect 10260 680 10270 740
rect 10330 690 10350 740
rect 10330 680 10340 690
rect 10720 630 10740 649
rect 10680 560 10690 630
rect 10760 560 10770 630
rect 10570 380 10580 440
rect 10640 380 10650 440
rect 10370 180 10380 250
rect 10450 180 10460 250
rect 10590 190 10620 380
rect 10170 60 10260 150
rect 10328 132 10388 142
rect 10436 132 10496 142
rect 10670 80 10780 110
rect 10328 62 10344 72
rect 10436 62 10496 72
rect 10170 -70 10176 60
rect 10270 -40 10280 20
rect 10340 -40 10350 20
rect 10110 -130 10120 -70
rect 10180 -130 10190 -70
rect 9730 -520 9740 -460
rect 9800 -520 9810 -460
rect 10124 -540 10130 -130
rect 10170 -270 10176 -130
rect 10290 -220 10340 -40
rect 10480 -170 10540 20
rect 10750 -70 10780 80
rect 10820 70 10830 130
rect 10890 70 10900 130
rect 10730 -130 10740 -70
rect 10800 -130 10810 -70
rect 10470 -230 10480 -170
rect 10540 -230 10550 -170
rect 10170 -360 10260 -270
rect 10328 -280 10388 -270
rect 10436 -280 10496 -270
rect 10750 -300 10780 -130
rect 10660 -330 10780 -300
rect 10328 -350 10344 -340
rect 10436 -350 10496 -340
rect 10170 -440 10176 -360
rect 10170 -540 10180 -440
rect 10370 -460 10380 -390
rect 10450 -460 10460 -390
rect 10124 -600 10180 -540
rect 10590 -580 10620 -410
rect 3780 -940 10180 -600
rect 10560 -640 10570 -580
rect 10630 -640 10640 -580
rect 10240 -670 10330 -660
rect 10240 -730 10260 -670
rect 10320 -730 10330 -670
rect 10730 -730 10740 -670
rect 10800 -730 10810 -670
rect 10240 -764 10330 -730
rect 10238 -770 10330 -764
rect 10238 -830 10250 -770
rect 10310 -830 10330 -770
rect 10580 -830 10590 -770
rect 10650 -830 10660 -770
rect 10238 -836 10330 -830
rect 10240 -840 10330 -836
rect 10390 -930 10400 -870
rect 10460 -930 10470 -870
rect 10600 -930 10630 -830
rect 3780 -1770 3800 -940
rect 10339 -986 10399 -976
rect 10447 -986 10507 -976
rect 10740 -1000 10780 -730
rect 10660 -1030 10780 -1000
rect 10339 -1056 10355 -1046
rect 10447 -1056 10507 -1046
rect 10490 -1180 10550 -1090
rect 10480 -1240 10490 -1180
rect 10550 -1240 10560 -1180
rect 10490 -1340 10550 -1240
rect 10339 -1386 10399 -1376
rect 10447 -1386 10507 -1376
rect 10740 -1400 10780 -1030
rect 10840 -990 10870 70
rect 10940 -160 10970 1790
rect 11030 870 11060 1900
rect 11010 810 11020 870
rect 11080 810 11090 870
rect 11020 520 11080 530
rect 11020 450 11080 460
rect 11030 250 11060 450
rect 11010 190 11020 250
rect 11080 190 11090 250
rect 10900 -220 10910 -160
rect 10970 -220 10980 -160
rect 10900 -340 10910 -280
rect 10970 -340 10980 -280
rect 10840 -1050 10850 -990
rect 10910 -1050 10920 -990
rect 10950 -1380 10980 -340
rect 11030 -400 11060 190
rect 11010 -460 11020 -400
rect 11080 -460 11090 -400
rect 11120 -580 11150 2430
rect 11190 2340 11200 2400
rect 11260 2340 11270 2400
rect 11200 430 11230 2340
rect 11270 2087 11280 2147
rect 11340 2087 11350 2147
rect 11290 740 11320 2087
rect 11630 1720 11700 2810
rect 11620 1650 11630 1720
rect 11700 1650 11710 1720
rect 11450 1540 11460 1600
rect 11520 1540 11530 1600
rect 11360 1370 11420 1380
rect 11360 1300 11420 1310
rect 11270 680 11280 740
rect 11340 680 11350 740
rect 11180 370 11190 430
rect 11250 370 11260 430
rect 11080 -640 11090 -580
rect 11150 -640 11160 -580
rect 11010 -910 11020 -850
rect 11080 -910 11090 -850
rect 10660 -1430 10780 -1400
rect 10920 -1440 10930 -1380
rect 10990 -1440 11000 -1380
rect 10339 -1456 10355 -1446
rect 10447 -1456 10507 -1446
rect 11030 -1490 11060 -910
rect 10380 -1560 10390 -1500
rect 10450 -1560 10460 -1500
rect 10600 -1630 10630 -1500
rect 11010 -1550 11020 -1490
rect 11080 -1550 11090 -1490
rect 11120 -1630 11150 -640
rect 11200 -760 11230 370
rect 11180 -820 11190 -760
rect 11250 -820 11260 -760
rect 11290 -1190 11320 680
rect 11380 40 11410 1300
rect 11470 520 11500 1540
rect 11540 1490 11600 1500
rect 11540 1420 11600 1430
rect 11440 460 11450 520
rect 11510 460 11520 520
rect 11550 140 11580 1420
rect 11630 630 11700 1650
rect 11620 560 11630 630
rect 11700 560 11710 630
rect 11530 130 11580 140
rect 11500 70 11510 130
rect 11570 70 11580 130
rect 11360 30 11420 40
rect 11360 -40 11420 -30
rect 11550 -860 11580 70
rect 11630 -670 11700 560
rect 11690 -730 11700 -670
rect 11630 -780 11700 -730
rect 11510 -920 11520 -860
rect 11580 -920 11590 -860
rect 11270 -1250 11280 -1190
rect 11340 -1250 11350 -1190
rect 10570 -1690 10580 -1630
rect 10640 -1690 10650 -1630
rect 11070 -1690 11080 -1630
rect 11140 -1690 11150 -1630
rect 3700 -1830 3800 -1770
rect 3890 -1780 6890 -1720
rect 6950 -1780 10030 -1720
rect 3700 -1840 10140 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1890 10140 -1840
rect 3700 -1900 10140 -1890
<< via1 >>
rect 6890 2690 6950 2750
rect 6890 560 6950 620
rect 6890 360 6950 420
rect 9740 70 9800 130
rect 10520 2562 10580 2570
rect 10520 2512 10577 2562
rect 10577 2512 10580 2562
rect 10520 2510 10580 2512
rect 10680 2566 10750 2580
rect 10680 2512 10747 2566
rect 10747 2512 10750 2566
rect 10680 2510 10750 2512
rect 11010 2520 11070 2580
rect 10260 2410 10280 2470
rect 10280 2410 10320 2470
rect 10590 2350 10600 2400
rect 10600 2350 10650 2400
rect 10590 2340 10650 2350
rect 10280 2127 10340 2137
rect 10280 2077 10330 2127
rect 10330 2077 10340 2127
rect 11110 2430 11170 2490
rect 10510 1954 10570 1960
rect 10510 1904 10511 1954
rect 10511 1904 10570 1954
rect 10510 1900 10570 1904
rect 10680 1954 10750 1960
rect 10680 1900 10747 1954
rect 10747 1900 10750 1954
rect 10680 1890 10750 1900
rect 11010 1900 11070 1960
rect 10520 1838 10580 1850
rect 10520 1790 10580 1838
rect 10930 1790 10990 1850
rect 10760 1650 10830 1720
rect 10280 1520 10340 1580
rect 10620 1570 10629 1600
rect 10629 1570 10663 1600
rect 10663 1570 10680 1600
rect 10620 1540 10680 1570
rect 10500 1340 10563 1406
rect 10550 1230 10610 1290
rect 10800 1240 10860 1300
rect 10360 1009 10420 1020
rect 10360 961 10420 1009
rect 10630 1025 10700 1030
rect 10630 977 10634 1025
rect 10634 977 10699 1025
rect 10699 977 10700 1025
rect 10630 970 10700 977
rect 10360 960 10420 961
rect 10550 864 10610 870
rect 10550 816 10554 864
rect 10554 816 10610 864
rect 10550 810 10610 816
rect 10270 680 10330 740
rect 10690 560 10760 630
rect 10580 380 10640 440
rect 10380 180 10450 250
rect 10328 72 10388 132
rect 10436 72 10496 132
rect 10280 -40 10340 20
rect 10120 -130 10130 -70
rect 10130 -130 10170 -70
rect 10170 -130 10180 -70
rect 9740 -520 9800 -460
rect 10830 70 10890 130
rect 10740 -130 10800 -70
rect 10480 -230 10540 -170
rect 10328 -340 10388 -280
rect 10436 -340 10496 -280
rect 10380 -460 10450 -390
rect 10570 -640 10630 -580
rect 10260 -730 10320 -670
rect 10740 -730 10800 -670
rect 10590 -830 10650 -770
rect 10400 -930 10460 -870
rect 10339 -1046 10399 -986
rect 10447 -1046 10507 -986
rect 10490 -1240 10550 -1180
rect 10339 -1446 10399 -1386
rect 10447 -1446 10507 -1386
rect 11020 810 11080 870
rect 11020 460 11080 520
rect 11020 190 11080 250
rect 10910 -220 10970 -160
rect 10910 -340 10970 -280
rect 10850 -1050 10910 -990
rect 11020 -460 11080 -400
rect 11200 2340 11260 2400
rect 11280 2087 11340 2147
rect 11630 1650 11700 1720
rect 11460 1540 11520 1600
rect 11360 1310 11420 1370
rect 11280 680 11340 740
rect 11190 370 11250 430
rect 11090 -640 11150 -580
rect 11020 -910 11080 -850
rect 10930 -1440 10990 -1380
rect 10390 -1560 10450 -1500
rect 11020 -1550 11080 -1490
rect 11190 -820 11250 -760
rect 11540 1430 11600 1490
rect 11450 460 11510 520
rect 11630 560 11700 630
rect 11510 70 11570 130
rect 11360 -30 11420 30
rect 11630 -730 11690 -670
rect 11520 -920 11580 -860
rect 11280 -1250 11340 -1190
rect 10580 -1690 10640 -1630
rect 11080 -1690 11140 -1630
rect 6890 -1780 6950 -1720
<< metal2 >>
rect 6890 2750 6950 2760
rect 6890 620 6950 2690
rect 10540 2625 11750 2655
rect 10540 2580 10570 2625
rect 10680 2580 10750 2590
rect 10520 2570 10580 2580
rect 10520 2500 10580 2510
rect 11010 2580 11070 2590
rect 10750 2530 11010 2560
rect 11070 2530 11750 2560
rect 11010 2510 11070 2520
rect 10680 2500 10750 2510
rect 11110 2490 11170 2500
rect 10260 2470 10320 2480
rect 10320 2440 11110 2470
rect 11110 2420 11170 2430
rect 10260 2400 10320 2410
rect 10590 2400 10650 2410
rect 11200 2400 11260 2410
rect 10650 2360 11200 2390
rect 10590 2330 10650 2340
rect 11200 2330 11260 2340
rect 11280 2147 11340 2157
rect 10280 2137 10340 2147
rect 10340 2087 11280 2117
rect 11280 2077 11340 2087
rect 10280 2067 10340 2077
rect 10530 2010 11750 2040
rect 10530 1970 10560 2010
rect 10510 1960 10570 1970
rect 10510 1890 10570 1900
rect 10680 1960 10750 1970
rect 11010 1960 11070 1970
rect 10750 1900 11010 1930
rect 11010 1890 11070 1900
rect 10680 1880 10750 1890
rect 10520 1850 10580 1860
rect 10930 1850 10990 1860
rect 10580 1810 10930 1840
rect 10520 1780 10580 1790
rect 10930 1780 10990 1790
rect 10760 1720 10830 1730
rect 11630 1720 11700 1730
rect 10830 1650 11630 1720
rect 10760 1640 10830 1650
rect 11630 1640 11700 1650
rect 10620 1600 10680 1610
rect 10280 1580 10340 1590
rect 11460 1600 11520 1610
rect 10680 1550 11460 1580
rect 10620 1530 10680 1540
rect 11460 1530 11520 1540
rect 10280 1510 10340 1520
rect 10290 1480 10320 1510
rect 11540 1490 11600 1500
rect 10290 1450 11540 1480
rect 11540 1420 11600 1430
rect 10500 1406 10563 1416
rect 10563 1370 10580 1380
rect 11360 1370 11420 1380
rect 10563 1340 11360 1370
rect 10500 1330 10563 1340
rect 10800 1300 10860 1310
rect 11360 1300 11420 1310
rect 10550 1290 10610 1300
rect 10800 1230 10860 1240
rect 10550 1220 10610 1230
rect 10360 1020 10420 1030
rect 10560 1020 10590 1220
rect 10420 980 10590 1020
rect 10630 1030 10700 1040
rect 10810 1020 10850 1230
rect 10700 980 10850 1020
rect 10630 960 10700 970
rect 10360 950 10420 960
rect 10550 870 10610 880
rect 11020 870 11080 880
rect 10610 820 11020 850
rect 10550 800 10610 810
rect 11020 800 11080 810
rect 10270 740 10330 750
rect 11280 740 11340 750
rect 10330 680 11280 720
rect 10270 670 10330 680
rect 11280 670 11340 680
rect 3610 560 6890 600
rect 10690 630 10760 640
rect 11630 630 11700 640
rect 6950 560 7610 600
rect 6890 550 6950 560
rect 6890 420 6950 430
rect 6890 -290 6950 360
rect 7570 120 7610 560
rect 10760 560 11630 630
rect 10690 550 10760 560
rect 11630 550 11700 560
rect 11020 520 11080 530
rect 11450 520 11510 530
rect 11080 470 11450 500
rect 11020 450 11080 460
rect 11450 450 11510 460
rect 10580 440 10640 450
rect 11190 430 11250 440
rect 10640 390 11190 420
rect 10580 370 10640 380
rect 11190 360 11250 370
rect 10380 250 10450 260
rect 11020 250 11080 260
rect 10450 200 11020 240
rect 11020 180 11080 190
rect 10380 170 10450 180
rect 9740 130 9800 140
rect 7570 80 9740 120
rect 10328 132 10388 142
rect 9800 80 10328 120
rect 9740 60 9800 70
rect 10328 62 10388 72
rect 10436 132 10496 142
rect 10830 130 10890 140
rect 10496 80 10830 120
rect 10436 62 10496 72
rect 10830 60 10890 70
rect 11510 130 11570 140
rect 11510 60 11570 70
rect 11360 30 11420 40
rect 10280 20 10340 30
rect 10340 -20 11360 10
rect 11420 -20 11750 10
rect 11360 -40 11420 -30
rect 10280 -50 10340 -40
rect 10120 -70 10180 -60
rect 10740 -70 10800 -60
rect 10180 -120 10740 -80
rect 10120 -140 10180 -130
rect 10740 -140 10800 -130
rect 10910 -160 10970 -150
rect 10480 -170 10540 -160
rect 10540 -210 10910 -180
rect 10910 -230 10970 -220
rect 10480 -240 10540 -230
rect 10328 -280 10388 -270
rect 3610 -330 10328 -290
rect 6890 -1720 6950 -330
rect 9600 -1400 9640 -330
rect 10328 -350 10388 -340
rect 10436 -280 10496 -270
rect 10910 -280 10970 -270
rect 10496 -330 10910 -300
rect 10436 -350 10496 -340
rect 10910 -350 10970 -340
rect 10380 -390 10450 -380
rect 9740 -460 9800 -450
rect 11020 -400 11080 -390
rect 10450 -450 11020 -410
rect 10380 -470 10450 -460
rect 11020 -470 11080 -460
rect 9740 -530 9800 -520
rect 9750 -1000 9790 -530
rect 10570 -580 10630 -570
rect 11090 -580 11150 -570
rect 10630 -630 11090 -600
rect 10570 -650 10630 -640
rect 11090 -650 11150 -640
rect 10260 -670 10320 -660
rect 10740 -670 10800 -660
rect 10320 -720 10740 -680
rect 10260 -740 10320 -730
rect 11630 -670 11690 -660
rect 10800 -720 11630 -680
rect 10740 -740 10800 -730
rect 11630 -740 11690 -730
rect 11190 -760 11250 -750
rect 10590 -770 10650 -760
rect 10650 -810 11190 -780
rect 11190 -830 11250 -820
rect 10590 -840 10650 -830
rect 11020 -850 11080 -840
rect 10400 -870 10460 -860
rect 10460 -900 11020 -870
rect 11520 -860 11580 -850
rect 11080 -900 11520 -870
rect 11020 -920 11080 -910
rect 11520 -930 11580 -920
rect 10400 -940 10460 -930
rect 10339 -986 10399 -976
rect 9750 -1040 10339 -1000
rect 10339 -1056 10399 -1046
rect 10447 -986 10507 -976
rect 10850 -990 10910 -980
rect 10507 -1030 10850 -1000
rect 10447 -1056 10507 -1046
rect 10850 -1060 10910 -1050
rect 10490 -1180 10550 -1170
rect 11280 -1190 11340 -1180
rect 10550 -1230 11280 -1200
rect 10490 -1250 10550 -1240
rect 11280 -1260 11340 -1250
rect 10339 -1386 10399 -1376
rect 9600 -1440 10339 -1400
rect 10339 -1456 10399 -1446
rect 10447 -1386 10507 -1376
rect 10930 -1380 10990 -1370
rect 10507 -1430 10930 -1390
rect 10447 -1456 10507 -1446
rect 10930 -1450 10990 -1440
rect 11020 -1490 11080 -1480
rect 10390 -1500 10450 -1490
rect 10450 -1550 11020 -1530
rect 10450 -1560 11080 -1550
rect 10390 -1570 10450 -1560
rect 10580 -1630 10640 -1620
rect 11080 -1630 11140 -1620
rect 10640 -1670 11080 -1640
rect 10580 -1700 10640 -1690
rect 11080 -1700 11140 -1690
rect 6890 -1790 6950 -1780
use sky130_fd_pr__pfet_01v8_lvt_B59788  sky130_fd_pr__pfet_01v8_lvt_B59788_0
timestamp 1711994487
transform 1 0 6954 0 1 -681
box -3254 -1219 3254 1219
use sky130_fd_pr__pfet_01v8_M4CK9Z  sky130_fd_pr__pfet_01v8_M4CK9Z_0
timestamp 1711995413
transform 1 0 10461 0 -1 -313
box -359 -261 359 261
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10766 0 -1 2777
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1710522493
transform -1 0 10766 0 1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10490 0 -1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1710522493
transform -1 0 10490 0 -1 2777
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1710522493
transform -1 0 10490 0 1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1710522493
transform 1 0 10214 0 1 601
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1710522493
transform 1 0 10490 0 1 601
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10858 0 -1 1689
box -38 -48 406 592
use sky130_fd_pr__pfet_01v8_lvt_B59788  XM24
timestamp 1711994487
transform 1 0 6954 0 1 1651
box -3254 -1219 3254 1219
use sky130_fd_pr__nfet_01v8_75Z3GH  XM27
timestamp 1711995063
transform 1 0 10521 0 1 -1416
box -311 -252 311 252
use sky130_fd_pr__pfet_01v8_M4CK9Z  XM29
timestamp 1711995413
transform 1 0 10461 0 1 103
box -359 -261 359 261
use sky130_fd_pr__nfet_01v8_75Z3GH  XM37
timestamp 1711995063
transform 1 0 10521 0 -1 -1018
box -311 -252 311 252
<< labels >>
flabel metal1 11030 305 11060 335 0 FreeSans 80 0 0 0 LOAD_CAL_Z
flabel metal1 10940 300 10970 330 0 FreeSans 80 0 0 0 EN_COMP_Z
flabel metal1 11120 310 11150 340 0 FreeSans 80 0 0 0 CAL_RESULTi
flabel metal1 11200 480 11230 510 0 FreeSans 80 0 0 0 CAL_RESULT_Z
flabel metal1 11290 460 11320 490 0 FreeSans 80 0 0 0 EN_COMPi
rlabel metal2 3610 -330 3650 -290 1 CAL_P
port 3 n
rlabel metal2 3610 560 3650 600 1 CAL_N
port 4 n
rlabel metal1 9980 2820 10140 2880 1 VDD
port 0 n
rlabel metal1 10280 2820 10440 2880 1 VSS
port 6 n
rlabel metal2 11720 2530 11750 2560 1 CAL_CYCLE
port 7 n
rlabel metal2 11720 2625 11750 2655 1 CAL_RESULT
port 1 n
rlabel metal2 11715 2010 11745 2040 1 EN_COMP
port 2 n
rlabel metal2 11715 -20 11745 10 1 EN
port 5 n
<< end >>
