* NGSPICE file created from state_machine.ext - technology: sky130A

.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_ef_sc_hd__decap_12.spice

* pin order for ef_sc_hd_decap_12 cell is different in the openlane generated netlist vs magic generated netlist, modified openlane generated netlist manually to match

.subckt state_machine VDD VSS clk clk_data comp_p data[0] data[1] data[2] data[3]
+ data[4] data[5] en_comp en_offset_cal en_offset_cal_o en_vcm_sw_o en_vcm_sw_o_i
+ offset_cal_cycle rst_z sample_o single_ended start vcm_dummy_o vcm_o[0] vcm_o[10]
+ vcm_o[1] vcm_o[2] vcm_o[3] vcm_o[4] vcm_o[5] vcm_o[6] vcm_o[7] vcm_o[8] vcm_o[9]
+ vcm_o_i[0] vcm_o_i[10] vcm_o_i[1] vcm_o_i[2] vcm_o_i[3] vcm_o_i[4] vcm_o_i[5] vcm_o_i[6]
+ vcm_o_i[7] vcm_o_i[8] vcm_o_i[9] vin_n_sw_on vin_p_sw_on vref_z_n_o[0] vref_z_n_o[10]
+ vref_z_n_o[1] vref_z_n_o[2] vref_z_n_o[3] vref_z_n_o[4] vref_z_n_o[5] vref_z_n_o[6]
+ vref_z_n_o[7] vref_z_n_o[8] vref_z_n_o[9] vref_z_p_o[0] vref_z_p_o[10] vref_z_p_o[1]
+ vref_z_p_o[2] vref_z_p_o[3] vref_z_p_o[4] vref_z_p_o[5] vref_z_p_o[6] vref_z_p_o[7]
+ vref_z_p_o[8] vref_z_p_o[9] vss_n_o[0] vss_n_o[10] vss_n_o[1] vss_n_o[2] vss_n_o[3]
+ vss_n_o[4] vss_n_o[5] vss_n_o[6] vss_n_o[7] vss_n_o[8] vss_n_o[9] vss_p_o[0] vss_p_o[10]
+ vss_p_o[1] vss_p_o[2] vss_p_o[3] vss_p_o[4] vss_p_o[5] vss_p_o[6] vss_p_o[7] vss_p_o[8]
+ vss_p_o[9]
XFILLER_0_2_7 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_294_ counter\[9\] _103_ VSS VSS VDD VDD net42 sky130_fd_sc_hd__nor2_1
X_363_ _026_ net107 net117 VSS VSS VDD VDD _020_ sky130_fd_sc_hd__o21a_1
Xfanout105 state\[1\] VSS VSS VDD VDD net105 sky130_fd_sc_hd__buf_2
XFILLER_0_9_274 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_346_ net1 _137_ _136_ VSS VSS VDD VDD _007_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_66 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_277_ _099_ _085_ VSS VSS VDD VDD net62 sky130_fd_sc_hd__nand2b_1
X_200_ net99 net11 net110 VSS VSS VDD VDD _059_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_4_82 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_329_ net1 _124_ _123_ VSS VSS VDD VDD _003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_228 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_114 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput20 net20 VSS VSS VDD VDD clk_data sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 VSS VSS VDD VDD vref_z_n_o[8] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VSS VSS VDD VDD vref_z_p_o[8] sky130_fd_sc_hd__buf_2
Xoutput42 net42 VSS VSS VDD VDD vcm_o[8] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VSS VSS VDD VDD sample_o sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_35 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput86 net86 VSS VSS VDD VDD vss_p_o[8] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VSS VSS VDD VDD vss_n_o[8] sky130_fd_sc_hd__buf_2
X_293_ counter\[8\] _103_ VSS VSS VDD VDD net41 sky130_fd_sc_hd__nor2_1
X_362_ net107 net92 _141_ net116 VSS VSS VDD VDD _019_ sky130_fd_sc_hd__a22o_1
Xfanout106 state\[0\] VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_253 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_9_242 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_67 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ result\[3\] net91 VSS VSS VDD VDD _137_ sky130_fd_sc_hd__and2_1
X_276_ result\[7\] result\[6\] net97 VSS VSS VDD VDD _099_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Left_14 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_328_ result\[9\] _104_ VSS VSS VDD VDD _124_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_19 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_259_ net103 net107 net32 _069_ VSS VSS VDD VDD _091_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_6_Right_6 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput54 net54 VSS VSS VDD VDD vref_z_n_o[9] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VSS VSS VDD VDD data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 VSS VSS VDD VDD vref_z_p_o[9] sky130_fd_sc_hd__buf_2
Xoutput43 net43 VSS VSS VDD VDD vcm_o[9] sky130_fd_sc_hd__buf_2
Xoutput32 net32 VSS VSS VDD VDD vcm_dummy_o sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_36 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 net87 VSS VSS VDD VDD vss_p_o[9] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VSS VSS VDD VDD vss_n_o[9] sky130_fd_sc_hd__buf_2
X_361_ net108 net92 net90 counter\[9\] VSS VSS VDD VDD _018_ sky130_fd_sc_hd__a22o_1
X_292_ counter\[7\] _103_ VSS VSS VDD VDD net40 sky130_fd_sc_hd__nor2_1
XFILLER_0_4_195 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xfanout107 counter\[11\] VSS VSS VDD VDD net107 sky130_fd_sc_hd__buf_2
XFILLER_0_1_198 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_68 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_275_ net100 _035_ _083_ _098_ VSS VSS VDD VDD net61 sky130_fd_sc_hd__o211ai_1
X_344_ _134_ _135_ _051_ VSS VSS VDD VDD _136_ sky130_fd_sc_hd__a21o_1
X_189_ net106 net18 net19 net105 VSS VSS VDD VDD _052_ sky130_fd_sc_hd__or4b_4
X_327_ _121_ _122_ _051_ VSS VSS VDD VDD _123_ sky130_fd_sc_hd__a21o_1
X_258_ result\[10\] _069_ VSS VSS VDD VDD net54 sky130_fd_sc_hd__nand2_1
XFILLER_0_6_19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput22 net22 VSS VSS VDD VDD data[1] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VSS VSS VDD VDD vss_p_o[0] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VSS VSS VDD VDD vcm_o[0] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VSS VSS VDD VDD vss_n_o[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_37 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput44 net44 VSS VSS VDD VDD vref_z_n_o[0] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VSS VSS VDD VDD vref_z_p_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_7_84 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_360_ counter\[9\] net92 net90 counter\[8\] VSS VSS VDD VDD _017_ sky130_fd_sc_hd__a22o_1
X_291_ counter\[6\] _103_ VSS VSS VDD VDD net39 sky130_fd_sc_hd__nor2_1
Xfanout108 counter\[10\] VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_166 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_69 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_274_ net100 result\[5\] VSS VSS VDD VDD _098_ sky130_fd_sc_hd__nand2_1
X_343_ net109 counter\[5\] net98 VSS VSS VDD VDD _135_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_4_85 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_326_ net102 counter\[9\] net108 VSS VSS VDD VDD _122_ sky130_fd_sc_hd__or3b_1
Xfanout90 _141_ VSS VSS VDD VDD net90 sky130_fd_sc_hd__buf_2
X_257_ net53 _090_ VSS VSS VDD VDD net86 sky130_fd_sc_hd__nand2_1
X_188_ net106 state\[1\] VSS VSS VDD VDD _051_ sky130_fd_sc_hd__nand2b_2
X_309_ _034_ _051_ VSS VSS VDD VDD net20 sky130_fd_sc_hd__nor2_1
XFILLER_0_8_139 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput45 net45 VSS VSS VDD VDD vref_z_n_o[10] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VSS VSS VDD VDD data[2] sky130_fd_sc_hd__clkbuf_4
Xoutput56 net56 VSS VSS VDD VDD vref_z_p_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_7_183 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput34 net34 VSS VSS VDD VDD vcm_o[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_38 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 net78 VSS VSS VDD VDD vss_p_o[10] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VSS VSS VDD VDD vss_n_o[10] sky130_fd_sc_hd__buf_2
X_290_ counter\[5\] _103_ VSS VSS VDD VDD net38 sky130_fd_sc_hd__nor2_1
XFILLER_0_9_201 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xfanout109 counter\[4\] VSS VSS VDD VDD net109 sky130_fd_sc_hd__buf_2
X_342_ net98 counter\[3\] net109 VSS VSS VDD VDD _134_ sky130_fd_sc_hd__or3b_1
X_273_ net94 result\[5\] _061_ _081_ _097_ VSS VSS VDD VDD net60 sky130_fd_sc_hd__a221o_1
XFILLER_0_5_270 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xfanout91 _104_ VSS VSS VDD VDD net91 sky130_fd_sc_hd__clkbuf_2
X_187_ state\[0\] net105 VSS VSS VDD VDD _050_ sky130_fd_sc_hd__and2b_1
X_256_ net108 _037_ _052_ net95 VSS VSS VDD VDD _090_ sky130_fd_sc_hd__a211o_1
X_325_ net108 net107 net102 VSS VSS VDD VDD _121_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_8_Left_18 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_239_ _052_ _080_ VSS VSS VDD VDD _081_ sky130_fd_sc_hd__or2_1
X_308_ _051_ _112_ _105_ net115 VSS VSS VDD VDD _156_ sky130_fd_sc_hd__a2bb2o_1
Xoutput24 net24 VSS VSS VDD VDD data[3] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 VSS VSS VDD VDD vref_z_n_o[1] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VSS VSS VDD VDD vcm_o[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_39 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput57 net57 VSS VSS VDD VDD vref_z_p_o[1] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VSS VSS VDD VDD vss_p_o[1] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VSS VSS VDD VDD vss_n_o[1] sky130_fd_sc_hd__buf_2
X_341_ _133_ _117_ _132_ VSS VSS VDD VDD _006_ sky130_fd_sc_hd__mux2_1
X_272_ net94 _040_ VSS VSS VDD VDD _097_ sky130_fd_sc_hd__nor2_1
X_324_ _117_ result\[10\] _120_ VSS VSS VDD VDD _002_ sky130_fd_sc_hd__mux2_1
X_186_ _033_ result\[5\] _049_ VSS VSS VDD VDD net26 sky130_fd_sc_hd__o21ai_1
Xfanout92 net93 VSS VSS VDD VDD net92 sky130_fd_sc_hd__buf_2
X_255_ net102 net108 net32 _068_ VSS VSS VDD VDD _089_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_9_70 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_238_ net99 counter\[6\] VSS VSS VDD VDD _080_ sky130_fd_sc_hd__nand2_1
X_307_ _107_ _109_ _110_ _111_ VSS VSS VDD VDD _112_ sky130_fd_sc_hd__and4_1
X_169_ result\[3\] VSS VSS VDD VDD _038_ sky130_fd_sc_hd__inv_2
Xoutput25 net25 VSS VSS VDD VDD data[4] sky130_fd_sc_hd__clkbuf_4
Xoutput36 net36 VSS VSS VDD VDD vcm_o[2] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VSS VSS VDD VDD vss_n_o[2] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VSS VSS VDD VDD vref_z_n_o[2] sky130_fd_sc_hd__buf_2
Xoutput58 net58 VSS VSS VDD VDD vref_z_p_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_7_54 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_340_ result\[7\] net91 VSS VSS VDD VDD _133_ sky130_fd_sc_hd__and2_1
X_271_ _078_ _096_ VSS VSS VDD VDD net59 sky130_fd_sc_hd__nand2_1
X_323_ _026_ _118_ _119_ _115_ VSS VSS VDD VDD _120_ sky130_fd_sc_hd__a31o_1
Xfanout93 _050_ VSS VSS VDD VDD net93 sky130_fd_sc_hd__buf_2
X_185_ net100 net110 result\[11\] VSS VSS VDD VDD _049_ sky130_fd_sc_hd__or3_1
X_254_ result\[9\] _068_ VSS VSS VDD VDD net53 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_71 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_168_ result\[8\] VSS VSS VDD VDD _037_ sky130_fd_sc_hd__inv_2
X_306_ counter\[7\] counter\[3\] counter\[2\] net109 VSS VSS VDD VDD _111_ sky130_fd_sc_hd__and4_1
X_237_ result\[5\] _060_ VSS VSS VDD VDD net49 sky130_fd_sc_hd__nand2_1
Xoutput26 net26 VSS VSS VDD VDD data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput48 net48 VSS VSS VDD VDD vref_z_n_o[3] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VSS VSS VDD VDD vcm_o[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput59 net59 VSS VSS VDD VDD vref_z_p_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_1_104 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_40 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_237 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_270_ _038_ _040_ net94 VSS VSS VDD VDD _096_ sky130_fd_sc_hd__mux2_1
X_399_ clknet_2_2__leaf_clk _018_ net113 VSS VSS VDD VDD counter\[9\] sky130_fd_sc_hd__dfrtp_4
X_322_ net107 net103 VSS VSS VDD VDD _119_ sky130_fd_sc_hd__nand2b_1
X_184_ _048_ VSS VSS VDD VDD net25 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_72 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout94 _027_ VSS VSS VDD VDD net94 sky130_fd_sc_hd__clkbuf_4
X_253_ net52 _088_ VSS VSS VDD VDD net85 sky130_fd_sc_hd__nand2_1
X_236_ net48 _079_ VSS VSS VDD VDD net81 sky130_fd_sc_hd__nand2_1
X_305_ counter\[6\] counter\[5\] counter\[1\] VSS VSS VDD VDD _110_ sky130_fd_sc_hd__and3_1
X_167_ result\[1\] VSS VSS VDD VDD _036_ sky130_fd_sc_hd__inv_2
X_219_ result\[11\] net8 _070_ VSS VSS VDD VDD _071_ sky130_fd_sc_hd__or3b_1
Xoutput49 net49 VSS VSS VDD VDD vref_z_n_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_7_154 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_132 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_110 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xoutput38 net38 VSS VSS VDD VDD vcm_o[4] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VSS VSS VDD VDD en_comp sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_clk clk VSS VSS VDD VDD clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_157 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_34 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_41 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_398_ clknet_2_2__leaf_clk _017_ net113 VSS VSS VDD VDD counter\[8\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_9_73 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_252_ _029_ result\[7\] net89 net101 VSS VSS VDD VDD _088_ sky130_fd_sc_hd__o211ai_1
X_183_ result\[10\] result\[4\] net110 VSS VSS VDD VDD _048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_20 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout95 _027_ VSS VSS VDD VDD net95 sky130_fd_sc_hd__dlymetal6s2s_1
X_321_ net103 net108 net107 VSS VSS VDD VDD _118_ sky130_fd_sc_hd__or3b_1
X_304_ net103 counter\[0\] VSS VSS VDD VDD _109_ sky130_fd_sc_hd__xor2_1
X_235_ counter\[5\] _038_ _052_ net94 VSS VSS VDD VDD _079_ sky130_fd_sc_hd__a211o_1
X_166_ result\[6\] VSS VSS VDD VDD _035_ sky130_fd_sc_hd__inv_2
X_218_ net103 net107 VSS VSS VDD VDD _070_ sky130_fd_sc_hd__and2b_1
Xoutput39 net39 VSS VSS VDD VDD vcm_o[5] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VSS VSS VDD VDD en_offset_cal_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_79 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_169 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_180 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_42 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_250 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_397_ clknet_2_2__leaf_clk _016_ net113 VSS VSS VDD VDD counter\[7\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_2_0__f_clk clknet_0_clk VSS VSS VDD VDD clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_182_ _047_ VSS VSS VDD VDD net24 sky130_fd_sc_hd__inv_2
X_251_ net101 counter\[9\] net89 _066_ VSS VSS VDD VDD _087_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_21 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 net98 VSS VSS VDD VDD net96 sky130_fd_sc_hd__clkbuf_2
X_320_ net94 _028_ net92 _117_ _116_ VSS VSS VDD VDD _001_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_9_74 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_13 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_234_ net98 counter\[5\] net88 _059_ VSS VSS VDD VDD _078_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_48 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_303_ net104 counter\[0\] VSS VSS VDD VDD _108_ sky130_fd_sc_hd__nor2_1
X_165_ counter\[5\] VSS VSS VDD VDD _034_ sky130_fd_sc_hd__inv_2
X_217_ net103 net89 _069_ _041_ VSS VSS VDD VDD net76 sky130_fd_sc_hd__a22o_1
XFILLER_0_7_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput29 net29 VSS VSS VDD VDD en_vcm_sw_o sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_43 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_195 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_396_ clknet_2_1__leaf_clk _015_ net111 VSS VSS VDD VDD counter\[6\] sky130_fd_sc_hd__dfrtp_4
X_181_ result\[9\] result\[3\] net109 VSS VSS VDD VDD _047_ sky130_fd_sc_hd__mux2_1
Xfanout97 net98 VSS VSS VDD VDD net97 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_22 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ result\[8\] _066_ VSS VSS VDD VDD net52 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_75 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_379_ counter\[2\] counter\[3\] net97 VSS VSS VDD VDD _153_ sky130_fd_sc_hd__nand3b_1
X_164_ net110 VSS VSS VDD VDD _033_ sky130_fd_sc_hd__inv_2
X_233_ result\[4\] _059_ VSS VSS VDD VDD net48 sky130_fd_sc_hd__nand2_1
X_302_ net107 net108 counter\[9\] counter\[8\] VSS VSS VDD VDD _107_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_113 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_216_ net103 net17 net108 VSS VSS VDD VDD _069_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_4_138 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_44 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_174__1 clknet_2_2__leaf_clk VSS VSS VDD VDD net114 sky130_fd_sc_hd__inv_2
X_395_ clknet_2_1__leaf_clk _014_ net111 VSS VSS VDD VDD counter\[5\] sky130_fd_sc_hd__dfrtp_4
X_180_ _046_ VSS VSS VDD VDD net23 sky130_fd_sc_hd__inv_2
Xfanout98 single_ended_reg VSS VSS VDD VDD net98 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_76 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_23 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ net96 counter\[1\] counter\[2\] VSS VSS VDD VDD _152_ sky130_fd_sc_hd__or3b_1
X_301_ net6 _106_ _000_ VSS VSS VDD VDD _155_ sky130_fd_sc_hd__a21o_1
X_232_ net47 _077_ VSS VSS VDD VDD net80 sky130_fd_sc_hd__nand2_1
X_163_ counter\[2\] VSS VSS VDD VDD _032_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_70 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_215_ net103 net89 _068_ _039_ VSS VSS VDD VDD net75 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_55 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_82 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_175 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_220 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_81 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_394_ clknet_2_0__leaf_clk _013_ net111 VSS VSS VDD VDD counter\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_201 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_256 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_77 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ net1 _151_ _150_ VSS VSS VDD VDD _024_ sky130_fd_sc_hd__mux2_1
Xfanout88 net89 VSS VSS VDD VDD net88 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_24 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 single_ended_reg VSS VSS VDD VDD net99 sky130_fd_sc_hd__buf_2
X_231_ _033_ result\[2\] net88 net98 VSS VSS VDD VDD _077_ sky130_fd_sc_hd__o211ai_1
X_300_ net106 net105 VSS VSS VDD VDD _106_ sky130_fd_sc_hd__nor2_1
X_162_ counter\[7\] VSS VSS VDD VDD _031_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_82 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xinput1 comp_p VSS VSS VDD VDD net1 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_56 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ net102 net16 counter\[9\] VSS VSS VDD VDD _068_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_7_137 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_110 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_243 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_393_ clknet_2_0__leaf_clk _012_ net111 VSS VSS VDD VDD counter\[3\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_9_78 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 net32 VSS VSS VDD VDD net89 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_25 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ result\[6\] net91 VSS VSS VDD VDD _151_ sky130_fd_sc_hd__and2_1
X_161_ counter\[8\] VSS VSS VDD VDD _030_ sky130_fd_sc_hd__inv_2
X_230_ net98 net109 net88 _058_ VSS VSS VDD VDD _076_ sky130_fd_sc_hd__a31o_1
X_359_ counter\[8\] net92 net90 counter\[7\] VSS VSS VDD VDD _016_ sky130_fd_sc_hd__a22o_1
Xinput2 en_offset_cal VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_57 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ net101 counter\[9\] VSS VSS VDD VDD _067_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_130 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_155 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_392_ clknet_2_0__leaf_clk _011_ net111 VSS VSS VDD VDD counter\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_0_26 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_79 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ counter\[6\] _051_ _063_ _149_ counter\[7\] VSS VSS VDD VDD _150_ sky130_fd_sc_hd__o32a_1
X_358_ counter\[7\] net93 net90 counter\[6\] VSS VSS VDD VDD _015_ sky130_fd_sc_hd__a22o_1
X_160_ counter\[9\] VSS VSS VDD VDD _029_ sky130_fd_sc_hd__inv_2
X_289_ net110 _103_ VSS VSS VDD VDD net37 sky130_fd_sc_hd__nor2_1
Xinput3 en_vcm_sw_o_i VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_58 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ net102 net89 _066_ _037_ VSS VSS VDD VDD net74 sky130_fd_sc_hd__a22o_1
XFILLER_0_2_63 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_189 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_391_ clknet_2_2__leaf_clk _010_ net112 VSS VSS VDD VDD counter\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_0_27 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ net106 net105 net101 counter\[8\] VSS VSS VDD VDD _149_ sky130_fd_sc_hd__nand4b_1
Xinput4 rst_z VSS VSS VDD VDD net4 sky130_fd_sc_hd__buf_1
X_357_ counter\[6\] net93 net90 counter\[5\] VSS VSS VDD VDD _014_ sky130_fd_sc_hd__a22o_1
X_288_ counter\[3\] _103_ VSS VSS VDD VDD net36 sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1__f_clk clknet_0_clk VSS VSS VDD VDD clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_6_59 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ net101 net15 counter\[8\] VSS VSS VDD VDD _066_ sky130_fd_sc_hd__nor3b_1
X_409_ clknet_2_0__leaf_clk _025_ net111 VSS VSS VDD VDD result\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_151 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_110 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_176 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_390_ clknet_2_2__leaf_clk _009_ net112 VSS VSS VDD VDD counter\[0\] sky130_fd_sc_hd__dfrtp_1
X_373_ net103 net5 _106_ VSS VSS VDD VDD _023_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_28 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_274 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_31 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_42 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
Xinput5 single_ended VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkbuf_1
X_287_ counter\[2\] _103_ VSS VSS VDD VDD net35 sky130_fd_sc_hd__nor2_1
X_356_ net109 net90 net20 VSS VSS VDD VDD _013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_193 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_408_ clknet_2_1__leaf_clk _024_ net4 VSS VSS VDD VDD result\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_119 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_210_ net100 counter\[8\] VSS VSS VDD VDD _065_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_141 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_339_ _031_ net92 _065_ _131_ _030_ VSS VSS VDD VDD _132_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_166 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_188 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_169 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_29 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _117_ result\[2\] _148_ VSS VSS VDD VDD _022_ sky130_fd_sc_hd__mux2_1
X_355_ net109 net93 net90 counter\[3\] VSS VSS VDD VDD _012_ sky130_fd_sc_hd__a22o_1
X_286_ counter\[1\] _103_ VSS VSS VDD VDD net33 sky130_fd_sc_hd__nor2_1
Xinput6 start VSS VSS VDD VDD net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_12 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_407_ clknet_2_3__leaf_clk _023_ net113 VSS VSS VDD VDD single_ended_reg sky130_fd_sc_hd__dfrtp_1
X_338_ net106 net105 net101 counter\[9\] VSS VSS VDD VDD _131_ sky130_fd_sc_hd__and4b_1
XFILLER_0_2_88 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_269_ net96 _038_ _076_ _095_ VSS VSS VDD VDD net58 sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_7_60 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_371_ net93 _146_ _147_ _115_ VSS VSS VDD VDD _148_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_210 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_22 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_77 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_285_ net94 net88 VSS VSS VDD VDD _103_ sky130_fd_sc_hd__nand2_4
X_354_ counter\[3\] net93 net90 counter\[2\] VSS VSS VDD VDD _011_ sky130_fd_sc_hd__a22o_1
Xinput7 vcm_o_i[0] VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkbuf_1
X_337_ net1 _130_ _129_ VSS VSS VDD VDD _005_ sky130_fd_sc_hd__mux2_1
X_268_ net97 result\[2\] VSS VSS VDD VDD _095_ sky130_fd_sc_hd__nand2_1
X_199_ net98 net88 _058_ _038_ VSS VSS VDD VDD net69 sky130_fd_sc_hd__a22o_1
X_406_ clknet_2_0__leaf_clk _022_ net111 VSS VSS VDD VDD result\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_7_61 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 vcm_o_i[2] VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_146 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_370_ counter\[3\] net109 net96 VSS VSS VDD VDD _147_ sky130_fd_sc_hd__nand3b_1
X_353_ counter\[1\] net90 _138_ VSS VSS VDD VDD _010_ sky130_fd_sc_hd__a21o_1
X_284_ net99 result\[10\] _053_ _071_ VSS VSS VDD VDD net56 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_30 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 vcm_o_i[10] VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkbuf_1
X_405_ clknet_2_1__leaf_clk _021_ net4 VSS VSS VDD VDD result\[5\] sky130_fd_sc_hd__dfrtp_2
X_336_ result\[4\] net91 VSS VSS VDD VDD _130_ sky130_fd_sc_hd__and2_1
X_198_ net98 net10 counter\[3\] VSS VSS VDD VDD _058_ sky130_fd_sc_hd__nor3b_1
X_267_ net94 result\[2\] _057_ _074_ _094_ VSS VSS VDD VDD net57 sky130_fd_sc_hd__a221o_1
X_319_ net1 net91 VSS VSS VDD VDD _117_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_62 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 vcm_o_i[3] VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_117 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_0_90 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_352_ counter\[1\] net93 net90 net118 VSS VSS VDD VDD _009_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_31 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 vcm_o_i[1] VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkbuf_1
X_283_ _091_ _102_ VSS VSS VDD VDD net65 sky130_fd_sc_hd__nand2_1
XFILLER_0_9_175 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_197_ result\[2\] _057_ _053_ VSS VSS VDD VDD net68 sky130_fd_sc_hd__o21ai_2
X_266_ net94 _036_ VSS VSS VDD VDD _094_ sky130_fd_sc_hd__nor2_1
X_404_ clknet_2_2__leaf_clk _156_ net112 VSS VSS VDD VDD state\[1\] sky130_fd_sc_hd__dfrtp_1
X_335_ net99 counter\[5\] _080_ _128_ _051_ VSS VSS VDD VDD _129_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_2_58 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_318_ _051_ _070_ net91 result\[11\] VSS VSS VDD VDD _116_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_7_63 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 vcm_o_i[4] VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkbuf_1
X_249_ net51 _086_ VSS VSS VDD VDD net84 sky130_fd_sc_hd__nand2_1
XFILLER_0_2_170 VSS VDD VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_8_207 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_276 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xhold1 counter_sample VSS VSS VDD VDD net115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_14 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_32 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_282_ _039_ _041_ net95 VSS VSS VDD VDD _102_ sky130_fd_sc_hd__mux2_1
X_351_ net106 net105 VSS VSS VDD VDD _141_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_165 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_403_ clknet_2_3__leaf_clk _155_ net112 VSS VSS VDD VDD state\[0\] sky130_fd_sc_hd__dfrtp_1
X_334_ net110 counter\[5\] VSS VSS VDD VDD _128_ sky130_fd_sc_hd__nand2b_1
X_196_ net96 _032_ net9 VSS VSS VDD VDD _057_ sky130_fd_sc_hd__or3_1
X_265_ net94 result\[1\] _054_ _055_ _093_ VSS VSS VDD VDD net55 sky130_fd_sc_hd__a221o_1
X_179_ result\[8\] result\[2\] net110 VSS VSS VDD VDD _046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_64 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 vcm_o_i[5] VSS VSS VDD VDD net13 sky130_fd_sc_hd__clkbuf_1
X_317_ net92 _114_ _105_ VSS VSS VDD VDD net29 sky130_fd_sc_hd__a21o_1
X_248_ counter\[8\] _035_ _052_ net95 VSS VSS VDD VDD _086_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_182 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk VSS VSS VDD VDD clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold2 counter\[10\] VSS VSS VDD VDD net116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_33 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _140_ net1 _139_ VSS VSS VDD VDD _008_ sky130_fd_sc_hd__mux2_1
X_281_ _089_ _101_ VSS VSS VDD VDD net64 sky130_fd_sc_hd__nand2_1
XFILLER_0_9_111 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_402_ clknet_2_3__leaf_clk _000_ net112 VSS VSS VDD VDD counter_sample sky130_fd_sc_hd__dfrtp_1
X_333_ _127_ net1 _126_ VSS VSS VDD VDD _004_ sky130_fd_sc_hd__mux2_1
X_195_ net96 _032_ net9 VSS VSS VDD VDD _056_ sky130_fd_sc_hd__nor3_1
X_264_ net96 result\[0\] VSS VSS VDD VDD _093_ sky130_fd_sc_hd__and2_1
X_316_ net106 net105 VSS VSS VDD VDD _115_ sky130_fd_sc_hd__xnor2_2
Xinput14 vcm_o_i[6] VSS VSS VDD VDD net14 sky130_fd_sc_hd__clkbuf_1
X_247_ net100 counter\[8\] net89 _064_ VSS VSS VDD VDD _085_ sky130_fd_sc_hd__a31o_1
X_178_ _045_ VSS VSS VDD VDD net22 sky130_fd_sc_hd__inv_2
XFILLER_0_8_15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
Xhold3 state\[1\] VSS VSS VDD VDD net117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_34 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_280_ _037_ _039_ net95 VSS VSS VDD VDD _101_ sky130_fd_sc_hd__mux2_1
X_332_ result\[8\] net91 VSS VSS VDD VDD _127_ sky130_fd_sc_hd__and2_1
X_401_ clknet_2_3__leaf_clk _020_ net112 VSS VSS VDD VDD counter\[11\] sky130_fd_sc_hd__dfrtp_1
X_194_ result\[1\] _055_ _053_ VSS VSS VDD VDD net66 sky130_fd_sc_hd__o21ai_2
X_263_ _041_ _053_ net45 VSS VSS VDD VDD net78 sky130_fd_sc_hd__o21ai_1
X_177_ result\[7\] result\[1\] net109 VSS VSS VDD VDD _045_ sky130_fd_sc_hd__mux2_1
Xinput15 vcm_o_i[7] VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkbuf_1
X_315_ net2 _114_ VSS VSS VDD VDD net30 sky130_fd_sc_hd__and2_1
X_246_ result\[7\] _064_ VSS VSS VDD VDD net51 sky130_fd_sc_hd__nand2_1
X_229_ result\[3\] _058_ VSS VSS VDD VDD net47 sky130_fd_sc_hd__nand2_1
Xhold4 counter\[0\] VSS VSS VDD VDD net118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_45 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_83 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_271 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_146 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_331_ _030_ net92 _067_ _125_ _029_ VSS VSS VDD VDD _126_ sky130_fd_sc_hd__a32o_1
X_193_ net96 net7 counter\[1\] VSS VSS VDD VDD _055_ sky130_fd_sc_hd__or3b_1
X_400_ clknet_2_2__leaf_clk _019_ net112 VSS VSS VDD VDD counter\[10\] sky130_fd_sc_hd__dfrtp_1
X_262_ net103 _028_ net8 result\[11\] VSS VSS VDD VDD net45 sky130_fd_sc_hd__or4b_1
XFILLER_0_6_138 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_160 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_176_ _044_ VSS VSS VDD VDD net21 sky130_fd_sc_hd__inv_2
Xinput16 vcm_o_i[8] VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkbuf_1
X_314_ net2 _108_ _113_ net114 net92 VSS VSS VDD VDD net27 sky130_fd_sc_hd__o311a_2
X_245_ net50 _084_ VSS VSS VDD VDD net83 sky130_fd_sc_hd__nand2_1
X_159_ counter\[11\] VSS VSS VDD VDD _028_ sky130_fd_sc_hd__inv_2
X_228_ result\[2\] _056_ _075_ VSS VSS VDD VDD net79 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_46 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_9_125 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_9_103 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_330_ net106 net105 net101 net108 VSS VSS VDD VDD _125_ sky130_fd_sc_hd__and4b_1
XFILLER_0_6_83 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_192_ net94 _032_ _052_ VSS VSS VDD VDD _054_ sky130_fd_sc_hd__or3_1
X_261_ net54 _092_ VSS VSS VDD VDD net87 sky130_fd_sc_hd__nand2_1
XFILLER_0_5_172 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_175_ result\[6\] result\[0\] net109 VSS VSS VDD VDD _044_ sky130_fd_sc_hd__mux2_1
Xinput17 vcm_o_i[9] VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_1_Left_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_244_ _031_ result\[5\] net89 net100 VSS VSS VDD VDD _084_ sky130_fd_sc_hd__o211ai_1
X_313_ _108_ _113_ VSS VSS VDD VDD _114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_164 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_227_ result\[1\] _073_ net88 net96 VSS VSS VDD VDD _075_ sky130_fd_sc_hd__o211a_1
X_158_ net97 VSS VSS VDD VDD _027_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_47 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_226 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_94 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_260_ net107 _039_ _052_ net95 VSS VSS VDD VDD _092_ sky130_fd_sc_hd__a211o_1
X_389_ clknet_2_0__leaf_clk _008_ net111 VSS VSS VDD VDD result\[0\] sky130_fd_sc_hd__dfrtp_1
X_191_ net98 net88 VSS VSS VDD VDD _053_ sky130_fd_sc_hd__nand2_2
Xinput18 vin_n_sw_on VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkbuf_1
X_243_ net100 counter\[7\] net89 _062_ VSS VSS VDD VDD _083_ sky130_fd_sc_hd__a31o_1
X_312_ counter\[1\] net104 VSS VSS VDD VDD _113_ sky130_fd_sc_hd__and2b_1
X_157_ net106 VSS VSS VDD VDD _026_ sky130_fd_sc_hd__inv_2
X_226_ _052_ _073_ VSS VSS VDD VDD _074_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_268 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_48 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ result\[7\] net14 _063_ _053_ VSS VSS VDD VDD net73 sky130_fd_sc_hd__o31ai_1
XFILLER_0_6_96 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_190_ _052_ VSS VSS VDD VDD net32 sky130_fd_sc_hd__inv_2
X_388_ clknet_2_0__leaf_clk _007_ net111 VSS VSS VDD VDD result\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_119 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xinput19 vin_p_sw_on VSS VSS VDD VDD net19 sky130_fd_sc_hd__buf_1
X_242_ result\[6\] _062_ VSS VSS VDD VDD net50 sky130_fd_sc_hd__nand2_1
X_311_ net112 net2 VSS VSS VDD VDD net28 sky130_fd_sc_hd__and2_1
X_173_ net3 VSS VSS VDD VDD _042_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_86 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_225_ net96 counter\[3\] VSS VSS VDD VDD _073_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_49 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ net101 net14 counter\[7\] VSS VSS VDD VDD _064_ sky130_fd_sc_hd__nor3b_1
Xclkbuf_2_3__f_clk clknet_0_clk VSS VSS VDD VDD clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_139 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_387_ clknet_2_3__leaf_clk _006_ net113 VSS VSS VDD VDD result\[7\] sky130_fd_sc_hd__dfrtp_2
X_310_ net105 _042_ _106_ net107 VSS VSS VDD VDD net31 sky130_fd_sc_hd__a211oi_2
X_241_ result\[5\] _060_ _082_ VSS VSS VDD VDD net82 sky130_fd_sc_hd__a21o_1
X_172_ result\[10\] VSS VSS VDD VDD _041_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_156 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3_54 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_224_ result\[2\] _056_ VSS VSS VDD VDD net46 sky130_fd_sc_hd__nand2_1
X_207_ net101 counter\[7\] VSS VSS VDD VDD _063_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_20 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_0_55 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_386_ clknet_2_1__leaf_clk _005_ net111 VSS VSS VDD VDD result\[4\] sky130_fd_sc_hd__dfrtp_1
X_171_ result\[4\] VSS VSS VDD VDD _040_ sky130_fd_sc_hd__inv_2
X_240_ result\[4\] _080_ net89 net99 VSS VSS VDD VDD _082_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_135 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_11 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_369_ net97 counter\[2\] counter\[3\] VSS VSS VDD VDD _146_ sky130_fd_sc_hd__or3b_1
Xfanout110 counter\[4\] VSS VSS VDD VDD net110 sky130_fd_sc_hd__clkbuf_2
X_223_ net44 _072_ VSS VSS VDD VDD net77 sky130_fd_sc_hd__nand2_1
X_206_ net99 net88 _062_ _035_ VSS VSS VDD VDD net72 sky130_fd_sc_hd__a22o_1
XFILLER_0_3_252 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_274 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_50 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_119 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_385_ clknet_2_3__leaf_clk _004_ net113 VSS VSS VDD VDD result\[8\] sky130_fd_sc_hd__dfrtp_1
Xoutput80 net80 VSS VSS VDD VDD vss_p_o[2] sky130_fd_sc_hd__buf_2
X_170_ result\[9\] VSS VSS VDD VDD _039_ sky130_fd_sc_hd__inv_2
X_368_ net1 _145_ _144_ VSS VSS VDD VDD _021_ sky130_fd_sc_hd__mux2_1
X_299_ net115 _104_ VSS VSS VDD VDD _000_ sky130_fd_sc_hd__nor2_1
Xfanout111 net4 VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkbuf_4
Xfanout100 single_ended_reg VSS VSS VDD VDD net100 sky130_fd_sc_hd__clkbuf_2
X_222_ _032_ result\[0\] net88 net96 VSS VSS VDD VDD _072_ sky130_fd_sc_hd__o211ai_1
X_205_ net100 net13 counter\[6\] VSS VSS VDD VDD _062_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_9_44 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_242 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_51 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_384_ clknet_2_3__leaf_clk _003_ net113 VSS VSS VDD VDD result\[9\] sky130_fd_sc_hd__dfrtp_1
Xoutput81 net81 VSS VSS VDD VDD vss_p_o[3] sky130_fd_sc_hd__buf_2
Xoutput70 net70 VSS VSS VDD VDD vss_n_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_2_148 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_298_ _104_ VSS VSS VDD VDD _105_ sky130_fd_sc_hd__inv_2
X_367_ result\[5\] net91 VSS VSS VDD VDD _145_ sky130_fd_sc_hd__and2_1
Xfanout112 net113 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkbuf_4
Xfanout101 net104 VSS VSS VDD VDD net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_35 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_221_ _036_ _055_ VSS VSS VDD VDD net44 sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_9_Left_19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_6_273 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_204_ result\[5\] _061_ _053_ VSS VSS VDD VDD net71 sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_257 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_52 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_383_ clknet_2_3__leaf_clk _002_ net112 VSS VSS VDD VDD result\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_7 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput82 net82 VSS VSS VDD VDD vss_p_o[4] sky130_fd_sc_hd__buf_2
Xoutput71 net71 VSS VSS VDD VDD vss_n_o[4] sky130_fd_sc_hd__buf_2
Xoutput60 net60 VSS VSS VDD VDD vref_z_p_o[4] sky130_fd_sc_hd__buf_2
X_297_ state\[1\] state\[0\] VSS VSS VDD VDD _104_ sky130_fd_sc_hd__nand2b_1
X_366_ _142_ _143_ _051_ VSS VSS VDD VDD _144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_190 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xfanout113 net4 VSS VSS VDD VDD net113 sky130_fd_sc_hd__buf_2
Xfanout102 net104 VSS VSS VDD VDD net102 sky130_fd_sc_hd__clkbuf_2
X_220_ _053_ _071_ VSS VSS VDD VDD net67 sky130_fd_sc_hd__nand2_1
X_349_ result\[0\] net91 VSS VSS VDD VDD _140_ sky130_fd_sc_hd__and2_1
X_203_ net99 _034_ net12 VSS VSS VDD VDD _061_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_24 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_53 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput61 net61 VSS VSS VDD VDD vref_z_p_o[5] sky130_fd_sc_hd__buf_2
Xoutput50 net50 VSS VSS VDD VDD vref_z_n_o[5] sky130_fd_sc_hd__buf_2
X_382_ clknet_2_3__leaf_clk _001_ net112 VSS VSS VDD VDD result\[11\] sky130_fd_sc_hd__dfrtp_1
Xoutput83 net83 VSS VSS VDD VDD vss_p_o[5] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VSS VSS VDD VDD vss_n_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_5_103 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_296_ counter\[11\] _103_ VSS VSS VDD VDD net34 sky130_fd_sc_hd__nor2_1
X_365_ net100 counter\[5\] counter\[6\] VSS VSS VDD VDD _143_ sky130_fd_sc_hd__or3b_1
Xfanout103 net104 VSS VSS VDD VDD net103 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_0_Left_10 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_279_ net102 _037_ _087_ _100_ VSS VSS VDD VDD net63 sky130_fd_sc_hd__o211ai_2
X_348_ counter\[1\] net92 _108_ _113_ _138_ VSS VSS VDD VDD _139_ sky130_fd_sc_hd__a32o_1
X_202_ net99 _034_ net12 VSS VSS VDD VDD _060_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_5_54 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput51 net51 VSS VSS VDD VDD vref_z_n_o[6] sky130_fd_sc_hd__buf_2
X_381_ _117_ result\[1\] _154_ VSS VSS VDD VDD _025_ sky130_fd_sc_hd__mux2_1
Xoutput40 net40 VSS VSS VDD VDD vcm_o[6] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VSS VSS VDD VDD vss_p_o[6] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VSS VSS VDD VDD vss_n_o[6] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VSS VSS VDD VDD vref_z_p_o[6] sky130_fd_sc_hd__buf_2
X_295_ net108 _103_ VSS VSS VDD VDD net43 sky130_fd_sc_hd__nor2_1
X_364_ counter\[6\] counter\[7\] net99 VSS VSS VDD VDD _142_ sky130_fd_sc_hd__nand3b_1
Xfanout104 single_ended_reg VSS VSS VDD VDD net104 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_8_65 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_278_ net101 result\[7\] VSS VSS VDD VDD _100_ sky130_fd_sc_hd__nand2_1
X_347_ net106 net105 counter\[2\] VSS VSS VDD VDD _138_ sky130_fd_sc_hd__and3b_1
X_201_ net99 net88 _059_ _040_ VSS VSS VDD VDD net70 sky130_fd_sc_hd__a22o_1
XFILLER_0_4_70 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput52 net52 VSS VSS VDD VDD vref_z_n_o[7] sky130_fd_sc_hd__buf_2
Xoutput41 net41 VSS VSS VDD VDD vcm_o[7] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VSS VSS VDD VDD offset_cal_cycle sky130_fd_sc_hd__buf_2
X_380_ net91 _152_ _153_ _115_ VSS VSS VDD VDD _154_ sky130_fd_sc_hd__a31o_1
Xoutput63 net63 VSS VSS VDD VDD vref_z_p_o[7] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VSS VSS VDD VDD vss_p_o[7] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VSS VSS VDD VDD vss_n_o[7] sky130_fd_sc_hd__buf_2
.ends

