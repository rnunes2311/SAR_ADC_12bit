magic
tech sky130A
magscale 1 2
timestamp 1711310191
<< metal3 >>
rect -886 1441 886 1469
rect -886 -1441 802 1441
rect 866 -1441 886 1441
rect -886 -1469 886 -1441
<< via3 >>
rect 802 -1441 866 1441
<< mimcap >>
rect -846 1389 554 1429
rect -846 -1389 -806 1389
rect 514 -1389 554 1389
rect -846 -1429 554 -1389
<< mimcapcontact >>
rect -806 -1389 514 1389
<< metal4 >>
rect 786 1441 882 1457
rect -807 1389 515 1390
rect -807 -1389 -806 1389
rect 514 -1389 515 1389
rect -807 -1390 515 -1389
rect 786 -1441 802 1441
rect 866 -1441 882 1441
rect 786 -1457 882 -1441
<< properties >>
string FIXED_BBOX -886 -1469 594 1469
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7 l 14.29 val 208.15 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
