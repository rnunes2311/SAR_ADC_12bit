magic
tech sky130A
magscale 1 2
timestamp 1715418002
<< nwell >>
rect 6802 -170 6990 -136
rect 6802 -252 7236 -170
<< pwell >>
rect 6560 -430 6620 -350
<< nsubdiff >>
rect 5560 323 5896 416
rect 6522 327 6858 420
<< locali >>
rect 5540 1070 7820 1100
rect 5540 1010 5600 1070
rect 7730 1010 7820 1070
rect 5540 940 7820 1010
rect 7090 610 7200 660
rect 5560 323 5896 416
rect 6522 327 6858 420
rect 7075 131 7291 181
rect 5540 -1030 5580 -290
rect 5890 -1020 6520 -810
rect 6850 -1020 6880 -290
rect 5540 -1520 5740 -1030
rect 6700 -1520 6880 -1020
rect 5540 -1630 7820 -1520
rect 5540 -1690 5600 -1630
rect 7730 -1690 7820 -1630
rect 5540 -1740 7820 -1690
<< viali >>
rect 5600 1010 7730 1070
rect 6959 611 7022 658
rect 7560 600 7620 660
rect 6958 133 7024 181
rect 7560 130 7620 190
rect 7240 -490 7300 -430
rect 7540 -477 7607 -429
rect 5600 -1690 7730 -1630
<< metal1 >>
rect 5540 1070 7820 1100
rect 5540 1010 5600 1070
rect 7730 1010 7820 1070
rect 5540 990 5650 1010
rect 5710 990 5900 1010
rect 5970 990 6040 1010
rect 6110 990 6320 1010
rect 6390 990 6450 1010
rect 6520 990 6710 1010
rect 6770 990 7320 1010
rect 7380 990 7420 1010
rect 7480 990 7820 1010
rect 5540 940 7820 990
rect 5560 810 5770 850
rect 5880 815 6075 845
rect 6355 815 6540 845
rect 5560 520 5600 810
rect 5640 680 5650 740
rect 5710 680 5720 740
rect 5775 565 5850 595
rect 5560 480 5770 520
rect 5560 250 5600 480
rect 5820 410 5850 565
rect 5770 350 5780 410
rect 5840 350 5850 410
rect 5560 210 5770 250
rect 5560 -80 5600 210
rect 5640 70 5650 130
rect 5710 70 5720 130
rect 5560 -120 5770 -80
rect 5560 -390 5600 -120
rect 5800 -350 5830 20
rect 5880 -85 5910 815
rect 5960 680 5970 740
rect 6030 680 6040 740
rect 6380 680 6390 740
rect 6450 680 6460 740
rect 5960 580 5970 640
rect 6030 580 6040 640
rect 6380 580 6390 640
rect 6450 580 6460 640
rect 5960 490 5970 550
rect 6030 490 6040 550
rect 6380 490 6390 550
rect 6450 490 6460 550
rect 6060 350 6070 410
rect 6130 350 6140 410
rect 6280 350 6290 410
rect 6350 350 6360 410
rect 6095 85 6180 115
rect 6150 -70 6180 85
rect 6240 85 6325 115
rect 5880 -115 6055 -85
rect 5880 -180 5910 -115
rect 6120 -130 6130 -70
rect 6190 -130 6200 -70
rect 5860 -240 5870 -180
rect 5930 -240 5940 -180
rect 5800 -360 5860 -350
rect 5560 -430 5750 -390
rect 5800 -430 5860 -420
rect 5900 -395 5930 -240
rect 5900 -425 6075 -395
rect 5560 -900 5590 -430
rect 5630 -540 5640 -480
rect 5700 -540 5710 -480
rect 5630 -700 5640 -640
rect 5700 -700 5710 -640
rect 5900 -705 5930 -425
rect 6150 -530 6180 -130
rect 6240 -180 6270 85
rect 6510 -70 6540 815
rect 6660 810 6860 850
rect 6700 680 6710 740
rect 6770 680 6780 740
rect 6570 565 6645 595
rect 6570 410 6600 565
rect 6820 530 6860 810
rect 6950 664 6960 670
rect 6947 658 6960 664
rect 7020 664 7030 670
rect 7020 658 7034 664
rect 6947 611 6959 658
rect 7022 611 7034 658
rect 6947 610 6960 611
rect 7020 610 7034 611
rect 6947 605 7034 610
rect 7548 660 7632 666
rect 7548 600 7560 660
rect 7620 600 7632 660
rect 7548 594 7632 600
rect 6660 490 6870 530
rect 6570 350 6580 410
rect 6640 350 6650 410
rect 6820 250 6860 490
rect 7540 340 7820 460
rect 6660 210 6870 250
rect 6700 70 6710 130
rect 6770 70 6780 130
rect 6480 -85 6490 -70
rect 6355 -115 6490 -85
rect 6480 -130 6490 -115
rect 6550 -130 6560 -70
rect 6220 -240 6230 -180
rect 6290 -240 6300 -180
rect 6100 -560 6180 -530
rect 6240 -530 6270 -240
rect 6490 -390 6520 -130
rect 6590 -350 6620 20
rect 6820 -80 6860 210
rect 7548 190 7632 196
rect 6950 187 6960 190
rect 6946 181 6960 187
rect 7020 187 7030 190
rect 7020 181 7036 187
rect 6946 133 6958 181
rect 7024 133 7036 181
rect 6946 130 6960 133
rect 7020 130 7036 133
rect 6946 127 7036 130
rect 7548 130 7560 190
rect 7620 130 7632 190
rect 7548 124 7632 130
rect 6650 -120 6860 -80
rect 6340 -430 6520 -390
rect 6560 -360 6620 -350
rect 6820 -380 6860 -120
rect 7310 -180 7320 -120
rect 7380 -180 7390 -120
rect 7410 -180 7420 -120
rect 7480 -180 7490 -120
rect 6650 -420 6860 -380
rect 6560 -430 6620 -420
rect 6240 -560 6320 -530
rect 5960 -590 6020 -580
rect 6020 -650 6030 -590
rect 6380 -650 6390 -590
rect 6450 -650 6460 -590
rect 5960 -660 6020 -650
rect 6490 -700 6520 -430
rect 6690 -540 6700 -480
rect 6760 -540 6770 -480
rect 6690 -700 6700 -640
rect 6760 -700 6770 -640
rect 5900 -735 6065 -705
rect 5900 -740 5930 -735
rect 6340 -740 6520 -700
rect 5770 -810 5780 -750
rect 5840 -810 5850 -750
rect 6580 -810 6590 -750
rect 6650 -810 6660 -750
rect 6820 -900 6854 -420
rect 7220 -424 7310 -420
rect 7220 -430 7312 -424
rect 7220 -490 7240 -430
rect 7300 -490 7312 -430
rect 7528 -429 7619 -423
rect 7528 -477 7540 -429
rect 7607 -430 7619 -429
rect 7528 -483 7550 -477
rect 7540 -490 7550 -483
rect 7610 -490 7620 -430
rect 7220 -496 7312 -490
rect 7220 -500 7310 -496
rect 7700 -640 7820 340
rect 7080 -740 7160 -660
rect 7540 -760 7820 -640
rect 7220 -900 7230 -880
rect 5560 -940 7230 -900
rect 7290 -940 7300 -880
rect 5630 -1040 5640 -980
rect 5700 -1040 5710 -980
rect 5630 -1520 5710 -1040
rect 5770 -1050 5780 -990
rect 5840 -1050 5850 -990
rect 5950 -1050 5960 -990
rect 6020 -1025 6030 -990
rect 6020 -1050 6040 -1025
rect 6380 -1050 6390 -990
rect 6450 -1050 6460 -990
rect 6580 -1050 6590 -990
rect 6650 -1050 6660 -990
rect 6690 -1040 6700 -980
rect 6760 -1040 6770 -980
rect 5820 -1240 5850 -1050
rect 6010 -1220 6040 -1050
rect 6070 -1140 6080 -1080
rect 6140 -1140 6150 -1080
rect 6390 -1220 6420 -1050
rect 6500 -1174 6560 -1100
rect 6590 -1174 6620 -1050
rect 6466 -1180 6620 -1174
rect 6500 -1202 6560 -1180
rect 6590 -1240 6620 -1180
rect 5860 -1370 5870 -1310
rect 5930 -1370 5940 -1310
rect 6180 -1370 6190 -1310
rect 6250 -1370 6260 -1310
rect 5870 -1460 5930 -1370
rect 6490 -1376 6500 -1316
rect 6560 -1376 6570 -1316
rect 6280 -1470 6290 -1410
rect 6350 -1470 6360 -1410
rect 6690 -1520 6770 -1040
rect 7700 -1520 7820 -760
rect 5540 -1630 7820 -1520
rect 5540 -1690 5600 -1630
rect 7730 -1690 7820 -1630
rect 5540 -1740 7820 -1690
<< via1 >>
rect 5650 1010 5710 1050
rect 5900 1010 5970 1050
rect 6040 1010 6110 1050
rect 6320 1010 6390 1050
rect 6450 1010 6520 1050
rect 6710 1010 6770 1050
rect 7320 1010 7380 1050
rect 7420 1010 7480 1050
rect 5650 990 5710 1010
rect 5900 990 5970 1010
rect 6040 990 6110 1010
rect 6320 990 6390 1010
rect 6450 990 6520 1010
rect 6710 990 6770 1010
rect 7320 990 7380 1010
rect 7420 990 7480 1010
rect 5650 680 5710 740
rect 5780 350 5840 410
rect 5650 70 5710 130
rect 5970 680 6030 740
rect 6390 680 6450 740
rect 5970 580 6030 640
rect 6390 580 6450 640
rect 5970 490 6030 550
rect 6390 490 6450 550
rect 6070 350 6130 410
rect 6290 350 6350 410
rect 6130 -130 6190 -70
rect 5870 -240 5930 -180
rect 5800 -420 5860 -360
rect 5640 -540 5700 -480
rect 5640 -700 5700 -640
rect 6710 680 6770 740
rect 6960 658 7020 670
rect 6960 611 7020 658
rect 6960 610 7020 611
rect 7560 600 7620 660
rect 6580 350 6640 410
rect 6710 70 6770 130
rect 6490 -130 6550 -70
rect 6230 -240 6290 -180
rect 6960 181 7020 190
rect 6960 133 7020 181
rect 6960 130 7020 133
rect 7560 130 7620 190
rect 6560 -420 6620 -360
rect 7320 -180 7380 -120
rect 7420 -180 7480 -120
rect 5960 -650 6020 -590
rect 6390 -650 6450 -590
rect 6700 -540 6760 -480
rect 6700 -700 6760 -640
rect 5780 -810 5840 -750
rect 6590 -810 6650 -750
rect 7240 -490 7300 -430
rect 7550 -477 7607 -430
rect 7607 -477 7610 -430
rect 7550 -490 7610 -477
rect 7230 -940 7290 -880
rect 5640 -1040 5700 -980
rect 5780 -1050 5840 -990
rect 5960 -1050 6020 -990
rect 6390 -1050 6450 -990
rect 6590 -1050 6650 -990
rect 6700 -1040 6760 -980
rect 6080 -1140 6140 -1080
rect 5870 -1370 5930 -1310
rect 6190 -1370 6250 -1310
rect 6500 -1376 6560 -1316
rect 6290 -1470 6350 -1410
<< metal2 >>
rect 5650 1050 5710 1060
rect 5650 740 5710 990
rect 5900 1050 6520 1060
rect 5970 990 6040 1050
rect 6110 990 6320 1050
rect 6390 990 6450 1050
rect 5900 980 6520 990
rect 6710 1050 6770 1060
rect 5650 130 5710 680
rect 5970 740 6040 980
rect 6030 680 6040 740
rect 5970 640 6040 680
rect 6030 580 6040 640
rect 5970 550 6040 580
rect 6030 490 6040 550
rect 5970 480 6040 490
rect 6390 740 6450 980
rect 6390 640 6450 680
rect 6390 550 6450 580
rect 6390 480 6450 490
rect 6710 740 6770 990
rect 7320 1050 7480 1060
rect 7380 990 7420 1050
rect 5780 410 5840 420
rect 6070 410 6130 420
rect 5840 360 6070 400
rect 5780 340 5840 350
rect 6070 340 6130 350
rect 6290 410 6350 420
rect 6580 410 6640 420
rect 6350 360 6580 400
rect 6290 340 6350 350
rect 6580 340 6640 350
rect 5650 60 5710 70
rect 6710 130 6770 680
rect 6960 670 7020 680
rect 7020 615 7115 645
rect 6960 600 7020 610
rect 6960 190 7020 200
rect 6960 120 7020 130
rect 6710 60 6770 70
rect 6130 -70 6190 -60
rect 6490 -70 6550 -60
rect 6190 -120 6490 -90
rect 6130 -140 6190 -130
rect 6975 -90 7005 120
rect 6550 -120 7005 -90
rect 6490 -140 6550 -130
rect 5870 -180 5930 -170
rect 6230 -180 6290 -170
rect 5930 -230 6230 -200
rect 5870 -250 5930 -240
rect 7085 -200 7115 615
rect 7320 -120 7480 990
rect 7560 660 7620 670
rect 7620 610 7860 650
rect 7560 590 7620 600
rect 7560 190 7620 200
rect 7620 140 7860 180
rect 7560 120 7620 130
rect 7380 -180 7420 -120
rect 7320 -190 7480 -180
rect 6290 -230 7115 -200
rect 6230 -250 6290 -240
rect 5800 -360 5860 -350
rect 6560 -360 6620 -350
rect 5860 -415 6000 -385
rect 5800 -430 5860 -420
rect 5640 -480 5700 -470
rect 5640 -640 5700 -540
rect 5970 -580 6000 -415
rect 6415 -420 6560 -390
rect 6415 -580 6445 -420
rect 6560 -430 6620 -420
rect 7240 -430 7300 -420
rect 6700 -480 6760 -470
rect 5960 -590 6020 -580
rect 5960 -660 6020 -650
rect 6390 -590 6450 -580
rect 6390 -660 6450 -650
rect 6700 -640 6760 -540
rect 5640 -980 5700 -700
rect 5780 -750 5840 -740
rect 5780 -820 5840 -810
rect 5790 -980 5820 -820
rect 5970 -980 6010 -660
rect 6400 -980 6440 -660
rect 6590 -750 6650 -740
rect 6590 -820 6650 -810
rect 6610 -980 6640 -820
rect 6700 -980 6760 -700
rect 7240 -500 7300 -490
rect 7550 -430 7610 -420
rect 7610 -480 7860 -440
rect 7550 -500 7610 -490
rect 7240 -870 7280 -500
rect 7230 -880 7290 -870
rect 7230 -950 7290 -940
rect 5640 -1050 5700 -1040
rect 5780 -990 5840 -980
rect 5780 -1060 5840 -1050
rect 5960 -990 6020 -980
rect 5960 -1060 6020 -1050
rect 6390 -990 6450 -980
rect 6390 -1060 6450 -1050
rect 6590 -990 6650 -980
rect 6700 -1050 6760 -1040
rect 6590 -1060 6650 -1050
rect 6080 -1080 6140 -1070
rect 5450 -1130 6080 -1090
rect 6080 -1150 6140 -1140
rect 5870 -1310 5930 -1300
rect 6190 -1310 6250 -1300
rect 5930 -1360 6190 -1320
rect 5870 -1380 5930 -1370
rect 6500 -1316 6560 -1306
rect 6250 -1366 6500 -1326
rect 6190 -1380 6250 -1370
rect 6500 -1386 6560 -1376
rect 6290 -1410 6350 -1400
rect 5450 -1460 6290 -1420
rect 6290 -1480 6350 -1470
use sky130_fd_pr__nfet_01v8_7XK7PK  sky130_fd_pr__nfet_01v8_7XK7PK_0
timestamp 1711976318
transform -1 0 6682 0 1 -662
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_0
timestamp 1711974973
transform 1 0 6050 0 1 -562
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KPCVAL  sky130_fd_pr__pfet_01v8_KPCVAL_0
timestamp 1711975452
transform 1 0 6683 0 1 67
box -211 -319 211 319
use sky130_fd_sc_hd__buf_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 7630 0 1 -692
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 6894 0 1 396
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1710522493
transform 1 0 6894 0 -1 396
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7170 0 -1 396
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x7
timestamp 1710522493
transform 1 0 7170 0 1 396
box -38 -48 498 592
use sky130_fd_pr__nfet_01v8_lvt_DTMSLK  XM1
timestamp 1711975147
transform 1 0 6216 0 1 -1276
box -530 -310 530 310
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1711974973
transform 1 0 6366 0 1 -562
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_UNYNRG  XM5
timestamp 1711975388
transform 1 0 5735 0 1 667
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGASDL  XM6
timestamp 1711974973
transform 1 0 6051 0 1 367
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGASDL  XM9
timestamp 1711974973
transform 1 0 6367 0 1 367
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_YRYNRG  XM10
timestamp 1711975601
transform 1 0 5735 0 1 67
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XG57AL  XM11
timestamp 1711975388
transform 1 0 6683 0 1 667
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_7XK7PK  XM18
timestamp 1711976318
transform 1 0 5734 0 1 -662
box -211 -410 211 410
<< labels >>
rlabel metal2 7820 -480 7860 -440 1 EN
port 3 n
rlabel metal2 5450 -1130 5490 -1090 1 VIN_P
port 1 n
rlabel metal2 5450 -1460 5490 -1420 1 VIN_N
port 2 n
rlabel metal2 7820 140 7860 180 1 OUT_N
port 5 n
rlabel metal2 7820 610 7860 650 1 OUT_P
port 4 n
rlabel locali 5570 970 5830 1080 1 VDD
port 0 n
rlabel metal1 5580 -1710 5840 -1600 1 VSS
port 6 n
<< end >>
