magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< nwell >>
rect -246 -2855 246 2855
<< pmos >>
rect -50 1036 50 2636
rect -50 -800 50 800
rect -50 -2636 50 -1036
<< pdiff >>
rect -108 2624 -50 2636
rect -108 1048 -96 2624
rect -62 1048 -50 2624
rect -108 1036 -50 1048
rect 50 2624 108 2636
rect 50 1048 62 2624
rect 96 1048 108 2624
rect 50 1036 108 1048
rect -108 788 -50 800
rect -108 -788 -96 788
rect -62 -788 -50 788
rect -108 -800 -50 -788
rect 50 788 108 800
rect 50 -788 62 788
rect 96 -788 108 788
rect 50 -800 108 -788
rect -108 -1048 -50 -1036
rect -108 -2624 -96 -1048
rect -62 -2624 -50 -1048
rect -108 -2636 -50 -2624
rect 50 -1048 108 -1036
rect 50 -2624 62 -1048
rect 96 -2624 108 -1048
rect 50 -2636 108 -2624
<< pdiffc >>
rect -96 1048 -62 2624
rect 62 1048 96 2624
rect -96 -788 -62 788
rect 62 -788 96 788
rect -96 -2624 -62 -1048
rect 62 -2624 96 -1048
<< nsubdiff >>
rect -210 2785 -114 2819
rect 114 2785 210 2819
rect -210 2723 -176 2785
rect 176 2723 210 2785
rect -210 -2785 -176 -2723
rect 176 -2785 210 -2723
rect -210 -2819 -114 -2785
rect 114 -2819 210 -2785
<< nsubdiffcont >>
rect -114 2785 114 2819
rect -210 -2723 -176 2723
rect 176 -2723 210 2723
rect -114 -2819 114 -2785
<< poly >>
rect -50 2717 50 2733
rect -50 2683 -34 2717
rect 34 2683 50 2717
rect -50 2636 50 2683
rect -50 989 50 1036
rect -50 955 -34 989
rect 34 955 50 989
rect -50 939 50 955
rect -50 881 50 897
rect -50 847 -34 881
rect 34 847 50 881
rect -50 800 50 847
rect -50 -847 50 -800
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect -50 -897 50 -881
rect -50 -955 50 -939
rect -50 -989 -34 -955
rect 34 -989 50 -955
rect -50 -1036 50 -989
rect -50 -2683 50 -2636
rect -50 -2717 -34 -2683
rect 34 -2717 50 -2683
rect -50 -2733 50 -2717
<< polycont >>
rect -34 2683 34 2717
rect -34 955 34 989
rect -34 847 34 881
rect -34 -881 34 -847
rect -34 -989 34 -955
rect -34 -2717 34 -2683
<< locali >>
rect -210 2785 -114 2819
rect 114 2785 210 2819
rect -210 2723 -176 2785
rect 176 2723 210 2785
rect -50 2683 -34 2717
rect 34 2683 50 2717
rect -96 2624 -62 2640
rect -96 1032 -62 1048
rect 62 2624 96 2640
rect 62 1032 96 1048
rect -50 955 -34 989
rect 34 955 50 989
rect -50 847 -34 881
rect 34 847 50 881
rect -96 788 -62 804
rect -96 -804 -62 -788
rect 62 788 96 804
rect 62 -804 96 -788
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect -50 -989 -34 -955
rect 34 -989 50 -955
rect -96 -1048 -62 -1032
rect -96 -2640 -62 -2624
rect 62 -1048 96 -1032
rect 62 -2640 96 -2624
rect -50 -2717 -34 -2683
rect 34 -2717 50 -2683
rect -210 -2785 -176 -2723
rect 176 -2785 210 -2723
rect -210 -2819 -114 -2785
rect 114 -2819 210 -2785
<< viali >>
rect -34 2683 34 2717
rect -96 1048 -62 2624
rect 62 1048 96 2624
rect -34 955 34 989
rect -34 847 34 881
rect -96 -788 -62 788
rect 62 -788 96 788
rect -34 -881 34 -847
rect -34 -989 34 -955
rect -96 -2624 -62 -1048
rect 62 -2624 96 -1048
rect -34 -2717 34 -2683
<< metal1 >>
rect -46 2717 46 2723
rect -46 2683 -34 2717
rect 34 2683 46 2717
rect -46 2677 46 2683
rect -102 2624 -56 2636
rect -102 1048 -96 2624
rect -62 1048 -56 2624
rect -102 1036 -56 1048
rect 56 2624 102 2636
rect 56 1048 62 2624
rect 96 1048 102 2624
rect 56 1036 102 1048
rect -46 989 46 995
rect -46 955 -34 989
rect 34 955 46 989
rect -46 949 46 955
rect -46 881 46 887
rect -46 847 -34 881
rect 34 847 46 881
rect -46 841 46 847
rect -102 788 -56 800
rect -102 -788 -96 788
rect -62 -788 -56 788
rect -102 -800 -56 -788
rect 56 788 102 800
rect 56 -788 62 788
rect 96 -788 102 788
rect 56 -800 102 -788
rect -46 -847 46 -841
rect -46 -881 -34 -847
rect 34 -881 46 -847
rect -46 -887 46 -881
rect -46 -955 46 -949
rect -46 -989 -34 -955
rect 34 -989 46 -955
rect -46 -995 46 -989
rect -102 -1048 -56 -1036
rect -102 -2624 -96 -1048
rect -62 -2624 -56 -1048
rect -102 -2636 -56 -2624
rect 56 -1048 102 -1036
rect 56 -2624 62 -1048
rect 96 -2624 102 -1048
rect 56 -2636 102 -2624
rect -46 -2683 46 -2677
rect -46 -2717 -34 -2683
rect 34 -2717 46 -2683
rect -46 -2723 46 -2717
<< properties >>
string FIXED_BBOX -193 -2802 193 2802
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
