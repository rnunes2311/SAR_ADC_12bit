magic
tech sky130A
magscale 1 2
timestamp 1711884628
<< error_p >>
rect -77 262 -19 268
rect 115 262 173 268
rect -77 228 -65 262
rect 115 228 127 262
rect -77 222 -19 228
rect 115 222 173 228
rect -173 -228 -115 -222
rect 19 -228 77 -222
rect -173 -262 -161 -228
rect 19 -262 31 -228
rect -173 -268 -115 -262
rect 19 -268 77 -262
<< pwell >>
rect -359 -400 359 400
<< nmoslvt >>
rect -159 -190 -129 190
rect -63 -190 -33 190
rect 33 -190 63 190
rect 129 -190 159 190
<< ndiff >>
rect -221 178 -159 190
rect -221 -178 -209 178
rect -175 -178 -159 178
rect -221 -190 -159 -178
rect -129 178 -63 190
rect -129 -178 -113 178
rect -79 -178 -63 178
rect -129 -190 -63 -178
rect -33 178 33 190
rect -33 -178 -17 178
rect 17 -178 33 178
rect -33 -190 33 -178
rect 63 178 129 190
rect 63 -178 79 178
rect 113 -178 129 178
rect 63 -190 129 -178
rect 159 178 221 190
rect 159 -178 175 178
rect 209 -178 221 178
rect 159 -190 221 -178
<< ndiffc >>
rect -209 -178 -175 178
rect -113 -178 -79 178
rect -17 -178 17 178
rect 79 -178 113 178
rect 175 -178 209 178
<< psubdiff >>
rect -323 330 -227 364
rect 227 330 323 364
rect -323 -330 -289 330
rect 289 268 323 330
rect 289 -330 323 -268
rect -323 -364 -227 -330
rect 227 -364 323 -330
<< psubdiffcont >>
rect -227 330 227 364
rect 289 -268 323 268
rect -227 -364 227 -330
<< poly >>
rect -81 262 -15 278
rect -81 228 -65 262
rect -31 228 -15 262
rect -159 190 -129 216
rect -81 212 -15 228
rect 111 262 177 278
rect 111 228 127 262
rect 161 228 177 262
rect -63 190 -33 212
rect 33 190 63 216
rect 111 212 177 228
rect 129 190 159 212
rect -159 -212 -129 -190
rect -177 -228 -111 -212
rect -63 -216 -33 -190
rect 33 -212 63 -190
rect -177 -262 -161 -228
rect -127 -262 -111 -228
rect -177 -278 -111 -262
rect 15 -228 81 -212
rect 129 -216 159 -190
rect 15 -262 31 -228
rect 65 -262 81 -228
rect 15 -278 81 -262
<< polycont >>
rect -65 228 -31 262
rect 127 228 161 262
rect -161 -262 -127 -228
rect 31 -262 65 -228
<< locali >>
rect -323 330 -227 364
rect 227 330 323 364
rect -323 -330 -289 330
rect 289 268 323 330
rect -81 228 -65 262
rect -31 228 -15 262
rect 111 228 127 262
rect 161 228 177 262
rect -209 178 -175 194
rect -209 -194 -175 -178
rect -113 178 -79 194
rect -113 -194 -79 -178
rect -17 178 17 194
rect -17 -194 17 -178
rect 79 178 113 194
rect 79 -194 113 -178
rect 175 178 209 194
rect 175 -194 209 -178
rect -177 -262 -161 -228
rect -127 -262 -111 -228
rect 15 -262 31 -228
rect 65 -262 81 -228
rect 289 -330 323 -268
rect -323 -364 -227 -330
rect 227 -364 323 -330
<< viali >>
rect -65 228 -31 262
rect 127 228 161 262
rect -209 -178 -175 178
rect -113 -178 -79 178
rect -17 -178 17 178
rect 79 -178 113 178
rect 175 -178 209 178
rect -161 -262 -127 -228
rect 31 -262 65 -228
<< metal1 >>
rect -77 262 -19 268
rect -77 228 -65 262
rect -31 228 -19 262
rect -77 222 -19 228
rect 115 262 173 268
rect 115 228 127 262
rect 161 228 173 262
rect 115 222 173 228
rect -215 178 -169 190
rect -215 -178 -209 178
rect -175 -178 -169 178
rect -215 -190 -169 -178
rect -119 178 -73 190
rect -119 -178 -113 178
rect -79 -178 -73 178
rect -119 -190 -73 -178
rect -23 178 23 190
rect -23 -178 -17 178
rect 17 -178 23 178
rect -23 -190 23 -178
rect 73 178 119 190
rect 73 -178 79 178
rect 113 -178 119 178
rect 73 -190 119 -178
rect 169 178 215 190
rect 169 -178 175 178
rect 209 -178 215 178
rect 169 -190 215 -178
rect -173 -228 -115 -222
rect -173 -262 -161 -228
rect -127 -262 -115 -228
rect -173 -268 -115 -262
rect 19 -228 77 -222
rect 19 -262 31 -228
rect 65 -262 77 -228
rect 19 -268 77 -262
<< properties >>
string FIXED_BBOX -306 -347 306 347
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.9 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
