magic
tech sky130A
magscale 1 2
timestamp 1714331631
<< viali >>
rect 2053 7497 2087 7531
rect 2881 7497 2915 7531
rect 3801 7497 3835 7531
rect 4169 7497 4203 7531
rect 6101 7497 6135 7531
rect 6377 7497 6411 7531
rect 8493 7497 8527 7531
rect 8953 7497 8987 7531
rect 11713 7497 11747 7531
rect 13553 7497 13587 7531
rect 19441 7497 19475 7531
rect 26709 7497 26743 7531
rect 26985 7497 27019 7531
rect 27445 7497 27479 7531
rect 1409 7429 1443 7463
rect 1777 7429 1811 7463
rect 5549 7429 5583 7463
rect 5825 7429 5859 7463
rect 7573 7429 7607 7463
rect 8125 7429 8159 7463
rect 8401 7429 8435 7463
rect 9413 7429 9447 7463
rect 13461 7429 13495 7463
rect 15853 7429 15887 7463
rect 2237 7361 2271 7395
rect 2605 7361 2639 7395
rect 2697 7361 2731 7395
rect 3617 7361 3651 7395
rect 4261 7361 4295 7395
rect 4721 7361 4755 7395
rect 5641 7361 5675 7395
rect 6745 7361 6779 7395
rect 8217 7361 8251 7395
rect 9321 7361 9355 7395
rect 10425 7361 10459 7395
rect 10977 7361 11011 7395
rect 11069 7361 11103 7395
rect 11161 7361 11195 7395
rect 11621 7361 11655 7395
rect 12357 7361 12391 7395
rect 14289 7361 14323 7395
rect 15485 7361 15519 7395
rect 17509 7361 17543 7395
rect 18613 7361 18647 7395
rect 19257 7361 19291 7395
rect 22201 7361 22235 7395
rect 22753 7361 22787 7395
rect 23305 7361 23339 7395
rect 23856 7361 23890 7395
rect 23949 7361 23983 7395
rect 24225 7361 24259 7395
rect 26249 7361 26283 7395
rect 26525 7361 26559 7395
rect 27169 7361 27203 7395
rect 27261 7361 27295 7395
rect 4445 7293 4479 7327
rect 6837 7293 6871 7327
rect 7021 7293 7055 7327
rect 7665 7293 7699 7327
rect 7757 7293 7791 7327
rect 9597 7293 9631 7327
rect 12173 7293 12207 7327
rect 14105 7293 14139 7327
rect 14473 7293 14507 7327
rect 15301 7293 15335 7327
rect 18153 7293 18187 7327
rect 19809 7293 19843 7327
rect 20085 7293 20119 7327
rect 21925 7293 21959 7327
rect 25697 7293 25731 7327
rect 25973 7293 26007 7327
rect 3525 7225 3559 7259
rect 17601 7225 17635 7259
rect 17969 7225 18003 7259
rect 18061 7225 18095 7259
rect 18797 7225 18831 7259
rect 23581 7225 23615 7259
rect 2421 7157 2455 7191
rect 4813 7157 4847 7191
rect 7205 7157 7239 7191
rect 10333 7157 10367 7191
rect 10885 7157 10919 7191
rect 12541 7157 12575 7191
rect 15669 7157 15703 7191
rect 15945 7157 15979 7191
rect 17417 7157 17451 7191
rect 18429 7157 18463 7191
rect 21557 7157 21591 7191
rect 22661 7157 22695 7191
rect 23121 7157 23155 7191
rect 24041 7157 24075 7191
rect 26065 7157 26099 7191
rect 1501 6953 1535 6987
rect 1869 6953 1903 6987
rect 6469 6953 6503 6987
rect 7008 6953 7042 6987
rect 9216 6953 9250 6987
rect 10793 6953 10827 6987
rect 14197 6953 14231 6987
rect 15681 6953 15715 6987
rect 17785 6953 17819 6987
rect 18245 6953 18279 6987
rect 20545 6953 20579 6987
rect 18337 6885 18371 6919
rect 4169 6817 4203 6851
rect 6745 6817 6779 6851
rect 8953 6817 8987 6851
rect 11437 6817 11471 6851
rect 13737 6817 13771 6851
rect 18797 6817 18831 6851
rect 18981 6817 19015 6851
rect 19257 6817 19291 6851
rect 21189 6817 21223 6851
rect 21833 6817 21867 6851
rect 22385 6817 22419 6851
rect 1685 6749 1719 6783
rect 2053 6749 2087 6783
rect 2421 6749 2455 6783
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 6285 6749 6319 6783
rect 6439 6749 6473 6783
rect 11713 6749 11747 6783
rect 13645 6749 13679 6783
rect 15945 6749 15979 6783
rect 16037 6749 16071 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 18705 6749 18739 6783
rect 19441 6749 19475 6783
rect 19717 6749 19751 6783
rect 21557 6749 21591 6783
rect 22661 6749 22695 6783
rect 23304 6749 23338 6783
rect 23397 6749 23431 6783
rect 23765 6749 23799 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 24409 6749 24443 6783
rect 26525 6749 26559 6783
rect 26801 6749 26835 6783
rect 26893 6749 26927 6783
rect 27261 6749 27295 6783
rect 4445 6681 4479 6715
rect 6193 6681 6227 6715
rect 11161 6681 11195 6715
rect 11989 6681 12023 6715
rect 16313 6681 16347 6715
rect 19809 6681 19843 6715
rect 19993 6681 20027 6715
rect 21649 6681 21683 6715
rect 24685 6681 24719 6715
rect 2237 6613 2271 6647
rect 3617 6613 3651 6647
rect 8493 6613 8527 6647
rect 10701 6613 10735 6647
rect 11253 6613 11287 6647
rect 13461 6613 13495 6647
rect 19625 6613 19659 6647
rect 20913 6613 20947 6647
rect 21005 6613 21039 6647
rect 23029 6613 23063 6647
rect 23581 6613 23615 6647
rect 26157 6613 26191 6647
rect 26341 6613 26375 6647
rect 26617 6613 26651 6647
rect 27077 6613 27111 6647
rect 27445 6613 27479 6647
rect 1501 6409 1535 6443
rect 4629 6409 4663 6443
rect 4997 6409 5031 6443
rect 7941 6409 7975 6443
rect 9321 6409 9355 6443
rect 10701 6409 10735 6443
rect 10793 6409 10827 6443
rect 11161 6409 11195 6443
rect 12173 6409 12207 6443
rect 12633 6409 12667 6443
rect 14197 6409 14231 6443
rect 14565 6409 14599 6443
rect 15761 6409 15795 6443
rect 16129 6409 16163 6443
rect 19809 6409 19843 6443
rect 22753 6409 22787 6443
rect 24961 6409 24995 6443
rect 25421 6409 25455 6443
rect 27445 6409 27479 6443
rect 7757 6341 7791 6375
rect 16773 6341 16807 6375
rect 17785 6341 17819 6375
rect 18337 6341 18371 6375
rect 23397 6341 23431 6375
rect 25329 6341 25363 6375
rect 1685 6273 1719 6307
rect 2053 6273 2087 6307
rect 2145 6273 2179 6307
rect 5641 6273 5675 6307
rect 5917 6273 5951 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 8769 6273 8803 6307
rect 9229 6273 9263 6307
rect 9689 6273 9723 6307
rect 10333 6273 10367 6307
rect 12541 6273 12575 6307
rect 13001 6273 13035 6307
rect 13185 6273 13219 6307
rect 13461 6273 13495 6307
rect 13645 6273 13679 6307
rect 14749 6273 14783 6307
rect 15209 6273 15243 6307
rect 15669 6273 15703 6307
rect 16221 6273 16255 6307
rect 16405 6273 16439 6307
rect 16957 6273 16991 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 19901 6273 19935 6307
rect 22017 6273 22051 6307
rect 22385 6273 22419 6307
rect 22569 6273 22603 6307
rect 23029 6273 23063 6307
rect 26525 6273 26559 6307
rect 27261 6273 27295 6307
rect 2421 6205 2455 6239
rect 4169 6205 4203 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 5457 6205 5491 6239
rect 5733 6205 5767 6239
rect 5825 6205 5859 6239
rect 6469 6205 6503 6239
rect 6745 6205 6779 6239
rect 9781 6205 9815 6239
rect 9873 6205 9907 6239
rect 10517 6205 10551 6239
rect 12817 6205 12851 6239
rect 14013 6205 14047 6239
rect 14105 6205 14139 6239
rect 15577 6205 15611 6239
rect 18061 6205 18095 6239
rect 21649 6205 21683 6239
rect 22293 6205 22327 6239
rect 22477 6205 22511 6239
rect 23121 6205 23155 6239
rect 25513 6205 25547 6239
rect 1869 6137 1903 6171
rect 10241 6137 10275 6171
rect 16313 6137 16347 6171
rect 16681 6137 16715 6171
rect 7665 6069 7699 6103
rect 8677 6069 8711 6103
rect 9045 6069 9079 6103
rect 13093 6069 13127 6103
rect 13553 6069 13587 6103
rect 14841 6069 14875 6103
rect 15117 6069 15151 6103
rect 17693 6069 17727 6103
rect 21925 6069 21959 6103
rect 22937 6069 22971 6103
rect 24869 6069 24903 6103
rect 26709 6069 26743 6103
rect 3801 5865 3835 5899
rect 5733 5865 5767 5899
rect 6101 5865 6135 5899
rect 7205 5865 7239 5899
rect 7941 5865 7975 5899
rect 8953 5865 8987 5899
rect 9321 5865 9355 5899
rect 9505 5865 9539 5899
rect 12541 5865 12575 5899
rect 13645 5865 13679 5899
rect 14289 5865 14323 5899
rect 15761 5865 15795 5899
rect 18153 5865 18187 5899
rect 19349 5865 19383 5899
rect 19809 5865 19843 5899
rect 27445 5865 27479 5899
rect 1501 5797 1535 5831
rect 3157 5797 3191 5831
rect 13553 5797 13587 5831
rect 17417 5797 17451 5831
rect 27077 5797 27111 5831
rect 4445 5729 4479 5763
rect 4629 5729 4663 5763
rect 4905 5729 4939 5763
rect 5089 5729 5123 5763
rect 6653 5729 6687 5763
rect 9045 5729 9079 5763
rect 9137 5729 9171 5763
rect 9873 5729 9907 5763
rect 11989 5729 12023 5763
rect 12357 5729 12391 5763
rect 12449 5729 12483 5763
rect 12633 5729 12667 5763
rect 13001 5729 13035 5763
rect 13737 5729 13771 5763
rect 14933 5729 14967 5763
rect 15301 5729 15335 5763
rect 15577 5729 15611 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 19533 5729 19567 5763
rect 22477 5729 22511 5763
rect 24409 5729 24443 5763
rect 24685 5729 24719 5763
rect 1685 5661 1719 5695
rect 2053 5661 2087 5695
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5365 5661 5399 5695
rect 5457 5661 5491 5695
rect 5549 5661 5583 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 6929 5661 6963 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8309 5661 8343 5695
rect 8401 5661 8435 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 12725 5661 12759 5695
rect 13093 5661 13127 5695
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 13461 5661 13495 5695
rect 14473 5661 14507 5695
rect 14565 5661 14599 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 15945 5661 15979 5695
rect 16037 5661 16071 5695
rect 16129 5661 16163 5695
rect 16247 5661 16281 5695
rect 16405 5661 16439 5695
rect 17325 5661 17359 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 18521 5661 18555 5695
rect 18613 5661 18647 5695
rect 18889 5661 18923 5695
rect 19257 5661 19291 5695
rect 19901 5661 19935 5695
rect 21741 5661 21775 5695
rect 21925 5661 21959 5695
rect 22017 5661 22051 5695
rect 22109 5661 22143 5695
rect 26525 5661 26559 5695
rect 26893 5661 26927 5695
rect 27261 5661 27295 5695
rect 6561 5593 6595 5627
rect 7021 5593 7055 5627
rect 11713 5593 11747 5627
rect 14657 5593 14691 5627
rect 14795 5593 14829 5627
rect 16840 5593 16874 5627
rect 16957 5593 16991 5627
rect 17576 5593 17610 5627
rect 19073 5593 19107 5627
rect 20177 5593 20211 5627
rect 22753 5593 22787 5627
rect 1869 5525 1903 5559
rect 4261 5525 4295 5559
rect 6009 5525 6043 5559
rect 6469 5525 6503 5559
rect 7573 5525 7607 5559
rect 7757 5525 7791 5559
rect 8585 5525 8619 5559
rect 10241 5525 10275 5559
rect 12817 5525 12851 5559
rect 15301 5525 15335 5559
rect 16681 5525 16715 5559
rect 17049 5525 17083 5559
rect 17693 5525 17727 5559
rect 21649 5525 21683 5559
rect 22385 5525 22419 5559
rect 24225 5525 24259 5559
rect 26157 5525 26191 5559
rect 26709 5525 26743 5559
rect 1501 5321 1535 5355
rect 8769 5321 8803 5355
rect 9873 5321 9907 5355
rect 9965 5321 9999 5355
rect 13645 5321 13679 5355
rect 18429 5321 18463 5355
rect 20269 5321 20303 5355
rect 20729 5321 20763 5355
rect 22569 5321 22603 5355
rect 24225 5321 24259 5355
rect 27445 5321 27479 5355
rect 9505 5253 9539 5287
rect 11253 5253 11287 5287
rect 11897 5253 11931 5287
rect 12449 5253 12483 5287
rect 12633 5253 12667 5287
rect 14933 5253 14967 5287
rect 16773 5253 16807 5287
rect 19533 5253 19567 5287
rect 23489 5253 23523 5287
rect 25237 5253 25271 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 3249 5185 3283 5219
rect 3433 5185 3467 5219
rect 3709 5185 3743 5219
rect 4077 5185 4111 5219
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 5357 5185 5391 5219
rect 5549 5175 5583 5209
rect 5665 5185 5699 5219
rect 6101 5185 6135 5219
rect 6469 5185 6503 5219
rect 6837 5185 6871 5219
rect 7205 5185 7239 5219
rect 7665 5185 7699 5219
rect 7849 5185 7883 5219
rect 7941 5185 7975 5219
rect 8033 5185 8067 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 9044 5185 9078 5219
rect 9137 5185 9171 5219
rect 9229 5185 9263 5219
rect 9322 5185 9356 5219
rect 9597 5185 9631 5219
rect 9694 5185 9728 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 10885 5185 10919 5219
rect 11161 5185 11195 5219
rect 11345 5185 11379 5219
rect 12357 5185 12391 5219
rect 12541 5185 12575 5219
rect 12725 5185 12759 5219
rect 13093 5185 13127 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 15761 5185 15795 5219
rect 16865 5185 16899 5219
rect 17325 5185 17359 5219
rect 17509 5185 17543 5219
rect 17969 5185 18003 5219
rect 18889 5185 18923 5219
rect 19165 5185 19199 5219
rect 19257 5185 19291 5219
rect 19349 5185 19383 5219
rect 20453 5185 20487 5219
rect 20913 5185 20947 5219
rect 21189 5185 21223 5219
rect 21557 5175 21591 5209
rect 21833 5185 21867 5219
rect 22293 5185 22327 5219
rect 22753 5185 22787 5219
rect 23121 5185 23155 5219
rect 23305 5185 23339 5219
rect 23765 5185 23799 5219
rect 23857 5185 23891 5219
rect 24133 5185 24167 5219
rect 24317 5185 24351 5219
rect 24409 5185 24443 5219
rect 24593 5185 24627 5219
rect 24869 5185 24903 5219
rect 25881 5185 25915 5219
rect 26525 5185 26559 5219
rect 27261 5185 27295 5219
rect 3525 5117 3559 5151
rect 4353 5117 4387 5151
rect 5917 5117 5951 5151
rect 6561 5117 6595 5151
rect 6929 5117 6963 5151
rect 7113 5117 7147 5151
rect 7297 5117 7331 5151
rect 7389 5117 7423 5151
rect 10701 5117 10735 5151
rect 11069 5117 11103 5151
rect 11989 5117 12023 5151
rect 12081 5117 12115 5151
rect 12817 5117 12851 5151
rect 15025 5117 15059 5151
rect 16037 5117 16071 5151
rect 16497 5117 16531 5151
rect 18061 5117 18095 5151
rect 18153 5117 18187 5151
rect 18613 5117 18647 5151
rect 18705 5117 18739 5151
rect 18797 5117 18831 5151
rect 19717 5117 19751 5151
rect 20545 5117 20579 5151
rect 20821 5117 20855 5151
rect 22109 5117 22143 5151
rect 6377 5049 6411 5083
rect 11529 5049 11563 5083
rect 15209 5049 15243 5083
rect 15669 5049 15703 5083
rect 16221 5049 16255 5083
rect 17417 5049 17451 5083
rect 17601 5049 17635 5083
rect 19993 5049 20027 5083
rect 20177 5049 20211 5083
rect 1869 4981 1903 5015
rect 2145 4981 2179 5015
rect 3433 4981 3467 5015
rect 3893 4981 3927 5015
rect 4445 4981 4479 5015
rect 4629 4981 4663 5015
rect 4813 4981 4847 5015
rect 5457 4981 5491 5015
rect 5733 4981 5767 5015
rect 6745 4981 6779 5015
rect 8493 4981 8527 5015
rect 13001 4981 13035 5015
rect 21005 4981 21039 5015
rect 21465 4981 21499 5015
rect 22293 4981 22327 5015
rect 22477 4981 22511 5015
rect 22753 4981 22787 5015
rect 23949 4981 23983 5015
rect 24593 4981 24627 5015
rect 25053 4981 25087 5015
rect 26709 4981 26743 5015
rect 2132 4777 2166 4811
rect 3801 4777 3835 4811
rect 4905 4777 4939 4811
rect 5641 4777 5675 4811
rect 11805 4777 11839 4811
rect 12541 4777 12575 4811
rect 13001 4777 13035 4811
rect 13369 4777 13403 4811
rect 15393 4777 15427 4811
rect 15945 4777 15979 4811
rect 22017 4777 22051 4811
rect 27445 4777 27479 4811
rect 1501 4709 1535 4743
rect 3617 4709 3651 4743
rect 4997 4709 5031 4743
rect 8401 4709 8435 4743
rect 9321 4709 9355 4743
rect 9689 4709 9723 4743
rect 15853 4709 15887 4743
rect 20361 4709 20395 4743
rect 21097 4709 21131 4743
rect 21833 4709 21867 4743
rect 24409 4709 24443 4743
rect 1869 4641 1903 4675
rect 4445 4641 4479 4675
rect 12633 4641 12667 4675
rect 13737 4641 13771 4675
rect 15117 4641 15151 4675
rect 15761 4641 15795 4675
rect 19809 4641 19843 4675
rect 20637 4641 20671 4675
rect 20729 4641 20763 4675
rect 20821 4641 20855 4675
rect 23765 4641 23799 4675
rect 1685 4573 1719 4607
rect 4169 4573 4203 4607
rect 4721 4573 4755 4607
rect 4813 4573 4847 4607
rect 5089 4573 5123 4607
rect 6929 4573 6963 4607
rect 7389 4573 7423 4607
rect 7665 4573 7699 4607
rect 7941 4573 7975 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 8585 4573 8619 4607
rect 9597 4573 9631 4607
rect 9689 4573 9723 4607
rect 9781 4573 9815 4607
rect 9965 4573 9999 4607
rect 10057 4573 10091 4607
rect 10149 4573 10183 4607
rect 10519 4573 10553 4607
rect 12909 4573 12943 4607
rect 13001 4573 13035 4607
rect 13185 4573 13219 4607
rect 13461 4573 13495 4607
rect 13553 4573 13587 4607
rect 14105 4573 14139 4607
rect 14381 4573 14415 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 15485 4573 15519 4607
rect 16037 4573 16071 4607
rect 16129 4573 16163 4607
rect 16313 4573 16347 4607
rect 16405 4573 16439 4607
rect 16589 4573 16623 4607
rect 16773 4573 16807 4607
rect 16957 4573 16991 4607
rect 17049 4573 17083 4607
rect 17233 4573 17267 4607
rect 17325 4573 17359 4607
rect 17509 4573 17543 4607
rect 17601 4573 17635 4607
rect 17785 4573 17819 4607
rect 17877 4573 17911 4607
rect 18153 4573 18187 4607
rect 18245 4573 18279 4607
rect 18429 4573 18463 4607
rect 18521 4573 18555 4607
rect 18797 4573 18831 4607
rect 18981 4573 19015 4607
rect 19717 4573 19751 4607
rect 20269 4573 20303 4607
rect 20545 4573 20579 4607
rect 21005 4573 21039 4607
rect 21189 4573 21223 4607
rect 21281 4573 21315 4607
rect 21649 4573 21683 4607
rect 24041 4573 24075 4607
rect 24225 4573 24259 4607
rect 26157 4573 26191 4607
rect 26249 4573 26283 4607
rect 26617 4573 26651 4607
rect 26893 4573 26927 4607
rect 27261 4573 27295 4607
rect 8033 4505 8067 4539
rect 8217 4505 8251 4539
rect 9137 4505 9171 4539
rect 9413 4505 9447 4539
rect 17969 4505 18003 4539
rect 19625 4505 19659 4539
rect 20177 4505 20211 4539
rect 21465 4505 21499 4539
rect 21557 4505 21591 4539
rect 23489 4505 23523 4539
rect 25881 4505 25915 4539
rect 4261 4437 4295 4471
rect 7113 4437 7147 4471
rect 10425 4437 10459 4471
rect 12357 4437 12391 4471
rect 13737 4437 13771 4471
rect 16221 4437 16255 4471
rect 16497 4437 16531 4471
rect 16773 4437 16807 4471
rect 17049 4437 17083 4471
rect 18981 4437 19015 4471
rect 19257 4437 19291 4471
rect 23857 4437 23891 4471
rect 26341 4437 26375 4471
rect 26801 4437 26835 4471
rect 27077 4437 27111 4471
rect 6377 4233 6411 4267
rect 7113 4233 7147 4267
rect 11069 4233 11103 4267
rect 11529 4233 11563 4267
rect 13001 4233 13035 4267
rect 23305 4233 23339 4267
rect 23581 4233 23615 4267
rect 4905 4165 4939 4199
rect 7297 4165 7331 4199
rect 9505 4165 9539 4199
rect 13277 4165 13311 4199
rect 16957 4165 16991 4199
rect 18061 4165 18095 4199
rect 19533 4165 19567 4199
rect 19901 4165 19935 4199
rect 21557 4165 21591 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2237 4097 2271 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5089 4097 5123 4131
rect 5503 4097 5537 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 5916 4097 5950 4131
rect 6009 4097 6043 4131
rect 6556 4097 6590 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 6928 4097 6962 4131
rect 7021 4097 7055 4131
rect 7481 4097 7515 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 8033 4097 8067 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8493 4097 8527 4131
rect 8769 4097 8803 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 9413 4097 9447 4131
rect 9689 4097 9723 4131
rect 9965 4097 9999 4131
rect 10058 4097 10092 4131
rect 10241 4097 10275 4131
rect 10333 4097 10367 4131
rect 10471 4097 10505 4131
rect 10885 4097 10919 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 11989 4097 12023 4131
rect 12265 4097 12299 4131
rect 12357 4097 12391 4131
rect 12449 4097 12483 4131
rect 12633 4097 12667 4131
rect 12817 4097 12851 4131
rect 13461 4097 13495 4131
rect 13553 4097 13587 4131
rect 13737 4097 13771 4131
rect 13829 4097 13863 4131
rect 14105 4097 14139 4131
rect 14381 4097 14415 4131
rect 14841 4097 14875 4131
rect 15301 4097 15335 4131
rect 15393 4097 15427 4131
rect 15853 4097 15887 4131
rect 16159 4097 16193 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 17049 4097 17083 4131
rect 17141 4097 17175 4131
rect 17785 4097 17819 4131
rect 17969 4097 18003 4131
rect 18153 4097 18187 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 18981 4097 19015 4131
rect 19158 4097 19192 4131
rect 19303 4097 19337 4131
rect 19441 4097 19475 4131
rect 19625 4097 19659 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 22753 4097 22787 4131
rect 22937 4097 22971 4131
rect 23029 4097 23063 4131
rect 23121 4097 23155 4131
rect 23857 4097 23891 4131
rect 24133 4097 24167 4131
rect 25789 4097 25823 4131
rect 26065 4097 26099 4131
rect 26249 4097 26283 4131
rect 26525 4097 26559 4131
rect 26985 4097 27019 4131
rect 27261 4097 27295 4131
rect 2513 4029 2547 4063
rect 4261 4029 4295 4063
rect 4813 4029 4847 4063
rect 7665 4029 7699 4063
rect 7849 4029 7883 4063
rect 8861 4029 8895 4063
rect 9873 4029 9907 4063
rect 10701 4029 10735 4063
rect 12081 4029 12115 4063
rect 13921 4029 13955 4063
rect 14197 4029 14231 4063
rect 14289 4029 14323 4063
rect 14657 4029 14691 4063
rect 15025 4029 15059 4063
rect 15117 4029 15151 4063
rect 16681 4029 16715 4063
rect 18797 4029 18831 4063
rect 23765 4029 23799 4063
rect 24225 4029 24259 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 1501 3961 1535 3995
rect 1869 3961 1903 3995
rect 5273 3961 5307 3995
rect 10609 3961 10643 3995
rect 14933 3961 14967 3995
rect 15669 3961 15703 3995
rect 15945 3961 15979 3995
rect 25513 3961 25547 3995
rect 26065 3961 26099 3995
rect 27445 3961 27479 3995
rect 5365 3893 5399 3927
rect 8585 3893 8619 3927
rect 12633 3893 12667 3927
rect 15531 3893 15565 3927
rect 15761 3893 15795 3927
rect 18337 3893 18371 3927
rect 19073 3893 19107 3927
rect 19809 3893 19843 3927
rect 24501 3893 24535 3927
rect 25697 3893 25731 3927
rect 25881 3893 25915 3927
rect 26709 3893 26743 3927
rect 27077 3893 27111 3927
rect 1501 3689 1535 3723
rect 6009 3689 6043 3723
rect 6193 3689 6227 3723
rect 6745 3689 6779 3723
rect 10149 3689 10183 3723
rect 13277 3689 13311 3723
rect 14933 3689 14967 3723
rect 19073 3689 19107 3723
rect 20269 3689 20303 3723
rect 27445 3689 27479 3723
rect 13461 3621 13495 3655
rect 19809 3621 19843 3655
rect 23489 3621 23523 3655
rect 1869 3553 1903 3587
rect 3617 3553 3651 3587
rect 5365 3553 5399 3587
rect 6285 3553 6319 3587
rect 8125 3553 8159 3587
rect 10333 3553 10367 3587
rect 12357 3553 12391 3587
rect 15117 3553 15151 3587
rect 17969 3553 18003 3587
rect 19901 3553 19935 3587
rect 23397 3553 23431 3587
rect 24593 3553 24627 3587
rect 24777 3553 24811 3587
rect 25421 3553 25455 3587
rect 1685 3485 1719 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4629 3485 4663 3519
rect 4721 3485 4755 3519
rect 4905 3485 4939 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6377 3485 6411 3519
rect 6653 3485 6687 3519
rect 6837 3485 6871 3519
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 7941 3485 7975 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9137 3485 9171 3519
rect 9689 3485 9723 3519
rect 9781 3485 9815 3519
rect 9965 3485 9999 3519
rect 10057 3485 10091 3519
rect 10241 3485 10275 3519
rect 12449 3485 12483 3519
rect 13921 3485 13955 3519
rect 14105 3485 14139 3519
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 15301 3485 15335 3519
rect 16497 3485 16531 3519
rect 16681 3485 16715 3519
rect 18705 3485 18739 3519
rect 18797 3485 18831 3519
rect 18889 3485 18923 3519
rect 19533 3485 19567 3519
rect 20545 3485 20579 3519
rect 23213 3485 23247 3519
rect 23673 3485 23707 3519
rect 24225 3485 24259 3519
rect 25053 3485 25087 3519
rect 25697 3485 25731 3519
rect 25789 3485 25823 3519
rect 26157 3485 26191 3519
rect 26525 3485 26559 3519
rect 26893 3485 26927 3519
rect 27261 3485 27295 3519
rect 2145 3417 2179 3451
rect 3801 3417 3835 3451
rect 7573 3417 7607 3451
rect 7665 3417 7699 3451
rect 8217 3417 8251 3451
rect 10609 3417 10643 3451
rect 13093 3417 13127 3451
rect 14289 3417 14323 3451
rect 14381 3417 14415 3451
rect 18153 3417 18187 3451
rect 18245 3417 18279 3451
rect 18521 3417 18555 3451
rect 19257 3417 19291 3451
rect 20269 3417 20303 3451
rect 20821 3417 20855 3451
rect 22569 3417 22603 3451
rect 4169 3349 4203 3383
rect 4445 3349 4479 3383
rect 5457 3349 5491 3383
rect 5825 3349 5859 3383
rect 8493 3349 8527 3383
rect 8953 3349 8987 3383
rect 9597 3349 9631 3383
rect 9873 3349 9907 3383
rect 12633 3349 12667 3383
rect 12725 3349 12759 3383
rect 12817 3349 12851 3383
rect 13001 3349 13035 3383
rect 13293 3349 13327 3383
rect 13737 3349 13771 3383
rect 14657 3349 14691 3383
rect 16589 3349 16623 3383
rect 18337 3349 18371 3383
rect 19441 3349 19475 3383
rect 19625 3349 19659 3383
rect 20453 3349 20487 3383
rect 22661 3349 22695 3383
rect 23857 3349 23891 3383
rect 24041 3349 24075 3383
rect 24685 3349 24719 3383
rect 25513 3349 25547 3383
rect 25973 3349 26007 3383
rect 26341 3349 26375 3383
rect 26709 3349 26743 3383
rect 27077 3349 27111 3383
rect 1869 3145 1903 3179
rect 4261 3145 4295 3179
rect 5457 3145 5491 3179
rect 5733 3145 5767 3179
rect 7573 3145 7607 3179
rect 8309 3145 8343 3179
rect 8677 3145 8711 3179
rect 8769 3145 8803 3179
rect 10609 3145 10643 3179
rect 21005 3145 21039 3179
rect 21833 3145 21867 3179
rect 24133 3145 24167 3179
rect 25697 3145 25731 3179
rect 27445 3145 27479 3179
rect 2421 3077 2455 3111
rect 4629 3077 4663 3111
rect 5917 3077 5951 3111
rect 9597 3077 9631 3111
rect 9689 3077 9723 3111
rect 10333 3077 10367 3111
rect 11805 3077 11839 3111
rect 14197 3077 14231 3111
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2145 3009 2179 3043
rect 4445 3009 4479 3043
rect 4537 3009 4571 3043
rect 4813 3009 4847 3043
rect 4905 3009 4939 3043
rect 5181 3009 5215 3043
rect 5641 3009 5675 3043
rect 6101 3009 6135 3043
rect 6193 3009 6227 3043
rect 6469 3009 6503 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 7849 3009 7883 3043
rect 8953 3009 8987 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 9781 3009 9815 3043
rect 10057 3009 10091 3043
rect 10241 3009 10275 3043
rect 10425 3009 10459 3043
rect 11529 3009 11563 3043
rect 11713 3009 11747 3043
rect 11897 3009 11931 3043
rect 12173 3009 12207 3043
rect 16313 3009 16347 3043
rect 16681 3009 16715 3043
rect 18981 3009 19015 3043
rect 19073 3009 19107 3043
rect 19257 3009 19291 3043
rect 19717 3009 19751 3043
rect 20177 3009 20211 3043
rect 20545 3009 20579 3043
rect 20637 3009 20671 3043
rect 20821 3009 20855 3043
rect 21097 3009 21131 3043
rect 21281 3009 21315 3043
rect 21373 3009 21407 3043
rect 21465 3009 21499 3043
rect 22385 3009 22419 3043
rect 24501 3009 24535 3043
rect 24685 3009 24719 3043
rect 24777 3009 24811 3043
rect 24961 3009 24995 3043
rect 25053 3009 25087 3043
rect 25145 3009 25179 3043
rect 25329 3009 25363 3043
rect 25881 3009 25915 3043
rect 25973 3009 26007 3043
rect 26525 3009 26559 3043
rect 26985 3009 27019 3043
rect 27169 3009 27203 3043
rect 27261 3009 27295 3043
rect 4169 2941 4203 2975
rect 7297 2941 7331 2975
rect 8033 2941 8067 2975
rect 8217 2941 8251 2975
rect 9137 2941 9171 2975
rect 12449 2941 12483 2975
rect 14289 2941 14323 2975
rect 16037 2941 16071 2975
rect 16957 2941 16991 2975
rect 18705 2941 18739 2975
rect 19809 2941 19843 2975
rect 20269 2941 20303 2975
rect 22017 2941 22051 2975
rect 22109 2941 22143 2975
rect 22201 2941 22235 2975
rect 22661 2941 22695 2975
rect 25513 2941 25547 2975
rect 1501 2873 1535 2907
rect 6193 2873 6227 2907
rect 12081 2873 12115 2907
rect 19533 2873 19567 2907
rect 21649 2873 21683 2907
rect 24593 2873 24627 2907
rect 26157 2873 26191 2907
rect 26985 2873 27019 2907
rect 4997 2805 5031 2839
rect 6469 2805 6503 2839
rect 7297 2805 7331 2839
rect 7757 2805 7791 2839
rect 9965 2805 9999 2839
rect 18797 2805 18831 2839
rect 19073 2805 19107 2839
rect 24317 2805 24351 2839
rect 26709 2805 26743 2839
rect 1501 2601 1535 2635
rect 1869 2601 1903 2635
rect 3801 2601 3835 2635
rect 5549 2601 5583 2635
rect 5733 2601 5767 2635
rect 5917 2601 5951 2635
rect 6837 2601 6871 2635
rect 9505 2601 9539 2635
rect 12449 2601 12483 2635
rect 13461 2601 13495 2635
rect 14657 2601 14691 2635
rect 15577 2601 15611 2635
rect 16405 2601 16439 2635
rect 17785 2601 17819 2635
rect 21465 2601 21499 2635
rect 22017 2601 22051 2635
rect 23673 2601 23707 2635
rect 24133 2601 24167 2635
rect 26525 2601 26559 2635
rect 2605 2533 2639 2567
rect 4905 2533 4939 2567
rect 6377 2533 6411 2567
rect 8033 2533 8067 2567
rect 13001 2533 13035 2567
rect 23397 2533 23431 2567
rect 23489 2533 23523 2567
rect 5457 2465 5491 2499
rect 7849 2465 7883 2499
rect 9781 2465 9815 2499
rect 9891 2465 9925 2499
rect 12633 2465 12667 2499
rect 13645 2465 13679 2499
rect 13829 2465 13863 2499
rect 14841 2465 14875 2499
rect 17509 2465 17543 2499
rect 17601 2465 17635 2499
rect 19257 2465 19291 2499
rect 21281 2465 21315 2499
rect 23029 2465 23063 2499
rect 25605 2465 25639 2499
rect 26157 2465 26191 2499
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 2421 2397 2455 2431
rect 2789 2397 2823 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4077 2397 4111 2431
rect 4169 2397 4203 2431
rect 4353 2397 4387 2431
rect 4721 2397 4755 2431
rect 5089 2397 5123 2431
rect 5181 2397 5215 2431
rect 6101 2397 6135 2431
rect 6561 2397 6595 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7113 2397 7147 2431
rect 7205 2397 7239 2431
rect 7665 2397 7699 2431
rect 7757 2397 7791 2431
rect 8125 2397 8159 2431
rect 8309 2397 8343 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 9696 2397 9730 2431
rect 10057 2397 10091 2431
rect 10609 2397 10643 2431
rect 10701 2397 10735 2431
rect 10885 2397 10919 2431
rect 10977 2397 11011 2431
rect 11161 2397 11195 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 12725 2397 12759 2431
rect 12817 2397 12851 2431
rect 13093 2397 13127 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 14381 2397 14415 2431
rect 14473 2397 14507 2431
rect 14749 2397 14783 2431
rect 14933 2397 14967 2431
rect 15025 2397 15059 2431
rect 15761 2397 15795 2431
rect 15853 2397 15887 2431
rect 16129 2397 16163 2431
rect 16221 2397 16255 2431
rect 16865 2397 16899 2431
rect 17417 2397 17451 2431
rect 17877 2397 17911 2431
rect 18245 2397 18279 2431
rect 18981 2397 19015 2431
rect 21649 2397 21683 2431
rect 21833 2397 21867 2431
rect 22477 2397 22511 2431
rect 22661 2397 22695 2431
rect 22937 2397 22971 2431
rect 23857 2397 23891 2431
rect 23949 2397 23983 2431
rect 24409 2397 24443 2431
rect 25237 2397 25271 2431
rect 25329 2397 25363 2431
rect 25513 2397 25547 2431
rect 25789 2397 25823 2431
rect 26341 2397 26375 2431
rect 26617 2397 26651 2431
rect 26801 2397 26835 2431
rect 3065 2329 3099 2363
rect 3249 2329 3283 2363
rect 7021 2329 7055 2363
rect 8401 2329 8435 2363
rect 11069 2329 11103 2363
rect 14289 2329 14323 2363
rect 16037 2329 16071 2363
rect 18061 2329 18095 2363
rect 18153 2329 18187 2363
rect 21005 2329 21039 2363
rect 22569 2329 22603 2363
rect 22799 2329 22833 2363
rect 25973 2329 26007 2363
rect 27169 2329 27203 2363
rect 27537 2329 27571 2363
rect 2237 2261 2271 2295
rect 3525 2261 3559 2295
rect 4537 2261 4571 2295
rect 7389 2261 7423 2295
rect 8677 2261 8711 2295
rect 9229 2261 9263 2295
rect 10241 2261 10275 2295
rect 10425 2261 10459 2295
rect 10793 2261 10827 2295
rect 11713 2261 11747 2295
rect 13277 2261 13311 2295
rect 15209 2261 15243 2295
rect 17049 2261 17083 2295
rect 18429 2261 18463 2295
rect 18797 2261 18831 2295
rect 22293 2261 22327 2295
rect 24593 2261 24627 2295
rect 25053 2261 25087 2295
rect 25421 2261 25455 2295
rect 26709 2261 26743 2295
<< metal1 >>
rect 18230 7964 18236 8016
rect 18288 8004 18294 8016
rect 26970 8004 26976 8016
rect 18288 7976 26976 8004
rect 18288 7964 18294 7976
rect 26970 7964 26976 7976
rect 27028 7964 27034 8016
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 27338 7936 27344 7948
rect 7524 7908 27344 7936
rect 7524 7896 7530 7908
rect 27338 7896 27344 7908
rect 27396 7896 27402 7948
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 25038 7868 25044 7880
rect 10376 7840 25044 7868
rect 10376 7828 10382 7840
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 8202 7800 8208 7812
rect 7064 7772 8208 7800
rect 7064 7760 7070 7772
rect 8202 7760 8208 7772
rect 8260 7800 8266 7812
rect 11330 7800 11336 7812
rect 8260 7772 11336 7800
rect 8260 7760 8266 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 20438 7800 20444 7812
rect 15252 7772 20444 7800
rect 15252 7760 15258 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 1210 7692 1216 7744
rect 1268 7732 1274 7744
rect 2682 7732 2688 7744
rect 1268 7704 2688 7732
rect 1268 7692 1274 7704
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 17954 7732 17960 7744
rect 2924 7704 17960 7732
rect 2924 7692 2930 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 26510 7732 26516 7744
rect 19024 7704 26516 7732
rect 19024 7692 19030 7704
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 1104 7642 27876 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 27876 7642
rect 1104 7568 27876 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1176 7500 2053 7528
rect 1176 7488 1182 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 2866 7488 2872 7540
rect 2924 7488 2930 7540
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7497 3847 7531
rect 3789 7491 3847 7497
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 4203 7500 6040 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 1397 7463 1455 7469
rect 1397 7460 1409 7463
rect 1360 7432 1409 7460
rect 1360 7420 1366 7432
rect 1397 7429 1409 7432
rect 1443 7429 1455 7463
rect 1397 7423 1455 7429
rect 1765 7463 1823 7469
rect 1765 7429 1777 7463
rect 1811 7460 1823 7463
rect 2774 7460 2780 7472
rect 1811 7432 2780 7460
rect 1811 7429 1823 7432
rect 1765 7423 1823 7429
rect 2774 7420 2780 7432
rect 2832 7420 2838 7472
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2240 7324 2268 7355
rect 2590 7352 2596 7404
rect 2648 7352 2654 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 3804 7392 3832 7491
rect 5537 7463 5595 7469
rect 3651 7364 3832 7392
rect 4172 7432 5488 7460
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4172 7324 4200 7432
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4614 7392 4620 7404
rect 4295 7364 4620 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 2240 7296 4200 7324
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4396 7296 4445 7324
rect 4396 7284 4402 7296
rect 4433 7293 4445 7296
rect 4479 7324 4491 7327
rect 4479 7296 5396 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 4706 7256 4712 7268
rect 3559 7228 4712 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 3752 7160 4813 7188
rect 3752 7148 3758 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 5368 7188 5396 7296
rect 5460 7256 5488 7432
rect 5537 7429 5549 7463
rect 5583 7460 5595 7463
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5583 7432 5825 7460
rect 5583 7429 5595 7432
rect 5537 7423 5595 7429
rect 5813 7429 5825 7432
rect 5859 7429 5871 7463
rect 6012 7460 6040 7500
rect 6086 7488 6092 7540
rect 6144 7488 6150 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6178 7460 6184 7472
rect 6012 7432 6184 7460
rect 5813 7423 5871 7429
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 6380 7392 6408 7491
rect 8478 7488 8484 7540
rect 8536 7488 8542 7540
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 7558 7420 7564 7472
rect 7616 7420 7622 7472
rect 8113 7463 8171 7469
rect 8113 7429 8125 7463
rect 8159 7460 8171 7463
rect 8389 7463 8447 7469
rect 8389 7460 8401 7463
rect 8159 7432 8401 7460
rect 8159 7429 8171 7432
rect 8113 7423 8171 7429
rect 8389 7429 8401 7432
rect 8435 7429 8447 7463
rect 8389 7423 8447 7429
rect 5675 7364 6408 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6696 7364 6745 7392
rect 6696 7352 6702 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8956 7392 8984 7491
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 10928 7500 11713 7528
rect 10928 7488 10934 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13320 7500 13553 7528
rect 13320 7488 13326 7500
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 13541 7491 13599 7497
rect 15286 7488 15292 7540
rect 15344 7528 15350 7540
rect 15344 7500 17540 7528
rect 15344 7488 15350 7500
rect 9030 7420 9036 7472
rect 9088 7460 9094 7472
rect 9401 7463 9459 7469
rect 9401 7460 9413 7463
rect 9088 7432 9413 7460
rect 9088 7420 9094 7432
rect 9401 7429 9413 7432
rect 9447 7429 9459 7463
rect 11238 7460 11244 7472
rect 9401 7423 9459 7429
rect 10980 7432 11244 7460
rect 8251 7364 8984 7392
rect 9309 7395 9367 7401
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10870 7392 10876 7404
rect 10459 7364 10876 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6328 7296 6837 7324
rect 6328 7284 6334 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7006 7284 7012 7336
rect 7064 7284 7070 7336
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7742 7284 7748 7336
rect 7800 7284 7806 7336
rect 9324 7256 9352 7355
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10980 7401 11008 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 12434 7420 12440 7472
rect 12492 7460 12498 7472
rect 13449 7463 13507 7469
rect 13449 7460 13461 7463
rect 12492 7432 13461 7460
rect 12492 7420 12498 7432
rect 13449 7429 13461 7432
rect 13495 7429 13507 7463
rect 13449 7423 13507 7429
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 15841 7463 15899 7469
rect 15841 7460 15853 7463
rect 13872 7432 15853 7460
rect 13872 7420 13878 7432
rect 15841 7429 15853 7432
rect 15887 7429 15899 7463
rect 15841 7423 15899 7429
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11195 7364 11621 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11609 7361 11621 7364
rect 11655 7361 11667 7395
rect 11609 7355 11667 7361
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 9766 7324 9772 7336
rect 9631 7296 9772 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11072 7324 11100 7355
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 17512 7401 17540 7500
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19484 7500 22232 7528
rect 19484 7488 19490 7500
rect 19058 7460 19064 7472
rect 17880 7432 19064 7460
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 12400 7364 14289 7392
rect 12400 7352 12406 7364
rect 14277 7361 14289 7364
rect 14323 7392 14335 7395
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 14323 7364 15485 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17770 7392 17776 7404
rect 17543 7364 17776 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 10836 7296 11100 7324
rect 10836 7284 10842 7296
rect 12158 7284 12164 7336
rect 12216 7284 12222 7336
rect 14090 7284 14096 7336
rect 14148 7284 14154 7336
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14240 7296 14473 7324
rect 14240 7284 14246 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 15286 7284 15292 7336
rect 15344 7284 15350 7336
rect 15488 7324 15516 7355
rect 17770 7352 17776 7364
rect 17828 7352 17834 7404
rect 17880 7324 17908 7432
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 18046 7352 18052 7404
rect 18104 7392 18110 7404
rect 22204 7401 22232 7500
rect 22756 7500 23428 7528
rect 22756 7401 22784 7500
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18104 7364 18613 7392
rect 18104 7352 18110 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7361 19303 7395
rect 22189 7395 22247 7401
rect 19245 7355 19303 7361
rect 15488 7296 17908 7324
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18874 7324 18880 7336
rect 18196 7296 18880 7324
rect 18196 7284 18202 7296
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 5460 7228 7328 7256
rect 9324 7228 13676 7256
rect 7006 7188 7012 7200
rect 5368 7160 7012 7188
rect 4801 7151 4859 7157
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7190 7148 7196 7200
rect 7248 7148 7254 7200
rect 7300 7188 7328 7228
rect 9950 7188 9956 7200
rect 7300 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 10502 7188 10508 7200
rect 10367 7160 10508 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10873 7191 10931 7197
rect 10873 7157 10885 7191
rect 10919 7188 10931 7191
rect 12434 7188 12440 7200
rect 10919 7160 12440 7188
rect 10919 7157 10931 7160
rect 10873 7151 10931 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12526 7148 12532 7200
rect 12584 7148 12590 7200
rect 13648 7188 13676 7228
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 17589 7259 17647 7265
rect 14332 7228 17540 7256
rect 14332 7216 14338 7228
rect 15286 7188 15292 7200
rect 13648 7160 15292 7188
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15654 7148 15660 7200
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15804 7160 15945 7188
rect 15804 7148 15810 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 17276 7160 17417 7188
rect 17276 7148 17282 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17512 7188 17540 7228
rect 17589 7225 17601 7259
rect 17635 7256 17647 7259
rect 17862 7256 17868 7268
rect 17635 7228 17868 7256
rect 17635 7225 17647 7228
rect 17589 7219 17647 7225
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 17954 7216 17960 7268
rect 18012 7216 18018 7268
rect 18049 7259 18107 7265
rect 18049 7225 18061 7259
rect 18095 7256 18107 7259
rect 18230 7256 18236 7268
rect 18095 7228 18236 7256
rect 18095 7225 18107 7228
rect 18049 7219 18107 7225
rect 18230 7216 18236 7228
rect 18288 7216 18294 7268
rect 18785 7259 18843 7265
rect 18785 7256 18797 7259
rect 18340 7228 18797 7256
rect 18340 7188 18368 7228
rect 18785 7225 18797 7228
rect 18831 7256 18843 7259
rect 19260 7256 19288 7355
rect 19794 7284 19800 7336
rect 19852 7284 19858 7336
rect 20070 7284 20076 7336
rect 20128 7284 20134 7336
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21192 7324 21220 7378
rect 22189 7361 22201 7395
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 20864 7296 21925 7324
rect 20864 7284 20870 7296
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 22204 7324 22232 7355
rect 23290 7352 23296 7404
rect 23348 7352 23354 7404
rect 23400 7392 23428 7500
rect 26694 7488 26700 7540
rect 26752 7488 26758 7540
rect 26970 7488 26976 7540
rect 27028 7488 27034 7540
rect 27430 7488 27436 7540
rect 27488 7488 27494 7540
rect 23474 7420 23480 7472
rect 23532 7460 23538 7472
rect 23532 7432 24256 7460
rect 23532 7420 23538 7432
rect 23842 7392 23848 7404
rect 23400 7364 23848 7392
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 24026 7392 24032 7404
rect 23983 7364 24032 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 24026 7352 24032 7364
rect 24084 7352 24090 7404
rect 24228 7401 24256 7432
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 25222 7352 25228 7404
rect 25280 7392 25286 7404
rect 26237 7395 26295 7401
rect 26237 7392 26249 7395
rect 25280 7364 26249 7392
rect 25280 7352 25286 7364
rect 26237 7361 26249 7364
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 26510 7352 26516 7404
rect 26568 7352 26574 7404
rect 27154 7352 27160 7404
rect 27212 7352 27218 7404
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 25130 7324 25136 7336
rect 22204 7296 25136 7324
rect 21913 7287 21971 7293
rect 25130 7284 25136 7296
rect 25188 7284 25194 7336
rect 25682 7284 25688 7336
rect 25740 7284 25746 7336
rect 25961 7327 26019 7333
rect 25961 7293 25973 7327
rect 26007 7324 26019 7327
rect 26142 7324 26148 7336
rect 26007 7296 26148 7324
rect 26007 7293 26019 7296
rect 25961 7287 26019 7293
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 26326 7284 26332 7336
rect 26384 7324 26390 7336
rect 27264 7324 27292 7355
rect 26384 7296 27292 7324
rect 26384 7284 26390 7296
rect 18831 7228 19288 7256
rect 18831 7225 18843 7228
rect 18785 7219 18843 7225
rect 23474 7216 23480 7268
rect 23532 7256 23538 7268
rect 23569 7259 23627 7265
rect 23569 7256 23581 7259
rect 23532 7228 23581 7256
rect 23532 7216 23538 7228
rect 23569 7225 23581 7228
rect 23615 7225 23627 7259
rect 23569 7219 23627 7225
rect 23842 7216 23848 7268
rect 23900 7256 23906 7268
rect 25222 7256 25228 7268
rect 23900 7228 25228 7256
rect 23900 7216 23906 7228
rect 25222 7216 25228 7228
rect 25280 7216 25286 7268
rect 17512 7160 18368 7188
rect 17405 7151 17463 7157
rect 18414 7148 18420 7200
rect 18472 7148 18478 7200
rect 21082 7148 21088 7200
rect 21140 7188 21146 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 21140 7160 21557 7188
rect 21140 7148 21146 7160
rect 21545 7157 21557 7160
rect 21591 7157 21603 7191
rect 21545 7151 21603 7157
rect 22649 7191 22707 7197
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 22922 7188 22928 7200
rect 22695 7160 22928 7188
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 22922 7148 22928 7160
rect 22980 7148 22986 7200
rect 23106 7148 23112 7200
rect 23164 7148 23170 7200
rect 23934 7148 23940 7200
rect 23992 7188 23998 7200
rect 24029 7191 24087 7197
rect 24029 7188 24041 7191
rect 23992 7160 24041 7188
rect 23992 7148 23998 7160
rect 24029 7157 24041 7160
rect 24075 7157 24087 7191
rect 24029 7151 24087 7157
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 1104 7098 27876 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 27876 7098
rect 1104 7024 27876 7046
rect 1486 6944 1492 6996
rect 1544 6944 1550 6996
rect 1854 6944 1860 6996
rect 1912 6944 1918 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4304 6956 5488 6984
rect 4304 6944 4310 6956
rect 2682 6916 2688 6928
rect 2056 6888 2688 6916
rect 2056 6848 2084 6888
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 5460 6916 5488 6956
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 5592 6956 6469 6984
rect 5592 6944 5598 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 6457 6947 6515 6953
rect 6996 6987 7054 6993
rect 6996 6953 7008 6987
rect 7042 6984 7054 6987
rect 7190 6984 7196 6996
rect 7042 6956 7196 6984
rect 7042 6953 7054 6956
rect 6996 6947 7054 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 9030 6984 9036 6996
rect 7432 6956 9036 6984
rect 7432 6944 7438 6956
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9204 6987 9262 6993
rect 9204 6953 9216 6987
rect 9250 6984 9262 6987
rect 9306 6984 9312 6996
rect 9250 6956 9312 6984
rect 9250 6953 9262 6956
rect 9204 6947 9262 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10502 6984 10508 6996
rect 9732 6956 10508 6984
rect 9732 6944 9738 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 10778 6944 10784 6996
rect 10836 6944 10842 6996
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 11146 6984 11152 6996
rect 10928 6956 11152 6984
rect 10928 6944 10934 6956
rect 11146 6944 11152 6956
rect 11204 6984 11210 6996
rect 11204 6956 13216 6984
rect 11204 6944 11210 6956
rect 5810 6916 5816 6928
rect 5460 6888 5816 6916
rect 5810 6876 5816 6888
rect 5868 6916 5874 6928
rect 5868 6888 6868 6916
rect 5868 6876 5874 6888
rect 1688 6820 2084 6848
rect 1688 6789 1716 6820
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 2188 6820 4169 6848
rect 2188 6808 2194 6820
rect 4157 6817 4169 6820
rect 4203 6848 4215 6851
rect 5626 6848 5632 6860
rect 4203 6820 5632 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 5626 6808 5632 6820
rect 5684 6848 5690 6860
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 5684 6820 6745 6848
rect 5684 6808 5690 6820
rect 6733 6817 6745 6820
rect 6779 6817 6791 6851
rect 6840 6848 6868 6888
rect 8941 6851 8999 6857
rect 6840 6820 8248 6848
rect 6733 6811 6791 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2222 6780 2228 6792
rect 2087 6752 2228 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 6144 6752 6285 6780
rect 6144 6740 6150 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6427 6783 6485 6789
rect 6427 6749 6439 6783
rect 6473 6780 6485 6783
rect 6546 6780 6552 6792
rect 6473 6752 6552 6780
rect 6473 6749 6485 6752
rect 6427 6743 6485 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 4430 6672 4436 6724
rect 4488 6672 4494 6724
rect 5810 6712 5816 6724
rect 5658 6684 5816 6712
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6681 6239 6715
rect 8220 6712 8248 6820
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 8987 6820 11192 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 10502 6780 10508 6792
rect 10350 6752 10508 6780
rect 10502 6740 10508 6752
rect 10560 6780 10566 6792
rect 11054 6780 11060 6792
rect 10560 6752 11060 6780
rect 10560 6740 10566 6752
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11164 6780 11192 6820
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 11388 6820 11437 6848
rect 11388 6808 11394 6820
rect 11425 6817 11437 6820
rect 11471 6848 11483 6851
rect 12710 6848 12716 6860
rect 11471 6820 12716 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 11698 6780 11704 6792
rect 11164 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 9674 6712 9680 6724
rect 8220 6698 9680 6712
rect 8234 6684 9680 6698
rect 6181 6675 6239 6681
rect 1210 6604 1216 6656
rect 1268 6644 1274 6656
rect 2225 6647 2283 6653
rect 2225 6644 2237 6647
rect 1268 6616 2237 6644
rect 1268 6604 1274 6616
rect 2225 6613 2237 6616
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 5718 6644 5724 6656
rect 3651 6616 5724 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6196 6644 6224 6675
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 11149 6715 11207 6721
rect 10520 6684 10824 6712
rect 6270 6644 6276 6656
rect 6196 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8352 6616 8493 6644
rect 8352 6604 8358 6616
rect 8481 6613 8493 6616
rect 8527 6644 8539 6647
rect 10520 6644 10548 6684
rect 8527 6616 10548 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10652 6616 10701 6644
rect 10652 6604 10658 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10796 6644 10824 6684
rect 11149 6681 11161 6715
rect 11195 6712 11207 6715
rect 11195 6684 11928 6712
rect 11195 6681 11207 6684
rect 11149 6675 11207 6681
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 10796 6616 11253 6644
rect 10689 6607 10747 6613
rect 11241 6613 11253 6616
rect 11287 6613 11299 6647
rect 11900 6644 11928 6684
rect 11974 6672 11980 6724
rect 12032 6672 12038 6724
rect 13188 6712 13216 6956
rect 14182 6944 14188 6996
rect 14240 6944 14246 6996
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 15669 6987 15727 6993
rect 15669 6984 15681 6987
rect 14608 6956 15681 6984
rect 14608 6944 14614 6956
rect 15669 6953 15681 6956
rect 15715 6953 15727 6987
rect 15669 6947 15727 6953
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 18233 6987 18291 6993
rect 18233 6953 18245 6987
rect 18279 6984 18291 6987
rect 18279 6956 18736 6984
rect 18279 6953 18291 6956
rect 18233 6947 18291 6953
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13320 6820 13737 6848
rect 13320 6808 13326 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 17788 6848 17816 6944
rect 18322 6876 18328 6928
rect 18380 6876 18386 6928
rect 18598 6848 18604 6860
rect 15620 6820 17540 6848
rect 17788 6820 18604 6848
rect 15620 6808 15626 6820
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13633 6783 13691 6789
rect 13633 6780 13645 6783
rect 13412 6752 13645 6780
rect 13412 6740 13418 6752
rect 13633 6749 13645 6752
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17512 6780 17540 6820
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18708 6848 18736 6956
rect 20070 6944 20076 6996
rect 20128 6984 20134 6996
rect 20533 6987 20591 6993
rect 20533 6984 20545 6987
rect 20128 6956 20545 6984
rect 20128 6944 20134 6956
rect 20533 6953 20545 6956
rect 20579 6953 20591 6987
rect 20533 6947 20591 6953
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 26326 6984 26332 6996
rect 22704 6956 26332 6984
rect 22704 6944 22710 6956
rect 26326 6944 26332 6956
rect 26384 6944 26390 6996
rect 18874 6876 18880 6928
rect 18932 6916 18938 6928
rect 18932 6888 19380 6916
rect 18932 6876 18938 6888
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 18708 6820 18797 6848
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 18969 6851 19027 6857
rect 18969 6817 18981 6851
rect 19015 6848 19027 6851
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19015 6820 19257 6848
rect 19015 6817 19027 6820
rect 18969 6811 19027 6817
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19352 6848 19380 6888
rect 19352 6820 19840 6848
rect 19245 6811 19303 6817
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17512 6752 17877 6780
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18506 6780 18512 6792
rect 18095 6752 18512 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 14274 6712 14280 6724
rect 13188 6698 14280 6712
rect 13202 6684 14280 6698
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 15378 6712 15384 6724
rect 15226 6684 15384 6712
rect 15378 6672 15384 6684
rect 15436 6712 15442 6724
rect 15436 6684 16252 6712
rect 15436 6672 15442 6684
rect 12802 6644 12808 6656
rect 11900 6616 12808 6644
rect 11241 6607 11299 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 13449 6647 13507 6653
rect 13449 6644 13461 6647
rect 13412 6616 13461 6644
rect 13412 6604 13418 6616
rect 13449 6613 13461 6616
rect 13495 6613 13507 6647
rect 16224 6644 16252 6684
rect 16298 6672 16304 6724
rect 16356 6672 16362 6724
rect 17880 6712 17908 6743
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18690 6740 18696 6792
rect 18748 6740 18754 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19610 6780 19616 6792
rect 19475 6752 19616 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 19702 6740 19708 6792
rect 19760 6740 19766 6792
rect 19812 6780 19840 6820
rect 21174 6808 21180 6860
rect 21232 6808 21238 6860
rect 21818 6808 21824 6860
rect 21876 6808 21882 6860
rect 22370 6808 22376 6860
rect 22428 6808 22434 6860
rect 22738 6808 22744 6860
rect 22796 6848 22802 6860
rect 23842 6848 23848 6860
rect 22796 6820 23848 6848
rect 22796 6808 22802 6820
rect 20070 6780 20076 6792
rect 19812 6752 20076 6780
rect 20070 6740 20076 6752
rect 20128 6780 20134 6792
rect 23308 6789 23336 6820
rect 23842 6808 23848 6820
rect 23900 6808 23906 6860
rect 24670 6808 24676 6860
rect 24728 6848 24734 6860
rect 27614 6848 27620 6860
rect 24728 6820 26740 6848
rect 24728 6808 24734 6820
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 20128 6752 21557 6780
rect 20128 6740 20134 6752
rect 21545 6749 21557 6752
rect 21591 6780 21603 6783
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 21591 6752 22661 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 23292 6783 23350 6789
rect 23292 6749 23304 6783
rect 23338 6749 23350 6783
rect 23292 6743 23350 6749
rect 23385 6783 23443 6789
rect 23385 6749 23397 6783
rect 23431 6749 23443 6783
rect 23385 6743 23443 6749
rect 17526 6684 17816 6712
rect 17880 6684 18092 6712
rect 17788 6644 17816 6684
rect 17954 6644 17960 6656
rect 16224 6616 17960 6644
rect 13449 6607 13507 6613
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 18064 6644 18092 6684
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 19797 6715 19855 6721
rect 19797 6712 19809 6715
rect 19208 6684 19809 6712
rect 19208 6672 19214 6684
rect 19797 6681 19809 6684
rect 19843 6681 19855 6715
rect 19797 6675 19855 6681
rect 19978 6672 19984 6724
rect 20036 6672 20042 6724
rect 21637 6715 21695 6721
rect 21637 6681 21649 6715
rect 21683 6712 21695 6715
rect 22370 6712 22376 6724
rect 21683 6684 22376 6712
rect 21683 6681 21695 6684
rect 21637 6675 21695 6681
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 22664 6712 22692 6743
rect 22922 6712 22928 6724
rect 22664 6684 22928 6712
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 23106 6672 23112 6724
rect 23164 6712 23170 6724
rect 23400 6712 23428 6743
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 23934 6740 23940 6792
rect 23992 6740 23998 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 23164 6684 23428 6712
rect 23164 6672 23170 6684
rect 19334 6644 19340 6656
rect 18064 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19518 6604 19524 6656
rect 19576 6644 19582 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19576 6616 19625 6644
rect 19576 6604 19582 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 20898 6604 20904 6656
rect 20956 6604 20962 6656
rect 20990 6604 20996 6656
rect 21048 6604 21054 6656
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22612 6616 23029 6644
rect 22612 6604 22618 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 23569 6647 23627 6653
rect 23569 6644 23581 6647
rect 23440 6616 23581 6644
rect 23440 6604 23446 6616
rect 23569 6613 23581 6616
rect 23615 6613 23627 6647
rect 24044 6644 24072 6743
rect 24394 6740 24400 6792
rect 24452 6740 24458 6792
rect 26510 6740 26516 6792
rect 26568 6740 26574 6792
rect 24673 6715 24731 6721
rect 24673 6681 24685 6715
rect 24719 6712 24731 6715
rect 24946 6712 24952 6724
rect 24719 6684 24952 6712
rect 24719 6681 24731 6684
rect 24673 6675 24731 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 25130 6672 25136 6724
rect 25188 6672 25194 6724
rect 25958 6672 25964 6724
rect 26016 6712 26022 6724
rect 26712 6712 26740 6820
rect 26804 6820 27620 6848
rect 26804 6789 26832 6820
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 26878 6740 26884 6792
rect 26936 6740 26942 6792
rect 27249 6783 27307 6789
rect 27249 6749 27261 6783
rect 27295 6749 27307 6783
rect 27249 6743 27307 6749
rect 27264 6712 27292 6743
rect 26016 6684 26648 6712
rect 26712 6684 27292 6712
rect 26016 6672 26022 6684
rect 25498 6644 25504 6656
rect 24044 6616 25504 6644
rect 23569 6607 23627 6613
rect 25498 6604 25504 6616
rect 25556 6604 25562 6656
rect 26142 6604 26148 6656
rect 26200 6604 26206 6656
rect 26326 6604 26332 6656
rect 26384 6604 26390 6656
rect 26620 6653 26648 6684
rect 26605 6647 26663 6653
rect 26605 6613 26617 6647
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 27062 6604 27068 6656
rect 27120 6604 27126 6656
rect 27433 6647 27491 6653
rect 27433 6613 27445 6647
rect 27479 6644 27491 6647
rect 27522 6644 27528 6656
rect 27479 6616 27528 6644
rect 27479 6613 27491 6616
rect 27433 6607 27491 6613
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 1104 6554 27876 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 27876 6554
rect 1104 6480 27876 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 1360 6412 1501 6440
rect 1360 6400 1366 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 1489 6403 1547 6409
rect 1964 6412 4384 6440
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1964 6304 1992 6412
rect 4246 6372 4252 6384
rect 3634 6344 4252 6372
rect 1719 6276 1992 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 2130 6264 2136 6316
rect 2188 6264 2194 6316
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 3786 6236 3792 6248
rect 2455 6208 3792 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 1234 6128 1240 6180
rect 1292 6168 1298 6180
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1292 6140 1869 6168
rect 1292 6128 1298 6140
rect 1857 6137 1869 6140
rect 1903 6137 1915 6171
rect 1857 6131 1915 6137
rect 3602 6128 3608 6180
rect 3660 6168 3666 6180
rect 3896 6168 3924 6344
rect 4246 6332 4252 6344
rect 4304 6332 4310 6384
rect 4356 6372 4384 6412
rect 4430 6400 4436 6452
rect 4488 6440 4494 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4488 6412 4629 6440
rect 4488 6400 4494 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 5718 6440 5724 6452
rect 5040 6412 5724 6440
rect 5040 6400 5046 6412
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7708 6412 7941 6440
rect 7708 6400 7714 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8168 6412 8800 6440
rect 8168 6400 8174 6412
rect 5534 6372 5540 6384
rect 4356 6344 5540 6372
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6372 7803 6375
rect 8662 6372 8668 6384
rect 7791 6344 8668 6372
rect 7791 6341 7803 6344
rect 7745 6335 7803 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 8772 6372 8800 6412
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 9674 6440 9680 6452
rect 9646 6400 9680 6440
rect 9732 6400 9738 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10652 6412 10701 6440
rect 10652 6400 10658 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 10689 6403 10747 6409
rect 10778 6400 10784 6452
rect 10836 6400 10842 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11238 6440 11244 6452
rect 11195 6412 11244 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12032 6412 12173 6440
rect 12032 6400 12038 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12621 6443 12679 6449
rect 12621 6440 12633 6443
rect 12584 6412 12633 6440
rect 12584 6400 12590 6412
rect 12621 6409 12633 6412
rect 12667 6409 12679 6443
rect 12621 6403 12679 6409
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 14148 6412 14197 6440
rect 14148 6400 14154 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 14550 6400 14556 6452
rect 14608 6400 14614 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 15378 6440 15384 6452
rect 14884 6412 15384 6440
rect 14884 6400 14890 6412
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 15712 6412 15761 6440
rect 15712 6400 15718 6412
rect 15749 6409 15761 6412
rect 15795 6409 15807 6443
rect 15749 6403 15807 6409
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 16298 6440 16304 6452
rect 16163 6412 16304 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 18046 6440 18052 6452
rect 17880 6412 18052 6440
rect 9646 6372 9674 6400
rect 8772 6344 9674 6372
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10502 6372 10508 6384
rect 9824 6344 10508 6372
rect 9824 6332 9830 6344
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5408 6276 5641 6304
rect 5408 6264 5414 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 8110 6304 8116 6316
rect 6104 6276 8116 6304
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4798 6236 4804 6248
rect 4203 6208 4804 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5307 6208 5457 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 3660 6140 3924 6168
rect 3660 6128 3666 6140
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 5092 6168 5120 6199
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5592 6208 5733 6236
rect 5592 6196 5598 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 6104 6236 6132 6276
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8536 6276 8585 6304
rect 8536 6264 8542 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 5868 6208 6132 6236
rect 5868 6196 5874 6208
rect 6362 6196 6368 6248
rect 6420 6236 6426 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6420 6208 6469 6236
rect 6420 6196 6426 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 6730 6196 6736 6248
rect 6788 6196 6794 6248
rect 9232 6236 9260 6267
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 10336 6313 10364 6344
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 11514 6372 11520 6384
rect 10560 6344 11520 6372
rect 10560 6332 10566 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 13354 6372 13360 6384
rect 12308 6344 13360 6372
rect 12308 6332 12314 6344
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9456 6276 9689 6304
rect 9456 6264 9462 6276
rect 9677 6273 9689 6276
rect 9723 6304 9735 6307
rect 10321 6307 10379 6313
rect 9723 6276 10272 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9306 6236 9312 6248
rect 9232 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9548 6208 9781 6236
rect 9548 6196 9554 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 10244 6236 10272 6276
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 11882 6304 11888 6316
rect 10321 6267 10379 6273
rect 10428 6276 11888 6304
rect 10428 6236 10456 6276
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 11940 6276 12541 6304
rect 11940 6264 11946 6276
rect 12529 6273 12541 6276
rect 12575 6304 12587 6307
rect 12989 6307 13047 6313
rect 12575 6276 12940 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 10244 6208 10456 6236
rect 10502 6196 10508 6248
rect 10560 6196 10566 6248
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 12342 6236 12348 6248
rect 11020 6208 12348 6236
rect 11020 6196 11026 6208
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6205 12863 6239
rect 12912 6236 12940 6276
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13078 6304 13084 6316
rect 13035 6276 13084 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13170 6264 13176 6316
rect 13228 6264 13234 6316
rect 13280 6304 13308 6344
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 13556 6344 15700 6372
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 13280 6276 13461 6304
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13556 6236 13584 6344
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 14734 6264 14740 6316
rect 14792 6264 14798 6316
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6304 15255 6307
rect 15286 6304 15292 6316
rect 15243 6276 15292 6304
rect 15243 6273 15255 6276
rect 15197 6267 15255 6273
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 15672 6313 15700 6344
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 16761 6375 16819 6381
rect 16761 6372 16773 6375
rect 16632 6344 16773 6372
rect 16632 6332 16638 6344
rect 16761 6341 16773 6344
rect 16807 6341 16819 6375
rect 17678 6372 17684 6384
rect 16761 6335 16819 6341
rect 17236 6344 17684 6372
rect 17236 6316 17264 6344
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 17770 6332 17776 6384
rect 17828 6332 17834 6384
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 15746 6304 15752 6316
rect 15703 6276 15752 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 15896 6276 16221 6304
rect 15896 6264 15902 6276
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16482 6304 16488 6316
rect 16439 6276 16488 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 17880 6304 17908 6412
rect 18046 6400 18052 6412
rect 18104 6440 18110 6452
rect 19150 6440 19156 6452
rect 18104 6412 19156 6440
rect 18104 6400 18110 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19797 6443 19855 6449
rect 19797 6440 19809 6443
rect 19392 6412 19809 6440
rect 19392 6400 19398 6412
rect 19797 6409 19809 6412
rect 19843 6440 19855 6443
rect 20254 6440 20260 6452
rect 19843 6412 20260 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 22741 6443 22799 6449
rect 22741 6440 22753 6443
rect 21232 6412 22753 6440
rect 21232 6400 21238 6412
rect 22741 6409 22753 6412
rect 22787 6409 22799 6443
rect 23290 6440 23296 6452
rect 22741 6403 22799 6409
rect 23032 6412 23296 6440
rect 18322 6332 18328 6384
rect 18380 6332 18386 6384
rect 22830 6372 22836 6384
rect 22480 6344 22836 6372
rect 17543 6276 17908 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 19426 6264 19432 6316
rect 19484 6264 19490 6316
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 19978 6304 19984 6316
rect 19935 6276 19984 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 22480 6304 22508 6344
rect 22830 6332 22836 6344
rect 22888 6332 22894 6384
rect 22428 6276 22508 6304
rect 22428 6264 22434 6276
rect 22554 6264 22560 6316
rect 22612 6264 22618 6316
rect 23032 6313 23060 6412
rect 23290 6400 23296 6412
rect 23348 6440 23354 6452
rect 24854 6440 24860 6452
rect 23348 6412 24860 6440
rect 23348 6400 23354 6412
rect 24854 6400 24860 6412
rect 24912 6400 24918 6452
rect 24946 6400 24952 6452
rect 25004 6400 25010 6452
rect 25409 6443 25467 6449
rect 25409 6409 25421 6443
rect 25455 6440 25467 6443
rect 26050 6440 26056 6452
rect 25455 6412 26056 6440
rect 25455 6409 25467 6412
rect 25409 6403 25467 6409
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 27430 6400 27436 6452
rect 27488 6400 27494 6452
rect 23382 6332 23388 6384
rect 23440 6332 23446 6384
rect 24118 6332 24124 6384
rect 24176 6332 24182 6384
rect 25317 6375 25375 6381
rect 25317 6341 25329 6375
rect 25363 6372 25375 6375
rect 26326 6372 26332 6384
rect 25363 6344 26332 6372
rect 25363 6341 25375 6344
rect 25317 6335 25375 6341
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 12912 6208 13584 6236
rect 12805 6199 12863 6205
rect 6270 6168 6276 6180
rect 4764 6140 6276 6168
rect 4764 6128 4770 6140
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 7484 6140 9353 6168
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 7484 6100 7512 6140
rect 6236 6072 7512 6100
rect 7653 6103 7711 6109
rect 6236 6060 6242 6072
rect 7653 6069 7665 6103
rect 7699 6100 7711 6103
rect 7834 6100 7840 6112
rect 7699 6072 7840 6100
rect 7699 6069 7711 6072
rect 7653 6063 7711 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 8628 6072 8677 6100
rect 8628 6060 8634 6072
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 8665 6063 8723 6069
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8996 6072 9045 6100
rect 8996 6060 9002 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9325 6100 9353 6140
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9456 6140 10241 6168
rect 9456 6128 9462 6140
rect 10229 6137 10241 6140
rect 10275 6168 10287 6171
rect 12710 6168 12716 6180
rect 10275 6140 12716 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 12820 6168 12848 6199
rect 13998 6196 14004 6248
rect 14056 6196 14062 6248
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 15562 6196 15568 6248
rect 15620 6196 15626 6248
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 16080 6208 18061 6236
rect 16080 6196 16086 6208
rect 14366 6168 14372 6180
rect 12820 6140 14372 6168
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 16114 6168 16120 6180
rect 14608 6140 16120 6168
rect 14608 6128 14614 6140
rect 16114 6128 16120 6140
rect 16172 6128 16178 6180
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16669 6171 16727 6177
rect 16669 6168 16681 6171
rect 16347 6140 16681 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16669 6137 16681 6140
rect 16715 6137 16727 6171
rect 16669 6131 16727 6137
rect 12158 6100 12164 6112
rect 9325 6072 12164 6100
rect 9033 6063 9091 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 12400 6072 13093 6100
rect 12400 6060 12406 6072
rect 13081 6069 13093 6072
rect 13127 6069 13139 6103
rect 13081 6063 13139 6069
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14792 6072 14841 6100
rect 14792 6060 14798 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 14976 6072 15117 6100
rect 14976 6060 14982 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 15654 6100 15660 6112
rect 15344 6072 15660 6100
rect 15344 6060 15350 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 17126 6100 17132 6112
rect 16540 6072 17132 6100
rect 16540 6060 16546 6072
rect 17126 6060 17132 6072
rect 17184 6100 17190 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 17184 6072 17693 6100
rect 17184 6060 17190 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17880 6100 17908 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 19444 6236 19472 6264
rect 18049 6199 18107 6205
rect 18156 6208 19472 6236
rect 21637 6239 21695 6245
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18156 6168 18184 6208
rect 21637 6205 21649 6239
rect 21683 6205 21695 6239
rect 21637 6199 21695 6205
rect 18012 6140 18184 6168
rect 18012 6128 18018 6140
rect 19886 6128 19892 6180
rect 19944 6168 19950 6180
rect 21652 6168 21680 6199
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 22281 6239 22339 6245
rect 22281 6236 22293 6239
rect 21876 6208 22293 6236
rect 21876 6196 21882 6208
rect 22281 6205 22293 6208
rect 22327 6205 22339 6239
rect 22281 6199 22339 6205
rect 22462 6196 22468 6248
rect 22520 6196 22526 6248
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6205 23167 6239
rect 23109 6199 23167 6205
rect 23124 6168 23152 6199
rect 23842 6196 23848 6248
rect 23900 6236 23906 6248
rect 25332 6236 25360 6335
rect 26326 6332 26332 6344
rect 26384 6332 26390 6384
rect 25406 6264 25412 6316
rect 25464 6304 25470 6316
rect 26513 6307 26571 6313
rect 26513 6304 26525 6307
rect 25464 6276 26525 6304
rect 25464 6264 25470 6276
rect 26513 6273 26525 6276
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 27246 6264 27252 6316
rect 27304 6264 27310 6316
rect 23900 6208 25360 6236
rect 23900 6196 23906 6208
rect 25498 6196 25504 6248
rect 25556 6236 25562 6248
rect 26326 6236 26332 6248
rect 25556 6208 26332 6236
rect 25556 6196 25562 6208
rect 26326 6196 26332 6208
rect 26384 6196 26390 6248
rect 19944 6140 23152 6168
rect 19944 6128 19950 6140
rect 19904 6100 19932 6128
rect 17880 6072 19932 6100
rect 21913 6103 21971 6109
rect 17681 6063 17739 6069
rect 21913 6069 21925 6103
rect 21959 6100 21971 6103
rect 22186 6100 22192 6112
rect 21959 6072 22192 6100
rect 21959 6069 21971 6072
rect 21913 6063 21971 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22278 6060 22284 6112
rect 22336 6100 22342 6112
rect 22925 6103 22983 6109
rect 22925 6100 22937 6103
rect 22336 6072 22937 6100
rect 22336 6060 22342 6072
rect 22925 6069 22937 6072
rect 22971 6069 22983 6103
rect 23124 6100 23152 6140
rect 24394 6100 24400 6112
rect 23124 6072 24400 6100
rect 22925 6063 22983 6069
rect 24394 6060 24400 6072
rect 24452 6060 24458 6112
rect 24857 6103 24915 6109
rect 24857 6069 24869 6103
rect 24903 6100 24915 6103
rect 25222 6100 25228 6112
rect 24903 6072 25228 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 25222 6060 25228 6072
rect 25280 6060 25286 6112
rect 26694 6060 26700 6112
rect 26752 6060 26758 6112
rect 1104 6010 27876 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 27876 6010
rect 1104 5936 27876 5958
rect 3786 5856 3792 5908
rect 3844 5856 3850 5908
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 5350 5896 5356 5908
rect 4488 5868 5356 5896
rect 4488 5856 4494 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5500 5868 5733 5896
rect 5500 5856 5506 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 5721 5859 5779 5865
rect 5810 5856 5816 5908
rect 5868 5896 5874 5908
rect 5868 5868 6040 5896
rect 5868 5856 5874 5868
rect 1166 5788 1172 5840
rect 1224 5828 1230 5840
rect 1489 5831 1547 5837
rect 1489 5828 1501 5831
rect 1224 5800 1501 5828
rect 1224 5788 1230 5800
rect 1489 5797 1501 5800
rect 1535 5797 1547 5831
rect 1489 5791 1547 5797
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 3878 5828 3884 5840
rect 3191 5800 3884 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 4982 5828 4988 5840
rect 4172 5800 4988 5828
rect 4062 5760 4068 5772
rect 3344 5732 4068 5760
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2866 5692 2872 5704
rect 2087 5664 2872 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 3344 5701 3372 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 3292 5664 3341 5692
rect 3292 5652 3298 5664
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 3970 5692 3976 5704
rect 3559 5664 3976 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 1854 5516 1860 5568
rect 1912 5516 1918 5568
rect 3436 5556 3464 5655
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4172 5701 4200 5800
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 5902 5828 5908 5840
rect 5092 5800 5908 5828
rect 5092 5769 5120 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 6012 5828 6040 5868
rect 6086 5856 6092 5908
rect 6144 5856 6150 5908
rect 7193 5899 7251 5905
rect 7193 5865 7205 5899
rect 7239 5896 7251 5899
rect 7742 5896 7748 5908
rect 7239 5868 7748 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7852 5868 7941 5896
rect 6914 5828 6920 5840
rect 6012 5800 6920 5828
rect 6914 5788 6920 5800
rect 6972 5828 6978 5840
rect 7282 5828 7288 5840
rect 6972 5800 7288 5828
rect 6972 5788 6978 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4479 5732 4629 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4617 5723 4675 5729
rect 4724 5732 4905 5760
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4724 5692 4752 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 5077 5723 5135 5729
rect 5460 5732 6653 5760
rect 5460 5704 5488 5732
rect 6012 5704 6040 5732
rect 6641 5729 6653 5732
rect 6687 5760 6699 5763
rect 6730 5760 6736 5772
rect 6687 5732 6736 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7852 5760 7880 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8812 5868 8953 5896
rect 8812 5856 8818 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 9088 5868 9321 5896
rect 9088 5856 9094 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 9490 5856 9496 5908
rect 9548 5856 9554 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 12066 5896 12072 5908
rect 9640 5868 12072 5896
rect 9640 5856 9646 5868
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 12618 5896 12624 5908
rect 12575 5868 12624 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 13446 5896 13452 5908
rect 12768 5868 13452 5896
rect 12768 5856 12774 5868
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 13814 5896 13820 5908
rect 13679 5868 13820 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14056 5868 14289 5896
rect 14056 5856 14062 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15620 5868 15761 5896
rect 15620 5856 15626 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 17000 5868 18153 5896
rect 17000 5856 17006 5868
rect 18141 5865 18153 5868
rect 18187 5865 18199 5899
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 18141 5859 18199 5865
rect 18432 5868 19349 5896
rect 10134 5828 10140 5840
rect 9876 5800 10140 5828
rect 8938 5760 8944 5772
rect 6840 5732 7880 5760
rect 7944 5732 8944 5760
rect 4580 5664 4752 5692
rect 4801 5695 4859 5701
rect 4580 5652 4586 5664
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5258 5692 5264 5704
rect 5031 5664 5264 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 4816 5624 4844 5655
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5350 5652 5356 5704
rect 5408 5652 5414 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 5718 5692 5724 5704
rect 5583 5664 5724 5692
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6840 5692 6868 5732
rect 7944 5704 7972 5732
rect 8938 5720 8944 5732
rect 8996 5760 9002 5772
rect 9876 5769 9904 5800
rect 10134 5788 10140 5800
rect 10192 5828 10198 5840
rect 10594 5828 10600 5840
rect 10192 5800 10600 5828
rect 10192 5788 10198 5800
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 13078 5828 13084 5840
rect 12912 5800 13084 5828
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8996 5732 9045 5760
rect 8996 5720 9002 5732
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 10962 5760 10968 5772
rect 9861 5723 9919 5729
rect 10520 5732 10968 5760
rect 6104 5664 6868 5692
rect 6917 5695 6975 5701
rect 3936 5596 4844 5624
rect 5736 5624 5764 5652
rect 6104 5624 6132 5664
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7190 5692 7196 5704
rect 6963 5664 7196 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 8260 5664 8309 5692
rect 8260 5652 8266 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 9140 5692 9168 5723
rect 8496 5664 9168 5692
rect 5736 5596 6132 5624
rect 3936 5584 3942 5596
rect 6178 5584 6184 5636
rect 6236 5624 6242 5636
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 6236 5596 6561 5624
rect 6236 5584 6242 5596
rect 6549 5593 6561 5596
rect 6595 5593 6607 5627
rect 6549 5587 6607 5593
rect 7009 5627 7067 5633
rect 7009 5593 7021 5627
rect 7055 5624 7067 5627
rect 8404 5624 8432 5652
rect 7055 5596 8432 5624
rect 7055 5593 7067 5596
rect 7009 5587 7067 5593
rect 4062 5556 4068 5568
rect 3436 5528 4068 5556
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4798 5556 4804 5568
rect 4295 5528 4804 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4798 5516 4804 5528
rect 4856 5556 4862 5568
rect 5810 5556 5816 5568
rect 4856 5528 5816 5556
rect 4856 5516 4862 5528
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 5997 5559 6055 5565
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6362 5556 6368 5568
rect 6043 5528 6368 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 6638 5556 6644 5568
rect 6503 5528 6644 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7607 5528 7757 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 8496 5556 8524 5664
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 10520 5692 10548 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11756 5732 11989 5760
rect 11756 5720 11762 5732
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 12342 5720 12348 5772
rect 12400 5720 12406 5772
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 12621 5763 12679 5769
rect 12483 5732 12572 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 9732 5664 10548 5692
rect 9732 5652 9738 5664
rect 11146 5584 11152 5636
rect 11204 5584 11210 5636
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 11701 5627 11759 5633
rect 11701 5624 11713 5627
rect 11664 5596 11713 5624
rect 11664 5584 11670 5596
rect 11701 5593 11713 5596
rect 11747 5593 11759 5627
rect 11701 5587 11759 5593
rect 7892 5528 8524 5556
rect 8573 5559 8631 5565
rect 7892 5516 7898 5528
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8662 5556 8668 5568
rect 8619 5528 8668 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 12544 5556 12572 5732
rect 12621 5729 12633 5763
rect 12667 5760 12679 5763
rect 12802 5760 12808 5772
rect 12667 5732 12808 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 12912 5692 12940 5800
rect 13078 5788 13084 5800
rect 13136 5788 13142 5840
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 13538 5828 13544 5840
rect 13228 5800 13544 5828
rect 13228 5788 13234 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 16482 5828 16488 5840
rect 15304 5800 16488 5828
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5760 13047 5763
rect 13035 5732 13676 5760
rect 13035 5729 13047 5732
rect 12989 5723 13047 5729
rect 12759 5664 12940 5692
rect 13081 5695 13139 5701
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13354 5692 13360 5704
rect 13311 5664 13360 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12544 5528 12817 5556
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13096 5556 13124 5655
rect 13188 5568 13216 5655
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 13648 5692 13676 5732
rect 13722 5720 13728 5772
rect 13780 5720 13786 5772
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 15304 5769 15332 5800
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 17405 5831 17463 5837
rect 17405 5797 17417 5831
rect 17451 5797 17463 5831
rect 17405 5791 17463 5797
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 15528 5732 15577 5760
rect 15528 5720 15534 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 17420 5760 17448 5791
rect 17494 5788 17500 5840
rect 17552 5828 17558 5840
rect 18046 5828 18052 5840
rect 17552 5800 18052 5828
rect 17552 5788 17558 5800
rect 18046 5788 18052 5800
rect 18104 5788 18110 5840
rect 18432 5828 18460 5868
rect 19337 5865 19349 5868
rect 19383 5865 19395 5899
rect 19337 5859 19395 5865
rect 19702 5856 19708 5908
rect 19760 5896 19766 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19760 5868 19809 5896
rect 19760 5856 19766 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 23474 5896 23480 5908
rect 19797 5859 19855 5865
rect 19996 5868 23480 5896
rect 18156 5800 18460 5828
rect 18156 5760 18184 5800
rect 15804 5732 16160 5760
rect 15804 5720 15810 5732
rect 14090 5692 14096 5704
rect 13648 5664 14096 5692
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15160 5664 15393 5692
rect 15160 5652 15166 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 15838 5692 15844 5704
rect 15703 5664 15844 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16022 5652 16028 5704
rect 16080 5652 16086 5704
rect 16132 5701 16160 5732
rect 16250 5732 16712 5760
rect 16250 5701 16278 5732
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16235 5695 16293 5701
rect 16235 5661 16247 5695
rect 16281 5661 16293 5695
rect 16235 5655 16293 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16574 5692 16580 5704
rect 16439 5664 16580 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16684 5692 16712 5732
rect 16960 5732 17448 5760
rect 17696 5732 18184 5760
rect 16960 5692 16988 5732
rect 16684 5664 16988 5692
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 17696 5692 17724 5732
rect 18322 5720 18328 5772
rect 18380 5720 18386 5772
rect 18432 5769 18460 5800
rect 18506 5788 18512 5840
rect 18564 5828 18570 5840
rect 19996 5828 20024 5868
rect 23474 5856 23480 5868
rect 23532 5896 23538 5908
rect 24302 5896 24308 5908
rect 23532 5868 24308 5896
rect 23532 5856 23538 5868
rect 24302 5856 24308 5868
rect 24360 5856 24366 5908
rect 27430 5856 27436 5908
rect 27488 5856 27494 5908
rect 18564 5800 20024 5828
rect 18564 5788 18570 5800
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 17420 5664 17724 5692
rect 17773 5695 17831 5701
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 14274 5624 14280 5636
rect 14056 5596 14280 5624
rect 14056 5584 14062 5596
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 14642 5584 14648 5636
rect 14700 5584 14706 5636
rect 16850 5633 16856 5636
rect 14783 5627 14841 5633
rect 14783 5593 14795 5627
rect 14829 5624 14841 5627
rect 16828 5627 16856 5633
rect 14829 5596 15792 5624
rect 14829 5593 14841 5596
rect 14783 5587 14841 5593
rect 13044 5528 13124 5556
rect 13044 5516 13050 5528
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 14182 5556 14188 5568
rect 13228 5528 14188 5556
rect 13228 5516 13234 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 15289 5559 15347 5565
rect 15289 5525 15301 5559
rect 15335 5556 15347 5559
rect 15562 5556 15568 5568
rect 15335 5528 15568 5556
rect 15335 5525 15347 5528
rect 15289 5519 15347 5525
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 15764 5556 15792 5596
rect 16828 5593 16840 5627
rect 16828 5587 16856 5593
rect 16850 5584 16856 5587
rect 16908 5584 16914 5636
rect 16945 5627 17003 5633
rect 16945 5593 16957 5627
rect 16991 5624 17003 5627
rect 17126 5624 17132 5636
rect 16991 5596 17132 5624
rect 16991 5593 17003 5596
rect 16945 5587 17003 5593
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 17218 5584 17224 5636
rect 17276 5624 17282 5636
rect 17420 5624 17448 5664
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 17862 5692 17868 5704
rect 17819 5664 17868 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18138 5692 18144 5704
rect 18095 5664 18144 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 18509 5695 18567 5701
rect 18509 5692 18521 5695
rect 18288 5664 18521 5692
rect 18288 5652 18294 5664
rect 18509 5661 18521 5664
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5692 18659 5695
rect 18782 5692 18788 5704
rect 18647 5664 18788 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 18892 5701 18920 5800
rect 23750 5788 23756 5840
rect 23808 5828 23814 5840
rect 24210 5828 24216 5840
rect 23808 5800 24216 5828
rect 23808 5788 23814 5800
rect 24210 5788 24216 5800
rect 24268 5828 24274 5840
rect 24268 5800 24532 5828
rect 24268 5788 24274 5800
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 19208 5732 19533 5760
rect 19208 5720 19214 5732
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 22465 5763 22523 5769
rect 19521 5723 19579 5729
rect 19628 5732 21956 5760
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19334 5692 19340 5704
rect 19291 5664 19340 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 17586 5633 17592 5636
rect 17276 5596 17448 5624
rect 17564 5627 17592 5633
rect 17276 5584 17282 5596
rect 17564 5593 17576 5627
rect 17564 5587 17592 5593
rect 17586 5584 17592 5587
rect 17644 5584 17650 5636
rect 19058 5584 19064 5636
rect 19116 5624 19122 5636
rect 19628 5624 19656 5732
rect 19886 5652 19892 5704
rect 19944 5652 19950 5704
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 21928 5701 21956 5732
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 24394 5760 24400 5772
rect 22511 5732 24400 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 24394 5720 24400 5732
rect 24452 5720 24458 5772
rect 24504 5760 24532 5800
rect 27062 5788 27068 5840
rect 27120 5788 27126 5840
rect 24673 5763 24731 5769
rect 24673 5760 24685 5763
rect 24504 5732 24685 5760
rect 24673 5729 24685 5732
rect 24719 5729 24731 5763
rect 24673 5723 24731 5729
rect 25038 5720 25044 5772
rect 25096 5760 25102 5772
rect 25096 5732 26924 5760
rect 25096 5720 25102 5732
rect 21729 5695 21787 5701
rect 21729 5692 21741 5695
rect 21692 5664 21741 5692
rect 21692 5652 21698 5664
rect 21729 5661 21741 5664
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 22005 5695 22063 5701
rect 22005 5661 22017 5695
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 19116 5596 19656 5624
rect 19116 5584 19122 5596
rect 20162 5584 20168 5636
rect 20220 5584 20226 5636
rect 21450 5624 21456 5636
rect 21390 5596 21456 5624
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 21560 5596 21772 5624
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 15764 5528 16681 5556
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 17034 5516 17040 5568
rect 17092 5516 17098 5568
rect 17144 5556 17172 5584
rect 17681 5559 17739 5565
rect 17681 5556 17693 5559
rect 17144 5528 17693 5556
rect 17681 5525 17693 5528
rect 17727 5556 17739 5559
rect 18230 5556 18236 5568
rect 17727 5528 18236 5556
rect 17727 5525 17739 5528
rect 17681 5519 17739 5525
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 19150 5516 19156 5568
rect 19208 5556 19214 5568
rect 19334 5556 19340 5568
rect 19208 5528 19340 5556
rect 19208 5516 19214 5528
rect 19334 5516 19340 5528
rect 19392 5556 19398 5568
rect 21560 5556 21588 5596
rect 19392 5528 21588 5556
rect 19392 5516 19398 5528
rect 21634 5516 21640 5568
rect 21692 5516 21698 5568
rect 21744 5556 21772 5596
rect 21818 5584 21824 5636
rect 21876 5624 21882 5636
rect 22020 5624 22048 5655
rect 22094 5652 22100 5704
rect 22152 5652 22158 5704
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26896 5701 26924 5732
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 26292 5664 26525 5692
rect 26292 5652 26298 5664
rect 26513 5661 26525 5664
rect 26559 5661 26571 5695
rect 26513 5655 26571 5661
rect 26881 5695 26939 5701
rect 26881 5661 26893 5695
rect 26927 5661 26939 5695
rect 26881 5655 26939 5661
rect 27246 5652 27252 5704
rect 27304 5652 27310 5704
rect 21876 5596 22048 5624
rect 22112 5624 22140 5652
rect 22646 5624 22652 5636
rect 22112 5596 22652 5624
rect 21876 5584 21882 5596
rect 22646 5584 22652 5596
rect 22704 5584 22710 5636
rect 22741 5627 22799 5633
rect 22741 5593 22753 5627
rect 22787 5593 22799 5627
rect 24118 5624 24124 5636
rect 23966 5596 24124 5624
rect 22741 5587 22799 5593
rect 22186 5556 22192 5568
rect 21744 5528 22192 5556
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 22370 5516 22376 5568
rect 22428 5516 22434 5568
rect 22756 5556 22784 5587
rect 24118 5584 24124 5596
rect 24176 5624 24182 5636
rect 25130 5624 25136 5636
rect 24176 5596 25136 5624
rect 24176 5584 24182 5596
rect 25130 5584 25136 5596
rect 25188 5584 25194 5636
rect 23750 5556 23756 5568
rect 22756 5528 23756 5556
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 24213 5559 24271 5565
rect 24213 5525 24225 5559
rect 24259 5556 24271 5559
rect 24854 5556 24860 5568
rect 24259 5528 24860 5556
rect 24259 5525 24271 5528
rect 24213 5519 24271 5525
rect 24854 5516 24860 5528
rect 24912 5556 24918 5568
rect 25406 5556 25412 5568
rect 24912 5528 25412 5556
rect 24912 5516 24918 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 26142 5516 26148 5568
rect 26200 5516 26206 5568
rect 26694 5516 26700 5568
rect 26752 5516 26758 5568
rect 1104 5466 27876 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 27876 5466
rect 1104 5392 27876 5414
rect 1150 5312 1156 5364
rect 1208 5352 1214 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 1208 5324 1501 5352
rect 1208 5312 1214 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 5718 5352 5724 5364
rect 1489 5315 1547 5321
rect 4080 5324 5724 5352
rect 3786 5284 3792 5296
rect 3252 5256 3792 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 1688 5080 1716 5179
rect 2056 5148 2084 5179
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 3252 5225 3280 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4080 5225 4108 5324
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4212 5256 5304 5284
rect 4212 5244 4218 5256
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 4028 5188 4077 5216
rect 4028 5176 4034 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4614 5216 4620 5228
rect 4065 5179 4123 5185
rect 4172 5188 4620 5216
rect 3142 5148 3148 5160
rect 2056 5120 3148 5148
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 4172 5148 4200 5188
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 4798 5216 4804 5228
rect 4755 5188 4804 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5166 5216 5172 5228
rect 4939 5188 5172 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5276 5216 5304 5256
rect 5345 5219 5403 5225
rect 5345 5216 5357 5219
rect 5276 5188 5357 5216
rect 5345 5185 5357 5188
rect 5391 5185 5403 5219
rect 5345 5179 5403 5185
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5552 5215 5580 5324
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 7208 5324 8064 5352
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 5960 5256 6868 5284
rect 5960 5244 5966 5256
rect 5653 5219 5711 5225
rect 5537 5209 5595 5215
rect 3559 5120 4200 5148
rect 4341 5151 4399 5157
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 5460 5148 5488 5176
rect 5537 5175 5549 5209
rect 5583 5175 5595 5209
rect 5653 5185 5665 5219
rect 5699 5216 5711 5219
rect 5994 5216 6000 5228
rect 5699 5188 6000 5216
rect 5699 5185 5711 5188
rect 5653 5179 5711 5185
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5216 6147 5219
rect 6270 5216 6276 5228
rect 6135 5188 6276 5216
rect 6135 5185 6147 5188
rect 6089 5179 6147 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 6840 5225 6868 5256
rect 7208 5225 7236 5324
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6420 5188 6469 5216
rect 6420 5176 6426 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7650 5176 7656 5228
rect 7708 5176 7714 5228
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 5537 5169 5595 5175
rect 4387 5120 5488 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6288 5148 6316 5176
rect 6549 5151 6607 5157
rect 6288 5120 6500 5148
rect 2682 5080 2688 5092
rect 1688 5052 2688 5080
rect 2682 5040 2688 5052
rect 2740 5040 2746 5092
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 2924 5052 6377 5080
rect 2924 5040 2930 5052
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6472 5080 6500 5120
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6595 5120 6929 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7098 5108 7104 5160
rect 7156 5108 7162 5160
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7742 5148 7748 5160
rect 7423 5120 7748 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7300 5080 7328 5111
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7852 5148 7880 5179
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8036 5225 8064 5324
rect 8294 5312 8300 5364
rect 8352 5312 8358 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 8110 5244 8116 5296
rect 8168 5284 8174 5296
rect 8312 5284 8340 5312
rect 8772 5284 8800 5315
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 9950 5312 9956 5364
rect 10008 5312 10014 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 13630 5352 13636 5364
rect 10560 5324 13636 5352
rect 10560 5312 10566 5324
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 15102 5352 15108 5364
rect 14148 5324 15108 5352
rect 14148 5312 14154 5324
rect 15102 5312 15108 5324
rect 15160 5352 15166 5364
rect 18138 5352 18144 5364
rect 15160 5324 18144 5352
rect 15160 5312 15166 5324
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18248 5324 18429 5352
rect 9493 5287 9551 5293
rect 8168 5256 8616 5284
rect 8772 5256 9353 5284
rect 8168 5244 8174 5256
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8202 5216 8208 5228
rect 8067 5188 8208 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8588 5225 8616 5256
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8352 5188 8401 5216
rect 8352 5176 8358 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 9030 5216 9036 5228
rect 8990 5188 9036 5216
rect 8573 5179 8631 5185
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9122 5176 9128 5228
rect 9180 5176 9186 5228
rect 9214 5176 9220 5228
rect 9272 5176 9278 5228
rect 9325 5225 9353 5256
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 10042 5284 10048 5296
rect 9539 5256 10048 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 10686 5284 10692 5296
rect 10152 5256 10692 5284
rect 9310 5219 9368 5225
rect 9310 5185 9322 5219
rect 9356 5185 9368 5219
rect 9310 5179 9368 5185
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 10152 5225 10180 5256
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 11241 5287 11299 5293
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 11422 5284 11428 5296
rect 11287 5256 11428 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 11882 5244 11888 5296
rect 11940 5244 11946 5296
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12437 5287 12495 5293
rect 12437 5284 12449 5287
rect 12308 5256 12449 5284
rect 12308 5244 12314 5256
rect 12437 5253 12449 5256
rect 12483 5253 12495 5287
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 12437 5247 12495 5253
rect 12544 5256 12633 5284
rect 9682 5219 9740 5225
rect 9682 5185 9694 5219
rect 9728 5185 9740 5219
rect 9682 5179 9740 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10778 5216 10784 5228
rect 10551 5188 10784 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 9047 5148 9075 5176
rect 9697 5148 9725 5179
rect 7852 5120 9725 5148
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10244 5148 10272 5179
rect 9824 5120 10272 5148
rect 10336 5148 10364 5179
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 10962 5216 10968 5228
rect 10919 5188 10968 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11146 5176 11152 5228
rect 11204 5176 11210 5228
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 11388 5188 12204 5216
rect 11388 5176 11394 5188
rect 10594 5148 10600 5160
rect 10336 5120 10600 5148
rect 9824 5108 9830 5120
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5148 11115 5151
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11103 5120 11989 5148
rect 11103 5117 11115 5120
rect 11057 5111 11115 5117
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 7926 5080 7932 5092
rect 6472 5052 7932 5080
rect 6365 5043 6423 5049
rect 7926 5040 7932 5052
rect 7984 5040 7990 5092
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 9950 5080 9956 5092
rect 8720 5052 9956 5080
rect 8720 5040 8726 5052
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10704 5080 10732 5111
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 11330 5080 11336 5092
rect 10284 5052 11336 5080
rect 10284 5040 10290 5052
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 11606 5080 11612 5092
rect 11563 5052 11612 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 12176 5080 12204 5188
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 12544 5225 12572 5256
rect 12621 5253 12633 5256
rect 12667 5253 12679 5287
rect 13170 5284 13176 5296
rect 12621 5247 12679 5253
rect 13004 5256 13176 5284
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 13004 5216 13032 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 14182 5244 14188 5296
rect 14240 5284 14246 5296
rect 14921 5287 14979 5293
rect 14240 5256 14780 5284
rect 14240 5244 14246 5256
rect 14752 5228 14780 5256
rect 14921 5253 14933 5287
rect 14967 5284 14979 5287
rect 15194 5284 15200 5296
rect 14967 5256 15200 5284
rect 14967 5253 14979 5256
rect 14921 5247 14979 5253
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 15838 5244 15844 5296
rect 15896 5284 15902 5296
rect 16574 5284 16580 5296
rect 15896 5256 16580 5284
rect 15896 5244 15902 5256
rect 16574 5244 16580 5256
rect 16632 5284 16638 5296
rect 16761 5287 16819 5293
rect 16761 5284 16773 5287
rect 16632 5256 16773 5284
rect 16632 5244 16638 5256
rect 16761 5253 16773 5256
rect 16807 5253 16819 5287
rect 18248 5284 18276 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 19978 5352 19984 5364
rect 18932 5324 19984 5352
rect 18932 5312 18938 5324
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20257 5355 20315 5361
rect 20257 5352 20269 5355
rect 20220 5324 20269 5352
rect 20220 5312 20226 5324
rect 20257 5321 20269 5324
rect 20303 5321 20315 5355
rect 20257 5315 20315 5321
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 22278 5352 22284 5364
rect 20763 5324 22284 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 22520 5324 22569 5352
rect 22520 5312 22526 5324
rect 22557 5321 22569 5324
rect 22603 5321 22615 5355
rect 22557 5315 22615 5321
rect 24210 5312 24216 5364
rect 24268 5312 24274 5364
rect 24302 5312 24308 5364
rect 24360 5352 24366 5364
rect 25774 5352 25780 5364
rect 24360 5324 25780 5352
rect 24360 5312 24366 5324
rect 25774 5312 25780 5324
rect 25832 5312 25838 5364
rect 27430 5312 27436 5364
rect 27488 5312 27494 5364
rect 19426 5284 19432 5296
rect 16761 5247 16819 5253
rect 17328 5256 18276 5284
rect 18892 5256 19432 5284
rect 12759 5188 13032 5216
rect 13081 5219 13139 5225
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 14642 5216 14648 5228
rect 13127 5188 14648 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12728 5148 12756 5179
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 14792 5188 15485 5216
rect 14792 5176 14798 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 15795 5188 16804 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 12676 5120 12756 5148
rect 12676 5108 12682 5120
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 14090 5148 14096 5160
rect 12860 5120 14096 5148
rect 12860 5108 12866 5120
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14516 5120 15025 5148
rect 14516 5108 14522 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15672 5148 15700 5176
rect 15013 5111 15071 5117
rect 15488 5120 15700 5148
rect 15488 5092 15516 5120
rect 15930 5108 15936 5160
rect 15988 5148 15994 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15988 5120 16037 5148
rect 15988 5108 15994 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 16776 5148 16804 5188
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 17218 5216 17224 5228
rect 16908 5188 17224 5216
rect 16908 5176 16914 5188
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17328 5225 17356 5256
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17543 5188 17632 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 16776 5120 17540 5148
rect 15197 5083 15255 5089
rect 12176 5052 13032 5080
rect 1144 4972 1150 5024
rect 1202 5012 1208 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1202 4984 1869 5012
rect 1202 4972 1208 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2133 5015 2191 5021
rect 2133 5012 2145 5015
rect 2096 4984 2145 5012
rect 2096 4972 2102 4984
rect 2133 4981 2145 4984
rect 2179 4981 2191 5015
rect 2133 4975 2191 4981
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3384 4984 3433 5012
rect 3384 4972 3390 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3421 4975 3479 4981
rect 3878 4972 3884 5024
rect 3936 4972 3942 5024
rect 4430 4972 4436 5024
rect 4488 4972 4494 5024
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4580 4984 4629 5012
rect 4580 4972 4586 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4764 4984 4813 5012
rect 4764 4972 4770 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 4801 4975 4859 4981
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 5316 4984 5457 5012
rect 5316 4972 5322 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 8202 5012 8208 5024
rect 6779 4984 8208 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 9122 5012 9128 5024
rect 8536 4984 9128 5012
rect 8536 4972 8542 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12710 5012 12716 5024
rect 11848 4984 12716 5012
rect 11848 4972 11854 4984
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 13004 5021 13032 5052
rect 15197 5049 15209 5083
rect 15243 5080 15255 5083
rect 15470 5080 15476 5092
rect 15243 5052 15476 5080
rect 15243 5049 15255 5052
rect 15197 5043 15255 5049
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 15654 5040 15660 5092
rect 15712 5040 15718 5092
rect 16209 5083 16267 5089
rect 16209 5049 16221 5083
rect 16255 5049 16267 5083
rect 16209 5043 16267 5049
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13538 5012 13544 5024
rect 13035 4984 13544 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 15102 4972 15108 5024
rect 15160 5012 15166 5024
rect 16114 5012 16120 5024
rect 15160 4984 16120 5012
rect 15160 4972 15166 4984
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16224 5012 16252 5043
rect 16390 5040 16396 5092
rect 16448 5080 16454 5092
rect 17405 5083 17463 5089
rect 17405 5080 17417 5083
rect 16448 5052 17417 5080
rect 16448 5040 16454 5052
rect 17405 5049 17417 5052
rect 17451 5049 17463 5083
rect 17405 5043 17463 5049
rect 16850 5012 16856 5024
rect 16224 4984 16856 5012
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17512 5012 17540 5120
rect 17604 5089 17632 5188
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17736 5188 17969 5216
rect 17736 5176 17742 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 18506 5214 18512 5228
rect 17957 5179 18015 5185
rect 18432 5186 18512 5214
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5117 18199 5151
rect 18432 5148 18460 5186
rect 18506 5176 18512 5186
rect 18564 5176 18570 5228
rect 18892 5225 18920 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19518 5244 19524 5296
rect 19576 5244 19582 5296
rect 22370 5284 22376 5296
rect 20456 5256 22376 5284
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 19150 5176 19156 5228
rect 19208 5176 19214 5228
rect 19242 5176 19248 5228
rect 19300 5176 19306 5228
rect 20456 5225 20484 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 22646 5244 22652 5296
rect 22704 5284 22710 5296
rect 23477 5287 23535 5293
rect 23477 5284 23489 5287
rect 22704 5256 23489 5284
rect 22704 5244 22710 5256
rect 23477 5253 23489 5256
rect 23523 5284 23535 5287
rect 23566 5284 23572 5296
rect 23523 5256 23572 5284
rect 23523 5253 23535 5256
rect 23477 5247 23535 5253
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 24026 5284 24032 5296
rect 23768 5256 24032 5284
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5185 19395 5219
rect 19337 5179 19395 5185
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 18432 5120 18613 5148
rect 18141 5111 18199 5117
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5148 18843 5151
rect 18831 5120 18920 5148
rect 18831 5117 18843 5120
rect 18785 5111 18843 5117
rect 17589 5083 17647 5089
rect 17589 5049 17601 5083
rect 17635 5049 17647 5083
rect 17589 5043 17647 5049
rect 17862 5040 17868 5092
rect 17920 5080 17926 5092
rect 18156 5080 18184 5111
rect 17920 5052 18184 5080
rect 17920 5040 17926 5052
rect 18230 5040 18236 5092
rect 18288 5080 18294 5092
rect 18708 5080 18736 5111
rect 18288 5052 18736 5080
rect 18892 5080 18920 5120
rect 19260 5080 19288 5176
rect 19352 5092 19380 5179
rect 20898 5176 20904 5228
rect 20956 5176 20962 5228
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 21545 5209 21603 5215
rect 21545 5175 21557 5209
rect 21591 5175 21603 5209
rect 21634 5176 21640 5228
rect 21692 5216 21698 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21692 5188 21833 5216
rect 21692 5176 21698 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 22281 5219 22339 5225
rect 22281 5216 22293 5219
rect 21821 5179 21879 5185
rect 21928 5188 22293 5216
rect 21545 5169 21603 5175
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 19794 5148 19800 5160
rect 19751 5120 19800 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 20530 5108 20536 5160
rect 20588 5108 20594 5160
rect 20809 5151 20867 5157
rect 20809 5117 20821 5151
rect 20855 5148 20867 5151
rect 21450 5148 21456 5160
rect 20855 5120 21456 5148
rect 20855 5117 20867 5120
rect 20809 5111 20867 5117
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 18892 5052 19288 5080
rect 18288 5040 18294 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 19886 5080 19892 5092
rect 19392 5052 19892 5080
rect 19392 5040 19398 5052
rect 19886 5040 19892 5052
rect 19944 5080 19950 5092
rect 19981 5083 20039 5089
rect 19981 5080 19993 5083
rect 19944 5052 19993 5080
rect 19944 5040 19950 5052
rect 19981 5049 19993 5052
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 20165 5083 20223 5089
rect 20165 5049 20177 5083
rect 20211 5080 20223 5083
rect 21560 5080 21588 5169
rect 21726 5108 21732 5160
rect 21784 5148 21790 5160
rect 21928 5148 21956 5188
rect 22281 5185 22293 5188
rect 22327 5216 22339 5219
rect 22738 5216 22744 5228
rect 22327 5188 22744 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 23014 5176 23020 5228
rect 23072 5216 23078 5228
rect 23109 5219 23167 5225
rect 23109 5216 23121 5219
rect 23072 5188 23121 5216
rect 23072 5176 23078 5188
rect 23109 5185 23121 5188
rect 23155 5185 23167 5219
rect 23109 5179 23167 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 23382 5216 23388 5228
rect 23339 5188 23388 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 23768 5225 23796 5256
rect 24026 5244 24032 5256
rect 24084 5244 24090 5296
rect 25225 5287 25283 5293
rect 25225 5284 25237 5287
rect 24136 5256 25237 5284
rect 24136 5228 24164 5256
rect 25225 5253 25237 5256
rect 25271 5253 25283 5287
rect 25225 5247 25283 5253
rect 23753 5219 23811 5225
rect 23753 5185 23765 5219
rect 23799 5185 23811 5219
rect 23753 5179 23811 5185
rect 23842 5176 23848 5228
rect 23900 5176 23906 5228
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 24394 5176 24400 5228
rect 24452 5176 24458 5228
rect 24578 5176 24584 5228
rect 24636 5176 24642 5228
rect 24857 5219 24915 5225
rect 24857 5185 24869 5219
rect 24903 5185 24915 5219
rect 24857 5179 24915 5185
rect 25869 5219 25927 5225
rect 25869 5185 25881 5219
rect 25915 5216 25927 5219
rect 26142 5216 26148 5228
rect 25915 5188 26148 5216
rect 25915 5185 25927 5188
rect 25869 5179 25927 5185
rect 21784 5120 21956 5148
rect 22097 5151 22155 5157
rect 21784 5108 21790 5120
rect 22097 5117 22109 5151
rect 22143 5148 22155 5151
rect 22143 5120 22876 5148
rect 22143 5117 22155 5120
rect 22097 5111 22155 5117
rect 21818 5080 21824 5092
rect 20211 5052 21824 5080
rect 20211 5049 20223 5052
rect 20165 5043 20223 5049
rect 21818 5040 21824 5052
rect 21876 5040 21882 5092
rect 19058 5012 19064 5024
rect 17512 4984 19064 5012
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 20990 4972 20996 5024
rect 21048 4972 21054 5024
rect 21453 5015 21511 5021
rect 21453 4981 21465 5015
rect 21499 5012 21511 5015
rect 22112 5012 22140 5111
rect 22186 5040 22192 5092
rect 22244 5080 22250 5092
rect 22848 5080 22876 5120
rect 24026 5108 24032 5160
rect 24084 5148 24090 5160
rect 24872 5148 24900 5179
rect 26142 5176 26148 5188
rect 26200 5176 26206 5228
rect 26510 5176 26516 5228
rect 26568 5176 26574 5228
rect 27154 5176 27160 5228
rect 27212 5216 27218 5228
rect 27249 5219 27307 5225
rect 27249 5216 27261 5219
rect 27212 5188 27261 5216
rect 27212 5176 27218 5188
rect 27249 5185 27261 5188
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 25038 5148 25044 5160
rect 24084 5120 25044 5148
rect 24084 5108 24090 5120
rect 25038 5108 25044 5120
rect 25096 5108 25102 5160
rect 24762 5080 24768 5092
rect 22244 5052 22784 5080
rect 22848 5052 24768 5080
rect 22244 5040 22250 5052
rect 21499 4984 22140 5012
rect 21499 4981 21511 4984
rect 21453 4975 21511 4981
rect 22278 4972 22284 5024
rect 22336 4972 22342 5024
rect 22465 5015 22523 5021
rect 22465 4981 22477 5015
rect 22511 5012 22523 5015
rect 22554 5012 22560 5024
rect 22511 4984 22560 5012
rect 22511 4981 22523 4984
rect 22465 4975 22523 4981
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 22756 5021 22784 5052
rect 24762 5040 24768 5052
rect 24820 5040 24826 5092
rect 24854 5040 24860 5092
rect 24912 5080 24918 5092
rect 24912 5052 25084 5080
rect 24912 5040 24918 5052
rect 22741 5015 22799 5021
rect 22741 4981 22753 5015
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 23198 4972 23204 5024
rect 23256 5012 23262 5024
rect 23937 5015 23995 5021
rect 23937 5012 23949 5015
rect 23256 4984 23949 5012
rect 23256 4972 23262 4984
rect 23937 4981 23949 4984
rect 23983 4981 23995 5015
rect 23937 4975 23995 4981
rect 24581 5015 24639 5021
rect 24581 4981 24593 5015
rect 24627 5012 24639 5015
rect 24946 5012 24952 5024
rect 24627 4984 24952 5012
rect 24627 4981 24639 4984
rect 24581 4975 24639 4981
rect 24946 4972 24952 4984
rect 25004 4972 25010 5024
rect 25056 5021 25084 5052
rect 25041 5015 25099 5021
rect 25041 4981 25053 5015
rect 25087 4981 25099 5015
rect 25041 4975 25099 4981
rect 26694 4972 26700 5024
rect 26752 4972 26758 5024
rect 1104 4922 27876 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 27876 4922
rect 1104 4848 27876 4870
rect 2120 4811 2178 4817
rect 2120 4777 2132 4811
rect 2166 4808 2178 4811
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2166 4780 3801 4808
rect 2166 4777 2178 4780
rect 2120 4771 2178 4777
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5166 4808 5172 4820
rect 4939 4780 5172 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5626 4768 5632 4820
rect 5684 4768 5690 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 7374 4808 7380 4820
rect 5776 4780 7380 4808
rect 5776 4768 5782 4780
rect 7374 4768 7380 4780
rect 7432 4808 7438 4820
rect 11606 4808 11612 4820
rect 7432 4780 11612 4808
rect 7432 4768 7438 4780
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11756 4780 11805 4808
rect 11756 4768 11762 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12526 4768 12532 4820
rect 12584 4768 12590 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4777 13047 4811
rect 12989 4771 13047 4777
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13722 4808 13728 4820
rect 13403 4780 13728 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 1118 4700 1124 4752
rect 1176 4740 1182 4752
rect 1489 4743 1547 4749
rect 1489 4740 1501 4743
rect 1176 4712 1501 4740
rect 1176 4700 1182 4712
rect 1489 4709 1501 4712
rect 1535 4709 1547 4743
rect 1489 4703 1547 4709
rect 3605 4743 3663 4749
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 4614 4740 4620 4752
rect 3651 4712 4620 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 4614 4700 4620 4712
rect 4672 4740 4678 4752
rect 4985 4743 5043 4749
rect 4985 4740 4997 4743
rect 4672 4712 4997 4740
rect 4672 4700 4678 4712
rect 4985 4709 4997 4712
rect 5031 4709 5043 4743
rect 4985 4703 5043 4709
rect 5810 4700 5816 4752
rect 5868 4740 5874 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 5868 4712 8401 4740
rect 5868 4700 5874 4712
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 8478 4700 8484 4752
rect 8536 4740 8542 4752
rect 9214 4740 9220 4752
rect 8536 4712 9220 4740
rect 8536 4700 8542 4712
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 9309 4743 9367 4749
rect 9309 4709 9321 4743
rect 9355 4740 9367 4743
rect 9490 4740 9496 4752
rect 9355 4712 9496 4740
rect 9355 4709 9367 4712
rect 9309 4703 9367 4709
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 11146 4740 11152 4752
rect 9723 4712 11152 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 13004 4740 13032 4771
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 14700 4780 15393 4808
rect 14700 4768 14706 4780
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 15930 4808 15936 4820
rect 15381 4771 15439 4777
rect 15488 4780 15936 4808
rect 15488 4740 15516 4780
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 19702 4808 19708 4820
rect 16040 4780 19708 4808
rect 11572 4712 13032 4740
rect 13740 4712 15516 4740
rect 11572 4700 11578 4712
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2130 4672 2136 4684
rect 1903 4644 2136 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2682 4632 2688 4684
rect 2740 4672 2746 4684
rect 4433 4675 4491 4681
rect 2740 4644 4292 4672
rect 2740 4632 2746 4644
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3936 4576 4169 4604
rect 3936 4564 3942 4576
rect 4157 4573 4169 4576
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 3602 4536 3608 4548
rect 3358 4508 3608 4536
rect 3602 4496 3608 4508
rect 3660 4496 3666 4548
rect 4264 4536 4292 4644
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 5350 4672 5356 4684
rect 4479 4644 5356 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 6932 4644 10548 4672
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4396 4576 4721 4604
rect 4396 4564 4402 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 4890 4604 4896 4616
rect 4847 4576 4896 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 6178 4604 6184 4616
rect 5123 4576 6184 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6932 4613 6960 4644
rect 10520 4616 10548 4644
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11664 4644 12296 4672
rect 11664 4632 11670 4644
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7374 4564 7380 4616
rect 7432 4564 7438 4616
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 7926 4564 7932 4616
rect 7984 4564 7990 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 8168 4576 8309 4604
rect 8168 4564 8174 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8478 4604 8484 4616
rect 8435 4576 8484 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9582 4604 9588 4616
rect 8619 4576 9588 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 6362 4536 6368 4548
rect 4264 4508 6368 4536
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 7116 4536 7144 4564
rect 7668 4536 7696 4564
rect 7116 4508 7696 4536
rect 8018 4496 8024 4548
rect 8076 4496 8082 4548
rect 8202 4496 8208 4548
rect 8260 4496 8266 4548
rect 9125 4539 9183 4545
rect 9125 4505 9137 4539
rect 9171 4505 9183 4539
rect 9125 4499 9183 4505
rect 9401 4539 9459 4545
rect 9401 4505 9413 4539
rect 9447 4505 9459 4539
rect 9692 4536 9720 4567
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10134 4564 10140 4616
rect 10192 4564 10198 4616
rect 10502 4604 10508 4616
rect 10465 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 11790 4604 11796 4616
rect 10652 4576 11796 4604
rect 10652 4564 10658 4576
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 12158 4536 12164 4548
rect 9692 4508 12164 4536
rect 9401 4499 9459 4505
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 3694 4468 3700 4480
rect 3568 4440 3700 4468
rect 3568 4428 3574 4440
rect 3694 4428 3700 4440
rect 3752 4468 3758 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 3752 4440 4261 4468
rect 3752 4428 3758 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 5994 4468 6000 4480
rect 4948 4440 6000 4468
rect 4948 4428 4954 4440
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 7098 4428 7104 4480
rect 7156 4428 7162 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 9140 4468 9168 4499
rect 7340 4440 9168 4468
rect 9416 4468 9444 4499
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 12268 4536 12296 4644
rect 12618 4632 12624 4684
rect 12676 4632 12682 4684
rect 12710 4632 12716 4684
rect 12768 4672 12774 4684
rect 13740 4681 13768 4712
rect 15838 4700 15844 4752
rect 15896 4700 15902 4752
rect 13004 4672 13216 4680
rect 13725 4675 13783 4681
rect 13725 4672 13737 4675
rect 12768 4652 13737 4672
rect 12768 4644 13032 4652
rect 13188 4644 13737 4652
rect 12768 4632 12774 4644
rect 13725 4641 13737 4644
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 13832 4644 14228 4672
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12492 4576 12909 4604
rect 12492 4564 12498 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13078 4604 13084 4616
rect 13035 4576 13084 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13538 4564 13544 4616
rect 13596 4564 13602 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 13832 4604 13860 4644
rect 13688 4576 13860 4604
rect 14093 4607 14151 4613
rect 13688 4564 13694 4576
rect 14093 4573 14105 4607
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14108 4536 14136 4567
rect 12268 4508 14136 4536
rect 14200 4536 14228 4644
rect 15102 4632 15108 4684
rect 15160 4632 15166 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 15344 4644 15516 4672
rect 15344 4632 15350 4644
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 14332 4576 14381 4604
rect 14332 4564 14338 4576
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 15010 4564 15016 4616
rect 15068 4564 15074 4616
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 15378 4604 15384 4616
rect 15243 4576 15384 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15488 4613 15516 4644
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16040 4613 16068 4780
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 20162 4808 20168 4820
rect 19852 4780 20168 4808
rect 19852 4768 19858 4780
rect 20162 4768 20168 4780
rect 20220 4808 20226 4820
rect 21726 4808 21732 4820
rect 20220 4780 21732 4808
rect 20220 4768 20226 4780
rect 16114 4700 16120 4752
rect 16172 4740 16178 4752
rect 17678 4740 17684 4752
rect 16172 4712 16620 4740
rect 16172 4700 16178 4712
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16114 4564 16120 4616
rect 16172 4564 16178 4616
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16592 4613 16620 4712
rect 17512 4712 17684 4740
rect 17126 4672 17132 4684
rect 16776 4644 17132 4672
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 16264 4576 16313 4604
rect 16264 4564 16270 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 16666 4604 16672 4616
rect 16623 4576 16672 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 16408 4536 16436 4567
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16776 4613 16804 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 14200 4508 16436 4536
rect 16960 4536 16988 4567
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 17512 4613 17540 4712
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 18230 4740 18236 4752
rect 17788 4712 18236 4740
rect 17788 4672 17816 4712
rect 18230 4700 18236 4712
rect 18288 4700 18294 4752
rect 18524 4712 19012 4740
rect 18524 4672 18552 4712
rect 17604 4644 17816 4672
rect 17880 4644 18552 4672
rect 17604 4616 17632 4644
rect 17880 4616 17908 4644
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4604 17279 4607
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17267 4576 17325 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 17586 4564 17592 4616
rect 17644 4564 17650 4616
rect 17770 4564 17776 4616
rect 17828 4564 17834 4616
rect 17862 4564 17868 4616
rect 17920 4564 17926 4616
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18141 4607 18199 4613
rect 18141 4604 18153 4607
rect 18104 4576 18153 4604
rect 18104 4564 18110 4576
rect 18141 4573 18153 4576
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 17957 4539 18015 4545
rect 17957 4536 17969 4539
rect 16960 4508 17969 4536
rect 17957 4505 17969 4508
rect 18003 4505 18015 4539
rect 18156 4536 18184 4567
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 18414 4564 18420 4616
rect 18472 4564 18478 4616
rect 18524 4613 18552 4644
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 18984 4672 19012 4712
rect 19150 4700 19156 4752
rect 19208 4740 19214 4752
rect 20349 4743 20407 4749
rect 20349 4740 20361 4743
rect 19208 4712 20361 4740
rect 19208 4700 19214 4712
rect 20349 4709 20361 4712
rect 20395 4709 20407 4743
rect 20349 4703 20407 4709
rect 19797 4675 19855 4681
rect 19797 4672 19809 4675
rect 18656 4644 18920 4672
rect 18984 4644 19809 4672
rect 18656 4632 18662 4644
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 18782 4564 18788 4616
rect 18840 4564 18846 4616
rect 18892 4604 18920 4644
rect 19797 4641 19809 4644
rect 19843 4641 19855 4675
rect 19797 4635 19855 4641
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 20622 4672 20628 4684
rect 19944 4644 20628 4672
rect 19944 4632 19950 4644
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 20732 4681 20760 4780
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 22002 4768 22008 4820
rect 22060 4768 22066 4820
rect 22480 4780 26924 4808
rect 21082 4700 21088 4752
rect 21140 4700 21146 4752
rect 21821 4743 21879 4749
rect 21821 4709 21833 4743
rect 21867 4740 21879 4743
rect 22480 4740 22508 4780
rect 21867 4712 22508 4740
rect 21867 4709 21879 4712
rect 21821 4703 21879 4709
rect 24026 4700 24032 4752
rect 24084 4740 24090 4752
rect 24397 4743 24455 4749
rect 24397 4740 24409 4743
rect 24084 4712 24409 4740
rect 24084 4700 24090 4712
rect 24397 4709 24409 4712
rect 24443 4709 24455 4743
rect 24397 4703 24455 4709
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4641 20775 4675
rect 20717 4635 20775 4641
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4672 20867 4675
rect 20855 4644 21496 4672
rect 20855 4641 20867 4644
rect 20809 4635 20867 4641
rect 18969 4607 19027 4613
rect 18969 4604 18981 4607
rect 18892 4576 18981 4604
rect 18969 4573 18981 4576
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19702 4564 19708 4616
rect 19760 4564 19766 4616
rect 20254 4564 20260 4616
rect 20312 4564 20318 4616
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20533 4607 20591 4613
rect 20533 4604 20545 4607
rect 20404 4576 20545 4604
rect 20404 4564 20410 4576
rect 20533 4573 20545 4576
rect 20579 4604 20591 4607
rect 20898 4604 20904 4616
rect 20579 4576 20904 4604
rect 20579 4573 20591 4576
rect 20533 4567 20591 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 19260 4536 19288 4564
rect 19613 4539 19671 4545
rect 19613 4536 19625 4539
rect 18156 4508 19625 4536
rect 17957 4499 18015 4505
rect 19613 4505 19625 4508
rect 19659 4536 19671 4539
rect 20165 4539 20223 4545
rect 20165 4536 20177 4539
rect 19659 4508 20177 4536
rect 19659 4505 19671 4508
rect 19613 4499 19671 4505
rect 20165 4505 20177 4508
rect 20211 4505 20223 4539
rect 20165 4499 20223 4505
rect 9766 4468 9772 4480
rect 9416 4440 9772 4468
rect 7340 4428 7346 4440
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10413 4471 10471 4477
rect 10413 4437 10425 4471
rect 10459 4468 10471 4471
rect 10870 4468 10876 4480
rect 10459 4440 10876 4468
rect 10459 4437 10471 4440
rect 10413 4431 10471 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 12032 4440 12357 4468
rect 12032 4428 12038 4440
rect 12345 4437 12357 4440
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 14826 4468 14832 4480
rect 13771 4440 14832 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15286 4428 15292 4480
rect 15344 4468 15350 4480
rect 16114 4468 16120 4480
rect 15344 4440 16120 4468
rect 15344 4428 15350 4440
rect 16114 4428 16120 4440
rect 16172 4428 16178 4480
rect 16206 4428 16212 4480
rect 16264 4428 16270 4480
rect 16482 4428 16488 4480
rect 16540 4428 16546 4480
rect 16758 4428 16764 4480
rect 16816 4428 16822 4480
rect 17034 4428 17040 4480
rect 17092 4428 17098 4480
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18414 4468 18420 4480
rect 17828 4440 18420 4468
rect 17828 4428 17834 4440
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 18598 4428 18604 4480
rect 18656 4468 18662 4480
rect 18874 4468 18880 4480
rect 18656 4440 18880 4468
rect 18656 4428 18662 4440
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 18969 4471 19027 4477
rect 18969 4437 18981 4471
rect 19015 4468 19027 4471
rect 19058 4468 19064 4480
rect 19015 4440 19064 4468
rect 19015 4437 19027 4440
rect 18969 4431 19027 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19150 4428 19156 4480
rect 19208 4468 19214 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 19208 4440 19257 4468
rect 19208 4428 19214 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 21008 4468 21036 4567
rect 21174 4564 21180 4616
rect 21232 4564 21238 4616
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 19484 4440 21036 4468
rect 21284 4468 21312 4564
rect 21468 4548 21496 4644
rect 22738 4632 22744 4684
rect 22796 4672 22802 4684
rect 23753 4675 23811 4681
rect 23753 4672 23765 4675
rect 22796 4644 23765 4672
rect 22796 4632 22802 4644
rect 23753 4641 23765 4644
rect 23799 4672 23811 4675
rect 23799 4644 26188 4672
rect 23799 4641 23811 4644
rect 23753 4635 23811 4641
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 24026 4564 24032 4616
rect 24084 4564 24090 4616
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4604 24271 4607
rect 24302 4604 24308 4616
rect 24259 4576 24308 4604
rect 24259 4573 24271 4576
rect 24213 4567 24271 4573
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 26160 4613 26188 4644
rect 26896 4613 26924 4780
rect 27430 4768 27436 4820
rect 27488 4768 27494 4820
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4604 26203 4607
rect 26237 4607 26295 4613
rect 26237 4604 26249 4607
rect 26191 4576 26249 4604
rect 26191 4573 26203 4576
rect 26145 4567 26203 4573
rect 26237 4573 26249 4576
rect 26283 4573 26295 4607
rect 26237 4567 26295 4573
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4573 26663 4607
rect 26605 4567 26663 4573
rect 26881 4607 26939 4613
rect 26881 4573 26893 4607
rect 26927 4573 26939 4607
rect 26881 4567 26939 4573
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27338 4604 27344 4616
rect 27295 4576 27344 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 21450 4496 21456 4548
rect 21508 4496 21514 4548
rect 21545 4539 21603 4545
rect 21545 4505 21557 4539
rect 21591 4536 21603 4539
rect 21726 4536 21732 4548
rect 21591 4508 21732 4536
rect 21591 4505 21603 4508
rect 21545 4499 21603 4505
rect 21726 4496 21732 4508
rect 21784 4536 21790 4548
rect 22094 4536 22100 4548
rect 21784 4508 22100 4536
rect 21784 4496 21790 4508
rect 22094 4496 22100 4508
rect 22152 4496 22158 4548
rect 23046 4508 23335 4536
rect 23198 4468 23204 4480
rect 21284 4440 23204 4468
rect 19484 4428 19490 4440
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23307 4468 23335 4508
rect 23474 4496 23480 4548
rect 23532 4496 23538 4548
rect 25130 4496 25136 4548
rect 25188 4496 25194 4548
rect 25869 4539 25927 4545
rect 25869 4505 25881 4539
rect 25915 4505 25927 4539
rect 26620 4536 26648 4567
rect 27338 4564 27344 4576
rect 27396 4564 27402 4616
rect 25869 4499 25927 4505
rect 26068 4508 26648 4536
rect 23658 4468 23664 4480
rect 23307 4440 23664 4468
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 23845 4471 23903 4477
rect 23845 4437 23857 4471
rect 23891 4468 23903 4471
rect 24210 4468 24216 4480
rect 23891 4440 24216 4468
rect 23891 4437 23903 4440
rect 23845 4431 23903 4437
rect 24210 4428 24216 4440
rect 24268 4428 24274 4480
rect 24486 4428 24492 4480
rect 24544 4468 24550 4480
rect 25884 4468 25912 4499
rect 26068 4480 26096 4508
rect 24544 4440 25912 4468
rect 24544 4428 24550 4440
rect 26050 4428 26056 4480
rect 26108 4428 26114 4480
rect 26326 4428 26332 4480
rect 26384 4428 26390 4480
rect 26789 4471 26847 4477
rect 26789 4437 26801 4471
rect 26835 4468 26847 4471
rect 26970 4468 26976 4480
rect 26835 4440 26976 4468
rect 26835 4437 26847 4440
rect 26789 4431 26847 4437
rect 26970 4428 26976 4440
rect 27028 4428 27034 4480
rect 27062 4428 27068 4480
rect 27120 4428 27126 4480
rect 1104 4378 27876 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 27876 4378
rect 1104 4304 27876 4326
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 5718 4264 5724 4276
rect 4120 4236 5724 4264
rect 4120 4224 4126 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6362 4224 6368 4276
rect 6420 4224 6426 4276
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 7466 4264 7472 4276
rect 7147 4236 7472 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 10594 4264 10600 4276
rect 8076 4236 10600 4264
rect 8076 4224 8082 4236
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10796 4236 11069 4264
rect 4893 4199 4951 4205
rect 4893 4165 4905 4199
rect 4939 4196 4951 4199
rect 4982 4196 4988 4208
rect 4939 4168 4988 4196
rect 4939 4165 4951 4168
rect 4893 4159 4951 4165
rect 4982 4156 4988 4168
rect 5040 4196 5046 4208
rect 5258 4196 5264 4208
rect 5040 4168 5264 4196
rect 5040 4156 5046 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 7285 4199 7343 4205
rect 5920 4168 7144 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1946 4128 1952 4140
rect 1719 4100 1952 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 1486 3952 1492 4004
rect 1544 3952 1550 4004
rect 1854 3952 1860 4004
rect 1912 3952 1918 4004
rect 2056 3992 2084 4091
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2225 4131 2283 4137
rect 2225 4128 2237 4131
rect 2188 4100 2237 4128
rect 2188 4088 2194 4100
rect 2225 4097 2237 4100
rect 2271 4097 2283 4131
rect 2225 4091 2283 4097
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4396 4100 4445 4128
rect 4396 4088 4402 4100
rect 4433 4097 4445 4100
rect 4479 4128 4491 4131
rect 4522 4128 4528 4140
rect 4479 4100 4528 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5166 4128 5172 4140
rect 5123 4100 5172 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5442 4088 5448 4140
rect 5500 4137 5506 4140
rect 5500 4131 5549 4137
rect 5500 4097 5503 4131
rect 5537 4097 5549 4131
rect 5500 4091 5549 4097
rect 5500 4088 5506 4091
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5718 4088 5724 4140
rect 5776 4088 5782 4140
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 5920 4137 5948 4168
rect 6546 4137 6552 4140
rect 5904 4131 5962 4137
rect 5904 4128 5916 4131
rect 5868 4100 5916 4128
rect 5868 4088 5874 4100
rect 5904 4097 5916 4100
rect 5950 4097 5962 4131
rect 5904 4091 5962 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6544 4128 6552 4137
rect 6507 4100 6552 4128
rect 5997 4091 6055 4097
rect 6544 4091 6552 4100
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 3786 4060 3792 4072
rect 2547 4032 3792 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4028 4032 4261 4060
rect 4028 4020 4034 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 6012 4060 6040 4091
rect 6546 4088 6552 4091
rect 6604 4088 6610 4140
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 4847 4032 6040 4060
rect 6748 4060 6776 4091
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 6916 4131 6974 4137
rect 6916 4128 6928 4131
rect 6880 4100 6928 4128
rect 6880 4088 6886 4100
rect 6916 4097 6928 4100
rect 6962 4097 6974 4131
rect 6916 4091 6974 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7116 4128 7144 4168
rect 7285 4165 7297 4199
rect 7331 4196 7343 4199
rect 7374 4196 7380 4208
rect 7331 4168 7380 4196
rect 7331 4165 7343 4168
rect 7285 4159 7343 4165
rect 7374 4156 7380 4168
rect 7432 4196 7438 4208
rect 9030 4196 9036 4208
rect 7432 4168 7604 4196
rect 7432 4156 7438 4168
rect 7466 4128 7472 4140
rect 7116 4100 7472 4128
rect 7009 4091 7067 4097
rect 7024 4060 7052 4091
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7576 4137 7604 4168
rect 8128 4168 9036 4196
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 6748 4032 6960 4060
rect 7024 4032 7665 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 2222 3992 2228 4004
rect 2056 3964 2228 3992
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 5261 3995 5319 4001
rect 5261 3961 5273 3995
rect 5307 3992 5319 3995
rect 6822 3992 6828 4004
rect 5307 3964 6828 3992
rect 5307 3961 5319 3964
rect 5261 3955 5319 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 6932 3992 6960 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 7006 3992 7012 4004
rect 6932 3964 7012 3992
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 7760 3992 7788 4091
rect 8018 4088 8024 4140
rect 8076 4088 8082 4140
rect 8128 4137 8156 4168
rect 8496 4137 8524 4168
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 9493 4199 9551 4205
rect 9493 4165 9505 4199
rect 9539 4196 9551 4199
rect 9858 4196 9864 4208
rect 9539 4168 9864 4196
rect 9539 4165 9551 4168
rect 9493 4159 9551 4165
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 10686 4196 10692 4208
rect 10244 4168 10692 4196
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8113 4091 8171 4097
rect 8220 4100 8309 4128
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8220 4060 8248 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 8128 4032 8248 4060
rect 8404 4060 8432 4091
rect 8404 4032 8524 4060
rect 7156 3964 7788 3992
rect 8128 3992 8156 4032
rect 8386 3992 8392 4004
rect 8128 3964 8392 3992
rect 7156 3952 7162 3964
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 3200 3896 5365 3924
rect 3200 3884 3206 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5353 3887 5411 3893
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6638 3924 6644 3936
rect 5684 3896 6644 3924
rect 5684 3884 5690 3896
rect 6638 3884 6644 3896
rect 6696 3924 6702 3936
rect 7116 3924 7144 3952
rect 6696 3896 7144 3924
rect 7760 3924 7788 3964
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 8496 3992 8524 4032
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 8772 4060 8800 4091
rect 8720 4032 8800 4060
rect 8720 4020 8726 4032
rect 8846 4020 8852 4072
rect 8904 4020 8910 4072
rect 9232 3992 9260 4091
rect 9324 4060 9352 4091
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 9674 4088 9680 4140
rect 9732 4088 9738 4140
rect 10244 4137 10272 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9784 4100 9965 4128
rect 9784 4060 9812 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10046 4131 10104 4137
rect 10046 4097 10058 4131
rect 10092 4097 10104 4131
rect 10046 4091 10104 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 9324 4032 9812 4060
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10060 4060 10088 4091
rect 10318 4088 10324 4140
rect 10376 4088 10382 4140
rect 10459 4131 10517 4137
rect 10459 4097 10471 4131
rect 10505 4128 10517 4131
rect 10796 4128 10824 4236
rect 11057 4233 11069 4236
rect 11103 4264 11115 4267
rect 11330 4264 11336 4276
rect 11103 4236 11336 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 11517 4267 11575 4273
rect 11517 4233 11529 4267
rect 11563 4264 11575 4267
rect 12066 4264 12072 4276
rect 11563 4236 12072 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 12526 4264 12532 4276
rect 12216 4236 12532 4264
rect 12216 4224 12222 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 12989 4267 13047 4273
rect 12989 4233 13001 4267
rect 13035 4264 13047 4267
rect 13538 4264 13544 4276
rect 13035 4236 13544 4264
rect 13035 4233 13047 4236
rect 12989 4227 13047 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 17862 4264 17868 4276
rect 14292 4236 17868 4264
rect 14292 4208 14320 4236
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18012 4236 18092 4264
rect 18012 4224 18018 4236
rect 13078 4196 13084 4208
rect 12452 4168 13084 4196
rect 12452 4140 12480 4168
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 13265 4199 13323 4205
rect 13265 4165 13277 4199
rect 13311 4196 13323 4199
rect 13630 4196 13636 4208
rect 13311 4168 13636 4196
rect 13311 4165 13323 4168
rect 13265 4159 13323 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 14274 4196 14280 4208
rect 13832 4168 14280 4196
rect 10505 4100 10824 4128
rect 10505 4097 10517 4100
rect 10459 4091 10517 4097
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 11146 4088 11152 4140
rect 11204 4088 11210 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11790 4128 11796 4140
rect 11747 4100 11796 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 9907 4032 10088 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11606 4060 11612 4072
rect 11112 4032 11612 4060
rect 11112 4020 11118 4032
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11900 4060 11928 4091
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11900 4032 12081 4060
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12360 4060 12388 4091
rect 12434 4088 12440 4140
rect 12492 4088 12498 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12584 4100 12633 4128
rect 12584 4088 12590 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12802 4088 12808 4140
rect 12860 4088 12866 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13280 4100 13461 4128
rect 12820 4060 12848 4088
rect 13280 4072 13308 4100
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13587 4100 13676 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 12360 4032 12848 4060
rect 12069 4023 12127 4029
rect 13262 4020 13268 4072
rect 13320 4020 13326 4072
rect 13648 4060 13676 4100
rect 13722 4088 13728 4140
rect 13780 4088 13786 4140
rect 13832 4137 13860 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 15010 4196 15016 4208
rect 14384 4168 15016 4196
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 14384 4137 14412 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 15194 4156 15200 4208
rect 15252 4196 15258 4208
rect 16390 4196 16396 4208
rect 15252 4168 16396 4196
rect 15252 4156 15258 4168
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 14829 4131 14887 4137
rect 14829 4128 14841 4131
rect 14608 4100 14841 4128
rect 14608 4088 14614 4100
rect 14829 4097 14841 4100
rect 14875 4097 14887 4131
rect 14829 4091 14887 4097
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 13648 4032 13860 4060
rect 9674 3992 9680 4004
rect 8496 3964 9680 3992
rect 7926 3924 7932 3936
rect 7760 3896 7932 3924
rect 6696 3884 6702 3896
rect 7926 3884 7932 3896
rect 7984 3924 7990 3936
rect 8496 3924 8524 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10597 3995 10655 4001
rect 10597 3992 10609 3995
rect 10008 3964 10609 3992
rect 10008 3952 10014 3964
rect 10597 3961 10609 3964
rect 10643 3961 10655 3995
rect 10597 3955 10655 3961
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 13280 3992 13308 4020
rect 13832 3992 13860 4032
rect 13906 4020 13912 4072
rect 13964 4020 13970 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14200 3992 14228 4023
rect 14274 4020 14280 4072
rect 14332 4020 14338 4072
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14516 4032 14657 4060
rect 14516 4020 14522 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 10836 3964 13032 3992
rect 13280 3964 13768 3992
rect 13832 3964 14412 3992
rect 10836 3952 10842 3964
rect 7984 3896 8524 3924
rect 8573 3927 8631 3933
rect 7984 3884 7990 3896
rect 8573 3893 8585 3927
rect 8619 3924 8631 3927
rect 9582 3924 9588 3936
rect 8619 3896 9588 3924
rect 8619 3893 8631 3896
rect 8573 3887 8631 3893
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 9640 3896 12633 3924
rect 9640 3884 9646 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 13004 3924 13032 3964
rect 13446 3924 13452 3936
rect 13004 3896 13452 3924
rect 12621 3887 12679 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13740 3924 13768 3964
rect 14384 3936 14412 3964
rect 14918 3952 14924 4004
rect 14976 3952 14982 4004
rect 15028 3992 15056 4023
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 15304 4060 15332 4091
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 15930 4128 15936 4140
rect 15887 4100 15936 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16114 4088 16120 4140
rect 16172 4137 16178 4140
rect 16316 4137 16344 4168
rect 16390 4156 16396 4168
rect 16448 4196 16454 4208
rect 16945 4199 17003 4205
rect 16945 4196 16957 4199
rect 16448 4168 16957 4196
rect 16448 4156 16454 4168
rect 16945 4165 16957 4168
rect 16991 4196 17003 4199
rect 17494 4196 17500 4208
rect 16991 4168 17500 4196
rect 16991 4165 17003 4168
rect 16945 4159 17003 4165
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 18064 4205 18092 4236
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 19334 4264 19340 4276
rect 18288 4236 19340 4264
rect 18288 4224 18294 4236
rect 19334 4224 19340 4236
rect 19392 4224 19398 4276
rect 20162 4264 20168 4276
rect 19812 4236 20168 4264
rect 18049 4199 18107 4205
rect 18049 4165 18061 4199
rect 18095 4165 18107 4199
rect 18049 4159 18107 4165
rect 18414 4156 18420 4208
rect 18472 4196 18478 4208
rect 18782 4196 18788 4208
rect 18472 4168 18788 4196
rect 18472 4156 18478 4168
rect 18782 4156 18788 4168
rect 18840 4156 18846 4208
rect 19058 4196 19064 4208
rect 18892 4168 19064 4196
rect 16172 4131 16205 4137
rect 16193 4097 16205 4131
rect 16172 4091 16205 4097
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16172 4088 16178 4091
rect 16850 4088 16856 4140
rect 16908 4088 16914 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17310 4128 17316 4140
rect 17175 4100 17316 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 15304 4032 16681 4060
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17052 4060 17080 4091
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17736 4100 17785 4128
rect 17736 4088 17742 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 17000 4032 17080 4060
rect 17972 4060 18000 4091
rect 18138 4088 18144 4140
rect 18196 4128 18202 4140
rect 18196 4100 18552 4128
rect 18196 4088 18202 4100
rect 18414 4060 18420 4072
rect 17972 4032 18420 4060
rect 17000 4020 17006 4032
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 15028 3964 15669 3992
rect 15657 3961 15669 3964
rect 15703 3992 15715 3995
rect 15933 3995 15991 4001
rect 15933 3992 15945 3995
rect 15703 3964 15945 3992
rect 15703 3961 15715 3964
rect 15657 3955 15715 3961
rect 15933 3961 15945 3964
rect 15979 3961 15991 3995
rect 15933 3955 15991 3961
rect 17678 3952 17684 4004
rect 17736 3992 17742 4004
rect 17972 3992 18000 4032
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 17736 3964 18000 3992
rect 18524 3992 18552 4100
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 18892 4137 18920 4168
rect 19058 4156 19064 4168
rect 19116 4156 19122 4208
rect 19521 4199 19579 4205
rect 19521 4165 19533 4199
rect 19567 4196 19579 4199
rect 19812 4196 19840 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 22738 4264 22744 4276
rect 22388 4236 22744 4264
rect 19567 4168 19840 4196
rect 19567 4165 19579 4168
rect 19521 4159 19579 4165
rect 19886 4156 19892 4208
rect 19944 4156 19950 4208
rect 21545 4199 21603 4205
rect 21545 4165 21557 4199
rect 21591 4196 21603 4199
rect 22388 4196 22416 4236
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 23290 4224 23296 4276
rect 23348 4224 23354 4276
rect 23569 4267 23627 4273
rect 23569 4233 23581 4267
rect 23615 4264 23627 4267
rect 24486 4264 24492 4276
rect 23615 4236 24492 4264
rect 23615 4233 23627 4236
rect 23569 4227 23627 4233
rect 24486 4224 24492 4236
rect 24544 4224 24550 4276
rect 24946 4224 24952 4276
rect 25004 4264 25010 4276
rect 26602 4264 26608 4276
rect 25004 4236 26608 4264
rect 25004 4224 25010 4236
rect 26602 4224 26608 4236
rect 26660 4224 26666 4276
rect 21591 4168 22416 4196
rect 21591 4165 21603 4168
rect 21545 4159 21603 4165
rect 22554 4156 22560 4208
rect 22612 4196 22618 4208
rect 24210 4196 24216 4208
rect 22612 4168 23152 4196
rect 22612 4156 22618 4168
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 19150 4137 19156 4140
rect 19146 4128 19156 4137
rect 19111 4100 19156 4128
rect 19146 4091 19156 4100
rect 19150 4088 19156 4091
rect 19208 4088 19214 4140
rect 19242 4088 19248 4140
rect 19300 4137 19306 4140
rect 19300 4131 19349 4137
rect 19300 4097 19303 4131
rect 19337 4097 19349 4131
rect 19300 4091 19349 4097
rect 19300 4088 19306 4091
rect 19426 4088 19432 4140
rect 19484 4088 19490 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19536 4100 19625 4128
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 18785 4063 18843 4069
rect 18785 4060 18797 4063
rect 18656 4032 18797 4060
rect 18656 4020 18662 4032
rect 18785 4029 18797 4032
rect 18831 4029 18843 4063
rect 19536 4060 19564 4100
rect 19613 4097 19625 4100
rect 19659 4128 19671 4131
rect 21634 4128 21640 4140
rect 19659 4100 21640 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22695 4100 22753 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 21450 4060 21456 4072
rect 18785 4023 18843 4029
rect 19260 4032 19564 4060
rect 19628 4032 21456 4060
rect 19260 3992 19288 4032
rect 18524 3964 19288 3992
rect 17736 3952 17742 3964
rect 19334 3952 19340 4004
rect 19392 3992 19398 4004
rect 19628 3992 19656 4032
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 21542 4020 21548 4072
rect 21600 4060 21606 4072
rect 22554 4060 22560 4072
rect 21600 4032 22560 4060
rect 21600 4020 21606 4032
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 22940 4060 22968 4091
rect 23014 4088 23020 4140
rect 23072 4088 23078 4140
rect 23124 4137 23152 4168
rect 23676 4168 24216 4196
rect 23109 4131 23167 4137
rect 23109 4097 23121 4131
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 23676 4060 23704 4168
rect 24210 4156 24216 4168
rect 24268 4156 24274 4208
rect 24302 4156 24308 4208
rect 24360 4196 24366 4208
rect 24360 4168 26280 4196
rect 24360 4156 24366 4168
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 24118 4088 24124 4140
rect 24176 4088 24182 4140
rect 25314 4128 25320 4140
rect 24228 4100 25320 4128
rect 24228 4069 24256 4100
rect 25314 4088 25320 4100
rect 25372 4128 25378 4140
rect 25590 4128 25596 4140
rect 25372 4100 25596 4128
rect 25372 4088 25378 4100
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 25774 4088 25780 4140
rect 25832 4088 25838 4140
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 26142 4128 26148 4140
rect 26099 4100 26148 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 26142 4088 26148 4100
rect 26200 4088 26206 4140
rect 26252 4137 26280 4168
rect 26237 4131 26295 4137
rect 26237 4097 26249 4131
rect 26283 4097 26295 4131
rect 26237 4091 26295 4097
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 27249 4131 27307 4137
rect 27249 4097 27261 4131
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 22940 4032 23704 4060
rect 23753 4063 23811 4069
rect 23753 4029 23765 4063
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 19392 3964 19656 3992
rect 19392 3952 19398 3964
rect 20438 3952 20444 4004
rect 20496 3992 20502 4004
rect 20496 3964 23520 3992
rect 20496 3952 20502 3964
rect 14090 3924 14096 3936
rect 13740 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 15562 3933 15568 3936
rect 15519 3927 15568 3933
rect 15519 3893 15531 3927
rect 15565 3893 15568 3927
rect 15519 3887 15568 3893
rect 15562 3884 15568 3887
rect 15620 3884 15626 3936
rect 15746 3884 15752 3936
rect 15804 3884 15810 3936
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 18138 3924 18144 3936
rect 17276 3896 18144 3924
rect 17276 3884 17282 3896
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 18506 3924 18512 3936
rect 18371 3896 18512 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 18932 3896 19073 3924
rect 18932 3884 18938 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 19794 3884 19800 3936
rect 19852 3884 19858 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23014 3924 23020 3936
rect 20680 3896 23020 3924
rect 20680 3884 20686 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23492 3924 23520 3964
rect 23566 3952 23572 4004
rect 23624 3992 23630 4004
rect 23768 3992 23796 4023
rect 25038 4020 25044 4072
rect 25096 4020 25102 4072
rect 25222 4020 25228 4072
rect 25280 4020 25286 4072
rect 27264 4060 27292 4091
rect 25424 4032 27292 4060
rect 25424 3992 25452 4032
rect 23624 3964 23796 3992
rect 23860 3964 25452 3992
rect 25501 3995 25559 4001
rect 23624 3952 23630 3964
rect 23860 3924 23888 3964
rect 25501 3961 25513 3995
rect 25547 3992 25559 3995
rect 26053 3995 26111 4001
rect 25547 3964 26004 3992
rect 25547 3961 25559 3964
rect 25501 3955 25559 3961
rect 23492 3896 23888 3924
rect 23934 3884 23940 3936
rect 23992 3924 23998 3936
rect 24489 3927 24547 3933
rect 24489 3924 24501 3927
rect 23992 3896 24501 3924
rect 23992 3884 23998 3896
rect 24489 3893 24501 3896
rect 24535 3893 24547 3927
rect 24489 3887 24547 3893
rect 24670 3884 24676 3936
rect 24728 3924 24734 3936
rect 25516 3924 25544 3955
rect 24728 3896 25544 3924
rect 24728 3884 24734 3896
rect 25682 3884 25688 3936
rect 25740 3884 25746 3936
rect 25774 3884 25780 3936
rect 25832 3924 25838 3936
rect 25869 3927 25927 3933
rect 25869 3924 25881 3927
rect 25832 3896 25881 3924
rect 25832 3884 25838 3896
rect 25869 3893 25881 3896
rect 25915 3893 25927 3927
rect 25976 3924 26004 3964
rect 26053 3961 26065 3995
rect 26099 3992 26111 3995
rect 26234 3992 26240 4004
rect 26099 3964 26240 3992
rect 26099 3961 26111 3964
rect 26053 3955 26111 3961
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 27430 3952 27436 4004
rect 27488 3952 27494 4004
rect 26142 3924 26148 3936
rect 25976 3896 26148 3924
rect 25869 3887 25927 3893
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 26694 3884 26700 3936
rect 26752 3884 26758 3936
rect 27062 3884 27068 3936
rect 27120 3884 27126 3936
rect 1104 3834 27876 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 27876 3834
rect 1104 3760 27876 3782
rect 1302 3680 1308 3732
rect 1360 3720 1366 3732
rect 1489 3723 1547 3729
rect 1489 3720 1501 3723
rect 1360 3692 1501 3720
rect 1360 3680 1366 3692
rect 1489 3689 1501 3692
rect 1535 3689 1547 3723
rect 1489 3683 1547 3689
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4430 3720 4436 3732
rect 4028 3692 4436 3720
rect 4028 3680 4034 3692
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5626 3720 5632 3732
rect 5408 3692 5632 3720
rect 5408 3680 5414 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5776 3692 6009 3720
rect 5776 3680 5782 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 6178 3680 6184 3732
rect 6236 3680 6242 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 6512 3692 6745 3720
rect 6512 3680 6518 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 6733 3683 6791 3689
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8662 3720 8668 3732
rect 8168 3692 8668 3720
rect 8168 3680 8174 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9950 3720 9956 3732
rect 9364 3692 9956 3720
rect 9364 3680 9370 3692
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 10100 3692 10149 3720
rect 10100 3680 10106 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10137 3683 10195 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 12618 3720 12624 3732
rect 11020 3692 12624 3720
rect 11020 3680 11026 3692
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 13265 3723 13323 3729
rect 13265 3720 13277 3723
rect 12676 3692 13277 3720
rect 12676 3680 12682 3692
rect 13265 3689 13277 3692
rect 13311 3689 13323 3723
rect 13265 3683 13323 3689
rect 14921 3723 14979 3729
rect 14921 3689 14933 3723
rect 14967 3720 14979 3723
rect 15010 3720 15016 3732
rect 14967 3692 15016 3720
rect 14967 3689 14979 3692
rect 14921 3683 14979 3689
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 17862 3680 17868 3732
rect 17920 3680 17926 3732
rect 19061 3723 19119 3729
rect 19061 3689 19073 3723
rect 19107 3720 19119 3723
rect 19426 3720 19432 3732
rect 19107 3692 19432 3720
rect 19107 3689 19119 3692
rect 19061 3683 19119 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 23842 3720 23848 3732
rect 20640 3692 23848 3720
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 3510 3652 3516 3664
rect 3292 3624 3516 3652
rect 3292 3612 3298 3624
rect 3510 3612 3516 3624
rect 3568 3612 3574 3664
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 4948 3624 5120 3652
rect 4948 3612 4954 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2130 3584 2136 3596
rect 1903 3556 2136 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 3605 3587 3663 3593
rect 2832 3556 3556 3584
rect 2832 3544 2838 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 3528 3516 3556 3556
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4798 3584 4804 3596
rect 3651 3556 4804 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3528 3488 3985 3516
rect 3973 3485 3985 3488
rect 4019 3516 4031 3519
rect 4062 3516 4068 3528
rect 4019 3488 4068 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4338 3516 4344 3528
rect 4295 3488 4344 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4632 3525 4660 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 2133 3451 2191 3457
rect 2133 3417 2145 3451
rect 2179 3417 2191 3451
rect 3789 3451 3847 3457
rect 3789 3448 3801 3451
rect 2133 3411 2191 3417
rect 3436 3420 3801 3448
rect 2148 3380 2176 3411
rect 3436 3380 3464 3420
rect 3789 3417 3801 3420
rect 3835 3417 3847 3451
rect 4724 3448 4752 3479
rect 3789 3411 3847 3417
rect 4632 3420 4752 3448
rect 4908 3448 4936 3479
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5092 3525 5120 3624
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5316 3624 9904 3652
rect 5316 3612 5322 3624
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5994 3584 6000 3596
rect 5399 3556 5672 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5442 3516 5448 3528
rect 5123 3488 5448 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5644 3525 5672 3556
rect 5828 3556 6000 3584
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5828 3448 5856 3556
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6546 3584 6552 3596
rect 6319 3556 6552 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 7064 3556 7328 3584
rect 7064 3544 7070 3556
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 4908 3420 5856 3448
rect 5920 3448 5948 3479
rect 6362 3476 6368 3528
rect 6420 3476 6426 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 6914 3516 6920 3528
rect 6871 3488 6920 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 6178 3448 6184 3460
rect 5920 3420 6184 3448
rect 4632 3392 4660 3420
rect 6178 3408 6184 3420
rect 6236 3448 6242 3460
rect 6656 3448 6684 3479
rect 6914 3476 6920 3488
rect 6972 3516 6978 3528
rect 7300 3525 7328 3556
rect 8110 3544 8116 3596
rect 8168 3544 8174 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8536 3556 9168 3584
rect 8536 3544 8542 3556
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6972 3488 7113 3516
rect 6972 3476 6978 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7524 3488 7941 3516
rect 7524 3476 7530 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 7929 3479 7987 3485
rect 8128 3488 8309 3516
rect 6236 3420 6684 3448
rect 7561 3451 7619 3457
rect 6236 3408 6242 3420
rect 7561 3417 7573 3451
rect 7607 3417 7619 3451
rect 7561 3411 7619 3417
rect 7653 3451 7711 3457
rect 7653 3417 7665 3451
rect 7699 3448 7711 3451
rect 7742 3448 7748 3460
rect 7699 3420 7748 3448
rect 7699 3417 7711 3420
rect 7653 3411 7711 3417
rect 2148 3352 3464 3380
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 3970 3380 3976 3392
rect 3660 3352 3976 3380
rect 3660 3340 3666 3352
rect 3970 3340 3976 3352
rect 4028 3380 4034 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 4028 3352 4169 3380
rect 4028 3340 4034 3352
rect 4157 3349 4169 3352
rect 4203 3380 4215 3383
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 4203 3352 4445 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 4433 3343 4491 3349
rect 4614 3340 4620 3392
rect 4672 3340 4678 3392
rect 4798 3340 4804 3392
rect 4856 3380 4862 3392
rect 5445 3383 5503 3389
rect 5445 3380 5457 3383
rect 4856 3352 5457 3380
rect 4856 3340 4862 3352
rect 5445 3349 5457 3352
rect 5491 3349 5503 3383
rect 5445 3343 5503 3349
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 6914 3380 6920 3392
rect 5859 3352 6920 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7576 3380 7604 3411
rect 7742 3408 7748 3420
rect 7800 3448 7806 3460
rect 8128 3448 8156 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8662 3516 8668 3528
rect 8619 3488 8668 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 7800 3420 8156 3448
rect 7800 3408 7806 3420
rect 8202 3408 8208 3460
rect 8260 3408 8266 3460
rect 8404 3448 8432 3479
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 8938 3516 8944 3528
rect 8864 3488 8944 3516
rect 8754 3448 8760 3460
rect 8404 3420 8760 3448
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 8110 3380 8116 3392
rect 7576 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8864 3380 8892 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9140 3525 9168 3556
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9876 3584 9904 3624
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11974 3652 11980 3664
rect 11756 3624 11980 3652
rect 11756 3612 11762 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12802 3652 12808 3664
rect 12176 3624 12808 3652
rect 10321 3587 10379 3593
rect 9640 3556 9812 3584
rect 9876 3556 10180 3584
rect 9640 3544 9646 3556
rect 9784 3525 9812 3556
rect 10152 3528 10180 3556
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 11716 3584 11744 3612
rect 10367 3556 11744 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 9692 3448 9720 3479
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 9968 3448 9996 3476
rect 9692 3420 9996 3448
rect 8527 3352 8892 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 9585 3383 9643 3389
rect 9585 3380 9597 3383
rect 9456 3352 9597 3380
rect 9456 3340 9462 3352
rect 9585 3349 9597 3352
rect 9631 3349 9643 3383
rect 9585 3343 9643 3349
rect 9858 3340 9864 3392
rect 9916 3340 9922 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10060 3380 10088 3479
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12066 3516 12072 3528
rect 11664 3488 12072 3516
rect 11664 3476 11670 3488
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 10594 3408 10600 3460
rect 10652 3408 10658 3460
rect 12176 3448 12204 3624
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 13449 3655 13507 3661
rect 13449 3621 13461 3655
rect 13495 3652 13507 3655
rect 17770 3652 17776 3664
rect 13495 3624 17776 3652
rect 13495 3621 13507 3624
rect 13449 3615 13507 3621
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 12345 3587 12403 3593
rect 12345 3553 12357 3587
rect 12391 3584 12403 3587
rect 12618 3584 12624 3596
rect 12391 3556 12624 3584
rect 12391 3553 12403 3556
rect 12345 3547 12403 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12986 3584 12992 3596
rect 12728 3556 12992 3584
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12308 3488 12449 3516
rect 12308 3476 12314 3488
rect 12437 3485 12449 3488
rect 12483 3516 12495 3519
rect 12728 3516 12756 3556
rect 12986 3544 12992 3556
rect 13044 3584 13050 3596
rect 13170 3584 13176 3596
rect 13044 3556 13176 3584
rect 13044 3544 13050 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 15105 3587 15163 3593
rect 13320 3556 14596 3584
rect 13320 3544 13326 3556
rect 12483 3488 12756 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 12860 3488 13768 3516
rect 12860 3476 12866 3488
rect 11900 3420 12204 3448
rect 11900 3380 11928 3420
rect 10008 3352 11928 3380
rect 10008 3340 10014 3352
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12268 3380 12296 3476
rect 13078 3408 13084 3460
rect 13136 3448 13142 3460
rect 13136 3420 13400 3448
rect 13136 3408 13142 3420
rect 12032 3352 12296 3380
rect 12032 3340 12038 3352
rect 12618 3340 12624 3392
rect 12676 3340 12682 3392
rect 12710 3340 12716 3392
rect 12768 3340 12774 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 12894 3380 12900 3392
rect 12851 3352 12900 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 12986 3340 12992 3392
rect 13044 3340 13050 3392
rect 13262 3340 13268 3392
rect 13320 3389 13326 3392
rect 13320 3383 13339 3389
rect 13327 3349 13339 3383
rect 13372 3380 13400 3420
rect 13630 3380 13636 3392
rect 13372 3352 13636 3380
rect 13320 3343 13339 3349
rect 13320 3340 13326 3343
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13740 3389 13768 3488
rect 13906 3476 13912 3528
rect 13964 3476 13970 3528
rect 14090 3476 14096 3528
rect 14148 3476 14154 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 14274 3408 14280 3460
rect 14332 3408 14338 3460
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3417 14427 3451
rect 14568 3448 14596 3556
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15562 3584 15568 3596
rect 15151 3556 15568 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 17402 3584 17408 3596
rect 15672 3556 17408 3584
rect 15194 3476 15200 3528
rect 15252 3476 15258 3528
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 15672 3448 15700 3556
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17880 3584 17908 3680
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 19150 3652 19156 3664
rect 18104 3624 19156 3652
rect 18104 3612 18110 3624
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 19242 3612 19248 3664
rect 19300 3652 19306 3664
rect 19610 3652 19616 3664
rect 19300 3624 19616 3652
rect 19300 3612 19306 3624
rect 19610 3612 19616 3624
rect 19668 3612 19674 3664
rect 19797 3655 19855 3661
rect 19797 3621 19809 3655
rect 19843 3652 19855 3655
rect 20640 3652 20668 3692
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 26234 3720 26240 3732
rect 24780 3692 26240 3720
rect 19843 3624 20668 3652
rect 19843 3621 19855 3624
rect 19797 3615 19855 3621
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 23477 3655 23535 3661
rect 23477 3652 23489 3655
rect 23072 3624 23489 3652
rect 23072 3612 23078 3624
rect 23477 3621 23489 3624
rect 23523 3652 23535 3655
rect 23523 3624 24624 3652
rect 23523 3621 23535 3624
rect 23477 3615 23535 3621
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 17880 3556 17969 3584
rect 17957 3553 17969 3556
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18414 3544 18420 3596
rect 18472 3584 18478 3596
rect 19889 3587 19947 3593
rect 18472 3556 19656 3584
rect 18472 3544 18478 3556
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 14568 3420 15700 3448
rect 14369 3411 14427 3417
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 14384 3380 14412 3411
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16298 3448 16304 3460
rect 15988 3420 16304 3448
rect 15988 3408 15994 3420
rect 16298 3408 16304 3420
rect 16356 3448 16362 3460
rect 16500 3448 16528 3479
rect 16666 3476 16672 3528
rect 16724 3476 16730 3528
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 17644 3488 18184 3516
rect 17644 3476 17650 3488
rect 18156 3460 18184 3488
rect 18432 3488 18705 3516
rect 16942 3448 16948 3460
rect 16356 3420 16948 3448
rect 16356 3408 16362 3420
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 18138 3408 18144 3460
rect 18196 3408 18202 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18432 3448 18460 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 18782 3476 18788 3528
rect 18840 3476 18846 3528
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19208 3488 19533 3516
rect 19208 3476 19214 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 18288 3420 18460 3448
rect 18509 3451 18567 3457
rect 18288 3408 18294 3420
rect 18509 3417 18521 3451
rect 18555 3448 18567 3451
rect 19245 3451 19303 3457
rect 19245 3448 19257 3451
rect 18555 3420 19257 3448
rect 18555 3417 18567 3420
rect 18509 3411 18567 3417
rect 19245 3417 19257 3420
rect 19291 3417 19303 3451
rect 19628 3448 19656 3556
rect 19889 3553 19901 3587
rect 19935 3584 19947 3587
rect 20070 3584 20076 3596
rect 19935 3556 20076 3584
rect 19935 3553 19947 3556
rect 19889 3547 19947 3553
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 20312 3556 22784 3584
rect 20312 3544 20318 3556
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 20438 3516 20444 3528
rect 19852 3488 20444 3516
rect 19852 3476 19858 3488
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 20530 3476 20536 3528
rect 20588 3476 20594 3528
rect 22756 3516 22784 3556
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 24596 3593 24624 3624
rect 24780 3593 24808 3692
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 27430 3680 27436 3732
rect 27488 3680 27494 3732
rect 24854 3612 24860 3664
rect 24912 3652 24918 3664
rect 24912 3624 27292 3652
rect 24912 3612 24918 3624
rect 23385 3587 23443 3593
rect 23385 3584 23397 3587
rect 22888 3556 23397 3584
rect 22888 3544 22894 3556
rect 23385 3553 23397 3556
rect 23431 3553 23443 3587
rect 23385 3547 23443 3553
rect 24581 3587 24639 3593
rect 24581 3553 24593 3587
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25409 3587 25467 3593
rect 25409 3553 25421 3587
rect 25455 3584 25467 3587
rect 27062 3584 27068 3596
rect 25455 3556 27068 3584
rect 25455 3553 25467 3556
rect 25409 3547 25467 3553
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 21942 3488 22692 3516
rect 22756 3488 23213 3516
rect 20257 3451 20315 3457
rect 20257 3448 20269 3451
rect 19628 3420 20269 3448
rect 19245 3411 19303 3417
rect 20257 3417 20269 3420
rect 20303 3417 20315 3451
rect 20257 3411 20315 3417
rect 20806 3408 20812 3460
rect 20864 3408 20870 3460
rect 22278 3408 22284 3460
rect 22336 3448 22342 3460
rect 22557 3451 22615 3457
rect 22557 3448 22569 3451
rect 22336 3420 22569 3448
rect 22336 3408 22342 3420
rect 22557 3417 22569 3420
rect 22603 3417 22615 3451
rect 22664 3448 22692 3488
rect 23201 3485 23213 3488
rect 23247 3516 23259 3519
rect 23566 3516 23572 3528
rect 23247 3488 23572 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3512 23719 3519
rect 23934 3512 23940 3528
rect 23707 3485 23940 3512
rect 23661 3484 23940 3485
rect 23661 3479 23719 3484
rect 23934 3476 23940 3484
rect 23992 3476 23998 3528
rect 24210 3476 24216 3528
rect 24268 3476 24274 3528
rect 24670 3476 24676 3528
rect 24728 3516 24734 3528
rect 25041 3519 25099 3525
rect 25041 3516 25053 3519
rect 24728 3488 25053 3516
rect 24728 3476 24734 3488
rect 25041 3485 25053 3488
rect 25087 3485 25099 3519
rect 25685 3519 25743 3525
rect 25685 3516 25697 3519
rect 25041 3479 25099 3485
rect 25148 3488 25697 3516
rect 23106 3448 23112 3460
rect 22664 3420 23112 3448
rect 22557 3411 22615 3417
rect 23106 3408 23112 3420
rect 23164 3408 23170 3460
rect 25148 3448 25176 3488
rect 25685 3485 25697 3488
rect 25731 3485 25743 3519
rect 25685 3479 25743 3485
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3485 25835 3519
rect 25777 3479 25835 3485
rect 26145 3519 26203 3525
rect 26145 3485 26157 3519
rect 26191 3485 26203 3519
rect 26145 3479 26203 3485
rect 23216 3420 25176 3448
rect 13771 3352 14412 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 16577 3383 16635 3389
rect 16577 3349 16589 3383
rect 16623 3380 16635 3383
rect 16850 3380 16856 3392
rect 16623 3352 16856 3380
rect 16623 3349 16635 3352
rect 16577 3343 16635 3349
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 16960 3380 16988 3408
rect 23216 3392 23244 3420
rect 25590 3408 25596 3460
rect 25648 3448 25654 3460
rect 25792 3448 25820 3479
rect 26160 3448 26188 3479
rect 26234 3476 26240 3528
rect 26292 3516 26298 3528
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 26292 3488 26525 3516
rect 26292 3476 26298 3488
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 26513 3479 26571 3485
rect 26878 3476 26884 3528
rect 26936 3476 26942 3528
rect 27264 3525 27292 3624
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3485 27307 3519
rect 27249 3479 27307 3485
rect 25648 3420 25820 3448
rect 25884 3420 26188 3448
rect 25648 3408 25654 3420
rect 18322 3380 18328 3392
rect 16960 3352 18328 3380
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 18414 3340 18420 3392
rect 18472 3380 18478 3392
rect 19334 3380 19340 3392
rect 18472 3352 19340 3380
rect 18472 3340 18478 3352
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 19426 3340 19432 3392
rect 19484 3340 19490 3392
rect 19610 3340 19616 3392
rect 19668 3340 19674 3392
rect 20441 3383 20499 3389
rect 20441 3349 20453 3383
rect 20487 3380 20499 3383
rect 20714 3380 20720 3392
rect 20487 3352 20720 3380
rect 20487 3349 20499 3352
rect 20441 3343 20499 3349
rect 20714 3340 20720 3352
rect 20772 3340 20778 3392
rect 21082 3340 21088 3392
rect 21140 3380 21146 3392
rect 22649 3383 22707 3389
rect 22649 3380 22661 3383
rect 21140 3352 22661 3380
rect 21140 3340 21146 3352
rect 22649 3349 22661 3352
rect 22695 3349 22707 3383
rect 22649 3343 22707 3349
rect 23198 3340 23204 3392
rect 23256 3340 23262 3392
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 23845 3383 23903 3389
rect 23845 3380 23857 3383
rect 23808 3352 23857 3380
rect 23808 3340 23814 3352
rect 23845 3349 23857 3352
rect 23891 3349 23903 3383
rect 23845 3343 23903 3349
rect 23934 3340 23940 3392
rect 23992 3380 23998 3392
rect 24029 3383 24087 3389
rect 24029 3380 24041 3383
rect 23992 3352 24041 3380
rect 23992 3340 23998 3352
rect 24029 3349 24041 3352
rect 24075 3349 24087 3383
rect 24029 3343 24087 3349
rect 24670 3340 24676 3392
rect 24728 3340 24734 3392
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 25501 3383 25559 3389
rect 25501 3380 25513 3383
rect 24820 3352 25513 3380
rect 24820 3340 24826 3352
rect 25501 3349 25513 3352
rect 25547 3349 25559 3383
rect 25501 3343 25559 3349
rect 25774 3340 25780 3392
rect 25832 3380 25838 3392
rect 25884 3380 25912 3420
rect 25832 3352 25912 3380
rect 25832 3340 25838 3352
rect 25958 3340 25964 3392
rect 26016 3340 26022 3392
rect 26142 3340 26148 3392
rect 26200 3380 26206 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 26200 3352 26341 3380
rect 26200 3340 26206 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 26694 3340 26700 3392
rect 26752 3340 26758 3392
rect 27062 3340 27068 3392
rect 27120 3340 27126 3392
rect 1104 3290 27876 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 27876 3290
rect 1104 3216 27876 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1360 3148 1869 3176
rect 1360 3136 1366 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 1857 3139 1915 3145
rect 2424 3148 4261 3176
rect 2424 3117 2452 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5445 3179 5503 3185
rect 4580 3148 5396 3176
rect 4580 3136 4586 3148
rect 2409 3111 2467 3117
rect 2409 3077 2421 3111
rect 2455 3077 2467 3111
rect 2409 3071 2467 3077
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 4338 3108 4344 3120
rect 4120 3080 4344 3108
rect 4120 3068 4126 3080
rect 4338 3068 4344 3080
rect 4396 3108 4402 3120
rect 4617 3111 4675 3117
rect 4617 3108 4629 3111
rect 4396 3080 4629 3108
rect 4396 3068 4402 3080
rect 4617 3077 4629 3080
rect 4663 3108 4675 3111
rect 5258 3108 5264 3120
rect 4663 3080 5264 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 5368 3108 5396 3148
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5534 3176 5540 3188
rect 5491 3148 5540 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6086 3176 6092 3188
rect 5767 3148 6092 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 7064 3148 7573 3176
rect 7064 3136 7070 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 7561 3139 7619 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8076 3148 8309 3176
rect 8076 3136 8082 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 8662 3136 8668 3188
rect 8720 3136 8726 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 9306 3176 9312 3188
rect 8956 3148 9312 3176
rect 5902 3108 5908 3120
rect 5368 3080 5908 3108
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 2004 3012 2053 3040
rect 2004 3000 2010 3012
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2130 3000 2136 3052
rect 2188 3000 2194 3052
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4304 3012 4445 3040
rect 4304 3000 4310 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4522 3000 4528 3052
rect 4580 3000 4586 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4847 3012 4905 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 4893 3009 4905 3012
rect 4939 3040 4951 3043
rect 5074 3040 5080 3052
rect 4939 3012 5080 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4816 2972 4844 3003
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5368 3040 5396 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 5215 3012 5396 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5500 3012 5641 3040
rect 5500 3000 5506 3012
rect 5629 3009 5641 3012
rect 5675 3040 5687 3043
rect 5718 3040 5724 3052
rect 5675 3012 5724 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6104 3049 6132 3136
rect 6638 3108 6644 3120
rect 6196 3080 6644 3108
rect 6196 3049 6224 3080
rect 6638 3068 6644 3080
rect 6696 3108 6702 3120
rect 8386 3108 8392 3120
rect 6696 3080 7236 3108
rect 6696 3068 6702 3080
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 4203 2944 4844 2972
rect 6104 2972 6132 3003
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 7208 3049 7236 3080
rect 7668 3080 8392 3108
rect 7668 3049 7696 3080
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6604 3012 6929 3040
rect 6604 3000 6610 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7834 3000 7840 3052
rect 7892 3000 7898 3052
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 8956 3049 8984 3148
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9548 3148 10088 3176
rect 9548 3136 9554 3148
rect 9582 3108 9588 3120
rect 9232 3080 9588 3108
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8812 3012 8953 3040
rect 8812 3000 8818 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9232 3049 9260 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3108 9735 3111
rect 9950 3108 9956 3120
rect 9723 3080 9956 3108
rect 9723 3077 9735 3080
rect 9677 3071 9735 3077
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 9398 3000 9404 3052
rect 9456 3000 9462 3052
rect 10060 3049 10088 3148
rect 10134 3136 10140 3188
rect 10192 3136 10198 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10284 3148 10364 3176
rect 10284 3136 10290 3148
rect 10152 3108 10180 3136
rect 10336 3117 10364 3148
rect 10594 3136 10600 3188
rect 10652 3136 10658 3188
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 14458 3176 14464 3188
rect 10836 3148 14464 3176
rect 10836 3136 10842 3148
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 15378 3176 15384 3188
rect 14660 3148 15384 3176
rect 10321 3111 10379 3117
rect 10152 3080 10272 3108
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10134 3040 10140 3052
rect 10091 3012 10140 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 6104 2944 6960 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 1210 2864 1216 2916
rect 1268 2904 1274 2916
rect 1489 2907 1547 2913
rect 1489 2904 1501 2907
rect 1268 2876 1501 2904
rect 1268 2864 1274 2876
rect 1489 2873 1501 2876
rect 1535 2873 1547 2907
rect 1489 2867 1547 2873
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 3476 2876 5488 2904
rect 3476 2864 3482 2876
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 4982 2836 4988 2848
rect 3936 2808 4988 2836
rect 3936 2796 3942 2808
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5460 2836 5488 2876
rect 6178 2864 6184 2916
rect 6236 2864 6242 2916
rect 6932 2904 6960 2944
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7064 2944 7297 2972
rect 7064 2932 7070 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7984 2944 8033 2972
rect 7984 2932 7990 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 8220 2904 8248 2935
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8904 2944 9137 2972
rect 8904 2932 8910 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9416 2972 9444 3000
rect 9125 2935 9183 2941
rect 9244 2944 9444 2972
rect 9784 2972 9812 3003
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10244 3049 10272 3080
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 11793 3111 11851 3117
rect 10367 3080 11560 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10244 2972 10272 3003
rect 10410 3000 10416 3052
rect 10468 3000 10474 3052
rect 11532 3049 11560 3080
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 11974 3108 11980 3120
rect 11839 3080 11980 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 12124 3080 12926 3108
rect 12124 3068 12130 3080
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 14185 3111 14243 3117
rect 14185 3108 14197 3111
rect 13780 3080 14197 3108
rect 13780 3068 13786 3080
rect 14185 3077 14197 3080
rect 14231 3108 14243 3111
rect 14550 3108 14556 3120
rect 14231 3080 14556 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 14550 3068 14556 3080
rect 14608 3068 14614 3120
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 11563 3012 11652 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 11422 2972 11428 2984
rect 9784 2944 10180 2972
rect 10244 2944 11428 2972
rect 9244 2904 9272 2944
rect 6932 2876 7328 2904
rect 8220 2876 9272 2904
rect 6454 2836 6460 2848
rect 5460 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7300 2845 7328 2876
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 9784 2904 9812 2944
rect 9364 2876 9812 2904
rect 9364 2864 9370 2876
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 7742 2796 7748 2848
rect 7800 2796 7806 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9490 2836 9496 2848
rect 9088 2808 9496 2836
rect 9088 2796 9094 2808
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9950 2796 9956 2848
rect 10008 2796 10014 2848
rect 10152 2836 10180 2944
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 10962 2904 10968 2916
rect 10284 2876 10968 2904
rect 10284 2864 10290 2876
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 10778 2836 10784 2848
rect 10152 2808 10784 2836
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11624 2836 11652 3012
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11882 3000 11888 3052
rect 11940 3000 11946 3052
rect 12158 3000 12164 3052
rect 12216 3000 12222 3052
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14660 3040 14688 3148
rect 15378 3136 15384 3148
rect 15436 3176 15442 3188
rect 15930 3176 15936 3188
rect 15436 3148 15936 3176
rect 15436 3136 15442 3148
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 20530 3176 20536 3188
rect 16684 3148 20536 3176
rect 14734 3068 14740 3120
rect 14792 3108 14798 3120
rect 14792 3080 14858 3108
rect 14792 3068 14798 3080
rect 16684 3049 16712 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20993 3179 21051 3185
rect 20993 3176 21005 3179
rect 20864 3148 21005 3176
rect 20864 3136 20870 3148
rect 20993 3145 21005 3148
rect 21039 3145 21051 3179
rect 20993 3139 21051 3145
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21508 3148 21833 3176
rect 21508 3136 21514 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 23566 3136 23572 3188
rect 23624 3176 23630 3188
rect 24118 3176 24124 3188
rect 23624 3148 24124 3176
rect 23624 3136 23630 3148
rect 24118 3136 24124 3148
rect 24176 3136 24182 3188
rect 25130 3176 25136 3188
rect 24228 3148 25136 3176
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 20548 3108 20576 3136
rect 21634 3108 21640 3120
rect 18288 3080 19288 3108
rect 20548 3080 21640 3108
rect 18288 3068 18294 3080
rect 19260 3052 19288 3080
rect 21634 3068 21640 3080
rect 21692 3108 21698 3120
rect 22738 3108 22744 3120
rect 21692 3080 22744 3108
rect 21692 3068 21698 3080
rect 14424 3012 14688 3040
rect 16301 3043 16359 3049
rect 14424 3000 14430 3012
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16347 3012 16681 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 18969 3043 19027 3049
rect 18969 3040 18981 3043
rect 18156 3012 18981 3040
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12084 2944 12449 2972
rect 12084 2913 12112 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 14090 2972 14096 2984
rect 13228 2944 14096 2972
rect 13228 2932 13234 2944
rect 14090 2932 14096 2944
rect 14148 2972 14154 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14148 2944 14289 2972
rect 14148 2932 14154 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15344 2944 16037 2972
rect 15344 2932 15350 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 16942 2932 16948 2984
rect 17000 2932 17006 2984
rect 17678 2932 17684 2984
rect 17736 2972 17742 2984
rect 18156 2972 18184 3012
rect 18969 3009 18981 3012
rect 19015 3009 19027 3043
rect 18969 3003 19027 3009
rect 19058 3000 19064 3052
rect 19116 3000 19122 3052
rect 19242 3000 19248 3052
rect 19300 3000 19306 3052
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19576 3012 19717 3040
rect 19576 3000 19582 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 20162 3000 20168 3052
rect 20220 3000 20226 3052
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 20496 3012 20545 3040
rect 20496 3000 20502 3012
rect 20533 3009 20545 3012
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 17736 2944 18184 2972
rect 17736 2932 17742 2944
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18380 2944 18705 2972
rect 18380 2932 18386 2944
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 19076 2972 19104 3000
rect 18693 2935 18751 2941
rect 18800 2944 19104 2972
rect 12069 2907 12127 2913
rect 12069 2873 12081 2907
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 18046 2864 18052 2916
rect 18104 2904 18110 2916
rect 18414 2904 18420 2916
rect 18104 2876 18420 2904
rect 18104 2864 18110 2876
rect 18414 2864 18420 2876
rect 18472 2864 18478 2916
rect 18800 2904 18828 2944
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19484 2944 19809 2972
rect 19484 2932 19490 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 20254 2932 20260 2984
rect 20312 2932 20318 2984
rect 20548 2972 20576 3003
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 20806 3000 20812 3052
rect 20864 3000 20870 3052
rect 21082 3000 21088 3052
rect 21140 3000 21146 3052
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 21192 3012 21281 3040
rect 21192 2972 21220 3012
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 20548 2944 21220 2972
rect 21376 2972 21404 3003
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 22278 3040 22284 3052
rect 21928 3012 22284 3040
rect 21928 2972 21956 3012
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 22388 3049 22416 3080
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 22373 3043 22431 3049
rect 22373 3009 22385 3043
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 23658 3000 23664 3052
rect 23716 3040 23722 3052
rect 23716 3026 23782 3040
rect 23716 3012 23796 3026
rect 23716 3000 23722 3012
rect 21376 2944 21956 2972
rect 18524 2876 18828 2904
rect 12434 2836 12440 2848
rect 11624 2808 12440 2836
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 14918 2836 14924 2848
rect 12860 2808 14924 2836
rect 12860 2796 12866 2808
rect 14918 2796 14924 2808
rect 14976 2836 14982 2848
rect 16666 2836 16672 2848
rect 14976 2808 16672 2836
rect 14976 2796 14982 2808
rect 16666 2796 16672 2808
rect 16724 2836 16730 2848
rect 18524 2836 18552 2876
rect 18874 2864 18880 2916
rect 18932 2904 18938 2916
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 18932 2876 19533 2904
rect 18932 2864 18938 2876
rect 19521 2873 19533 2876
rect 19567 2873 19579 2907
rect 21376 2904 21404 2944
rect 22002 2932 22008 2984
rect 22060 2932 22066 2984
rect 22094 2932 22100 2984
rect 22152 2932 22158 2984
rect 22186 2932 22192 2984
rect 22244 2932 22250 2984
rect 22649 2975 22707 2981
rect 22649 2972 22661 2975
rect 22388 2944 22661 2972
rect 19521 2867 19579 2873
rect 20640 2876 21404 2904
rect 21637 2907 21695 2913
rect 20640 2848 20668 2876
rect 21637 2873 21649 2907
rect 21683 2904 21695 2907
rect 22388 2904 22416 2944
rect 22649 2941 22661 2944
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 23106 2932 23112 2984
rect 23164 2972 23170 2984
rect 23768 2972 23796 3012
rect 24228 2972 24256 3148
rect 25130 3136 25136 3148
rect 25188 3136 25194 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 25685 3179 25743 3185
rect 25685 3176 25697 3179
rect 25280 3148 25697 3176
rect 25280 3136 25286 3148
rect 25685 3145 25697 3148
rect 25731 3145 25743 3179
rect 25685 3139 25743 3145
rect 27430 3136 27436 3188
rect 27488 3136 27494 3188
rect 24854 3068 24860 3120
rect 24912 3068 24918 3120
rect 24489 3043 24547 3049
rect 24489 3009 24501 3043
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 23164 2944 24256 2972
rect 24504 2972 24532 3003
rect 24578 3000 24584 3052
rect 24636 3040 24642 3052
rect 24673 3043 24731 3049
rect 24673 3040 24685 3043
rect 24636 3012 24685 3040
rect 24636 3000 24642 3012
rect 24673 3009 24685 3012
rect 24719 3009 24731 3043
rect 24673 3003 24731 3009
rect 24765 3043 24823 3049
rect 24765 3009 24777 3043
rect 24811 3040 24823 3043
rect 24872 3040 24900 3068
rect 24811 3012 24900 3040
rect 24811 3009 24823 3012
rect 24765 3003 24823 3009
rect 24946 3000 24952 3052
rect 25004 3000 25010 3052
rect 25038 3000 25044 3052
rect 25096 3000 25102 3052
rect 25133 3043 25191 3049
rect 25133 3009 25145 3043
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 24854 2972 24860 2984
rect 24504 2944 24860 2972
rect 23164 2932 23170 2944
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 24964 2972 24992 3000
rect 25148 2972 25176 3003
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 25682 3000 25688 3052
rect 25740 3040 25746 3052
rect 25869 3043 25927 3049
rect 25869 3040 25881 3043
rect 25740 3012 25881 3040
rect 25740 3000 25746 3012
rect 25869 3009 25881 3012
rect 25915 3009 25927 3043
rect 25869 3003 25927 3009
rect 25961 3043 26019 3049
rect 25961 3009 25973 3043
rect 26007 3009 26019 3043
rect 25961 3003 26019 3009
rect 24964 2944 25176 2972
rect 25501 2975 25559 2981
rect 25501 2941 25513 2975
rect 25547 2972 25559 2975
rect 25976 2972 26004 3003
rect 26510 3000 26516 3052
rect 26568 3000 26574 3052
rect 26970 3000 26976 3052
rect 27028 3000 27034 3052
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 25547 2944 26004 2972
rect 25547 2941 25559 2944
rect 25501 2935 25559 2941
rect 26418 2932 26424 2984
rect 26476 2972 26482 2984
rect 27062 2972 27068 2984
rect 26476 2944 27068 2972
rect 26476 2932 26482 2944
rect 27062 2932 27068 2944
rect 27120 2972 27126 2984
rect 27172 2972 27200 3003
rect 27246 3000 27252 3052
rect 27304 3000 27310 3052
rect 27120 2944 27200 2972
rect 27120 2932 27126 2944
rect 21683 2876 22416 2904
rect 21683 2873 21695 2876
rect 21637 2867 21695 2873
rect 24118 2864 24124 2916
rect 24176 2904 24182 2916
rect 24394 2904 24400 2916
rect 24176 2876 24400 2904
rect 24176 2864 24182 2876
rect 24394 2864 24400 2876
rect 24452 2904 24458 2916
rect 24581 2907 24639 2913
rect 24581 2904 24593 2907
rect 24452 2876 24593 2904
rect 24452 2864 24458 2876
rect 24581 2873 24593 2876
rect 24627 2873 24639 2907
rect 24581 2867 24639 2873
rect 16724 2808 18552 2836
rect 16724 2796 16730 2808
rect 18782 2796 18788 2848
rect 18840 2796 18846 2848
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 19024 2808 19073 2836
rect 19024 2796 19030 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 19061 2799 19119 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 20622 2836 20628 2848
rect 19208 2808 20628 2836
rect 19208 2796 19214 2808
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 21910 2796 21916 2848
rect 21968 2836 21974 2848
rect 24305 2839 24363 2845
rect 24305 2836 24317 2839
rect 21968 2808 24317 2836
rect 21968 2796 21974 2808
rect 24305 2805 24317 2808
rect 24351 2805 24363 2839
rect 24596 2836 24624 2867
rect 25038 2864 25044 2916
rect 25096 2904 25102 2916
rect 26145 2907 26203 2913
rect 26145 2904 26157 2907
rect 25096 2876 26157 2904
rect 25096 2864 25102 2876
rect 26145 2873 26157 2876
rect 26191 2873 26203 2907
rect 26973 2907 27031 2913
rect 26973 2904 26985 2907
rect 26145 2867 26203 2873
rect 26252 2876 26985 2904
rect 26252 2836 26280 2876
rect 26973 2873 26985 2876
rect 27019 2873 27031 2907
rect 26973 2867 27031 2873
rect 24596 2808 26280 2836
rect 26697 2839 26755 2845
rect 24305 2799 24363 2805
rect 26697 2805 26709 2839
rect 26743 2836 26755 2839
rect 26878 2836 26884 2848
rect 26743 2808 26884 2836
rect 26743 2805 26755 2808
rect 26697 2799 26755 2805
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 1104 2746 27876 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 27876 2746
rect 1104 2672 27876 2694
rect 1486 2592 1492 2644
rect 1544 2592 1550 2644
rect 1854 2592 1860 2644
rect 1912 2592 1918 2644
rect 2746 2604 3556 2632
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 2593 2567 2651 2573
rect 2593 2564 2605 2567
rect 1360 2536 2605 2564
rect 1360 2524 1366 2536
rect 2593 2533 2605 2536
rect 2639 2533 2651 2567
rect 2593 2527 2651 2533
rect 1118 2456 1124 2508
rect 1176 2496 1182 2508
rect 2746 2496 2774 2604
rect 3528 2564 3556 2604
rect 3786 2592 3792 2644
rect 3844 2592 3850 2644
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2601 5595 2635
rect 5537 2595 5595 2601
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 5810 2632 5816 2644
rect 5767 2604 5816 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 4893 2567 4951 2573
rect 4893 2564 4905 2567
rect 3528 2536 4905 2564
rect 4893 2533 4905 2536
rect 4939 2533 4951 2567
rect 5552 2564 5580 2595
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 5994 2632 6000 2644
rect 5951 2604 6000 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 6825 2635 6883 2641
rect 6825 2632 6837 2635
rect 6696 2604 6837 2632
rect 6696 2592 6702 2604
rect 6825 2601 6837 2604
rect 6871 2601 6883 2635
rect 6825 2595 6883 2601
rect 7116 2604 9352 2632
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5552 2536 6377 2564
rect 4893 2527 4951 2533
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 7116 2564 7144 2604
rect 6512 2536 7144 2564
rect 6512 2524 6518 2536
rect 4798 2496 4804 2508
rect 1176 2468 2774 2496
rect 3252 2468 4804 2496
rect 1176 2456 1182 2468
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2314 2428 2320 2440
rect 2087 2400 2320 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2406 2388 2412 2440
rect 2464 2388 2470 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3252 2428 3280 2468
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5445 2499 5503 2505
rect 5040 2468 5212 2496
rect 5040 2456 5046 2468
rect 2823 2400 3280 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 3016 2332 3065 2360
rect 3016 2320 3022 2332
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 3694 2360 3700 2372
rect 3283 2332 3700 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 3988 2360 4016 2391
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4614 2428 4620 2440
rect 4387 2400 4620 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5184 2437 5212 2468
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 5902 2496 5908 2508
rect 5491 2468 5908 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5902 2456 5908 2468
rect 5960 2496 5966 2508
rect 7006 2496 7012 2508
rect 5960 2468 7012 2496
rect 5960 2456 5966 2468
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 6086 2388 6092 2440
rect 6144 2388 6150 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 4908 2360 4936 2388
rect 3988 2332 4936 2360
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 6564 2360 6592 2391
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7116 2437 7144 2536
rect 8021 2567 8079 2573
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 8294 2564 8300 2576
rect 8067 2536 8300 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8938 2564 8944 2576
rect 8588 2536 8944 2564
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8588 2496 8616 2536
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 7883 2468 8616 2496
rect 9324 2496 9352 2604
rect 9490 2592 9496 2644
rect 9548 2592 9554 2644
rect 12437 2635 12495 2641
rect 9692 2604 10732 2632
rect 9692 2496 9720 2604
rect 9324 2468 9720 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 5316 2332 6592 2360
rect 5316 2320 5322 2332
rect 1026 2252 1032 2304
rect 1084 2292 1090 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 1084 2264 2237 2292
rect 1084 2252 1090 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3878 2292 3884 2304
rect 3559 2264 3884 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 4525 2295 4583 2301
rect 4525 2292 4537 2295
rect 4028 2264 4537 2292
rect 4028 2252 4034 2264
rect 4525 2261 4537 2264
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 6932 2292 6960 2391
rect 7009 2363 7067 2369
rect 7009 2329 7021 2363
rect 7055 2360 7067 2363
rect 7208 2360 7236 2391
rect 7668 2360 7696 2391
rect 7055 2332 7236 2360
rect 7300 2332 7696 2360
rect 7760 2360 7788 2391
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 8076 2400 8125 2428
rect 8076 2388 8082 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8754 2428 8760 2440
rect 8527 2400 8760 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9324 2437 9352 2468
rect 9766 2456 9772 2508
rect 9824 2456 9830 2508
rect 9879 2499 9937 2505
rect 9879 2496 9891 2499
rect 9876 2474 9891 2496
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 7760 2332 8401 2360
rect 7055 2329 7067 2332
rect 7009 2323 7067 2329
rect 7300 2292 7328 2332
rect 4672 2264 7328 2292
rect 7377 2295 7435 2301
rect 4672 2252 4678 2264
rect 7377 2261 7389 2295
rect 7423 2292 7435 2295
rect 7558 2292 7564 2304
rect 7423 2264 7564 2292
rect 7423 2261 7435 2264
rect 7377 2255 7435 2261
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 7668 2292 7696 2332
rect 8389 2329 8401 2332
rect 8435 2360 8447 2363
rect 8846 2360 8852 2372
rect 8435 2332 8852 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 9140 2360 9168 2391
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9684 2431 9742 2437
rect 9684 2428 9696 2431
rect 9548 2400 9696 2428
rect 9548 2388 9554 2400
rect 9684 2397 9696 2400
rect 9730 2397 9742 2431
rect 9858 2422 9864 2474
rect 9925 2465 9937 2499
rect 9916 2459 9937 2465
rect 10704 2496 10732 2604
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12526 2632 12532 2644
rect 12483 2604 12532 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13412 2604 13461 2632
rect 13412 2592 13418 2604
rect 13449 2601 13461 2604
rect 13495 2632 13507 2635
rect 14274 2632 14280 2644
rect 13495 2604 14280 2632
rect 13495 2601 13507 2604
rect 13449 2595 13507 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14645 2635 14703 2641
rect 14645 2601 14657 2635
rect 14691 2632 14703 2635
rect 15286 2632 15292 2644
rect 14691 2604 15292 2632
rect 14691 2601 14703 2604
rect 14645 2595 14703 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 15562 2592 15568 2644
rect 15620 2592 15626 2644
rect 16393 2635 16451 2641
rect 16393 2601 16405 2635
rect 16439 2632 16451 2635
rect 16942 2632 16948 2644
rect 16439 2604 16948 2632
rect 16439 2601 16451 2604
rect 16393 2595 16451 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 17770 2592 17776 2644
rect 17828 2592 17834 2644
rect 20346 2632 20352 2644
rect 19306 2604 20352 2632
rect 12989 2567 13047 2573
rect 12989 2533 13001 2567
rect 13035 2564 13047 2567
rect 13035 2536 13676 2564
rect 13035 2533 13047 2536
rect 12989 2527 13047 2533
rect 13648 2505 13676 2536
rect 13722 2524 13728 2576
rect 13780 2524 13786 2576
rect 15102 2564 15108 2576
rect 14752 2536 15108 2564
rect 12621 2499 12679 2505
rect 10704 2468 12112 2496
rect 9916 2422 9922 2459
rect 9684 2391 9742 2397
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10704 2437 10732 2468
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 10870 2388 10876 2440
rect 10928 2388 10934 2440
rect 10962 2388 10968 2440
rect 11020 2388 11026 2440
rect 11164 2437 11192 2468
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 9582 2360 9588 2372
rect 9140 2332 9588 2360
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11532 2360 11560 2391
rect 11103 2332 11560 2360
rect 12084 2360 12112 2468
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13633 2499 13691 2505
rect 12667 2468 13124 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 12216 2400 12265 2428
rect 12216 2388 12222 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12492 2400 12541 2428
rect 12492 2388 12498 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 12710 2388 12716 2440
rect 12768 2388 12774 2440
rect 13096 2437 13124 2468
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 13740 2496 13768 2524
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13740 2468 13829 2496
rect 13633 2459 13691 2465
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 14182 2496 14188 2508
rect 13817 2459 13875 2465
rect 13924 2468 14188 2496
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 13924 2428 13952 2468
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14752 2496 14780 2536
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 17218 2564 17224 2576
rect 16132 2536 17224 2564
rect 14292 2468 14780 2496
rect 13771 2400 13952 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 12728 2360 12756 2388
rect 12084 2332 12756 2360
rect 12820 2360 12848 2391
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14292 2428 14320 2468
rect 14148 2400 14320 2428
rect 14148 2388 14154 2400
rect 14366 2388 14372 2440
rect 14424 2388 14430 2440
rect 14752 2437 14780 2468
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 14875 2468 15056 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 13998 2360 14004 2372
rect 12820 2332 14004 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 13998 2320 14004 2332
rect 14056 2320 14062 2372
rect 14274 2320 14280 2372
rect 14332 2320 14338 2372
rect 14476 2360 14504 2391
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15028 2437 15056 2468
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15746 2388 15752 2440
rect 15804 2388 15810 2440
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 15930 2428 15936 2440
rect 15887 2400 15936 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 16132 2437 16160 2536
rect 17218 2524 17224 2536
rect 17276 2564 17282 2576
rect 17862 2564 17868 2576
rect 17276 2536 17868 2564
rect 17276 2524 17282 2536
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 19306 2564 19334 2604
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 21453 2635 21511 2641
rect 21453 2632 21465 2635
rect 20496 2604 21465 2632
rect 20496 2592 20502 2604
rect 21453 2601 21465 2604
rect 21499 2601 21511 2635
rect 21453 2595 21511 2601
rect 22002 2592 22008 2644
rect 22060 2592 22066 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 22336 2604 23673 2632
rect 22336 2592 22342 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 24121 2635 24179 2641
rect 24121 2601 24133 2635
rect 24167 2632 24179 2635
rect 25958 2632 25964 2644
rect 24167 2604 25964 2632
rect 24167 2601 24179 2604
rect 24121 2595 24179 2601
rect 25958 2592 25964 2604
rect 26016 2592 26022 2644
rect 26510 2592 26516 2644
rect 26568 2592 26574 2644
rect 21634 2564 21640 2576
rect 18892 2536 19334 2564
rect 21284 2536 21640 2564
rect 17494 2456 17500 2508
rect 17552 2456 17558 2508
rect 17589 2499 17647 2505
rect 17589 2465 17601 2499
rect 17635 2496 17647 2499
rect 18782 2496 18788 2508
rect 17635 2468 18788 2496
rect 17635 2465 17647 2468
rect 17589 2459 17647 2465
rect 18782 2456 18788 2468
rect 18840 2456 18846 2508
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 17405 2431 17463 2437
rect 17405 2397 17417 2431
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 14476 2332 15332 2360
rect 7834 2292 7840 2304
rect 7668 2264 7840 2292
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 8662 2252 8668 2304
rect 8720 2252 8726 2304
rect 9214 2252 9220 2304
rect 9272 2252 9278 2304
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 10229 2295 10287 2301
rect 10229 2292 10241 2295
rect 9456 2264 10241 2292
rect 9456 2252 9462 2264
rect 10229 2261 10241 2264
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 10410 2252 10416 2304
rect 10468 2252 10474 2304
rect 10778 2252 10784 2304
rect 10836 2252 10842 2304
rect 11238 2252 11244 2304
rect 11296 2292 11302 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11296 2264 11713 2292
rect 11296 2252 11302 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13136 2264 13277 2292
rect 13136 2252 13142 2264
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 14976 2264 15209 2292
rect 14976 2252 14982 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15304 2292 15332 2332
rect 16022 2320 16028 2372
rect 16080 2320 16086 2372
rect 16298 2320 16304 2372
rect 16356 2360 16362 2372
rect 17420 2360 17448 2391
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 18230 2388 18236 2440
rect 18288 2388 18294 2440
rect 18892 2428 18920 2536
rect 19242 2456 19248 2508
rect 19300 2456 19306 2508
rect 21284 2505 21312 2536
rect 21634 2524 21640 2536
rect 21692 2524 21698 2576
rect 22296 2536 23244 2564
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2465 21327 2499
rect 22186 2496 22192 2508
rect 21269 2459 21327 2465
rect 21652 2468 22192 2496
rect 18340 2400 18920 2428
rect 16356 2332 17448 2360
rect 18049 2363 18107 2369
rect 16356 2320 16362 2332
rect 18049 2329 18061 2363
rect 18095 2329 18107 2363
rect 18049 2323 18107 2329
rect 16206 2292 16212 2304
rect 15304 2264 16212 2292
rect 15197 2255 15255 2261
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 18064 2292 18092 2323
rect 18138 2320 18144 2372
rect 18196 2320 18202 2372
rect 18340 2292 18368 2400
rect 18966 2388 18972 2440
rect 19024 2388 19030 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 21652 2437 21680 2468
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 21637 2431 21695 2437
rect 19392 2400 19918 2428
rect 19392 2388 19398 2400
rect 21637 2397 21649 2431
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 22296 2428 22324 2536
rect 22370 2456 22376 2508
rect 22428 2496 22434 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22428 2468 23029 2496
rect 22428 2456 22434 2468
rect 22664 2437 22692 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23216 2496 23244 2536
rect 23382 2524 23388 2576
rect 23440 2524 23446 2576
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 24578 2564 24584 2576
rect 23532 2536 24584 2564
rect 23532 2524 23538 2536
rect 24578 2524 24584 2536
rect 24636 2524 24642 2576
rect 24854 2524 24860 2576
rect 24912 2564 24918 2576
rect 25866 2564 25872 2576
rect 24912 2536 25872 2564
rect 24912 2524 24918 2536
rect 24118 2496 24124 2508
rect 23216 2468 24124 2496
rect 23017 2459 23075 2465
rect 24118 2456 24124 2468
rect 24176 2456 24182 2508
rect 25130 2456 25136 2508
rect 25188 2496 25194 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 25188 2468 25605 2496
rect 25188 2456 25194 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 25792 2496 25820 2536
rect 25866 2524 25872 2536
rect 25924 2524 25930 2576
rect 26145 2499 26203 2505
rect 26145 2496 26157 2499
rect 25792 2468 26157 2496
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 22296 2400 22477 2428
rect 21821 2391 21879 2397
rect 22465 2397 22477 2400
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 20993 2363 21051 2369
rect 18432 2332 19656 2360
rect 18432 2301 18460 2332
rect 17184 2264 18368 2292
rect 18417 2295 18475 2301
rect 17184 2252 17190 2264
rect 18417 2261 18429 2295
rect 18463 2261 18475 2295
rect 18417 2255 18475 2261
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18656 2264 18797 2292
rect 18656 2252 18662 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 19628 2292 19656 2332
rect 20993 2329 21005 2363
rect 21039 2329 21051 2363
rect 20993 2323 21051 2329
rect 21008 2292 21036 2323
rect 21358 2320 21364 2372
rect 21416 2360 21422 2372
rect 21836 2360 21864 2391
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 21416 2332 21864 2360
rect 21416 2320 21422 2332
rect 22554 2320 22560 2372
rect 22612 2320 22618 2372
rect 22787 2363 22845 2369
rect 22787 2329 22799 2363
rect 22833 2329 22845 2363
rect 23860 2360 23888 2391
rect 23934 2388 23940 2440
rect 23992 2388 23998 2440
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 24084 2400 24409 2428
rect 24084 2388 24090 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 25317 2431 25375 2437
rect 25317 2397 25329 2431
rect 25363 2428 25375 2431
rect 25406 2428 25412 2440
rect 25363 2400 25412 2428
rect 25363 2397 25375 2400
rect 25317 2391 25375 2397
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 25792 2437 25820 2468
rect 26145 2465 26157 2468
rect 26191 2465 26203 2499
rect 26145 2459 26203 2465
rect 26252 2468 26648 2496
rect 25777 2431 25835 2437
rect 25777 2397 25789 2431
rect 25823 2397 25835 2431
rect 26252 2428 26280 2468
rect 25777 2391 25835 2397
rect 25884 2400 26280 2428
rect 26329 2431 26387 2437
rect 25516 2360 25544 2388
rect 25884 2360 25912 2400
rect 26329 2397 26341 2431
rect 26375 2428 26387 2431
rect 26510 2428 26516 2440
rect 26375 2400 26516 2428
rect 26375 2397 26387 2400
rect 26329 2391 26387 2397
rect 26510 2388 26516 2400
rect 26568 2388 26574 2440
rect 26620 2437 26648 2468
rect 26605 2431 26663 2437
rect 26605 2397 26617 2431
rect 26651 2397 26663 2431
rect 26605 2391 26663 2397
rect 26786 2388 26792 2440
rect 26844 2388 26850 2440
rect 23860 2332 25452 2360
rect 25516 2332 25912 2360
rect 25961 2363 26019 2369
rect 22787 2323 22845 2329
rect 19628 2264 21036 2292
rect 18785 2255 18843 2261
rect 21082 2252 21088 2304
rect 21140 2292 21146 2304
rect 22281 2295 22339 2301
rect 22281 2292 22293 2295
rect 21140 2264 22293 2292
rect 21140 2252 21146 2264
rect 22281 2261 22293 2264
rect 22327 2261 22339 2295
rect 22802 2292 22830 2323
rect 23474 2292 23480 2304
rect 22802 2264 23480 2292
rect 22281 2255 22339 2261
rect 23474 2252 23480 2264
rect 23532 2252 23538 2304
rect 24210 2252 24216 2304
rect 24268 2292 24274 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24268 2264 24593 2292
rect 24268 2252 24274 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24946 2252 24952 2304
rect 25004 2292 25010 2304
rect 25424 2301 25452 2332
rect 25961 2329 25973 2363
rect 26007 2360 26019 2363
rect 27157 2363 27215 2369
rect 27157 2360 27169 2363
rect 26007 2332 27169 2360
rect 26007 2329 26019 2332
rect 25961 2323 26019 2329
rect 27157 2329 27169 2332
rect 27203 2329 27215 2363
rect 27157 2323 27215 2329
rect 27525 2363 27583 2369
rect 27525 2329 27537 2363
rect 27571 2360 27583 2363
rect 27798 2360 27804 2372
rect 27571 2332 27804 2360
rect 27571 2329 27583 2332
rect 27525 2323 27583 2329
rect 27798 2320 27804 2332
rect 27856 2320 27862 2372
rect 25041 2295 25099 2301
rect 25041 2292 25053 2295
rect 25004 2264 25053 2292
rect 25004 2252 25010 2264
rect 25041 2261 25053 2264
rect 25087 2261 25099 2295
rect 25041 2255 25099 2261
rect 25409 2295 25467 2301
rect 25409 2261 25421 2295
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 26694 2252 26700 2304
rect 26752 2252 26758 2304
rect 1104 2202 27876 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 27876 2202
rect 1104 2128 27876 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 2372 2060 5304 2088
rect 2372 2048 2378 2060
rect 1670 1980 1676 2032
rect 1728 2020 1734 2032
rect 5276 2020 5304 2060
rect 6086 2048 6092 2100
rect 6144 2088 6150 2100
rect 10778 2088 10784 2100
rect 6144 2060 10784 2088
rect 6144 2048 6150 2060
rect 10778 2048 10784 2060
rect 10836 2048 10842 2100
rect 11698 2048 11704 2100
rect 11756 2088 11762 2100
rect 14274 2088 14280 2100
rect 11756 2060 14280 2088
rect 11756 2048 11762 2060
rect 14274 2048 14280 2060
rect 14332 2088 14338 2100
rect 16022 2088 16028 2100
rect 14332 2060 16028 2088
rect 14332 2048 14338 2060
rect 16022 2048 16028 2060
rect 16080 2088 16086 2100
rect 17126 2088 17132 2100
rect 16080 2060 17132 2088
rect 16080 2048 16086 2060
rect 17126 2048 17132 2060
rect 17184 2048 17190 2100
rect 19058 2048 19064 2100
rect 19116 2088 19122 2100
rect 19116 2060 22094 2088
rect 19116 2048 19122 2060
rect 7742 2020 7748 2032
rect 1728 1992 2774 2020
rect 5276 1992 7748 2020
rect 1728 1980 1734 1992
rect 2746 1952 2774 1992
rect 7742 1980 7748 1992
rect 7800 1980 7806 2032
rect 7834 1980 7840 2032
rect 7892 2020 7898 2032
rect 12618 2020 12624 2032
rect 7892 1992 12624 2020
rect 7892 1980 7898 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 2746 1924 5304 1952
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 5276 1884 5304 1924
rect 5626 1912 5632 1964
rect 5684 1952 5690 1964
rect 21082 1952 21088 1964
rect 5684 1924 21088 1952
rect 5684 1912 5690 1924
rect 21082 1912 21088 1924
rect 21140 1912 21146 1964
rect 22066 1952 22094 2060
rect 23382 2048 23388 2100
rect 23440 2088 23446 2100
rect 27062 2088 27068 2100
rect 23440 2060 27068 2088
rect 23440 2048 23446 2060
rect 27062 2048 27068 2060
rect 27120 2048 27126 2100
rect 22186 1980 22192 2032
rect 22244 2020 22250 2032
rect 26694 2020 26700 2032
rect 22244 1992 26700 2020
rect 22244 1980 22250 1992
rect 26694 1980 26700 1992
rect 26752 1980 26758 2032
rect 25498 1952 25504 1964
rect 22066 1924 25504 1952
rect 25498 1912 25504 1924
rect 25556 1912 25562 1964
rect 10686 1884 10692 1896
rect 2464 1856 5120 1884
rect 5276 1856 10692 1884
rect 2464 1844 2470 1856
rect 2222 1774 2228 1826
rect 2280 1814 2286 1826
rect 2280 1786 4704 1814
rect 2280 1774 2286 1786
rect 4676 1604 4704 1786
rect 5092 1748 5120 1856
rect 10686 1844 10692 1856
rect 10744 1844 10750 1896
rect 16206 1844 16212 1896
rect 16264 1884 16270 1896
rect 18230 1884 18236 1896
rect 16264 1856 18236 1884
rect 16264 1844 16270 1856
rect 18230 1844 18236 1856
rect 18288 1884 18294 1896
rect 22554 1884 22560 1896
rect 18288 1856 22560 1884
rect 18288 1844 18294 1856
rect 22554 1844 22560 1856
rect 22612 1844 22618 1896
rect 9122 1776 9128 1828
rect 9180 1816 9186 1828
rect 27154 1816 27160 1828
rect 9180 1788 27160 1816
rect 9180 1776 9186 1788
rect 27154 1776 27160 1788
rect 27212 1776 27218 1828
rect 8570 1748 8576 1760
rect 5092 1720 8576 1748
rect 8570 1708 8576 1720
rect 8628 1708 8634 1760
rect 9950 1708 9956 1760
rect 10008 1748 10014 1760
rect 26234 1748 26240 1750
rect 10008 1720 26240 1748
rect 10008 1708 10014 1720
rect 26234 1698 26240 1720
rect 26292 1698 26298 1750
rect 4798 1636 4804 1688
rect 4856 1676 4862 1688
rect 5258 1676 5264 1688
rect 4856 1648 5264 1676
rect 4856 1636 4862 1648
rect 5258 1636 5264 1648
rect 5316 1636 5322 1688
rect 9490 1640 9496 1692
rect 9548 1680 9554 1692
rect 10410 1680 10416 1692
rect 9548 1652 10416 1680
rect 9548 1640 9554 1652
rect 10410 1640 10416 1652
rect 10468 1640 10474 1692
rect 22094 1630 22100 1682
rect 22152 1670 22158 1682
rect 26786 1670 26792 1682
rect 22152 1642 26792 1670
rect 22152 1630 22158 1642
rect 26786 1630 26792 1642
rect 26844 1630 26850 1682
rect 17034 1604 17040 1616
rect 4676 1576 17040 1604
rect 17034 1564 17040 1576
rect 17092 1564 17098 1616
<< via1 >>
rect 18236 7964 18288 8016
rect 26976 7964 27028 8016
rect 7472 7896 7524 7948
rect 27344 7896 27396 7948
rect 10324 7828 10376 7880
rect 25044 7828 25096 7880
rect 7012 7760 7064 7812
rect 8208 7760 8260 7812
rect 11336 7760 11388 7812
rect 15200 7760 15252 7812
rect 20444 7760 20496 7812
rect 1216 7692 1268 7744
rect 2688 7692 2740 7744
rect 2872 7692 2924 7744
rect 17960 7692 18012 7744
rect 18972 7692 19024 7744
rect 26516 7692 26568 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1124 7488 1176 7540
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 1308 7420 1360 7472
rect 2780 7420 2832 7472
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 4620 7352 4672 7404
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 4344 7284 4396 7336
rect 4712 7216 4764 7268
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 3700 7148 3752 7200
rect 6092 7531 6144 7540
rect 6092 7497 6101 7531
rect 6101 7497 6135 7531
rect 6135 7497 6144 7531
rect 6092 7488 6144 7497
rect 6184 7420 6236 7472
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 7564 7463 7616 7472
rect 7564 7429 7573 7463
rect 7573 7429 7607 7463
rect 7607 7429 7616 7463
rect 7564 7420 7616 7429
rect 6644 7352 6696 7404
rect 10876 7488 10928 7540
rect 13268 7488 13320 7540
rect 15292 7488 15344 7540
rect 9036 7420 9088 7472
rect 6276 7284 6328 7336
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 10876 7352 10928 7404
rect 11244 7420 11296 7472
rect 12440 7420 12492 7472
rect 13820 7420 13872 7472
rect 9772 7284 9824 7336
rect 10784 7284 10836 7336
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 12348 7352 12400 7361
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 14188 7284 14240 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 17776 7352 17828 7404
rect 19064 7420 19116 7472
rect 18052 7352 18104 7404
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18880 7284 18932 7336
rect 7012 7148 7064 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 9956 7148 10008 7200
rect 10508 7148 10560 7200
rect 12440 7148 12492 7200
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 14280 7216 14332 7268
rect 15292 7148 15344 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 15752 7148 15804 7200
rect 17224 7148 17276 7200
rect 17868 7216 17920 7268
rect 17960 7259 18012 7268
rect 17960 7225 17969 7259
rect 17969 7225 18003 7259
rect 18003 7225 18012 7259
rect 17960 7216 18012 7225
rect 18236 7216 18288 7268
rect 19800 7327 19852 7336
rect 19800 7293 19809 7327
rect 19809 7293 19843 7327
rect 19843 7293 19852 7327
rect 19800 7284 19852 7293
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 20812 7284 20864 7336
rect 23296 7395 23348 7404
rect 23296 7361 23305 7395
rect 23305 7361 23339 7395
rect 23339 7361 23348 7395
rect 23296 7352 23348 7361
rect 26700 7531 26752 7540
rect 26700 7497 26709 7531
rect 26709 7497 26743 7531
rect 26743 7497 26752 7531
rect 26700 7488 26752 7497
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 27436 7531 27488 7540
rect 27436 7497 27445 7531
rect 27445 7497 27479 7531
rect 27479 7497 27488 7531
rect 27436 7488 27488 7497
rect 23480 7420 23532 7472
rect 23848 7395 23900 7404
rect 23848 7361 23856 7395
rect 23856 7361 23890 7395
rect 23890 7361 23900 7395
rect 23848 7352 23900 7361
rect 24032 7352 24084 7404
rect 25228 7352 25280 7404
rect 26516 7395 26568 7404
rect 26516 7361 26525 7395
rect 26525 7361 26559 7395
rect 26559 7361 26568 7395
rect 26516 7352 26568 7361
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 25136 7284 25188 7336
rect 25688 7327 25740 7336
rect 25688 7293 25697 7327
rect 25697 7293 25731 7327
rect 25731 7293 25740 7327
rect 25688 7284 25740 7293
rect 26148 7284 26200 7336
rect 26332 7284 26384 7336
rect 23480 7216 23532 7268
rect 23848 7216 23900 7268
rect 25228 7216 25280 7268
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 21088 7148 21140 7200
rect 22928 7148 22980 7200
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 23940 7148 23992 7200
rect 26056 7191 26108 7200
rect 26056 7157 26065 7191
rect 26065 7157 26099 7191
rect 26099 7157 26108 7191
rect 26056 7148 26108 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1860 6987 1912 6996
rect 1860 6953 1869 6987
rect 1869 6953 1903 6987
rect 1903 6953 1912 6987
rect 1860 6944 1912 6953
rect 4252 6944 4304 6996
rect 2688 6876 2740 6928
rect 5540 6944 5592 6996
rect 7196 6944 7248 6996
rect 7380 6944 7432 6996
rect 9036 6944 9088 6996
rect 9312 6944 9364 6996
rect 9680 6944 9732 6996
rect 10508 6944 10560 6996
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 10876 6944 10928 6996
rect 11152 6944 11204 6996
rect 5816 6876 5868 6928
rect 2136 6808 2188 6860
rect 5632 6808 5684 6860
rect 2228 6740 2280 6792
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 6092 6740 6144 6792
rect 6552 6740 6604 6792
rect 4436 6715 4488 6724
rect 4436 6681 4445 6715
rect 4445 6681 4479 6715
rect 4479 6681 4488 6715
rect 4436 6672 4488 6681
rect 5816 6672 5868 6724
rect 10508 6740 10560 6792
rect 11060 6740 11112 6792
rect 11336 6808 11388 6860
rect 12716 6808 12768 6860
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 1216 6604 1268 6656
rect 5724 6604 5776 6656
rect 9680 6672 9732 6724
rect 6276 6604 6328 6656
rect 8300 6604 8352 6656
rect 10600 6604 10652 6656
rect 11980 6715 12032 6724
rect 11980 6681 11989 6715
rect 11989 6681 12023 6715
rect 12023 6681 12032 6715
rect 11980 6672 12032 6681
rect 14188 6987 14240 6996
rect 14188 6953 14197 6987
rect 14197 6953 14231 6987
rect 14231 6953 14240 6987
rect 14188 6944 14240 6953
rect 14556 6944 14608 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 13268 6808 13320 6860
rect 15568 6808 15620 6860
rect 18328 6919 18380 6928
rect 18328 6885 18337 6919
rect 18337 6885 18371 6919
rect 18371 6885 18380 6919
rect 18328 6876 18380 6885
rect 13360 6740 13412 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 18604 6808 18656 6860
rect 20076 6944 20128 6996
rect 22652 6944 22704 6996
rect 26332 6944 26384 6996
rect 18880 6876 18932 6928
rect 14280 6672 14332 6724
rect 15384 6672 15436 6724
rect 12808 6604 12860 6656
rect 13360 6604 13412 6656
rect 16304 6715 16356 6724
rect 16304 6681 16313 6715
rect 16313 6681 16347 6715
rect 16347 6681 16356 6715
rect 16304 6672 16356 6681
rect 18512 6740 18564 6792
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 19616 6740 19668 6792
rect 19708 6783 19760 6792
rect 19708 6749 19717 6783
rect 19717 6749 19751 6783
rect 19751 6749 19760 6783
rect 19708 6740 19760 6749
rect 21180 6851 21232 6860
rect 21180 6817 21189 6851
rect 21189 6817 21223 6851
rect 21223 6817 21232 6851
rect 21180 6808 21232 6817
rect 21824 6851 21876 6860
rect 21824 6817 21833 6851
rect 21833 6817 21867 6851
rect 21867 6817 21876 6851
rect 21824 6808 21876 6817
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 22744 6808 22796 6860
rect 20076 6740 20128 6792
rect 23848 6808 23900 6860
rect 24676 6808 24728 6860
rect 17960 6604 18012 6656
rect 19156 6672 19208 6724
rect 19984 6715 20036 6724
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 22376 6672 22428 6724
rect 22928 6672 22980 6724
rect 23112 6672 23164 6724
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 19340 6604 19392 6656
rect 19524 6604 19576 6656
rect 20904 6647 20956 6656
rect 20904 6613 20913 6647
rect 20913 6613 20947 6647
rect 20947 6613 20956 6647
rect 20904 6604 20956 6613
rect 20996 6647 21048 6656
rect 20996 6613 21005 6647
rect 21005 6613 21039 6647
rect 21039 6613 21048 6647
rect 20996 6604 21048 6613
rect 22560 6604 22612 6656
rect 23388 6604 23440 6656
rect 24400 6783 24452 6792
rect 24400 6749 24409 6783
rect 24409 6749 24443 6783
rect 24443 6749 24452 6783
rect 24400 6740 24452 6749
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 24952 6672 25004 6724
rect 25136 6672 25188 6724
rect 25964 6672 26016 6724
rect 27620 6808 27672 6860
rect 26884 6783 26936 6792
rect 26884 6749 26893 6783
rect 26893 6749 26927 6783
rect 26927 6749 26936 6783
rect 26884 6740 26936 6749
rect 25504 6604 25556 6656
rect 26148 6647 26200 6656
rect 26148 6613 26157 6647
rect 26157 6613 26191 6647
rect 26191 6613 26200 6647
rect 26148 6604 26200 6613
rect 26332 6647 26384 6656
rect 26332 6613 26341 6647
rect 26341 6613 26375 6647
rect 26375 6613 26384 6647
rect 26332 6604 26384 6613
rect 27068 6647 27120 6656
rect 27068 6613 27077 6647
rect 27077 6613 27111 6647
rect 27111 6613 27120 6647
rect 27068 6604 27120 6613
rect 27528 6604 27580 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1308 6400 1360 6452
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 3792 6196 3844 6248
rect 1240 6128 1292 6180
rect 3608 6128 3660 6180
rect 4252 6332 4304 6384
rect 4436 6400 4488 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5724 6400 5776 6452
rect 7656 6400 7708 6452
rect 8116 6400 8168 6452
rect 5540 6332 5592 6384
rect 8668 6332 8720 6384
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 9680 6400 9732 6452
rect 10600 6400 10652 6452
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 11244 6400 11296 6452
rect 11980 6400 12032 6452
rect 12532 6400 12584 6452
rect 14096 6400 14148 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 14832 6400 14884 6452
rect 15384 6400 15436 6452
rect 15660 6400 15712 6452
rect 16304 6400 16356 6452
rect 9772 6332 9824 6384
rect 5356 6264 5408 6316
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 8116 6307 8168 6316
rect 4804 6196 4856 6248
rect 4712 6128 4764 6180
rect 5540 6196 5592 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8484 6264 8536 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 5816 6196 5868 6205
rect 6368 6196 6420 6248
rect 6736 6239 6788 6248
rect 6736 6205 6745 6239
rect 6745 6205 6779 6239
rect 6779 6205 6788 6239
rect 6736 6196 6788 6205
rect 9404 6264 9456 6316
rect 10508 6332 10560 6384
rect 11520 6332 11572 6384
rect 12256 6332 12308 6384
rect 9312 6196 9364 6248
rect 9496 6196 9548 6248
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 11888 6264 11940 6316
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 10968 6196 11020 6248
rect 12348 6196 12400 6248
rect 13084 6264 13136 6316
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13360 6332 13412 6384
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 15292 6264 15344 6316
rect 16580 6332 16632 6384
rect 17684 6332 17736 6384
rect 17776 6375 17828 6384
rect 17776 6341 17785 6375
rect 17785 6341 17819 6375
rect 17819 6341 17828 6375
rect 17776 6332 17828 6341
rect 15752 6264 15804 6316
rect 15844 6264 15896 6316
rect 16488 6264 16540 6316
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 18052 6400 18104 6452
rect 19156 6400 19208 6452
rect 19340 6400 19392 6452
rect 20260 6400 20312 6452
rect 21180 6400 21232 6452
rect 18328 6375 18380 6384
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 19432 6264 19484 6316
rect 19984 6264 20036 6316
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22836 6332 22888 6384
rect 22376 6264 22428 6273
rect 22560 6307 22612 6316
rect 22560 6273 22569 6307
rect 22569 6273 22603 6307
rect 22603 6273 22612 6307
rect 22560 6264 22612 6273
rect 23296 6400 23348 6452
rect 24860 6400 24912 6452
rect 24952 6443 25004 6452
rect 24952 6409 24961 6443
rect 24961 6409 24995 6443
rect 24995 6409 25004 6443
rect 24952 6400 25004 6409
rect 26056 6400 26108 6452
rect 27436 6443 27488 6452
rect 27436 6409 27445 6443
rect 27445 6409 27479 6443
rect 27479 6409 27488 6443
rect 27436 6400 27488 6409
rect 23388 6375 23440 6384
rect 23388 6341 23397 6375
rect 23397 6341 23431 6375
rect 23431 6341 23440 6375
rect 23388 6332 23440 6341
rect 24124 6332 24176 6384
rect 6276 6128 6328 6180
rect 6184 6060 6236 6112
rect 7840 6060 7892 6112
rect 8576 6060 8628 6112
rect 8944 6060 8996 6112
rect 9404 6128 9456 6180
rect 12716 6128 12768 6180
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 16028 6196 16080 6248
rect 14372 6128 14424 6180
rect 14556 6128 14608 6180
rect 16120 6128 16172 6180
rect 12164 6060 12216 6112
rect 12348 6060 12400 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 14740 6060 14792 6112
rect 14924 6060 14976 6112
rect 15292 6060 15344 6112
rect 15660 6060 15712 6112
rect 16488 6060 16540 6112
rect 17132 6060 17184 6112
rect 17960 6128 18012 6180
rect 19892 6128 19944 6180
rect 21824 6196 21876 6248
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 23848 6196 23900 6248
rect 26332 6332 26384 6384
rect 25412 6264 25464 6316
rect 27252 6307 27304 6316
rect 27252 6273 27261 6307
rect 27261 6273 27295 6307
rect 27295 6273 27304 6307
rect 27252 6264 27304 6273
rect 25504 6239 25556 6248
rect 25504 6205 25513 6239
rect 25513 6205 25547 6239
rect 25547 6205 25556 6239
rect 25504 6196 25556 6205
rect 26332 6196 26384 6248
rect 22192 6060 22244 6112
rect 22284 6060 22336 6112
rect 24400 6060 24452 6112
rect 25228 6060 25280 6112
rect 26700 6103 26752 6112
rect 26700 6069 26709 6103
rect 26709 6069 26743 6103
rect 26743 6069 26752 6103
rect 26700 6060 26752 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 4436 5856 4488 5908
rect 5356 5856 5408 5908
rect 5448 5856 5500 5908
rect 5816 5856 5868 5908
rect 1172 5788 1224 5840
rect 3884 5788 3936 5840
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2872 5652 2924 5704
rect 3240 5652 3292 5704
rect 4068 5720 4120 5772
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 3976 5652 4028 5704
rect 4988 5788 5040 5840
rect 5908 5788 5960 5840
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7748 5856 7800 5908
rect 6920 5788 6972 5840
rect 7288 5788 7340 5840
rect 4528 5652 4580 5704
rect 6736 5720 6788 5772
rect 8760 5856 8812 5908
rect 9036 5856 9088 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 9588 5856 9640 5908
rect 12072 5856 12124 5908
rect 12624 5856 12676 5908
rect 12716 5856 12768 5908
rect 13452 5856 13504 5908
rect 13820 5856 13872 5908
rect 14004 5856 14056 5908
rect 15568 5856 15620 5908
rect 16948 5856 17000 5908
rect 3884 5584 3936 5636
rect 5264 5652 5316 5704
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 5724 5652 5776 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 8944 5720 8996 5772
rect 10140 5788 10192 5840
rect 10600 5788 10652 5840
rect 7196 5652 7248 5704
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8208 5652 8260 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 6184 5584 6236 5636
rect 4068 5516 4120 5568
rect 4804 5516 4856 5568
rect 5816 5516 5868 5568
rect 6368 5516 6420 5568
rect 6644 5516 6696 5568
rect 7840 5516 7892 5568
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 10968 5720 11020 5772
rect 11704 5720 11756 5772
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 9680 5652 9732 5661
rect 11152 5584 11204 5636
rect 11612 5584 11664 5636
rect 8668 5516 8720 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 12808 5720 12860 5772
rect 13084 5788 13136 5840
rect 13176 5788 13228 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 12992 5516 13044 5568
rect 13360 5652 13412 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 16488 5788 16540 5840
rect 15476 5720 15528 5772
rect 15752 5720 15804 5772
rect 17500 5788 17552 5840
rect 18052 5788 18104 5840
rect 19708 5856 19760 5908
rect 14096 5652 14148 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 15108 5652 15160 5704
rect 15844 5652 15896 5704
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16580 5652 16632 5704
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 18328 5763 18380 5772
rect 18328 5729 18337 5763
rect 18337 5729 18371 5763
rect 18371 5729 18380 5763
rect 18328 5720 18380 5729
rect 18512 5788 18564 5840
rect 23480 5856 23532 5908
rect 24308 5856 24360 5908
rect 27436 5899 27488 5908
rect 27436 5865 27445 5899
rect 27445 5865 27479 5899
rect 27479 5865 27488 5899
rect 27436 5856 27488 5865
rect 14004 5584 14056 5636
rect 14280 5584 14332 5636
rect 14648 5627 14700 5636
rect 14648 5593 14657 5627
rect 14657 5593 14691 5627
rect 14691 5593 14700 5627
rect 14648 5584 14700 5593
rect 16856 5627 16908 5636
rect 13176 5516 13228 5568
rect 14188 5516 14240 5568
rect 15568 5516 15620 5568
rect 16856 5593 16874 5627
rect 16874 5593 16908 5627
rect 16856 5584 16908 5593
rect 17132 5584 17184 5636
rect 17224 5584 17276 5636
rect 17868 5652 17920 5704
rect 18144 5652 18196 5704
rect 18236 5652 18288 5704
rect 18788 5652 18840 5704
rect 23756 5788 23808 5840
rect 24216 5788 24268 5840
rect 19156 5720 19208 5772
rect 19340 5652 19392 5704
rect 17592 5627 17644 5636
rect 17592 5593 17610 5627
rect 17610 5593 17644 5627
rect 17592 5584 17644 5593
rect 19064 5627 19116 5636
rect 19064 5593 19073 5627
rect 19073 5593 19107 5627
rect 19107 5593 19116 5627
rect 19892 5695 19944 5704
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 21640 5652 21692 5704
rect 24400 5763 24452 5772
rect 24400 5729 24409 5763
rect 24409 5729 24443 5763
rect 24443 5729 24452 5763
rect 24400 5720 24452 5729
rect 27068 5831 27120 5840
rect 27068 5797 27077 5831
rect 27077 5797 27111 5831
rect 27111 5797 27120 5831
rect 27068 5788 27120 5797
rect 25044 5720 25096 5772
rect 19064 5584 19116 5593
rect 20168 5627 20220 5636
rect 20168 5593 20177 5627
rect 20177 5593 20211 5627
rect 20211 5593 20220 5627
rect 20168 5584 20220 5593
rect 21456 5584 21508 5636
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 18236 5516 18288 5568
rect 19156 5516 19208 5568
rect 19340 5516 19392 5568
rect 21640 5559 21692 5568
rect 21640 5525 21649 5559
rect 21649 5525 21683 5559
rect 21683 5525 21692 5559
rect 21640 5516 21692 5525
rect 21824 5584 21876 5636
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 26240 5652 26292 5704
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 22652 5584 22704 5636
rect 22192 5516 22244 5568
rect 22376 5559 22428 5568
rect 22376 5525 22385 5559
rect 22385 5525 22419 5559
rect 22419 5525 22428 5559
rect 22376 5516 22428 5525
rect 24124 5584 24176 5636
rect 25136 5584 25188 5636
rect 23756 5516 23808 5568
rect 24860 5516 24912 5568
rect 25412 5516 25464 5568
rect 26148 5559 26200 5568
rect 26148 5525 26157 5559
rect 26157 5525 26191 5559
rect 26191 5525 26200 5559
rect 26148 5516 26200 5525
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1156 5312 1208 5364
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3792 5244 3844 5296
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3976 5176 4028 5228
rect 4160 5244 4212 5296
rect 3148 5108 3200 5160
rect 4620 5176 4672 5228
rect 4804 5176 4856 5228
rect 5172 5176 5224 5228
rect 5448 5176 5500 5228
rect 5724 5312 5776 5364
rect 5908 5244 5960 5296
rect 6000 5176 6052 5228
rect 6276 5176 6328 5228
rect 6368 5176 6420 5228
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 2688 5040 2740 5092
rect 2872 5040 2924 5092
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7748 5108 7800 5160
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8300 5312 8352 5364
rect 8116 5244 8168 5296
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10508 5312 10560 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 14096 5312 14148 5364
rect 15108 5312 15160 5364
rect 18144 5312 18196 5364
rect 8208 5176 8260 5228
rect 8300 5176 8352 5228
rect 9036 5219 9088 5228
rect 9036 5185 9044 5219
rect 9044 5185 9078 5219
rect 9078 5185 9088 5219
rect 9036 5176 9088 5185
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 10048 5244 10100 5296
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 10692 5244 10744 5296
rect 11428 5244 11480 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 12256 5244 12308 5296
rect 9772 5108 9824 5160
rect 10784 5176 10836 5228
rect 10968 5176 11020 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 10600 5108 10652 5160
rect 7932 5040 7984 5092
rect 8668 5040 8720 5092
rect 9956 5040 10008 5092
rect 10232 5040 10284 5092
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 11336 5040 11388 5092
rect 11612 5040 11664 5092
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 13176 5244 13228 5296
rect 14188 5244 14240 5296
rect 15200 5244 15252 5296
rect 15844 5244 15896 5296
rect 16580 5244 16632 5296
rect 18880 5312 18932 5364
rect 19984 5312 20036 5364
rect 20168 5312 20220 5364
rect 22284 5312 22336 5364
rect 22468 5312 22520 5364
rect 24216 5355 24268 5364
rect 24216 5321 24225 5355
rect 24225 5321 24259 5355
rect 24259 5321 24268 5355
rect 24216 5312 24268 5321
rect 24308 5312 24360 5364
rect 25780 5312 25832 5364
rect 27436 5355 27488 5364
rect 27436 5321 27445 5355
rect 27445 5321 27479 5355
rect 27479 5321 27488 5355
rect 27436 5312 27488 5321
rect 12624 5108 12676 5160
rect 14648 5176 14700 5228
rect 14740 5176 14792 5228
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 15660 5176 15712 5228
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 14096 5108 14148 5160
rect 14464 5108 14516 5160
rect 15936 5108 15988 5160
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17224 5176 17276 5228
rect 1150 4972 1202 5024
rect 2044 4972 2096 5024
rect 3332 4972 3384 5024
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 4528 4972 4580 5024
rect 4712 4972 4764 5024
rect 5264 4972 5316 5024
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 8208 4972 8260 5024
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 9128 4972 9180 5024
rect 11796 4972 11848 5024
rect 12716 4972 12768 5024
rect 15476 5040 15528 5092
rect 15660 5083 15712 5092
rect 15660 5049 15669 5083
rect 15669 5049 15703 5083
rect 15703 5049 15712 5083
rect 15660 5040 15712 5049
rect 13544 4972 13596 5024
rect 15108 4972 15160 5024
rect 16120 4972 16172 5024
rect 16396 5040 16448 5092
rect 16856 4972 16908 5024
rect 17684 5176 17736 5228
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 18512 5176 18564 5228
rect 19432 5244 19484 5296
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 22376 5244 22428 5296
rect 22652 5244 22704 5296
rect 23572 5244 23624 5296
rect 17868 5040 17920 5092
rect 18236 5040 18288 5092
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 21640 5176 21692 5228
rect 19800 5108 19852 5160
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 21456 5108 21508 5160
rect 19340 5040 19392 5092
rect 19892 5040 19944 5092
rect 21732 5108 21784 5160
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 23020 5176 23072 5228
rect 23388 5176 23440 5228
rect 24032 5244 24084 5296
rect 23848 5219 23900 5228
rect 23848 5185 23857 5219
rect 23857 5185 23891 5219
rect 23891 5185 23900 5219
rect 23848 5176 23900 5185
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 24584 5219 24636 5228
rect 24584 5185 24593 5219
rect 24593 5185 24627 5219
rect 24627 5185 24636 5219
rect 24584 5176 24636 5185
rect 21824 5040 21876 5092
rect 19064 4972 19116 5024
rect 20996 5015 21048 5024
rect 20996 4981 21005 5015
rect 21005 4981 21039 5015
rect 21039 4981 21048 5015
rect 20996 4972 21048 4981
rect 22192 5040 22244 5092
rect 24032 5108 24084 5160
rect 26148 5176 26200 5228
rect 26516 5219 26568 5228
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 27160 5176 27212 5228
rect 25044 5108 25096 5160
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 22560 4972 22612 5024
rect 24768 5040 24820 5092
rect 24860 5040 24912 5092
rect 23204 4972 23256 5024
rect 24952 4972 25004 5024
rect 26700 5015 26752 5024
rect 26700 4981 26709 5015
rect 26709 4981 26743 5015
rect 26743 4981 26752 5015
rect 26700 4972 26752 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5172 4768 5224 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 5724 4768 5776 4820
rect 7380 4768 7432 4820
rect 11612 4768 11664 4820
rect 11704 4768 11756 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 1124 4700 1176 4752
rect 4620 4700 4672 4752
rect 5816 4700 5868 4752
rect 8484 4700 8536 4752
rect 9220 4700 9272 4752
rect 9496 4700 9548 4752
rect 11152 4700 11204 4752
rect 11520 4700 11572 4752
rect 13728 4768 13780 4820
rect 14648 4768 14700 4820
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 2136 4632 2188 4684
rect 2688 4632 2740 4684
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 3884 4564 3936 4616
rect 3608 4496 3660 4548
rect 5356 4632 5408 4684
rect 4344 4564 4396 4616
rect 4896 4564 4948 4616
rect 6184 4564 6236 4616
rect 11612 4632 11664 4684
rect 7104 4564 7156 4616
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8116 4564 8168 4616
rect 8484 4564 8536 4616
rect 9588 4607 9640 4616
rect 9588 4573 9597 4607
rect 9597 4573 9631 4607
rect 9631 4573 9640 4607
rect 9588 4564 9640 4573
rect 6368 4496 6420 4548
rect 8024 4539 8076 4548
rect 8024 4505 8033 4539
rect 8033 4505 8067 4539
rect 8067 4505 8076 4539
rect 8024 4496 8076 4505
rect 8208 4539 8260 4548
rect 8208 4505 8217 4539
rect 8217 4505 8251 4539
rect 8251 4505 8260 4539
rect 8208 4496 8260 4505
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10508 4607 10560 4616
rect 10508 4573 10519 4607
rect 10519 4573 10553 4607
rect 10553 4573 10560 4607
rect 10508 4564 10560 4573
rect 10600 4564 10652 4616
rect 11796 4564 11848 4616
rect 3516 4428 3568 4480
rect 3700 4428 3752 4480
rect 4896 4428 4948 4480
rect 6000 4428 6052 4480
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7288 4428 7340 4480
rect 12164 4496 12216 4548
rect 12624 4675 12676 4684
rect 12624 4641 12633 4675
rect 12633 4641 12667 4675
rect 12667 4641 12676 4675
rect 12624 4632 12676 4641
rect 12716 4632 12768 4684
rect 15844 4743 15896 4752
rect 15844 4709 15853 4743
rect 15853 4709 15887 4743
rect 15887 4709 15896 4743
rect 15844 4700 15896 4709
rect 12440 4564 12492 4616
rect 13084 4564 13136 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 13636 4564 13688 4616
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 15292 4632 15344 4684
rect 14280 4564 14332 4616
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 15384 4564 15436 4616
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 19708 4768 19760 4820
rect 19800 4768 19852 4820
rect 20168 4768 20220 4820
rect 16120 4700 16172 4752
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16212 4564 16264 4616
rect 16672 4564 16724 4616
rect 17132 4632 17184 4684
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17684 4700 17736 4752
rect 18236 4700 18288 4752
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 18052 4564 18104 4616
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 18604 4632 18656 4684
rect 19156 4700 19208 4752
rect 18788 4607 18840 4616
rect 18788 4573 18797 4607
rect 18797 4573 18831 4607
rect 18831 4573 18840 4607
rect 18788 4564 18840 4573
rect 19892 4632 19944 4684
rect 20628 4675 20680 4684
rect 20628 4641 20637 4675
rect 20637 4641 20671 4675
rect 20671 4641 20680 4675
rect 20628 4632 20680 4641
rect 21732 4768 21784 4820
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 21088 4743 21140 4752
rect 21088 4709 21097 4743
rect 21097 4709 21131 4743
rect 21131 4709 21140 4743
rect 21088 4700 21140 4709
rect 24032 4700 24084 4752
rect 19248 4564 19300 4616
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20352 4564 20404 4616
rect 20904 4564 20956 4616
rect 9772 4428 9824 4480
rect 10876 4428 10928 4480
rect 11980 4428 12032 4480
rect 14832 4428 14884 4480
rect 15292 4428 15344 4480
rect 16120 4428 16172 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 16764 4471 16816 4480
rect 16764 4437 16773 4471
rect 16773 4437 16807 4471
rect 16807 4437 16816 4471
rect 16764 4428 16816 4437
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 17776 4428 17828 4480
rect 18420 4428 18472 4480
rect 18604 4428 18656 4480
rect 18880 4428 18932 4480
rect 19064 4428 19116 4480
rect 19156 4428 19208 4480
rect 19432 4428 19484 4480
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22744 4632 22796 4684
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 24308 4564 24360 4616
rect 27436 4811 27488 4820
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 21456 4539 21508 4548
rect 21456 4505 21465 4539
rect 21465 4505 21499 4539
rect 21499 4505 21508 4539
rect 21456 4496 21508 4505
rect 21732 4496 21784 4548
rect 22100 4496 22152 4548
rect 23204 4428 23256 4480
rect 23480 4539 23532 4548
rect 23480 4505 23489 4539
rect 23489 4505 23523 4539
rect 23523 4505 23532 4539
rect 23480 4496 23532 4505
rect 25136 4496 25188 4548
rect 27344 4564 27396 4616
rect 23664 4428 23716 4480
rect 24216 4428 24268 4480
rect 24492 4428 24544 4480
rect 26056 4428 26108 4480
rect 26332 4471 26384 4480
rect 26332 4437 26341 4471
rect 26341 4437 26375 4471
rect 26375 4437 26384 4471
rect 26332 4428 26384 4437
rect 26976 4428 27028 4480
rect 27068 4471 27120 4480
rect 27068 4437 27077 4471
rect 27077 4437 27111 4471
rect 27111 4437 27120 4471
rect 27068 4428 27120 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4068 4224 4120 4276
rect 5724 4224 5776 4276
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7472 4224 7524 4276
rect 8024 4224 8076 4276
rect 10600 4224 10652 4276
rect 4988 4156 5040 4208
rect 5264 4156 5316 4208
rect 1952 4088 2004 4140
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 2136 4088 2188 4140
rect 3608 4088 3660 4140
rect 4344 4088 4396 4140
rect 4528 4088 4580 4140
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5172 4088 5224 4140
rect 5448 4088 5500 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5724 4131 5776 4140
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 5816 4088 5868 4140
rect 6552 4131 6604 4140
rect 6552 4097 6556 4131
rect 6556 4097 6590 4131
rect 6590 4097 6604 4131
rect 3792 4020 3844 4072
rect 3976 4020 4028 4072
rect 6552 4088 6604 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6828 4088 6880 4140
rect 7380 4156 7432 4208
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 2228 3952 2280 4004
rect 6828 3952 6880 4004
rect 7012 3952 7064 4004
rect 7104 3952 7156 4004
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 9036 4156 9088 4208
rect 9864 4156 9916 4208
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 3148 3884 3200 3936
rect 5632 3884 5684 3936
rect 6644 3884 6696 3936
rect 8392 3952 8444 4004
rect 8668 4020 8720 4072
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 10692 4156 10744 4208
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 11336 4224 11388 4276
rect 12072 4224 12124 4276
rect 12164 4224 12216 4276
rect 12532 4224 12584 4276
rect 13544 4224 13596 4276
rect 17868 4224 17920 4276
rect 17960 4224 18012 4276
rect 13084 4156 13136 4208
rect 13636 4156 13688 4208
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 11796 4088 11848 4140
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 11060 4020 11112 4072
rect 11612 4020 11664 4072
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 12532 4088 12584 4140
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 13268 4020 13320 4072
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 14280 4156 14332 4208
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 15016 4156 15068 4208
rect 15200 4156 15252 4208
rect 14556 4088 14608 4140
rect 7932 3884 7984 3936
rect 9680 3952 9732 4004
rect 9956 3952 10008 4004
rect 10784 3952 10836 4004
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14280 4063 14332 4072
rect 14280 4029 14289 4063
rect 14289 4029 14323 4063
rect 14323 4029 14332 4063
rect 14280 4020 14332 4029
rect 14464 4020 14516 4072
rect 9588 3884 9640 3936
rect 13452 3884 13504 3936
rect 14924 3995 14976 4004
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 15936 4088 15988 4140
rect 16120 4131 16172 4140
rect 16396 4156 16448 4208
rect 17500 4156 17552 4208
rect 18236 4224 18288 4276
rect 19340 4224 19392 4276
rect 18420 4156 18472 4208
rect 18788 4156 18840 4208
rect 16120 4097 16159 4131
rect 16159 4097 16172 4131
rect 16120 4088 16172 4097
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 16948 4020 17000 4072
rect 17316 4088 17368 4140
rect 17684 4088 17736 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 17684 3952 17736 4004
rect 18420 4020 18472 4072
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 19064 4156 19116 4208
rect 20168 4224 20220 4276
rect 19892 4199 19944 4208
rect 19892 4165 19901 4199
rect 19901 4165 19935 4199
rect 19935 4165 19944 4199
rect 19892 4156 19944 4165
rect 22744 4224 22796 4276
rect 23296 4267 23348 4276
rect 23296 4233 23305 4267
rect 23305 4233 23339 4267
rect 23339 4233 23348 4267
rect 23296 4224 23348 4233
rect 24492 4224 24544 4276
rect 24952 4224 25004 4276
rect 26608 4224 26660 4276
rect 22560 4156 22612 4208
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19156 4131 19208 4140
rect 19156 4097 19158 4131
rect 19158 4097 19192 4131
rect 19192 4097 19208 4131
rect 19156 4088 19208 4097
rect 19248 4088 19300 4140
rect 19432 4131 19484 4140
rect 19432 4097 19441 4131
rect 19441 4097 19475 4131
rect 19475 4097 19484 4131
rect 19432 4088 19484 4097
rect 18604 4020 18656 4072
rect 21640 4088 21692 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 19340 3952 19392 4004
rect 21456 4020 21508 4072
rect 21548 4020 21600 4072
rect 22560 4020 22612 4072
rect 23020 4131 23072 4140
rect 23020 4097 23029 4131
rect 23029 4097 23063 4131
rect 23063 4097 23072 4131
rect 23020 4088 23072 4097
rect 24216 4156 24268 4208
rect 24308 4156 24360 4208
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 25320 4088 25372 4140
rect 25596 4088 25648 4140
rect 25780 4131 25832 4140
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 26148 4088 26200 4140
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 20444 3952 20496 4004
rect 14096 3884 14148 3936
rect 14372 3884 14424 3936
rect 15568 3884 15620 3936
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 17224 3884 17276 3936
rect 18144 3884 18196 3936
rect 18512 3884 18564 3936
rect 18880 3884 18932 3936
rect 19800 3927 19852 3936
rect 19800 3893 19809 3927
rect 19809 3893 19843 3927
rect 19843 3893 19852 3927
rect 19800 3884 19852 3893
rect 20628 3884 20680 3936
rect 23020 3884 23072 3936
rect 23572 3952 23624 4004
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 23940 3884 23992 3936
rect 24676 3884 24728 3936
rect 25688 3927 25740 3936
rect 25688 3893 25697 3927
rect 25697 3893 25731 3927
rect 25731 3893 25740 3927
rect 25688 3884 25740 3893
rect 25780 3884 25832 3936
rect 26240 3952 26292 4004
rect 27436 3995 27488 4004
rect 27436 3961 27445 3995
rect 27445 3961 27479 3995
rect 27479 3961 27488 3995
rect 27436 3952 27488 3961
rect 26148 3884 26200 3936
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 27068 3927 27120 3936
rect 27068 3893 27077 3927
rect 27077 3893 27111 3927
rect 27111 3893 27120 3927
rect 27068 3884 27120 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1308 3680 1360 3732
rect 3976 3680 4028 3732
rect 4436 3680 4488 3732
rect 5356 3680 5408 3732
rect 5632 3680 5684 3732
rect 5724 3680 5776 3732
rect 6184 3723 6236 3732
rect 6184 3689 6193 3723
rect 6193 3689 6227 3723
rect 6227 3689 6236 3723
rect 6184 3680 6236 3689
rect 6460 3680 6512 3732
rect 8116 3680 8168 3732
rect 8668 3680 8720 3732
rect 9312 3680 9364 3732
rect 9956 3680 10008 3732
rect 10048 3680 10100 3732
rect 10968 3680 11020 3732
rect 12624 3680 12676 3732
rect 15016 3680 15068 3732
rect 17868 3680 17920 3732
rect 19432 3680 19484 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 3240 3612 3292 3664
rect 3516 3612 3568 3664
rect 4896 3612 4948 3664
rect 2136 3544 2188 3596
rect 2780 3544 2832 3596
rect 1768 3476 1820 3528
rect 3240 3476 3292 3528
rect 4068 3476 4120 3528
rect 4344 3476 4396 3528
rect 4804 3544 4856 3596
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5264 3612 5316 3664
rect 5448 3476 5500 3528
rect 6000 3544 6052 3596
rect 6552 3544 6604 3596
rect 7012 3544 7064 3596
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 6184 3408 6236 3460
rect 6920 3476 6972 3528
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8484 3544 8536 3596
rect 7472 3476 7524 3528
rect 3608 3340 3660 3392
rect 3976 3340 4028 3392
rect 4620 3340 4672 3392
rect 4804 3340 4856 3392
rect 6920 3340 6972 3392
rect 7748 3408 7800 3460
rect 8208 3451 8260 3460
rect 8208 3417 8217 3451
rect 8217 3417 8251 3451
rect 8251 3417 8260 3451
rect 8208 3408 8260 3417
rect 8668 3476 8720 3528
rect 8760 3408 8812 3460
rect 8116 3340 8168 3392
rect 8944 3476 8996 3528
rect 9588 3544 9640 3596
rect 11704 3612 11756 3664
rect 11980 3612 12032 3664
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 9404 3340 9456 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 9956 3340 10008 3392
rect 10140 3476 10192 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 11612 3476 11664 3528
rect 12072 3476 12124 3528
rect 10600 3451 10652 3460
rect 10600 3417 10609 3451
rect 10609 3417 10643 3451
rect 10643 3417 10652 3451
rect 10600 3408 10652 3417
rect 12808 3612 12860 3664
rect 17776 3612 17828 3664
rect 12624 3544 12676 3596
rect 12256 3476 12308 3528
rect 12992 3544 13044 3596
rect 13176 3544 13228 3596
rect 13268 3544 13320 3596
rect 12808 3476 12860 3528
rect 11980 3340 12032 3392
rect 13084 3451 13136 3460
rect 13084 3417 13093 3451
rect 13093 3417 13127 3451
rect 13127 3417 13136 3451
rect 13084 3408 13136 3417
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 12716 3383 12768 3392
rect 12716 3349 12725 3383
rect 12725 3349 12759 3383
rect 12759 3349 12768 3383
rect 12716 3340 12768 3349
rect 12900 3340 12952 3392
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13268 3383 13320 3392
rect 13268 3349 13293 3383
rect 13293 3349 13320 3383
rect 13268 3340 13320 3349
rect 13636 3340 13688 3392
rect 13912 3519 13964 3528
rect 13912 3485 13921 3519
rect 13921 3485 13955 3519
rect 13955 3485 13964 3519
rect 13912 3476 13964 3485
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 15568 3544 15620 3596
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 17408 3544 17460 3596
rect 18052 3612 18104 3664
rect 19156 3612 19208 3664
rect 19248 3612 19300 3664
rect 19616 3612 19668 3664
rect 23848 3680 23900 3732
rect 23020 3612 23072 3664
rect 18420 3544 18472 3596
rect 15936 3408 15988 3460
rect 16304 3408 16356 3460
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 17592 3476 17644 3528
rect 16948 3408 17000 3460
rect 18144 3451 18196 3460
rect 18144 3417 18153 3451
rect 18153 3417 18187 3451
rect 18187 3417 18196 3451
rect 18144 3408 18196 3417
rect 18236 3451 18288 3460
rect 18236 3417 18245 3451
rect 18245 3417 18279 3451
rect 18279 3417 18288 3451
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19156 3476 19208 3528
rect 18236 3408 18288 3417
rect 20076 3544 20128 3596
rect 20260 3544 20312 3596
rect 19800 3476 19852 3528
rect 20444 3476 20496 3528
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 22836 3544 22888 3596
rect 26240 3680 26292 3732
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 24860 3612 24912 3664
rect 27068 3544 27120 3596
rect 20812 3451 20864 3460
rect 20812 3417 20821 3451
rect 20821 3417 20855 3451
rect 20855 3417 20864 3451
rect 20812 3408 20864 3417
rect 22284 3408 22336 3460
rect 23572 3476 23624 3528
rect 23940 3476 23992 3528
rect 24216 3519 24268 3528
rect 24216 3485 24225 3519
rect 24225 3485 24259 3519
rect 24259 3485 24268 3519
rect 24216 3476 24268 3485
rect 24676 3476 24728 3528
rect 23112 3408 23164 3460
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 16856 3340 16908 3392
rect 25596 3408 25648 3460
rect 26240 3476 26292 3528
rect 26884 3519 26936 3528
rect 26884 3485 26893 3519
rect 26893 3485 26927 3519
rect 26927 3485 26936 3519
rect 26884 3476 26936 3485
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 18420 3340 18472 3392
rect 19340 3340 19392 3392
rect 19432 3383 19484 3392
rect 19432 3349 19441 3383
rect 19441 3349 19475 3383
rect 19475 3349 19484 3383
rect 19432 3340 19484 3349
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 20720 3340 20772 3392
rect 21088 3340 21140 3392
rect 23204 3340 23256 3392
rect 23756 3340 23808 3392
rect 23940 3340 23992 3392
rect 24676 3383 24728 3392
rect 24676 3349 24685 3383
rect 24685 3349 24719 3383
rect 24719 3349 24728 3383
rect 24676 3340 24728 3349
rect 24768 3340 24820 3392
rect 25780 3340 25832 3392
rect 25964 3383 26016 3392
rect 25964 3349 25973 3383
rect 25973 3349 26007 3383
rect 26007 3349 26016 3383
rect 25964 3340 26016 3349
rect 26148 3340 26200 3392
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 27068 3383 27120 3392
rect 27068 3349 27077 3383
rect 27077 3349 27111 3383
rect 27111 3349 27120 3383
rect 27068 3340 27120 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1308 3136 1360 3188
rect 4528 3136 4580 3188
rect 4068 3068 4120 3120
rect 4344 3068 4396 3120
rect 5264 3068 5316 3120
rect 5540 3136 5592 3188
rect 6092 3136 6144 3188
rect 7012 3136 7064 3188
rect 8024 3136 8076 3188
rect 8668 3179 8720 3188
rect 8668 3145 8677 3179
rect 8677 3145 8711 3179
rect 8711 3145 8720 3179
rect 8668 3136 8720 3145
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 5908 3111 5960 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 1952 3000 2004 3052
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 3516 3000 3568 3052
rect 4252 3000 4304 3052
rect 4528 3043 4580 3052
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 5080 3000 5132 3052
rect 5908 3077 5917 3111
rect 5917 3077 5951 3111
rect 5951 3077 5960 3111
rect 5908 3068 5960 3077
rect 5448 3000 5500 3052
rect 5724 3000 5776 3052
rect 6644 3068 6696 3120
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 6552 3000 6604 3052
rect 8392 3068 8444 3120
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8760 3000 8812 3052
rect 9312 3136 9364 3188
rect 9496 3136 9548 3188
rect 9588 3111 9640 3120
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9588 3077 9597 3111
rect 9597 3077 9631 3111
rect 9631 3077 9640 3111
rect 9588 3068 9640 3077
rect 9956 3068 10008 3120
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 10140 3136 10192 3188
rect 10232 3136 10284 3188
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 10784 3136 10836 3188
rect 14464 3136 14516 3188
rect 1216 2864 1268 2916
rect 3424 2864 3476 2916
rect 3884 2796 3936 2848
rect 4988 2839 5040 2848
rect 4988 2805 4997 2839
rect 4997 2805 5031 2839
rect 5031 2805 5040 2839
rect 4988 2796 5040 2805
rect 6184 2907 6236 2916
rect 6184 2873 6193 2907
rect 6193 2873 6227 2907
rect 6227 2873 6236 2907
rect 6184 2864 6236 2873
rect 7012 2932 7064 2984
rect 7932 2932 7984 2984
rect 8852 2932 8904 2984
rect 10140 3000 10192 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 11980 3068 12032 3120
rect 12072 3068 12124 3120
rect 13728 3068 13780 3120
rect 14556 3068 14608 3120
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 9312 2864 9364 2916
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 9036 2796 9088 2848
rect 9496 2796 9548 2848
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 11428 2932 11480 2984
rect 10232 2864 10284 2916
rect 10968 2864 11020 2916
rect 10784 2796 10836 2848
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 14372 3000 14424 3052
rect 15384 3136 15436 3188
rect 15936 3136 15988 3188
rect 14740 3068 14792 3120
rect 20536 3136 20588 3188
rect 20812 3136 20864 3188
rect 21456 3136 21508 3188
rect 23572 3136 23624 3188
rect 24124 3179 24176 3188
rect 24124 3145 24133 3179
rect 24133 3145 24167 3179
rect 24167 3145 24176 3179
rect 24124 3136 24176 3145
rect 18236 3068 18288 3120
rect 21640 3068 21692 3120
rect 18052 3000 18104 3052
rect 13176 2932 13228 2984
rect 14096 2932 14148 2984
rect 15292 2932 15344 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 17684 2932 17736 2984
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19248 3043 19300 3052
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 19524 3000 19576 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 20444 3000 20496 3052
rect 18328 2932 18380 2984
rect 18052 2864 18104 2916
rect 18420 2864 18472 2916
rect 19432 2932 19484 2984
rect 20260 2975 20312 2984
rect 20260 2941 20269 2975
rect 20269 2941 20303 2975
rect 20303 2941 20312 2975
rect 20260 2932 20312 2941
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 21088 3043 21140 3052
rect 21088 3009 21097 3043
rect 21097 3009 21131 3043
rect 21131 3009 21140 3043
rect 21088 3000 21140 3009
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 22284 3000 22336 3052
rect 22744 3068 22796 3120
rect 23664 3000 23716 3052
rect 12440 2796 12492 2848
rect 12808 2796 12860 2848
rect 14924 2796 14976 2848
rect 16672 2796 16724 2848
rect 18880 2864 18932 2916
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 22100 2975 22152 2984
rect 22100 2941 22109 2975
rect 22109 2941 22143 2975
rect 22143 2941 22152 2975
rect 22100 2932 22152 2941
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 23112 2932 23164 2984
rect 25136 3136 25188 3188
rect 25228 3136 25280 3188
rect 27436 3179 27488 3188
rect 27436 3145 27445 3179
rect 27445 3145 27479 3179
rect 27479 3145 27488 3179
rect 27436 3136 27488 3145
rect 24860 3068 24912 3120
rect 24584 3000 24636 3052
rect 24952 3043 25004 3052
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 24860 2932 24912 2984
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 25688 3000 25740 3052
rect 26516 3043 26568 3052
rect 26516 3009 26525 3043
rect 26525 3009 26559 3043
rect 26559 3009 26568 3043
rect 26516 3000 26568 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 26424 2932 26476 2984
rect 27068 2932 27120 2984
rect 27252 3043 27304 3052
rect 27252 3009 27261 3043
rect 27261 3009 27295 3043
rect 27295 3009 27304 3043
rect 27252 3000 27304 3009
rect 24124 2864 24176 2916
rect 24400 2864 24452 2916
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 18972 2796 19024 2848
rect 19156 2796 19208 2848
rect 20628 2796 20680 2848
rect 21916 2796 21968 2848
rect 25044 2864 25096 2916
rect 26884 2796 26936 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 1308 2524 1360 2576
rect 1124 2456 1176 2508
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 5816 2592 5868 2644
rect 6000 2592 6052 2644
rect 6644 2592 6696 2644
rect 6460 2524 6512 2576
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2320 2388 2372 2440
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 4804 2456 4856 2508
rect 4988 2456 5040 2508
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 2964 2320 3016 2372
rect 3700 2320 3752 2372
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4620 2388 4672 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 4896 2388 4948 2440
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5908 2456 5960 2508
rect 7012 2456 7064 2508
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 5264 2320 5316 2372
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 8300 2524 8352 2576
rect 8944 2524 8996 2576
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 1032 2252 1084 2304
rect 3884 2252 3936 2304
rect 3976 2252 4028 2304
rect 4620 2252 4672 2304
rect 8024 2388 8076 2440
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8760 2388 8812 2440
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 7564 2252 7616 2304
rect 8852 2320 8904 2372
rect 9496 2388 9548 2440
rect 9864 2465 9891 2474
rect 9891 2465 9916 2474
rect 9864 2422 9916 2465
rect 12532 2592 12584 2644
rect 13360 2592 13412 2644
rect 14280 2592 14332 2644
rect 15292 2592 15344 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 16948 2592 17000 2644
rect 17776 2635 17828 2644
rect 17776 2601 17785 2635
rect 17785 2601 17819 2635
rect 17819 2601 17828 2635
rect 17776 2592 17828 2601
rect 13728 2524 13780 2576
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10324 2388 10376 2440
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 9588 2320 9640 2372
rect 12164 2388 12216 2440
rect 12440 2388 12492 2440
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 14188 2456 14240 2508
rect 15108 2524 15160 2576
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 14004 2320 14056 2372
rect 14280 2363 14332 2372
rect 14280 2329 14289 2363
rect 14289 2329 14323 2363
rect 14323 2329 14332 2363
rect 14280 2320 14332 2329
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 15936 2388 15988 2440
rect 17224 2524 17276 2576
rect 17868 2524 17920 2576
rect 20352 2592 20404 2644
rect 20444 2592 20496 2644
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 22284 2592 22336 2644
rect 25964 2592 26016 2644
rect 26516 2635 26568 2644
rect 26516 2601 26525 2635
rect 26525 2601 26559 2635
rect 26559 2601 26568 2635
rect 26516 2592 26568 2601
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 18788 2456 18840 2508
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 7840 2252 7892 2304
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 9404 2252 9456 2304
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 11244 2252 11296 2304
rect 13084 2252 13136 2304
rect 14924 2252 14976 2304
rect 16028 2363 16080 2372
rect 16028 2329 16037 2363
rect 16037 2329 16071 2363
rect 16071 2329 16080 2363
rect 16028 2320 16080 2329
rect 16304 2320 16356 2372
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 19248 2499 19300 2508
rect 19248 2465 19257 2499
rect 19257 2465 19291 2499
rect 19291 2465 19300 2499
rect 19248 2456 19300 2465
rect 21640 2524 21692 2576
rect 16212 2252 16264 2304
rect 16764 2252 16816 2304
rect 17132 2252 17184 2304
rect 18144 2363 18196 2372
rect 18144 2329 18153 2363
rect 18153 2329 18187 2363
rect 18187 2329 18196 2363
rect 18144 2320 18196 2329
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19340 2388 19392 2440
rect 22192 2456 22244 2508
rect 22376 2456 22428 2508
rect 23388 2567 23440 2576
rect 23388 2533 23397 2567
rect 23397 2533 23431 2567
rect 23431 2533 23440 2567
rect 23388 2524 23440 2533
rect 23480 2567 23532 2576
rect 23480 2533 23489 2567
rect 23489 2533 23523 2567
rect 23523 2533 23532 2567
rect 23480 2524 23532 2533
rect 24584 2524 24636 2576
rect 24860 2524 24912 2576
rect 24124 2456 24176 2508
rect 25136 2456 25188 2508
rect 25872 2524 25924 2576
rect 18604 2252 18656 2304
rect 21364 2320 21416 2372
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 22560 2363 22612 2372
rect 22560 2329 22569 2363
rect 22569 2329 22603 2363
rect 22603 2329 22612 2363
rect 22560 2320 22612 2329
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 24032 2388 24084 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 25412 2388 25464 2440
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 26516 2388 26568 2440
rect 26792 2431 26844 2440
rect 26792 2397 26801 2431
rect 26801 2397 26835 2431
rect 26835 2397 26844 2431
rect 26792 2388 26844 2397
rect 21088 2252 21140 2304
rect 23480 2252 23532 2304
rect 24216 2252 24268 2304
rect 24952 2252 25004 2304
rect 27804 2320 27856 2372
rect 26700 2295 26752 2304
rect 26700 2261 26709 2295
rect 26709 2261 26743 2295
rect 26743 2261 26752 2295
rect 26700 2252 26752 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 2320 2048 2372 2100
rect 1676 1980 1728 2032
rect 6092 2048 6144 2100
rect 10784 2048 10836 2100
rect 11704 2048 11756 2100
rect 14280 2048 14332 2100
rect 16028 2048 16080 2100
rect 17132 2048 17184 2100
rect 19064 2048 19116 2100
rect 7748 1980 7800 2032
rect 7840 1980 7892 2032
rect 12624 1980 12676 2032
rect 2412 1844 2464 1896
rect 5632 1912 5684 1964
rect 21088 1912 21140 1964
rect 23388 2048 23440 2100
rect 27068 2048 27120 2100
rect 22192 1980 22244 2032
rect 26700 1980 26752 2032
rect 25504 1912 25556 1964
rect 2228 1774 2280 1826
rect 10692 1844 10744 1896
rect 16212 1844 16264 1896
rect 18236 1844 18288 1896
rect 22560 1844 22612 1896
rect 9128 1776 9180 1828
rect 27160 1776 27212 1828
rect 8576 1708 8628 1760
rect 9956 1708 10008 1760
rect 26240 1698 26292 1750
rect 4804 1636 4856 1688
rect 5264 1636 5316 1688
rect 9496 1640 9548 1692
rect 10416 1640 10468 1692
rect 22100 1630 22152 1682
rect 26792 1630 26844 1682
rect 17040 1564 17092 1616
<< metal2 >>
rect 1214 7984 1270 7993
rect 1214 7919 1270 7928
rect 1228 7750 1256 7919
rect 1216 7744 1268 7750
rect 1122 7712 1178 7721
rect 1306 7710 1362 8110
rect 2688 7744 2740 7750
rect 1216 7686 1268 7692
rect 1122 7647 1178 7656
rect 1136 7546 1164 7647
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 1320 7478 1348 7710
rect 2688 7686 2740 7692
rect 2872 7744 2924 7750
rect 3698 7710 3754 8110
rect 6090 7710 6146 8110
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 2872 7686 2924 7692
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 2594 7440 2650 7449
rect 2700 7410 2728 7686
rect 2884 7546 2912 7686
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2594 7375 2596 7384
rect 1490 7168 1546 7177
rect 1490 7103 1546 7112
rect 1504 7002 1532 7103
rect 1872 7002 1900 7375
rect 2648 7375 2650 7384
rect 2688 7404 2740 7410
rect 2596 7346 2648 7352
rect 2688 7346 2740 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 2424 6905 2452 7142
rect 2688 6928 2740 6934
rect 2410 6896 2466 6905
rect 2136 6860 2188 6866
rect 2410 6831 2466 6840
rect 2686 6896 2688 6905
rect 2740 6896 2742 6905
rect 2686 6831 2742 6840
rect 2136 6802 2188 6808
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 1306 6624 1362 6633
rect 1228 6361 1256 6598
rect 1306 6559 1362 6568
rect 1320 6458 1348 6559
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1214 6352 1270 6361
rect 2148 6322 2176 6802
rect 2228 6792 2280 6798
rect 2412 6792 2464 6798
rect 2228 6734 2280 6740
rect 2410 6760 2412 6769
rect 2464 6760 2466 6769
rect 1214 6287 1270 6296
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1240 6180 1292 6186
rect 1240 6122 1292 6128
rect 1252 6089 1280 6122
rect 1238 6080 1294 6089
rect 1238 6015 1294 6024
rect 1172 5840 1224 5846
rect 1170 5808 1172 5817
rect 2056 5817 2084 6258
rect 1224 5808 1226 5817
rect 1170 5743 1226 5752
rect 2042 5808 2098 5817
rect 2042 5743 2098 5752
rect 1676 5704 1728 5710
rect 1674 5672 1676 5681
rect 1728 5672 1730 5681
rect 1674 5607 1730 5616
rect 1860 5568 1912 5574
rect 1858 5536 1860 5545
rect 1912 5536 1914 5545
rect 1858 5471 1914 5480
rect 1156 5364 1208 5370
rect 1156 5306 1208 5312
rect 1168 5273 1196 5306
rect 1154 5264 1210 5273
rect 1154 5199 1210 5208
rect 1766 5128 1822 5137
rect 1766 5063 1822 5072
rect 1150 5024 1202 5030
rect 1148 4992 1150 5001
rect 1202 4992 1204 5001
rect 1148 4927 1204 4936
rect 1124 4752 1176 4758
rect 1122 4720 1124 4729
rect 1176 4720 1178 4729
rect 1122 4655 1178 4664
rect 1674 4720 1730 4729
rect 1674 4655 1730 4664
rect 1688 4622 1716 4655
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1490 4448 1546 4457
rect 1490 4383 1546 4392
rect 1504 4010 1532 4383
rect 1674 4040 1730 4049
rect 1492 4004 1544 4010
rect 1674 3975 1730 3984
rect 1492 3946 1544 3952
rect 1306 3904 1362 3913
rect 1306 3839 1362 3848
rect 1320 3738 1348 3839
rect 1308 3732 1360 3738
rect 1308 3674 1360 3680
rect 1214 3632 1270 3641
rect 1214 3567 1270 3576
rect 1228 2922 1256 3567
rect 1306 3360 1362 3369
rect 1306 3295 1362 3304
rect 1320 3194 1348 3295
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 1490 3088 1546 3097
rect 1688 3058 1716 3975
rect 1780 3534 1808 5063
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1950 4584 2006 4593
rect 1950 4519 2006 4528
rect 1858 4176 1914 4185
rect 1964 4146 1992 4519
rect 1858 4111 1914 4120
rect 1952 4140 2004 4146
rect 1872 4010 1900 4111
rect 1952 4082 2004 4088
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1950 3088 2006 3097
rect 1490 3023 1546 3032
rect 1676 3052 1728 3058
rect 1216 2916 1268 2922
rect 1216 2858 1268 2864
rect 1504 2650 1532 3023
rect 1950 3023 1952 3032
rect 1676 2994 1728 3000
rect 2004 3023 2006 3032
rect 1952 2994 2004 3000
rect 1858 2816 1914 2825
rect 1858 2751 1914 2760
rect 1872 2650 1900 2751
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 1308 2576 1360 2582
rect 1030 2544 1086 2553
rect 1308 2518 1360 2524
rect 1030 2479 1086 2488
rect 1124 2508 1176 2514
rect 1044 2310 1072 2479
rect 1124 2450 1176 2456
rect 1032 2304 1084 2310
rect 1032 2246 1084 2252
rect 1136 1600 1164 2450
rect 1320 2281 1348 2518
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1306 2272 1362 2281
rect 1306 2207 1362 2216
rect 1688 2038 1716 2382
rect 1676 2032 1728 2038
rect 1676 1974 1728 1980
rect 2056 1600 2084 4966
rect 2148 4690 2176 6258
rect 2240 5273 2268 6734
rect 2410 6695 2466 6704
rect 2226 5264 2282 5273
rect 2226 5199 2282 5208
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2148 4146 2176 4626
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2148 3602 2176 4082
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2148 3058 2176 3538
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2240 1832 2268 3946
rect 2332 2553 2360 5170
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2700 4690 2728 5034
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2792 3602 2820 7414
rect 3330 7304 3386 7313
rect 3330 7239 3386 7248
rect 3344 6798 3372 7239
rect 3712 7206 3740 7710
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 6104 7546 6132 7710
rect 6458 7576 6514 7585
rect 6092 7540 6144 7546
rect 6458 7511 6514 7520
rect 6092 7482 6144 7488
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4344 7336 4396 7342
rect 4080 7296 4344 7324
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2884 5098 2912 5646
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 3160 3942 3188 5102
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3252 3777 3280 5646
rect 3344 5556 3372 6734
rect 3436 6361 3464 6734
rect 3422 6352 3478 6361
rect 3422 6287 3478 6296
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3344 5528 3556 5556
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3238 3768 3294 3777
rect 3238 3703 3294 3712
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 3252 3534 3280 3606
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2318 2544 2374 2553
rect 2318 2479 2374 2488
rect 3344 2446 3372 4966
rect 3436 2922 3464 5170
rect 3528 4486 3556 5528
rect 3620 4554 3648 6122
rect 3712 5234 3740 6287
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3804 5914 3832 6190
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3896 5642 3924 5782
rect 4080 5778 4108 7296
rect 4344 7278 4396 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4264 6390 4292 6938
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 6458 4476 6666
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3620 4146 3648 4490
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3804 4434 3832 5238
rect 3988 5234 4016 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5284 4108 5510
rect 4448 5409 4476 5850
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4434 5400 4490 5409
rect 4434 5335 4490 5344
rect 4160 5296 4212 5302
rect 4080 5256 4160 5284
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4622 3924 4966
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3608 4140 3660 4146
rect 3528 4100 3608 4128
rect 3528 3670 3556 4100
rect 3608 4082 3660 4088
rect 3606 3768 3662 3777
rect 3606 3703 3662 3712
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 3528 3058 3556 3606
rect 3620 3398 3648 3703
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 2332 2106 2360 2382
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2424 1902 2452 2382
rect 3712 2378 3740 4422
rect 3804 4406 3924 4434
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3804 2650 3832 4014
rect 3896 2854 3924 4406
rect 3988 4078 4016 5170
rect 4080 4604 4108 5256
rect 4160 5238 4212 5244
rect 4448 5030 4476 5335
rect 4540 5030 4568 5646
rect 4632 5234 4660 7346
rect 4724 7274 4752 7346
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 5906 7168 5962 7177
rect 5906 7103 5962 7112
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4758 4660 5170
rect 4724 5114 4752 6122
rect 4816 5574 4844 6190
rect 5000 5846 5028 6394
rect 5552 6390 5580 6938
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5356 6316 5408 6322
rect 5408 6276 5488 6304
rect 5356 6258 5408 6264
rect 5460 5914 5488 6276
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5368 5710 5396 5850
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 5228 4856 5234
rect 5172 5228 5224 5234
rect 4856 5188 4936 5216
rect 4804 5170 4856 5176
rect 4724 5086 4844 5114
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4344 4616 4396 4622
rect 4080 4576 4344 4604
rect 4344 4558 4396 4564
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3738 4016 4014
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3534 4108 4218
rect 4356 4146 4384 4558
rect 4632 4146 4660 4694
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4540 3924 4568 4082
rect 4540 3896 4660 3924
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4068 3528 4120 3534
rect 4344 3528 4396 3534
rect 4068 3470 4120 3476
rect 4250 3496 4306 3505
rect 4344 3470 4396 3476
rect 4250 3431 4306 3440
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3988 2428 4016 3334
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4080 2632 4108 3062
rect 4264 3058 4292 3431
rect 4356 3126 4384 3470
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4252 3052 4304 3058
rect 4448 3040 4476 3674
rect 4632 3398 4660 3896
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4528 3188 4580 3194
rect 4632 3176 4660 3334
rect 4580 3148 4660 3176
rect 4528 3130 4580 3136
rect 4528 3052 4580 3058
rect 4448 3012 4528 3040
rect 4252 2994 4304 3000
rect 4580 3012 4660 3040
rect 4528 2994 4580 3000
rect 4264 2961 4292 2994
rect 4250 2952 4306 2961
rect 4250 2887 4306 2896
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4080 2604 4200 2632
rect 4172 2446 4200 2604
rect 4632 2446 4660 3012
rect 4724 2446 4752 4966
rect 4816 4264 4844 5086
rect 4908 5001 4936 5188
rect 5172 5170 5224 5176
rect 4894 4992 4950 5001
rect 4894 4927 4950 4936
rect 5184 4826 5212 5170
rect 5276 5114 5304 5646
rect 5460 5234 5488 5646
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5276 5086 5396 5114
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4908 4486 4936 4558
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4816 4236 4936 4264
rect 4802 3768 4858 3777
rect 4802 3703 4858 3712
rect 4816 3602 4844 3703
rect 4908 3670 4936 4236
rect 5276 4214 5304 4966
rect 5368 4808 5396 5086
rect 5368 4780 5488 4808
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4988 4208 5040 4214
rect 5264 4208 5316 4214
rect 4988 4150 5040 4156
rect 5078 4176 5134 4185
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5000 3534 5028 4150
rect 5264 4150 5316 4156
rect 5078 4111 5134 4120
rect 5172 4140 5224 4146
rect 4988 3528 5040 3534
rect 5092 3505 5120 4111
rect 5172 4082 5224 4088
rect 5184 3913 5212 4082
rect 5170 3904 5226 3913
rect 5170 3839 5226 3848
rect 5368 3738 5396 4626
rect 5460 4321 5488 4780
rect 5446 4312 5502 4321
rect 5446 4247 5502 4256
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5354 3632 5410 3641
rect 4988 3470 5040 3476
rect 5078 3496 5134 3505
rect 5078 3431 5134 3440
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4816 2514 4844 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5276 3126 5304 3606
rect 5354 3567 5410 3576
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5080 3052 5132 3058
rect 5368 3040 5396 3567
rect 5460 3534 5488 4082
rect 5448 3528 5500 3534
rect 5446 3496 5448 3505
rect 5500 3496 5502 3505
rect 5446 3431 5502 3440
rect 5552 3194 5580 6190
rect 5644 4826 5672 6802
rect 5828 6730 5856 6870
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5736 6225 5764 6394
rect 5814 6352 5870 6361
rect 5920 6322 5948 7103
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5814 6287 5870 6296
rect 5908 6316 5960 6322
rect 5828 6254 5856 6287
rect 5908 6258 5960 6264
rect 5816 6248 5868 6254
rect 5722 6216 5778 6225
rect 5816 6190 5868 6196
rect 5722 6151 5778 6160
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5828 5710 5856 5850
rect 5920 5846 5948 6258
rect 6104 5914 6132 6734
rect 6196 6118 6224 7414
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6288 6662 6316 7278
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6186 6316 6598
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5736 5370 5764 5646
rect 5828 5574 5856 5646
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5920 5166 5948 5238
rect 6012 5234 6040 5646
rect 6196 5642 6224 6054
rect 6380 5658 6408 6190
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6288 5630 6408 5658
rect 6288 5234 6316 5630
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 5234 6408 5510
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4826 5764 4966
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5816 4752 5868 4758
rect 5736 4700 5816 4706
rect 5736 4694 5868 4700
rect 5736 4678 5856 4694
rect 5736 4282 5764 4678
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5644 3942 5672 4082
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5736 3738 5764 4082
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3052 5500 3058
rect 5132 3012 5212 3040
rect 5080 2994 5132 3000
rect 5184 2972 5212 3012
rect 5368 3012 5448 3040
rect 5368 2972 5396 3012
rect 5448 2994 5500 3000
rect 4894 2952 4950 2961
rect 5184 2944 5396 2972
rect 4894 2887 4950 2896
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4908 2446 4936 2887
rect 4988 2848 5040 2854
rect 4986 2816 4988 2825
rect 5040 2816 5042 2825
rect 4986 2751 5042 2760
rect 5000 2514 5028 2751
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4068 2440 4120 2446
rect 3988 2400 4068 2428
rect 4068 2382 4120 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4896 2440 4948 2446
rect 5080 2440 5132 2446
rect 4896 2382 4948 2388
rect 5078 2408 5080 2417
rect 5132 2408 5134 2417
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2228 1826 2280 1832
rect 2228 1768 2280 1774
rect 2976 1600 3004 2314
rect 4632 2310 4660 2382
rect 5078 2343 5134 2352
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 3896 1600 3924 2246
rect 3988 2009 4016 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 3974 2000 4030 2009
rect 3974 1935 4030 1944
rect 5276 1694 5304 2314
rect 5644 1970 5672 3674
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5736 3058 5764 3295
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5828 2650 5856 4082
rect 5920 3126 5948 5102
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6012 3602 6040 4422
rect 6196 3738 6224 4558
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4282 6408 4490
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6366 3904 6422 3913
rect 6366 3839 6422 3848
rect 6184 3732 6236 3738
rect 6104 3692 6184 3720
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 3233 6040 3538
rect 5998 3224 6054 3233
rect 6104 3194 6132 3692
rect 6184 3674 6236 3680
rect 6380 3534 6408 3839
rect 6472 3738 6500 7511
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 6497 6592 6734
rect 6550 6488 6606 6497
rect 6550 6423 6606 6432
rect 6656 6089 6684 7346
rect 7024 7342 7052 7754
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7206 7052 7278
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 7002 7236 7142
rect 7196 6996 7248 7002
rect 7380 6996 7432 7002
rect 7196 6938 7248 6944
rect 7300 6956 7380 6984
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6642 6080 6698 6089
rect 6642 6015 6698 6024
rect 6656 5574 6684 6015
rect 6748 5778 6776 6190
rect 7300 5846 7328 6956
rect 7380 6938 7432 6944
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6932 4264 6960 5782
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4622 7144 5102
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6564 4236 6960 4264
rect 6564 4146 6592 4236
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6656 3942 6684 4082
rect 6840 4010 6868 4082
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6552 3596 6604 3602
rect 6656 3584 6684 3878
rect 6604 3556 6684 3584
rect 6552 3538 6604 3544
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 5998 3159 6054 3168
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2514 5948 3062
rect 6196 2922 6224 3402
rect 6458 3224 6514 3233
rect 6458 3159 6514 3168
rect 6472 3058 6500 3159
rect 6564 3058 6592 3538
rect 6932 3534 6960 4236
rect 7116 4010 7144 4422
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7024 3602 7052 3946
rect 7208 3913 7236 5646
rect 7392 5545 7420 5646
rect 7378 5536 7434 5545
rect 7378 5471 7434 5480
rect 7484 5001 7512 7890
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7576 7313 7604 7414
rect 7656 7336 7708 7342
rect 7562 7304 7618 7313
rect 7656 7278 7708 7284
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7562 7239 7618 7248
rect 7668 6458 7696 7278
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7760 5914 7788 7278
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6322 8156 6394
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7562 5264 7618 5273
rect 7668 5234 7696 5646
rect 7852 5574 7880 6054
rect 8220 5710 8248 7754
rect 8482 7710 8538 8110
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 8496 7546 8524 7710
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 9048 7002 9076 7414
rect 9772 7336 9824 7342
rect 9402 7304 9458 7313
rect 9772 7278 9824 7284
rect 9402 7239 9458 7248
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6322 8340 6598
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7746 5264 7802 5273
rect 7562 5199 7618 5208
rect 7656 5228 7708 5234
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7392 4622 7420 4762
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7194 3904 7250 3913
rect 7194 3839 7250 3848
rect 7300 3777 7328 4422
rect 7484 4282 7512 4927
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7392 4049 7420 4150
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7378 4040 7434 4049
rect 7378 3975 7434 3984
rect 7286 3768 7342 3777
rect 7286 3703 7342 3712
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3398 6960 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7024 3194 7052 3538
rect 7484 3534 7512 4082
rect 7576 3641 7604 5199
rect 7746 5199 7802 5208
rect 7656 5170 7708 5176
rect 7760 5166 7788 5199
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7656 4616 7708 4622
rect 7852 4604 7880 5510
rect 7944 5234 7972 5646
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7944 5098 7972 5170
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7944 4622 7972 5034
rect 8128 4622 8156 5238
rect 8220 5234 8248 5646
rect 8312 5370 8340 6258
rect 8390 5808 8446 5817
rect 8390 5743 8446 5752
rect 8404 5710 8432 5743
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8390 5536 8446 5545
rect 8390 5471 8446 5480
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8298 5264 8354 5273
rect 8208 5228 8260 5234
rect 8298 5199 8300 5208
rect 8208 5170 8260 5176
rect 8352 5199 8354 5208
rect 8300 5170 8352 5176
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7708 4576 7880 4604
rect 7932 4616 7984 4622
rect 7656 4558 7708 4564
rect 7932 4558 7984 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7562 3632 7618 3641
rect 7562 3567 7618 3576
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7668 3233 7696 4558
rect 7944 4457 7972 4558
rect 8220 4554 8248 4966
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 7930 4448 7986 4457
rect 7930 4383 7986 4392
rect 8036 4282 8064 4490
rect 8024 4276 8076 4282
rect 7944 4236 8024 4264
rect 7944 4162 7972 4236
rect 8024 4218 8076 4224
rect 7760 4134 7972 4162
rect 8024 4140 8076 4146
rect 7760 3466 7788 4134
rect 8220 4128 8248 4490
rect 8076 4100 8248 4128
rect 8024 4082 8076 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7654 3224 7710 3233
rect 7012 3188 7064 3194
rect 7654 3159 7710 3168
rect 7012 3130 7064 3136
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6012 2094 6040 2586
rect 6472 2582 6500 2790
rect 6656 2650 6684 3062
rect 7852 3058 7880 4014
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7944 2990 7972 3878
rect 8036 3194 8064 4082
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8128 3602 8156 3674
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3505 8156 3538
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 7024 2514 7052 2926
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6104 2106 6132 2382
rect 5736 2066 6040 2094
rect 6092 2100 6144 2106
rect 5632 1964 5684 1970
rect 5632 1906 5684 1912
rect 4804 1688 4856 1694
rect 4804 1630 4856 1636
rect 5264 1688 5316 1694
rect 5264 1630 5316 1636
rect 4816 1600 4844 1630
rect 5736 1600 5764 2066
rect 6092 2042 6144 2048
rect 6656 1600 6684 2382
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 1600 7604 2246
rect 7760 2038 7788 2790
rect 8036 2446 8064 3130
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 2038 7880 2246
rect 7748 2032 7800 2038
rect 7748 1974 7800 1980
rect 7840 2032 7892 2038
rect 8128 2009 8156 3334
rect 8220 2145 8248 3402
rect 8312 2582 8340 5170
rect 8404 4740 8432 5471
rect 8496 5030 8524 6258
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8484 4752 8536 4758
rect 8404 4712 8484 4740
rect 8484 4694 8536 4700
rect 8496 4622 8524 4694
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8390 4312 8446 4321
rect 8390 4247 8446 4256
rect 8404 4010 8432 4247
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8404 3913 8432 3946
rect 8390 3904 8446 3913
rect 8390 3839 8446 3848
rect 8390 3768 8446 3777
rect 8390 3703 8446 3712
rect 8404 3126 8432 3703
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8312 2446 8340 2518
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8206 2136 8262 2145
rect 8206 2071 8262 2080
rect 7840 1974 7892 1980
rect 8114 2000 8170 2009
rect 8114 1935 8170 1944
rect 8496 1600 8524 3538
rect 8588 1766 8616 6054
rect 8680 5574 8708 6326
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8772 5914 8800 6258
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 5778 8984 6054
rect 9048 5914 9076 6938
rect 9324 6458 9352 6938
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9310 6352 9366 6361
rect 9416 6322 9444 7239
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9692 6730 9720 6938
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9310 6287 9366 6296
rect 9404 6316 9456 6322
rect 9324 6254 9352 6287
rect 9404 6258 9456 6264
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9310 5944 9366 5953
rect 9036 5908 9088 5914
rect 9310 5879 9366 5888
rect 9036 5850 9088 5856
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8942 5672 8998 5681
rect 8942 5607 8998 5616
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5098 8708 5510
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8668 4072 8720 4078
rect 8852 4072 8904 4078
rect 8668 4014 8720 4020
rect 8850 4040 8852 4049
rect 8904 4040 8906 4049
rect 8680 3738 8708 4014
rect 8850 3975 8906 3984
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8956 3534 8984 5607
rect 9126 5264 9182 5273
rect 9036 5228 9088 5234
rect 9126 5199 9128 5208
rect 9036 5170 9088 5176
rect 9180 5199 9182 5208
rect 9220 5228 9272 5234
rect 9128 5170 9180 5176
rect 9220 5170 9272 5176
rect 9048 4214 9076 5170
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8668 3528 8720 3534
rect 8944 3528 8996 3534
rect 8668 3470 8720 3476
rect 8850 3496 8906 3505
rect 8680 3194 8708 3470
rect 8760 3460 8812 3466
rect 8944 3470 8996 3476
rect 8850 3431 8906 3440
rect 8760 3402 8812 3408
rect 8772 3194 8800 3402
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8772 2446 8800 2994
rect 8864 2990 8892 3431
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8760 2440 8812 2446
rect 8666 2408 8722 2417
rect 8760 2382 8812 2388
rect 8864 2378 8892 2926
rect 8956 2582 8984 3334
rect 9048 3058 9076 4150
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9048 2854 9076 2994
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 8666 2343 8722 2352
rect 8852 2372 8904 2378
rect 8680 2310 8708 2343
rect 8852 2314 8904 2320
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 9140 1834 9168 4966
rect 9232 4758 9260 5170
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9232 3913 9260 4694
rect 9218 3904 9274 3913
rect 9218 3839 9274 3848
rect 9324 3738 9352 5879
rect 9416 5710 9444 6122
rect 9508 5914 9536 6190
rect 9586 6080 9642 6089
rect 9586 6015 9642 6024
rect 9600 5914 9628 6015
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9692 5710 9720 6394
rect 9784 6390 9812 7278
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9784 5273 9812 6326
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5370 9904 6190
rect 9968 5370 9996 7142
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5296 10100 5302
rect 9494 5264 9550 5273
rect 9770 5264 9826 5273
rect 9494 5199 9550 5208
rect 9588 5228 9640 5234
rect 9508 4758 9536 5199
rect 9640 5188 9720 5216
rect 10048 5238 10100 5244
rect 9770 5199 9826 5208
rect 9588 5170 9640 5176
rect 9692 5148 9720 5188
rect 9772 5160 9824 5166
rect 9692 5120 9772 5148
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3398 9444 4082
rect 9508 3754 9536 4694
rect 9588 4616 9640 4622
rect 9692 4604 9720 5120
rect 9772 5102 9824 5108
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9968 4865 9996 5034
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9968 4622 9996 4791
rect 10060 4622 10088 5238
rect 10152 4622 10180 5782
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5098 10272 5510
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 9772 4616 9824 4622
rect 9692 4576 9772 4604
rect 9588 4558 9640 4564
rect 9772 4558 9824 4564
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9600 3942 9628 4558
rect 9784 4486 9812 4558
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9678 4312 9734 4321
rect 9678 4247 9734 4256
rect 9692 4146 9720 4247
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9678 4040 9734 4049
rect 9678 3975 9680 3984
rect 9732 3975 9734 3984
rect 9680 3946 9732 3952
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9508 3726 9720 3754
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9310 3224 9366 3233
rect 9310 3159 9312 3168
rect 9364 3159 9366 3168
rect 9312 3130 9364 3136
rect 9324 2922 9352 3130
rect 9416 3058 9444 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9508 2854 9536 3130
rect 9600 3126 9628 3538
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9496 2644 9548 2650
rect 9600 2632 9628 3062
rect 9548 2604 9628 2632
rect 9496 2586 9548 2592
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9220 2304 9272 2310
rect 9218 2272 9220 2281
rect 9404 2304 9456 2310
rect 9272 2272 9274 2281
rect 9404 2246 9456 2252
rect 9218 2207 9274 2216
rect 9128 1828 9180 1834
rect 9128 1770 9180 1776
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 9416 1600 9444 2246
rect 9508 1698 9536 2382
rect 9588 2372 9640 2378
rect 9692 2360 9720 3726
rect 9784 3210 9812 4422
rect 9864 4208 9916 4214
rect 10060 4162 10088 4558
rect 9916 4156 10088 4162
rect 9864 4150 10088 4156
rect 9876 4134 10088 4150
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9862 3768 9918 3777
rect 9968 3738 9996 3946
rect 10060 3738 10088 4134
rect 9862 3703 9918 3712
rect 9956 3732 10008 3738
rect 9876 3398 9904 3703
rect 9956 3674 10008 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10152 3618 10180 4558
rect 10336 4264 10364 7822
rect 10874 7710 10930 8110
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10888 7546 10916 7710
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 7002 10548 7142
rect 10796 7002 10824 7278
rect 10888 7002 10916 7346
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 10520 6798 10548 6938
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10782 6624 10838 6633
rect 10612 6458 10640 6598
rect 10782 6559 10838 6568
rect 10796 6458 10824 6559
rect 10600 6452 10652 6458
rect 10784 6452 10836 6458
rect 10600 6394 10652 6400
rect 10704 6412 10784 6440
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10520 6254 10548 6326
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10612 5846 10640 6394
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10520 4622 10548 5306
rect 10704 5302 10732 6412
rect 10784 6394 10836 6400
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5778 11008 6190
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10782 5264 10838 5273
rect 10980 5234 11008 5714
rect 10782 5199 10784 5208
rect 10836 5199 10838 5208
rect 10968 5228 11020 5234
rect 10784 5170 10836 5176
rect 10968 5170 11020 5176
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10612 4622 10640 5102
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10612 4282 10640 4558
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10244 4236 10364 4264
rect 10600 4276 10652 4282
rect 10244 3777 10272 4236
rect 10600 4218 10652 4224
rect 10692 4208 10744 4214
rect 10744 4156 10824 4162
rect 10692 4150 10824 4156
rect 10324 4140 10376 4146
rect 10704 4134 10824 4150
rect 10888 4146 10916 4422
rect 10324 4082 10376 4088
rect 10336 4049 10364 4082
rect 10692 4072 10744 4078
rect 10322 4040 10378 4049
rect 10692 4014 10744 4020
rect 10322 3975 10378 3984
rect 10230 3768 10286 3777
rect 10230 3703 10286 3712
rect 9968 3590 10180 3618
rect 9968 3534 9996 3590
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3210 9996 3334
rect 9784 3182 9996 3210
rect 10152 3194 10180 3470
rect 10244 3194 10272 3470
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 3194 10640 3402
rect 9784 2514 9812 3182
rect 9968 3126 9996 3182
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10140 3052 10192 3058
rect 10416 3052 10468 3058
rect 10192 3012 10272 3040
rect 10140 2994 10192 3000
rect 10244 2922 10272 3012
rect 10416 2994 10468 3000
rect 10428 2961 10456 2994
rect 10414 2952 10470 2961
rect 10232 2916 10284 2922
rect 10414 2887 10470 2896
rect 10232 2858 10284 2864
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9864 2474 9916 2480
rect 9864 2416 9916 2422
rect 9876 2360 9904 2416
rect 9640 2332 9904 2360
rect 9588 2314 9640 2320
rect 9968 1766 9996 2790
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10060 2281 10088 2382
rect 10046 2272 10102 2281
rect 10046 2207 10102 2216
rect 9956 1760 10008 1766
rect 9956 1702 10008 1708
rect 9496 1692 9548 1698
rect 9496 1634 9548 1640
rect 10336 1600 10364 2382
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10428 1698 10456 2246
rect 10704 1902 10732 4014
rect 10796 4010 10824 4134
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 11072 4078 11100 6734
rect 11164 5642 11192 6938
rect 11256 6458 11284 7414
rect 11348 6866 11376 7754
rect 13266 7710 13322 8110
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 13280 7546 13308 7710
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12164 7336 12216 7342
rect 11426 7304 11482 7313
rect 12164 7278 12216 7284
rect 11426 7239 11482 7248
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11440 5302 11468 7239
rect 12070 7032 12126 7041
rect 12070 6967 12126 6976
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11164 4758 11192 5170
rect 11348 5098 11376 5170
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11164 4146 11192 4694
rect 11348 4282 11376 5034
rect 11532 4758 11560 6326
rect 11716 5778 11744 6734
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11992 6458 12020 6666
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11624 5098 11652 5578
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11716 4826 11744 5714
rect 11900 5302 11928 6258
rect 12084 5914 12112 6967
rect 12176 6372 12204 7278
rect 12256 6384 12308 6390
rect 12176 6344 12256 6372
rect 12176 6118 12204 6344
rect 12256 6326 12308 6332
rect 12360 6254 12388 7346
rect 12452 7206 12480 7414
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6458 12572 7142
rect 12716 6860 12768 6866
rect 13268 6860 13320 6866
rect 12768 6820 12940 6848
rect 12716 6802 12768 6808
rect 12622 6760 12678 6769
rect 12622 6695 12678 6704
rect 12806 6760 12862 6769
rect 12806 6695 12862 6704
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12360 5778 12388 6054
rect 12438 5944 12494 5953
rect 12636 5914 12664 6695
rect 12820 6662 12848 6695
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5914 12756 6122
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12438 5879 12494 5888
rect 12624 5908 12676 5914
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11624 4690 11652 4762
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10874 3224 10930 3233
rect 10784 3188 10836 3194
rect 10874 3159 10930 3168
rect 10784 3130 10836 3136
rect 10796 2854 10824 3130
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10888 2446 10916 3159
rect 10980 2922 11008 3674
rect 11624 3534 11652 4014
rect 11716 3670 11744 4762
rect 11808 4622 11836 4966
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4146 12020 4422
rect 12084 4282 12112 5102
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12176 4282 12204 4490
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12164 4276 12216 4282
rect 12268 4264 12296 5238
rect 12348 5228 12400 5234
rect 12452 5216 12480 5879
rect 12624 5850 12676 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5778 12848 6015
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12400 5188 12480 5216
rect 12348 5170 12400 5176
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12268 4236 12388 4264
rect 12164 4218 12216 4224
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 11808 3913 11836 4082
rect 11794 3904 11850 3913
rect 11794 3839 11850 3848
rect 11992 3726 12204 3754
rect 11992 3670 12020 3726
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3126 12020 3334
rect 12084 3126 12112 3470
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12176 3058 12204 3726
rect 12268 3534 12296 4082
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12360 3097 12388 4236
rect 12452 4146 12480 4558
rect 12544 4434 12572 4762
rect 12636 4690 12664 5102
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4690 12756 4966
rect 12820 4865 12848 5102
rect 12806 4856 12862 4865
rect 12806 4791 12862 4800
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12544 4406 12664 4434
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12544 4146 12572 4218
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12346 3088 12402 3097
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12164 3052 12216 3058
rect 12346 3023 12402 3032
rect 12164 2994 12216 3000
rect 11428 2984 11480 2990
rect 11716 2938 11744 2994
rect 11900 2961 11928 2994
rect 11480 2932 11744 2938
rect 11428 2926 11744 2932
rect 10968 2916 11020 2922
rect 11440 2910 11744 2926
rect 10968 2858 11020 2864
rect 10980 2446 11008 2858
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 10796 2106 10824 2246
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10692 1896 10744 1902
rect 10692 1838 10744 1844
rect 10416 1692 10468 1698
rect 10416 1634 10468 1640
rect 11256 1600 11284 2246
rect 11716 2106 11744 2910
rect 11886 2952 11942 2961
rect 11886 2887 11942 2896
rect 12452 2854 12480 4082
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2446 12480 2790
rect 12544 2650 12572 4082
rect 12636 3738 12664 4406
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12636 3602 12664 3674
rect 12820 3670 12848 4082
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12820 3534 12848 3606
rect 12808 3528 12860 3534
rect 12714 3496 12770 3505
rect 12808 3470 12860 3476
rect 12714 3431 12770 3440
rect 12728 3398 12756 3431
rect 12912 3398 12940 6820
rect 13268 6802 13320 6808
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13096 5846 13124 6258
rect 13188 5846 13216 6258
rect 13280 6089 13308 6802
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6662 13400 6734
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6390 13400 6598
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13636 6316 13688 6322
rect 13556 6276 13636 6304
rect 13556 6236 13584 6276
rect 13636 6258 13688 6264
rect 13372 6208 13584 6236
rect 13266 6080 13322 6089
rect 13266 6015 13322 6024
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12992 5568 13044 5574
rect 13096 5556 13124 5782
rect 13176 5568 13228 5574
rect 13096 5528 13176 5556
rect 12992 5510 13044 5516
rect 13176 5510 13228 5516
rect 13004 3602 13032 5510
rect 13188 5302 13216 5510
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13082 4856 13138 4865
rect 13082 4791 13138 4800
rect 13096 4622 13124 4791
rect 13188 4622 13216 5238
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13096 3466 13124 4150
rect 13280 4078 13308 6015
rect 13372 5710 13400 6208
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5953 13584 6054
rect 13542 5944 13598 5953
rect 13452 5908 13504 5914
rect 13832 5914 13860 7414
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 13910 6488 13966 6497
rect 14108 6458 14136 7278
rect 14200 7041 14228 7278
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14186 7032 14242 7041
rect 14186 6967 14188 6976
rect 14240 6967 14242 6976
rect 14188 6938 14240 6944
rect 14292 6730 14320 7210
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14568 6458 14596 6938
rect 13910 6423 13966 6432
rect 14096 6452 14148 6458
rect 13542 5879 13598 5888
rect 13820 5908 13872 5914
rect 13452 5850 13504 5856
rect 13820 5850 13872 5856
rect 13464 5710 13492 5850
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12900 3392 12952 3398
rect 12992 3392 13044 3398
rect 12900 3334 12952 3340
rect 12990 3360 12992 3369
rect 13044 3360 13046 3369
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 11704 2100 11756 2106
rect 11704 2042 11756 2048
rect 12176 1600 12204 2382
rect 12636 2038 12664 3334
rect 12728 3233 12756 3334
rect 12990 3295 13046 3304
rect 12714 3224 12770 3233
rect 12714 3159 12770 3168
rect 13188 2990 13216 3538
rect 13280 3505 13308 3538
rect 13266 3496 13322 3505
rect 13266 3431 13322 3440
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 12808 2848 12860 2854
rect 13280 2825 13308 3334
rect 12808 2790 12860 2796
rect 13266 2816 13322 2825
rect 12716 2440 12768 2446
rect 12820 2428 12848 2790
rect 13266 2751 13322 2760
rect 13372 2650 13400 5646
rect 13556 5030 13584 5782
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13634 5400 13690 5409
rect 13634 5335 13636 5344
rect 13688 5335 13690 5344
rect 13636 5306 13688 5312
rect 13544 5024 13596 5030
rect 13464 4984 13544 5012
rect 13464 4622 13492 4984
rect 13544 4966 13596 4972
rect 13740 4826 13768 5714
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13556 4282 13584 4558
rect 13544 4276 13596 4282
rect 13464 4236 13544 4264
rect 13464 3942 13492 4236
rect 13544 4218 13596 4224
rect 13648 4214 13676 4558
rect 13726 4312 13782 4321
rect 13726 4247 13782 4256
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13740 4146 13768 4247
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13924 4078 13952 6423
rect 14096 6394 14148 6400
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14278 6352 14334 6361
rect 14278 6287 14334 6296
rect 14738 6352 14794 6361
rect 14738 6287 14740 6296
rect 14004 6248 14056 6254
rect 14096 6248 14148 6254
rect 14004 6190 14056 6196
rect 14094 6216 14096 6225
rect 14148 6216 14150 6225
rect 14016 5914 14044 6190
rect 14094 6151 14150 6160
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13912 3528 13964 3534
rect 14016 3516 14044 5578
rect 14108 5370 14136 5646
rect 14292 5642 14320 6287
rect 14792 6287 14794 6296
rect 14740 6258 14792 6264
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14108 5166 14136 5306
rect 14200 5302 14228 5510
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4146 14136 5102
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14200 4060 14228 5238
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14292 4214 14320 4558
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14280 4072 14332 4078
rect 14200 4032 14280 4060
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3534 14136 3878
rect 13964 3488 14044 3516
rect 14096 3528 14148 3534
rect 13912 3470 13964 3476
rect 14096 3470 14148 3476
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3108 13676 3334
rect 13728 3120 13780 3126
rect 13648 3080 13728 3108
rect 13728 3062 13780 3068
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13740 2582 13768 3062
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14108 2446 14136 2926
rect 14200 2514 14228 4032
rect 14384 4060 14412 6122
rect 14568 5710 14596 6122
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14476 5166 14504 5646
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 5234 14688 5578
rect 14752 5234 14780 6054
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14660 4826 14688 5170
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14844 4570 14872 6394
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5778 14964 6054
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14936 5545 14964 5714
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 14922 5536 14978 5545
rect 14922 5471 14978 5480
rect 15120 5370 15148 5646
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15212 5302 15240 7754
rect 15658 7710 15714 8110
rect 17960 7744 18012 7750
rect 15672 7634 15700 7710
rect 18050 7710 18106 8110
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 17960 7686 18012 7692
rect 15672 7606 15792 7634
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15304 7342 15332 7482
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 7206 15332 7278
rect 15764 7206 15792 7606
rect 16578 7440 16634 7449
rect 16578 7375 16634 7384
rect 17776 7404 17828 7410
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15474 7032 15530 7041
rect 15474 6967 15530 6976
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15396 6458 15424 6666
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6338 15516 6967
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15580 6769 15608 6802
rect 15566 6760 15622 6769
rect 15566 6695 15622 6704
rect 15672 6458 15700 7142
rect 16394 6896 16450 6905
rect 16394 6831 16450 6840
rect 16028 6792 16080 6798
rect 15750 6760 15806 6769
rect 16028 6734 16080 6740
rect 15750 6695 15806 6704
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15488 6310 15700 6338
rect 15764 6322 15792 6695
rect 15304 6118 15332 6258
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15488 5778 15516 6310
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15672 6202 15700 6310
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15856 6202 15884 6258
rect 16040 6254 16068 6734
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16316 6458 16344 6666
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 15580 5914 15608 6190
rect 15672 6174 15884 6202
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 5772 15528 5778
rect 15396 5732 15476 5760
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15120 4690 15148 4966
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14752 4542 14872 4570
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14464 4072 14516 4078
rect 14384 4032 14464 4060
rect 14280 4014 14332 4020
rect 14464 4014 14516 4020
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14292 2650 14320 3402
rect 14384 3058 14412 3878
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14476 3194 14504 3470
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14568 3126 14596 4082
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14660 3398 14688 3431
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14752 3126 14780 4542
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 14740 3120 14792 3126
rect 14844 3097 14872 4422
rect 15028 4214 15056 4558
rect 15304 4486 15332 4626
rect 15396 4622 15424 5732
rect 15476 5714 15528 5720
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15580 5234 15608 5510
rect 15672 5234 15700 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5545 15792 5714
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 16028 5704 16080 5710
rect 16132 5692 16160 6122
rect 16080 5664 16344 5692
rect 16028 5646 16080 5652
rect 15750 5536 15806 5545
rect 15750 5471 15806 5480
rect 15856 5302 15884 5646
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15948 5166 15976 5646
rect 16210 5264 16266 5273
rect 16210 5199 16266 5208
rect 15936 5160 15988 5166
rect 15658 5128 15714 5137
rect 15476 5092 15528 5098
rect 15936 5102 15988 5108
rect 15658 5063 15660 5072
rect 15476 5034 15528 5040
rect 15712 5063 15714 5072
rect 15660 5034 15712 5040
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14936 3913 14964 3946
rect 14922 3904 14978 3913
rect 14922 3839 14978 3848
rect 14936 3233 14964 3839
rect 15028 3738 15056 4150
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15120 3380 15148 4014
rect 15212 3534 15240 4150
rect 15304 3534 15332 4422
rect 15396 4146 15424 4558
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15488 4026 15516 5034
rect 16120 5024 16172 5030
rect 15750 4992 15806 5001
rect 16120 4966 16172 4972
rect 15750 4927 15806 4936
rect 15764 4690 15792 4927
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15844 4752 15896 4758
rect 15842 4720 15844 4729
rect 15896 4720 15898 4729
rect 15752 4684 15804 4690
rect 15842 4655 15898 4664
rect 15752 4626 15804 4632
rect 15948 4570 15976 4762
rect 16132 4758 16160 4966
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16224 4622 16252 5199
rect 16120 4616 16172 4622
rect 15948 4564 16120 4570
rect 15948 4558 16172 4564
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15948 4542 16160 4558
rect 15948 4146 15976 4542
rect 16120 4480 16172 4486
rect 16212 4480 16264 4486
rect 16120 4422 16172 4428
rect 16210 4448 16212 4457
rect 16264 4448 16266 4457
rect 16132 4146 16160 4422
rect 16210 4383 16266 4392
rect 16316 4298 16344 5664
rect 16408 5098 16436 6831
rect 16592 6390 16620 7375
rect 17776 7346 17828 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 16670 7032 16726 7041
rect 16670 6967 16726 6976
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 6118 16528 6258
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 5846 16528 6054
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16500 5166 16528 5782
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5302 16620 5646
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16500 4978 16528 5102
rect 16224 4270 16344 4298
rect 16408 4950 16528 4978
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 15396 3998 15516 4026
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15304 3380 15332 3470
rect 15120 3352 15332 3380
rect 14922 3224 14978 3233
rect 14922 3159 14978 3168
rect 14740 3062 14792 3068
rect 14830 3088 14886 3097
rect 14372 3052 14424 3058
rect 14830 3023 14886 3032
rect 14372 2994 14424 3000
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14384 2446 14412 2994
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2446 14964 2790
rect 15120 2582 15148 3352
rect 15396 3194 15424 3998
rect 15568 3936 15620 3942
rect 15752 3936 15804 3942
rect 15568 3878 15620 3884
rect 15750 3904 15752 3913
rect 15804 3904 15806 3913
rect 15580 3602 15608 3878
rect 15750 3839 15806 3848
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15304 2650 15332 2926
rect 15580 2650 15608 3538
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 3194 15976 3402
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15948 2446 15976 3130
rect 16224 2446 16252 4270
rect 16408 4214 16436 4950
rect 16684 4622 16712 6967
rect 17236 6322 17264 7142
rect 17788 7002 17816 7346
rect 17972 7274 18000 7686
rect 18064 7410 18092 7710
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17880 6905 17908 7210
rect 17866 6896 17922 6905
rect 17866 6831 17922 6840
rect 17774 6488 17830 6497
rect 17774 6423 17830 6432
rect 17788 6390 17816 6423
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16960 5914 16988 6258
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17144 5642 17172 6054
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17590 5808 17646 5817
rect 17316 5704 17368 5710
rect 17512 5692 17540 5782
rect 17590 5743 17646 5752
rect 17368 5664 17540 5692
rect 17316 5646 17368 5652
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 16868 5234 16896 5578
rect 17040 5568 17092 5574
rect 17038 5536 17040 5545
rect 17092 5536 17094 5545
rect 16960 5494 17038 5522
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16868 5030 16896 5170
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16762 4584 16818 4593
rect 16762 4519 16818 4528
rect 16776 4486 16804 4519
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16396 4208 16448 4214
rect 16500 4185 16528 4422
rect 16960 4185 16988 5494
rect 17038 5471 17094 5480
rect 17236 5234 17264 5578
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17038 4720 17094 4729
rect 17038 4655 17094 4664
rect 17132 4684 17184 4690
rect 17052 4622 17080 4655
rect 17132 4626 17184 4632
rect 17040 4616 17092 4622
rect 17144 4593 17172 4626
rect 17040 4558 17092 4564
rect 17130 4584 17186 4593
rect 17130 4519 17186 4528
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16396 4150 16448 4156
rect 16486 4176 16542 4185
rect 16946 4176 17002 4185
rect 16868 4146 16946 4162
rect 16486 4111 16542 4120
rect 16856 4140 16946 4146
rect 16908 4134 16946 4140
rect 16946 4111 17002 4120
rect 16856 4082 16908 4088
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 12768 2400 12848 2428
rect 14096 2440 14148 2446
rect 12716 2382 12768 2388
rect 14096 2382 14148 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15752 2440 15804 2446
rect 15936 2440 15988 2446
rect 15804 2400 15884 2428
rect 15752 2382 15804 2388
rect 14004 2372 14056 2378
rect 14004 2314 14056 2320
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 13096 1600 13124 2246
rect 14016 1600 14044 2314
rect 14292 2106 14320 2314
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14936 1600 14964 2246
rect 15856 1600 15884 2400
rect 15936 2382 15988 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 16040 2106 16068 2314
rect 16224 2310 16252 2382
rect 16316 2378 16344 3402
rect 16684 2854 16712 3470
rect 16960 3466 16988 4014
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16868 2446 16896 3334
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16960 2650 16988 2926
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16028 2100 16080 2106
rect 16028 2042 16080 2048
rect 16224 1902 16252 2246
rect 16212 1896 16264 1902
rect 16212 1838 16264 1844
rect 16776 1600 16804 2246
rect 17052 1622 17080 4422
rect 17236 3942 17264 5170
rect 17328 4146 17356 5646
rect 17604 5642 17632 5743
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17604 4622 17632 5578
rect 17696 5234 17724 6326
rect 17880 5710 17908 6831
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6186 18000 6598
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18064 5930 18092 6394
rect 17972 5902 18092 5930
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 5545 17908 5646
rect 17866 5536 17922 5545
rect 17866 5471 17922 5480
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4758 17724 5170
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17236 2582 17264 3878
rect 17406 3768 17462 3777
rect 17406 3703 17462 3712
rect 17420 3602 17448 3703
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17512 2514 17540 4150
rect 17604 3534 17632 4558
rect 17696 4146 17724 4694
rect 17880 4622 17908 5034
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17788 4486 17816 4558
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4321 17816 4422
rect 17774 4312 17830 4321
rect 17880 4282 17908 4558
rect 17972 4321 18000 5902
rect 18052 5840 18104 5846
rect 18156 5794 18184 7278
rect 18248 7274 18276 7958
rect 20442 7812 20498 8110
rect 20442 7760 20444 7812
rect 20496 7760 20498 7812
rect 18972 7744 19024 7750
rect 20442 7710 20498 7760
rect 22834 7710 22890 8110
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 18972 7686 19024 7692
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18340 6390 18368 6870
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18104 5788 18184 5794
rect 18052 5782 18184 5788
rect 18064 5766 18184 5782
rect 18156 5710 18184 5766
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5574 18276 5646
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18144 5364 18196 5370
rect 18340 5352 18368 5714
rect 18196 5324 18368 5352
rect 18144 5306 18196 5312
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4622 18092 5102
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17958 4312 18014 4321
rect 17774 4247 17830 4256
rect 17868 4276 17920 4282
rect 17958 4247 17960 4256
rect 17868 4218 17920 4224
rect 18012 4247 18014 4256
rect 17960 4218 18012 4224
rect 18156 4146 18184 5306
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18248 4758 18276 5034
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 18432 4622 18460 7142
rect 18892 6934 18920 7278
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18524 5846 18552 6734
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 18510 5672 18566 5681
rect 18510 5607 18566 5616
rect 18524 5234 18552 5607
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18616 4690 18644 6802
rect 18696 6792 18748 6798
rect 18694 6760 18696 6769
rect 18748 6760 18750 6769
rect 18694 6695 18750 6704
rect 18786 6624 18842 6633
rect 18786 6559 18842 6568
rect 18800 6100 18828 6559
rect 18708 6072 18828 6100
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18602 4584 18658 4593
rect 18248 4282 18276 4558
rect 18432 4486 18460 4558
rect 18602 4519 18658 4528
rect 18616 4486 18644 4519
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18248 4026 18276 4218
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18432 4078 18460 4150
rect 18616 4078 18644 4422
rect 18708 4146 18736 6072
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18800 4622 18828 5646
rect 18878 5400 18934 5409
rect 18878 5335 18880 5344
rect 18932 5335 18934 5344
rect 18880 5306 18932 5312
rect 18984 4842 19012 7686
rect 20456 7670 20484 7710
rect 22847 7666 22875 7710
rect 22847 7638 23428 7666
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19076 5642 19104 7414
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19168 6458 19196 6666
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6458 19380 6598
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19168 5778 19196 6394
rect 19444 6322 19472 7482
rect 23400 7426 23428 7638
rect 23480 7472 23532 7478
rect 23400 7420 23480 7426
rect 23400 7414 23532 7420
rect 23296 7404 23348 7410
rect 23400 7398 23520 7414
rect 23848 7404 23900 7410
rect 23296 7346 23348 7352
rect 23848 7346 23900 7352
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 19800 7336 19852 7342
rect 20076 7336 20128 7342
rect 19852 7296 19932 7324
rect 19800 7278 19852 7284
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19338 5808 19394 5817
rect 19156 5772 19208 5778
rect 19208 5732 19288 5760
rect 19338 5743 19394 5752
rect 19156 5714 19208 5720
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19062 5400 19118 5409
rect 19062 5335 19118 5344
rect 19076 5030 19104 5335
rect 19168 5234 19196 5510
rect 19260 5234 19288 5732
rect 19352 5710 19380 5743
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5574 19380 5646
rect 19340 5568 19392 5574
rect 19444 5545 19472 6258
rect 19340 5510 19392 5516
rect 19430 5536 19486 5545
rect 19430 5471 19486 5480
rect 19536 5302 19564 6598
rect 19628 5817 19656 6734
rect 19720 5914 19748 6734
rect 19904 6186 19932 7296
rect 20076 7278 20128 7284
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20088 7002 20116 7278
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19996 6497 20024 6666
rect 19982 6488 20038 6497
rect 19982 6423 20038 6432
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19614 5808 19670 5817
rect 19614 5743 19670 5752
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 18892 4814 19012 4842
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18800 4214 18828 4558
rect 18892 4486 18920 4814
rect 18970 4584 19026 4593
rect 18970 4519 19026 4528
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18878 4312 18934 4321
rect 18878 4247 18934 4256
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17880 3998 18276 4026
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18604 4072 18656 4078
rect 18892 4060 18920 4247
rect 18984 4146 19012 4519
rect 19076 4486 19104 4966
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19168 4593 19196 4694
rect 19248 4616 19300 4622
rect 19154 4584 19210 4593
rect 19248 4558 19300 4564
rect 19154 4519 19210 4528
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18604 4014 18656 4020
rect 18800 4032 18920 4060
rect 17592 3528 17644 3534
rect 17696 3516 17724 3946
rect 17880 3738 17908 3998
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18512 3936 18564 3942
rect 18564 3884 18644 3890
rect 18512 3878 18644 3884
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 3664 17828 3670
rect 18052 3664 18104 3670
rect 17828 3612 18052 3618
rect 17776 3606 18104 3612
rect 18156 3618 18184 3878
rect 18524 3862 18644 3878
rect 18616 3777 18644 3862
rect 18418 3768 18474 3777
rect 18418 3703 18474 3712
rect 18602 3768 18658 3777
rect 18602 3703 18658 3712
rect 17788 3590 18092 3606
rect 18156 3590 18276 3618
rect 18432 3602 18460 3703
rect 17696 3488 17816 3516
rect 17592 3470 17644 3476
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17144 2106 17172 2246
rect 17132 2100 17184 2106
rect 17132 2042 17184 2048
rect 17040 1616 17092 1622
rect 1122 1200 1178 1600
rect 2042 1200 2098 1600
rect 2962 1200 3018 1600
rect 3882 1200 3938 1600
rect 4802 1200 4858 1600
rect 5722 1200 5778 1600
rect 6642 1200 6698 1600
rect 7562 1200 7618 1600
rect 8482 1200 8538 1600
rect 9402 1200 9458 1600
rect 10322 1200 10378 1600
rect 11242 1200 11298 1600
rect 12162 1200 12218 1600
rect 13082 1200 13138 1600
rect 14002 1200 14058 1600
rect 14922 1200 14978 1600
rect 15842 1200 15898 1600
rect 16762 1200 16818 1600
rect 17696 1600 17724 2926
rect 17788 2650 17816 3488
rect 18248 3466 18276 3590
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18800 3534 18828 4032
rect 19076 3992 19104 4150
rect 19168 4146 19196 4422
rect 19260 4146 19288 4558
rect 19352 4282 19380 5034
rect 19444 4486 19472 5238
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19444 4146 19472 4422
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 4004 19392 4010
rect 19076 3964 19340 3992
rect 19340 3946 19392 3952
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18892 3641 18920 3878
rect 19444 3738 19472 4082
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19628 3670 19656 5743
rect 19904 5710 19932 6122
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19996 5370 20024 6258
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19812 4826 19840 5102
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19720 4622 19748 4762
rect 19904 4690 19932 5034
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19708 4616 19760 4622
rect 19706 4584 19708 4593
rect 19760 4584 19762 4593
rect 19706 4519 19762 4528
rect 19892 4208 19944 4214
rect 19996 4196 20024 5306
rect 19944 4168 20024 4196
rect 19892 4150 19944 4156
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19156 3664 19208 3670
rect 18878 3632 18934 3641
rect 19156 3606 19208 3612
rect 19248 3664 19300 3670
rect 19248 3606 19300 3612
rect 19616 3664 19668 3670
rect 19616 3606 19668 3612
rect 18878 3567 18934 3576
rect 19168 3534 19196 3606
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18064 2922 18092 2994
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17880 2446 17908 2518
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18156 2378 18184 3402
rect 18248 3126 18276 3402
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18432 2922 18460 3334
rect 18892 2922 18920 3470
rect 19154 3224 19210 3233
rect 19260 3210 19288 3606
rect 19812 3534 19840 3878
rect 20088 3602 20116 6734
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20180 5370 20208 5578
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20180 4282 20208 4762
rect 20272 4622 20300 6394
rect 20824 5681 20852 7278
rect 21088 7200 21140 7206
rect 21008 7148 21088 7154
rect 22928 7200 22980 7206
rect 21008 7142 21140 7148
rect 21822 7168 21878 7177
rect 21008 7126 21128 7142
rect 21008 6662 21036 7126
rect 22928 7142 22980 7148
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 21822 7103 21878 7112
rect 21836 6866 21864 7103
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22374 6896 22430 6905
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21824 6860 21876 6866
rect 22374 6831 22376 6840
rect 21824 6802 21876 6808
rect 22428 6831 22430 6840
rect 22376 6802 22428 6808
rect 20904 6656 20956 6662
rect 20996 6656 21048 6662
rect 20904 6598 20956 6604
rect 20994 6624 20996 6633
rect 21048 6624 21050 6633
rect 20916 6225 20944 6598
rect 20994 6559 21050 6568
rect 20902 6216 20958 6225
rect 20902 6151 20958 6160
rect 20350 5672 20406 5681
rect 20350 5607 20406 5616
rect 20810 5672 20866 5681
rect 20810 5607 20866 5616
rect 20364 4622 20392 5607
rect 20916 5234 20944 6151
rect 21008 6066 21036 6559
rect 21192 6458 21220 6802
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21836 6254 21864 6802
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22388 6322 22416 6666
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22572 6322 22600 6598
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21178 6080 21234 6089
rect 21008 6038 21178 6066
rect 21178 6015 21234 6024
rect 21640 5704 21692 5710
rect 21454 5672 21510 5681
rect 21640 5646 21692 5652
rect 21454 5607 21456 5616
rect 21508 5607 21510 5616
rect 21456 5578 21508 5584
rect 21652 5574 21680 5646
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 20994 5264 21050 5273
rect 20904 5228 20956 5234
rect 21652 5250 21680 5510
rect 21284 5234 21680 5250
rect 20994 5199 21050 5208
rect 21180 5228 21232 5234
rect 20904 5170 20956 5176
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20272 4321 20300 4558
rect 20258 4312 20314 4321
rect 20168 4276 20220 4282
rect 20258 4247 20314 4256
rect 20168 4218 20220 4224
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19432 3392 19484 3398
rect 19616 3392 19668 3398
rect 19432 3334 19484 3340
rect 19614 3360 19616 3369
rect 19668 3360 19670 3369
rect 19352 3233 19380 3334
rect 19210 3182 19288 3210
rect 19338 3224 19394 3233
rect 19154 3159 19210 3168
rect 19338 3159 19394 3168
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18800 2514 18828 2790
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 18984 2446 19012 2790
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18248 1902 18276 2382
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18236 1896 18288 1902
rect 18236 1838 18288 1844
rect 18616 1600 18644 2246
rect 19076 2106 19104 2994
rect 19156 2848 19208 2854
rect 19154 2816 19156 2825
rect 19208 2816 19210 2825
rect 19154 2751 19210 2760
rect 19260 2514 19288 2994
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19352 2446 19380 3159
rect 19444 2990 19472 3334
rect 19614 3295 19670 3304
rect 20180 3058 20208 4218
rect 20258 4176 20314 4185
rect 20258 4111 20314 4120
rect 20272 3738 20300 4111
rect 20548 4049 20576 5102
rect 21008 5030 21036 5199
rect 21284 5228 21692 5234
rect 21284 5222 21640 5228
rect 21284 5216 21312 5222
rect 21232 5188 21312 5216
rect 21180 5170 21232 5176
rect 21640 5170 21692 5176
rect 21086 5128 21142 5137
rect 21086 5063 21142 5072
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 21100 4758 21128 5063
rect 21192 4865 21220 5170
rect 21456 5160 21508 5166
rect 21732 5160 21784 5166
rect 21508 5120 21588 5148
rect 21456 5102 21508 5108
rect 21178 4856 21234 4865
rect 21178 4791 21234 4800
rect 21088 4752 21140 4758
rect 21086 4720 21088 4729
rect 21140 4720 21142 4729
rect 20628 4684 20680 4690
rect 21086 4655 21142 4664
rect 20628 4626 20680 4632
rect 20534 4040 20590 4049
rect 20444 4004 20496 4010
rect 20534 3975 20590 3984
rect 20444 3946 20496 3952
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19064 2100 19116 2106
rect 19064 2042 19116 2048
rect 19536 1600 19564 2994
rect 20272 2990 20300 3538
rect 20456 3534 20484 3946
rect 20640 3942 20668 4626
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 21180 4616 21232 4622
rect 21272 4616 21324 4622
rect 21180 4558 21232 4564
rect 21270 4584 21272 4593
rect 21324 4584 21326 4593
rect 20916 4049 20944 4558
rect 21192 4321 21220 4558
rect 21270 4519 21326 4528
rect 21456 4548 21508 4554
rect 21456 4490 21508 4496
rect 21178 4312 21234 4321
rect 21178 4247 21234 4256
rect 21468 4078 21496 4490
rect 21560 4078 21588 5120
rect 21732 5102 21784 5108
rect 21744 4826 21772 5102
rect 21836 5098 21864 5578
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 22020 4826 22048 6258
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22098 5808 22154 5817
rect 22098 5743 22154 5752
rect 22112 5710 22140 5743
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22204 5574 22232 6054
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22204 5098 22232 5510
rect 22296 5370 22324 6054
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4146 21680 4558
rect 21744 4554 21772 4762
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 22020 4146 22048 4762
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21456 4072 21508 4078
rect 20902 4040 20958 4049
rect 21456 4014 21508 4020
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 20902 3975 20958 3984
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20442 3224 20498 3233
rect 20548 3194 20576 3470
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20442 3159 20498 3168
rect 20536 3188 20588 3194
rect 20456 3058 20484 3159
rect 20536 3130 20588 3136
rect 20444 3052 20496 3058
rect 20364 3012 20444 3040
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20364 2650 20392 3012
rect 20444 2994 20496 3000
rect 20628 3052 20680 3058
rect 20732 3040 20760 3334
rect 20824 3194 20852 3402
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21100 3058 21128 3334
rect 21468 3194 21496 4014
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 20812 3052 20864 3058
rect 20732 3012 20812 3040
rect 20628 2994 20680 3000
rect 20812 2994 20864 3000
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 20640 2854 20668 2994
rect 20628 2848 20680 2854
rect 20824 2825 20852 2994
rect 21468 2961 21496 2994
rect 21454 2952 21510 2961
rect 21454 2887 21510 2896
rect 20628 2790 20680 2796
rect 20810 2816 20866 2825
rect 20810 2751 20866 2760
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20456 1600 20484 2586
rect 21652 2582 21680 3062
rect 22112 2990 22140 4490
rect 22204 2990 22232 5034
rect 22296 5030 22324 5306
rect 22388 5302 22416 5510
rect 22480 5370 22508 6190
rect 22664 5794 22692 6938
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22572 5766 22692 5794
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22572 5030 22600 5766
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22664 5302 22692 5578
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22756 5234 22784 6802
rect 22940 6730 22968 7142
rect 23124 6730 23152 7142
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22284 5024 22336 5030
rect 22560 5024 22612 5030
rect 22284 4966 22336 4972
rect 22558 4992 22560 5001
rect 22612 4992 22614 5001
rect 22558 4927 22614 4936
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22756 4282 22784 4626
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22572 4078 22600 4150
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22296 3058 22324 3402
rect 22284 3052 22336 3058
rect 22336 3012 22416 3040
rect 22284 2994 22336 3000
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21928 2689 21956 2790
rect 21914 2680 21970 2689
rect 22020 2650 22048 2926
rect 22204 2836 22232 2926
rect 22112 2808 22232 2836
rect 21914 2615 21970 2624
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21100 1970 21128 2246
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 21376 1600 21404 2314
rect 22112 1688 22140 2808
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22204 2038 22232 2450
rect 22192 2032 22244 2038
rect 22192 1974 22244 1980
rect 22100 1682 22152 1688
rect 22100 1624 22152 1630
rect 22296 1600 22324 2586
rect 22388 2514 22416 3012
rect 22572 2689 22600 4014
rect 22756 3126 22784 4218
rect 22848 3602 22876 6326
rect 22940 4729 22968 6666
rect 23020 5228 23072 5234
rect 23124 5216 23152 6666
rect 23308 6458 23336 7346
rect 23860 7274 23888 7346
rect 23480 7268 23532 7274
rect 23480 7210 23532 7216
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23400 6390 23428 6598
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23492 5914 23520 7210
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23768 5846 23796 6734
rect 23860 6254 23888 6802
rect 23952 6798 23980 7142
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23846 6080 23902 6089
rect 23846 6015 23902 6024
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23072 5188 23152 5216
rect 23388 5228 23440 5234
rect 23020 5170 23072 5176
rect 23388 5170 23440 5176
rect 22926 4720 22982 4729
rect 22926 4655 22982 4664
rect 23032 4146 23060 5170
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4486 23244 4966
rect 23400 4729 23428 5170
rect 23386 4720 23442 4729
rect 23386 4655 23442 4664
rect 23308 4554 23520 4570
rect 23308 4548 23532 4554
rect 23308 4542 23480 4548
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23308 4282 23336 4542
rect 23480 4490 23532 4496
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 23032 3942 23060 4082
rect 23584 4010 23612 5238
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23032 3670 23060 3878
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 23124 2990 23152 3402
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 22926 2816 22982 2825
rect 22926 2751 22982 2760
rect 22558 2680 22614 2689
rect 22558 2615 22614 2624
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22572 2378 22600 2615
rect 22940 2446 22968 2751
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 22572 1902 22600 2314
rect 22560 1896 22612 1902
rect 22560 1838 22612 1844
rect 23216 1600 23244 3334
rect 23584 3194 23612 3470
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23676 3058 23704 4422
rect 23768 3398 23796 5510
rect 23860 5234 23888 6015
rect 24044 5302 24072 7346
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24136 5681 24164 6326
rect 24412 6118 24440 6734
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 24122 5672 24178 5681
rect 24122 5607 24124 5616
rect 24176 5607 24178 5616
rect 24124 5578 24176 5584
rect 24228 5370 24256 5782
rect 24320 5370 24348 5850
rect 24412 5778 24440 6054
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 24032 5296 24084 5302
rect 24032 5238 24084 5244
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 24044 5166 24072 5238
rect 24320 5234 24348 5306
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4758 24072 5102
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24044 4185 24072 4558
rect 24030 4176 24086 4185
rect 23848 4140 23900 4146
rect 24136 4146 24164 5170
rect 24306 4720 24362 4729
rect 24306 4655 24362 4664
rect 24320 4622 24348 4655
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 4214 24256 4422
rect 24320 4214 24348 4558
rect 24216 4208 24268 4214
rect 24216 4150 24268 4156
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24030 4111 24086 4120
rect 24124 4140 24176 4146
rect 23848 4082 23900 4088
rect 24124 4082 24176 4088
rect 23860 3738 23888 4082
rect 24030 4040 24086 4049
rect 24030 3975 24086 3984
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23952 3534 23980 3878
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23952 3233 23980 3334
rect 23938 3224 23994 3233
rect 23938 3159 23994 3168
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23400 2106 23428 2518
rect 23492 2310 23520 2518
rect 24044 2446 24072 3975
rect 24228 3534 24256 4150
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24122 3224 24178 3233
rect 24122 3159 24124 3168
rect 24176 3159 24178 3168
rect 24124 3130 24176 3136
rect 24412 2922 24440 5170
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24504 4282 24532 4422
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24596 3058 24624 5170
rect 24688 5137 24716 6802
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6458 24992 6666
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24872 5574 24900 6394
rect 25056 5778 25084 7822
rect 25226 7710 25282 8110
rect 26976 8016 27028 8022
rect 26976 7958 27028 7964
rect 27158 7984 27214 7993
rect 26516 7744 26568 7750
rect 25240 7410 25268 7710
rect 26516 7686 26568 7692
rect 26238 7576 26294 7585
rect 26238 7511 26294 7520
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25136 7336 25188 7342
rect 25688 7336 25740 7342
rect 25136 7278 25188 7284
rect 25410 7304 25466 7313
rect 25148 6730 25176 7278
rect 25228 7268 25280 7274
rect 25688 7278 25740 7284
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 25410 7239 25466 7248
rect 25228 7210 25280 7216
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25240 6118 25268 7210
rect 25424 6322 25452 7239
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25516 6254 25544 6598
rect 25700 6497 25728 7278
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 25964 6724 26016 6730
rect 25964 6666 26016 6672
rect 25686 6488 25742 6497
rect 25686 6423 25742 6432
rect 25504 6248 25556 6254
rect 25504 6190 25556 6196
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 25044 5160 25096 5166
rect 24674 5128 24730 5137
rect 25044 5102 25096 5108
rect 24674 5063 24730 5072
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 24860 5092 24912 5098
rect 24860 5034 24912 5040
rect 24674 4176 24730 4185
rect 24674 4111 24730 4120
rect 24688 3942 24716 4111
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24688 3534 24716 3878
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24780 3398 24808 5034
rect 24872 4185 24900 5034
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4282 24992 4966
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 24858 4176 24914 4185
rect 24858 4111 24914 4120
rect 24858 3768 24914 3777
rect 24858 3703 24914 3712
rect 24872 3670 24900 3703
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24858 3360 24914 3369
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24124 2916 24176 2922
rect 24124 2858 24176 2864
rect 24400 2916 24452 2922
rect 24400 2858 24452 2864
rect 24136 2514 24164 2858
rect 24596 2582 24624 2994
rect 24584 2576 24636 2582
rect 24688 2553 24716 3334
rect 24858 3295 24914 3304
rect 24872 3126 24900 3295
rect 24964 3176 24992 4218
rect 25056 4078 25084 5102
rect 25148 4554 25176 5578
rect 25136 4548 25188 4554
rect 25136 4490 25188 4496
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 25148 3194 25176 4490
rect 25240 4078 25268 6054
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25136 3188 25188 3194
rect 24964 3148 25084 3176
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25056 3058 25084 3148
rect 25136 3130 25188 3136
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24872 2582 24900 2926
rect 24964 2689 24992 2994
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 24950 2680 25006 2689
rect 24950 2615 25006 2624
rect 24860 2576 24912 2582
rect 24584 2518 24636 2524
rect 24674 2544 24730 2553
rect 24124 2508 24176 2514
rect 24860 2518 24912 2524
rect 24674 2479 24730 2488
rect 24124 2450 24176 2456
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23480 2304 23532 2310
rect 23952 2281 23980 2382
rect 24964 2310 24992 2615
rect 24216 2304 24268 2310
rect 23480 2246 23532 2252
rect 23938 2272 23994 2281
rect 24216 2246 24268 2252
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 23938 2207 23994 2216
rect 24228 2150 24256 2246
rect 24136 2122 24256 2150
rect 23388 2100 23440 2106
rect 23388 2042 23440 2048
rect 24136 1600 24164 2122
rect 25056 1600 25084 2858
rect 25148 2514 25176 3130
rect 25240 2961 25268 3130
rect 25332 3058 25360 4082
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25226 2952 25282 2961
rect 25226 2887 25282 2896
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25240 2446 25268 2887
rect 25424 2446 25452 5510
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25792 4146 25820 5306
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25608 4026 25636 4082
rect 25608 3998 25820 4026
rect 25792 3942 25820 3998
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25516 1970 25544 2382
rect 25608 2009 25636 3402
rect 25700 3058 25728 3878
rect 25976 3482 26004 6666
rect 26068 6458 26096 7142
rect 26160 6662 26188 7278
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 26160 6361 26188 6598
rect 26146 6352 26202 6361
rect 26146 6287 26202 6296
rect 26252 5710 26280 7511
rect 26528 7410 26556 7686
rect 26988 7546 27016 7958
rect 27158 7919 27214 7928
rect 27344 7948 27396 7954
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 26712 7449 26740 7482
rect 26698 7440 26754 7449
rect 26516 7404 26568 7410
rect 27172 7410 27200 7919
rect 27344 7890 27396 7896
rect 26698 7375 26754 7384
rect 27160 7404 27212 7410
rect 26516 7346 26568 7352
rect 27160 7346 27212 7352
rect 26332 7336 26384 7342
rect 26332 7278 26384 7284
rect 26344 7002 26372 7278
rect 27250 7032 27306 7041
rect 26332 6996 26384 7002
rect 27250 6967 27306 6976
rect 26332 6938 26384 6944
rect 27066 6896 27122 6905
rect 27066 6831 27122 6840
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26344 6390 26372 6598
rect 26528 6497 26556 6734
rect 26514 6488 26570 6497
rect 26436 6446 26514 6474
rect 26332 6384 26384 6390
rect 26332 6326 26384 6332
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26160 5234 26188 5510
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26344 4570 26372 6190
rect 26252 4542 26372 4570
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 25884 3454 26004 3482
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25792 2417 25820 3334
rect 25884 2582 25912 3454
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 25976 2825 26004 3334
rect 25962 2816 26018 2825
rect 25962 2751 26018 2760
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25778 2408 25834 2417
rect 25778 2343 25834 2352
rect 25976 2009 26004 2586
rect 25594 2000 25650 2009
rect 25504 1964 25556 1970
rect 25594 1935 25650 1944
rect 25962 2000 26018 2009
rect 25962 1935 26018 1944
rect 25504 1906 25556 1912
rect 26068 1890 26096 4422
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 26160 3942 26188 4082
rect 26252 4010 26280 4542
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 26252 3738 26280 3946
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26160 2553 26188 3334
rect 26146 2544 26202 2553
rect 26146 2479 26202 2488
rect 25976 1862 26096 1890
rect 25976 1600 26004 1862
rect 26252 1756 26280 3470
rect 26344 3369 26372 4422
rect 26330 3360 26386 3369
rect 26330 3295 26386 3304
rect 26436 2990 26464 6446
rect 26514 6423 26570 6432
rect 26700 6112 26752 6118
rect 26698 6080 26700 6089
rect 26752 6080 26754 6089
rect 26698 6015 26754 6024
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26712 5273 26740 5510
rect 26896 5409 26924 6734
rect 27080 6662 27108 6831
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 27264 6322 27292 6967
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27250 5944 27306 5953
rect 27250 5879 27306 5888
rect 27068 5840 27120 5846
rect 27066 5808 27068 5817
rect 27120 5808 27122 5817
rect 27066 5743 27122 5752
rect 27264 5710 27292 5879
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 26882 5400 26938 5409
rect 26882 5335 26938 5344
rect 26698 5264 26754 5273
rect 26516 5228 26568 5234
rect 26698 5199 26754 5208
rect 27160 5228 27212 5234
rect 26516 5170 26568 5176
rect 27160 5170 27212 5176
rect 26528 4457 26556 5170
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26712 4729 26740 4966
rect 26698 4720 26754 4729
rect 26698 4655 26754 4664
rect 26976 4480 27028 4486
rect 26514 4448 26570 4457
rect 27068 4480 27120 4486
rect 26976 4422 27028 4428
rect 27066 4448 27068 4457
rect 27120 4448 27122 4457
rect 26514 4383 26570 4392
rect 26608 4276 26660 4282
rect 26608 4218 26660 4224
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26528 3913 26556 4082
rect 26514 3904 26570 3913
rect 26514 3839 26570 3848
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26528 2650 26556 2994
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26620 2530 26648 4218
rect 26988 4146 27016 4422
rect 27066 4383 27122 4392
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26712 3641 26740 3878
rect 26698 3632 26754 3641
rect 27080 3602 27108 3878
rect 26698 3567 26754 3576
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 26884 3528 26936 3534
rect 26882 3496 26884 3505
rect 26936 3496 26938 3505
rect 26882 3431 26938 3440
rect 26700 3392 26752 3398
rect 27068 3392 27120 3398
rect 26700 3334 26752 3340
rect 27066 3360 27068 3369
rect 27120 3360 27122 3369
rect 26712 2825 26740 3334
rect 27066 3295 27122 3304
rect 26974 3224 27030 3233
rect 26974 3159 27030 3168
rect 26988 3058 27016 3159
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 26884 2848 26936 2854
rect 26698 2816 26754 2825
rect 26884 2790 26936 2796
rect 26698 2751 26754 2760
rect 26528 2502 26648 2530
rect 26528 2446 26556 2502
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 26700 2304 26752 2310
rect 26700 2246 26752 2252
rect 26712 2038 26740 2246
rect 26700 2032 26752 2038
rect 26700 1974 26752 1980
rect 26240 1750 26292 1756
rect 26240 1692 26292 1698
rect 26804 1688 26832 2382
rect 26792 1682 26844 1688
rect 26792 1624 26844 1630
rect 26896 1600 26924 2790
rect 27080 2106 27108 2926
rect 27068 2100 27120 2106
rect 27068 2042 27120 2048
rect 27172 1834 27200 5170
rect 27356 4622 27384 7890
rect 27434 7712 27490 7721
rect 27618 7710 27674 8110
rect 27434 7647 27490 7656
rect 27448 7546 27476 7647
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27526 7168 27582 7177
rect 27526 7103 27582 7112
rect 27540 6662 27568 7103
rect 27632 6866 27660 7710
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27528 6656 27580 6662
rect 27434 6624 27490 6633
rect 27528 6598 27580 6604
rect 27434 6559 27490 6568
rect 27448 6458 27476 6559
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27434 6352 27490 6361
rect 27434 6287 27490 6296
rect 27448 5914 27476 6287
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27434 5536 27490 5545
rect 27434 5471 27490 5480
rect 27448 5370 27476 5471
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27434 4992 27490 5001
rect 27434 4927 27490 4936
rect 27448 4826 27476 4927
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27344 4616 27396 4622
rect 27344 4558 27396 4564
rect 27434 4176 27490 4185
rect 27434 4111 27490 4120
rect 27448 4010 27476 4111
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27434 3904 27490 3913
rect 27434 3839 27490 3848
rect 27448 3738 27476 3839
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27448 3097 27476 3130
rect 27250 3088 27306 3097
rect 27250 3023 27252 3032
rect 27304 3023 27306 3032
rect 27434 3088 27490 3097
rect 27434 3023 27490 3032
rect 27252 2994 27304 3000
rect 27804 2372 27856 2378
rect 27804 2314 27856 2320
rect 27160 1828 27212 1834
rect 27160 1770 27212 1776
rect 27816 1600 27844 2314
rect 17040 1558 17092 1564
rect 17682 1200 17738 1600
rect 18602 1200 18658 1600
rect 19522 1200 19578 1600
rect 20442 1200 20498 1600
rect 21362 1200 21418 1600
rect 22282 1200 22338 1600
rect 23202 1200 23258 1600
rect 24122 1200 24178 1600
rect 25042 1200 25098 1600
rect 25962 1200 26018 1600
rect 26882 1200 26938 1600
rect 27802 1200 27858 1600
<< via2 >>
rect 1214 7928 1270 7984
rect 1122 7656 1178 7712
rect 1858 7384 1914 7440
rect 2594 7404 2650 7440
rect 2594 7384 2596 7404
rect 2596 7384 2648 7404
rect 2648 7384 2650 7404
rect 1490 7112 1546 7168
rect 2410 6840 2466 6896
rect 2686 6876 2688 6896
rect 2688 6876 2740 6896
rect 2740 6876 2742 6896
rect 2686 6840 2742 6876
rect 1306 6568 1362 6624
rect 1214 6296 1270 6352
rect 2410 6740 2412 6760
rect 2412 6740 2464 6760
rect 2464 6740 2466 6760
rect 1238 6024 1294 6080
rect 1170 5788 1172 5808
rect 1172 5788 1224 5808
rect 1224 5788 1226 5808
rect 1170 5752 1226 5788
rect 2042 5752 2098 5808
rect 1674 5652 1676 5672
rect 1676 5652 1728 5672
rect 1728 5652 1730 5672
rect 1674 5616 1730 5652
rect 1858 5516 1860 5536
rect 1860 5516 1912 5536
rect 1912 5516 1914 5536
rect 1858 5480 1914 5516
rect 1154 5208 1210 5264
rect 1766 5072 1822 5128
rect 1148 4972 1150 4992
rect 1150 4972 1202 4992
rect 1202 4972 1204 4992
rect 1148 4936 1204 4972
rect 1122 4700 1124 4720
rect 1124 4700 1176 4720
rect 1176 4700 1178 4720
rect 1122 4664 1178 4700
rect 1674 4664 1730 4720
rect 1490 4392 1546 4448
rect 1674 3984 1730 4040
rect 1306 3848 1362 3904
rect 1214 3576 1270 3632
rect 1306 3304 1362 3360
rect 1490 3032 1546 3088
rect 1950 4528 2006 4584
rect 1858 4120 1914 4176
rect 1950 3052 2006 3088
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 1858 2760 1914 2816
rect 1030 2488 1086 2544
rect 1306 2216 1362 2272
rect 2410 6704 2466 6740
rect 2226 5208 2282 5264
rect 3330 7248 3386 7304
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 6458 7520 6514 7576
rect 3422 6296 3478 6352
rect 3698 6296 3754 6352
rect 3238 3712 3294 3768
rect 2318 2488 2374 2544
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4434 5344 4490 5400
rect 3606 3712 3662 3768
rect 5906 7112 5962 7168
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3440 4306 3496
rect 4250 2896 4306 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4894 4936 4950 4992
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4802 3712 4858 3768
rect 5078 4120 5134 4176
rect 5170 3848 5226 3904
rect 5446 4256 5502 4312
rect 5078 3440 5134 3496
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 5354 3576 5410 3632
rect 5446 3476 5448 3496
rect 5448 3476 5500 3496
rect 5500 3476 5502 3496
rect 5446 3440 5502 3476
rect 5814 6296 5870 6352
rect 5722 6160 5778 6216
rect 4894 2896 4950 2952
rect 4986 2796 4988 2816
rect 4988 2796 5040 2816
rect 5040 2796 5042 2816
rect 4986 2760 5042 2796
rect 5078 2388 5080 2408
rect 5080 2388 5132 2408
rect 5132 2388 5134 2408
rect 5078 2352 5134 2388
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 3974 1944 4030 2000
rect 5722 3304 5778 3360
rect 6366 3848 6422 3904
rect 5998 3168 6054 3224
rect 6550 6432 6606 6488
rect 6642 6024 6698 6080
rect 6458 3168 6514 3224
rect 7378 5480 7434 5536
rect 7562 7248 7618 7304
rect 7562 5208 7618 5264
rect 9402 7248 9458 7304
rect 7470 4936 7526 4992
rect 7194 3848 7250 3904
rect 7378 3984 7434 4040
rect 7286 3712 7342 3768
rect 7746 5208 7802 5264
rect 8390 5752 8446 5808
rect 8390 5480 8446 5536
rect 8298 5228 8354 5264
rect 8298 5208 8300 5228
rect 8300 5208 8352 5228
rect 8352 5208 8354 5228
rect 7562 3576 7618 3632
rect 7930 4392 7986 4448
rect 7654 3168 7710 3224
rect 8114 3440 8170 3496
rect 8390 4256 8446 4312
rect 8390 3848 8446 3904
rect 8390 3712 8446 3768
rect 8206 2080 8262 2136
rect 8114 1944 8170 2000
rect 9310 6296 9366 6352
rect 9310 5888 9366 5944
rect 8942 5616 8998 5672
rect 8850 4020 8852 4040
rect 8852 4020 8904 4040
rect 8904 4020 8906 4040
rect 8850 3984 8906 4020
rect 9126 5228 9182 5264
rect 9126 5208 9128 5228
rect 9128 5208 9180 5228
rect 9180 5208 9182 5228
rect 8850 3440 8906 3496
rect 8666 2352 8722 2408
rect 9218 3848 9274 3904
rect 9586 6024 9642 6080
rect 9494 5208 9550 5264
rect 9770 5208 9826 5264
rect 9954 4800 10010 4856
rect 9678 4256 9734 4312
rect 9678 4004 9734 4040
rect 9678 3984 9680 4004
rect 9680 3984 9732 4004
rect 9732 3984 9734 4004
rect 9310 3188 9366 3224
rect 9310 3168 9312 3188
rect 9312 3168 9364 3188
rect 9364 3168 9366 3188
rect 9218 2252 9220 2272
rect 9220 2252 9272 2272
rect 9272 2252 9274 2272
rect 9218 2216 9274 2252
rect 9862 3712 9918 3768
rect 10782 6568 10838 6624
rect 10782 5228 10838 5264
rect 10782 5208 10784 5228
rect 10784 5208 10836 5228
rect 10836 5208 10838 5228
rect 10322 3984 10378 4040
rect 10230 3712 10286 3768
rect 10414 2896 10470 2952
rect 10046 2216 10102 2272
rect 11426 7248 11482 7304
rect 12070 6976 12126 7032
rect 12622 6704 12678 6760
rect 12806 6704 12862 6760
rect 12438 5888 12494 5944
rect 12806 6024 12862 6080
rect 10874 3168 10930 3224
rect 11794 3848 11850 3904
rect 12806 4800 12862 4856
rect 12346 3032 12402 3088
rect 11886 2896 11942 2952
rect 12714 3440 12770 3496
rect 13266 6024 13322 6080
rect 13082 4800 13138 4856
rect 13542 5888 13598 5944
rect 13910 6432 13966 6488
rect 14186 6996 14242 7032
rect 14186 6976 14188 6996
rect 14188 6976 14240 6996
rect 14240 6976 14242 6996
rect 12990 3340 12992 3360
rect 12992 3340 13044 3360
rect 13044 3340 13046 3360
rect 12990 3304 13046 3340
rect 12714 3168 12770 3224
rect 13266 3440 13322 3496
rect 13266 2760 13322 2816
rect 13634 5364 13690 5400
rect 13634 5344 13636 5364
rect 13636 5344 13688 5364
rect 13688 5344 13690 5364
rect 13726 4256 13782 4312
rect 14278 6296 14334 6352
rect 14738 6316 14794 6352
rect 14738 6296 14740 6316
rect 14740 6296 14792 6316
rect 14792 6296 14794 6316
rect 14094 6196 14096 6216
rect 14096 6196 14148 6216
rect 14148 6196 14150 6216
rect 14094 6160 14150 6196
rect 14922 5480 14978 5536
rect 16578 7384 16634 7440
rect 15474 6976 15530 7032
rect 15566 6704 15622 6760
rect 16394 6840 16450 6896
rect 15750 6704 15806 6760
rect 14646 3440 14702 3496
rect 15750 5480 15806 5536
rect 16210 5208 16266 5264
rect 15658 5092 15714 5128
rect 15658 5072 15660 5092
rect 15660 5072 15712 5092
rect 15712 5072 15714 5092
rect 14922 3848 14978 3904
rect 15750 4936 15806 4992
rect 15842 4700 15844 4720
rect 15844 4700 15896 4720
rect 15896 4700 15898 4720
rect 15842 4664 15898 4700
rect 16210 4428 16212 4448
rect 16212 4428 16264 4448
rect 16264 4428 16266 4448
rect 16210 4392 16266 4428
rect 16670 6976 16726 7032
rect 14922 3168 14978 3224
rect 14830 3032 14886 3088
rect 15750 3884 15752 3904
rect 15752 3884 15804 3904
rect 15804 3884 15806 3904
rect 15750 3848 15806 3884
rect 17866 6840 17922 6896
rect 17774 6432 17830 6488
rect 17590 5752 17646 5808
rect 17038 5516 17040 5536
rect 17040 5516 17092 5536
rect 17092 5516 17094 5536
rect 16762 4528 16818 4584
rect 17038 5480 17094 5516
rect 17038 4664 17094 4720
rect 17130 4528 17186 4584
rect 16486 4120 16542 4176
rect 16946 4120 17002 4176
rect 17866 5480 17922 5536
rect 17406 3712 17462 3768
rect 17774 4256 17830 4312
rect 17958 4276 18014 4312
rect 17958 4256 17960 4276
rect 17960 4256 18012 4276
rect 18012 4256 18014 4276
rect 18510 5616 18566 5672
rect 18694 6740 18696 6760
rect 18696 6740 18748 6760
rect 18748 6740 18750 6760
rect 18694 6704 18750 6740
rect 18786 6568 18842 6624
rect 18602 4528 18658 4584
rect 18878 5364 18934 5400
rect 18878 5344 18880 5364
rect 18880 5344 18932 5364
rect 18932 5344 18934 5364
rect 19338 5752 19394 5808
rect 19062 5344 19118 5400
rect 19430 5480 19486 5536
rect 19982 6432 20038 6488
rect 19614 5752 19670 5808
rect 18970 4528 19026 4584
rect 18878 4256 18934 4312
rect 19154 4528 19210 4584
rect 18418 3712 18474 3768
rect 18602 3712 18658 3768
rect 19706 4564 19708 4584
rect 19708 4564 19760 4584
rect 19760 4564 19762 4584
rect 19706 4528 19762 4564
rect 18878 3576 18934 3632
rect 19154 3168 19210 3224
rect 21822 7112 21878 7168
rect 22374 6860 22430 6896
rect 22374 6840 22376 6860
rect 22376 6840 22428 6860
rect 22428 6840 22430 6860
rect 20994 6604 20996 6624
rect 20996 6604 21048 6624
rect 21048 6604 21050 6624
rect 20994 6568 21050 6604
rect 20902 6160 20958 6216
rect 20350 5616 20406 5672
rect 20810 5616 20866 5672
rect 21178 6024 21234 6080
rect 21454 5636 21510 5672
rect 21454 5616 21456 5636
rect 21456 5616 21508 5636
rect 21508 5616 21510 5636
rect 20994 5208 21050 5264
rect 20258 4256 20314 4312
rect 19614 3340 19616 3360
rect 19616 3340 19668 3360
rect 19668 3340 19670 3360
rect 19338 3168 19394 3224
rect 19154 2796 19156 2816
rect 19156 2796 19208 2816
rect 19208 2796 19210 2816
rect 19154 2760 19210 2796
rect 19614 3304 19670 3340
rect 20258 4120 20314 4176
rect 21086 5072 21142 5128
rect 21178 4800 21234 4856
rect 21086 4700 21088 4720
rect 21088 4700 21140 4720
rect 21140 4700 21142 4720
rect 21086 4664 21142 4700
rect 20534 3984 20590 4040
rect 21270 4564 21272 4584
rect 21272 4564 21324 4584
rect 21324 4564 21326 4584
rect 21270 4528 21326 4564
rect 21178 4256 21234 4312
rect 22098 5752 22154 5808
rect 20902 3984 20958 4040
rect 20442 3168 20498 3224
rect 21454 2896 21510 2952
rect 20810 2760 20866 2816
rect 22558 4972 22560 4992
rect 22560 4972 22612 4992
rect 22612 4972 22614 4992
rect 22558 4936 22614 4972
rect 21914 2624 21970 2680
rect 23846 6024 23902 6080
rect 22926 4664 22982 4720
rect 23386 4664 23442 4720
rect 22926 2760 22982 2816
rect 22558 2624 22614 2680
rect 24122 5636 24178 5672
rect 24122 5616 24124 5636
rect 24124 5616 24176 5636
rect 24176 5616 24178 5636
rect 24030 4120 24086 4176
rect 24306 4664 24362 4720
rect 24030 3984 24086 4040
rect 23938 3168 23994 3224
rect 24122 3188 24178 3224
rect 24122 3168 24124 3188
rect 24124 3168 24176 3188
rect 24176 3168 24178 3188
rect 26238 7520 26294 7576
rect 25410 7248 25466 7304
rect 25686 6432 25742 6488
rect 24674 5072 24730 5128
rect 24674 4120 24730 4176
rect 24858 4120 24914 4176
rect 24858 3712 24914 3768
rect 24858 3304 24914 3360
rect 24950 2624 25006 2680
rect 24674 2488 24730 2544
rect 23938 2216 23994 2272
rect 25226 2896 25282 2952
rect 26146 6296 26202 6352
rect 27158 7928 27214 7984
rect 26698 7384 26754 7440
rect 27250 6976 27306 7032
rect 27066 6840 27122 6896
rect 25962 2760 26018 2816
rect 25778 2352 25834 2408
rect 25594 1944 25650 2000
rect 25962 1944 26018 2000
rect 26146 2488 26202 2544
rect 26330 3304 26386 3360
rect 26514 6432 26570 6488
rect 26698 6060 26700 6080
rect 26700 6060 26752 6080
rect 26752 6060 26754 6080
rect 26698 6024 26754 6060
rect 27250 5888 27306 5944
rect 27066 5788 27068 5808
rect 27068 5788 27120 5808
rect 27120 5788 27122 5808
rect 27066 5752 27122 5788
rect 26882 5344 26938 5400
rect 26698 5208 26754 5264
rect 26698 4664 26754 4720
rect 26514 4392 26570 4448
rect 27066 4428 27068 4448
rect 27068 4428 27120 4448
rect 27120 4428 27122 4448
rect 26514 3848 26570 3904
rect 27066 4392 27122 4428
rect 26698 3576 26754 3632
rect 26882 3476 26884 3496
rect 26884 3476 26936 3496
rect 26936 3476 26938 3496
rect 26882 3440 26938 3476
rect 27066 3340 27068 3360
rect 27068 3340 27120 3360
rect 27120 3340 27122 3360
rect 27066 3304 27122 3340
rect 26974 3168 27030 3224
rect 26698 2760 26754 2816
rect 27434 7656 27490 7712
rect 27526 7112 27582 7168
rect 27434 6568 27490 6624
rect 27434 6296 27490 6352
rect 27434 5480 27490 5536
rect 27434 4936 27490 4992
rect 27434 4120 27490 4176
rect 27434 3848 27490 3904
rect 27250 3052 27306 3088
rect 27250 3032 27252 3052
rect 27252 3032 27304 3052
rect 27304 3032 27306 3052
rect 27434 3032 27490 3088
<< metal3 >>
rect 560 7986 960 8016
rect 1209 7986 1275 7989
rect 560 7984 1275 7986
rect 560 7928 1214 7984
rect 1270 7928 1275 7984
rect 560 7926 1275 7928
rect 560 7896 960 7926
rect 1209 7923 1275 7926
rect 27153 7986 27219 7989
rect 28020 7986 28420 8016
rect 27153 7984 28420 7986
rect 27153 7928 27158 7984
rect 27214 7928 28420 7984
rect 27153 7926 28420 7928
rect 27153 7923 27219 7926
rect 28020 7896 28420 7926
rect 560 7714 960 7744
rect 1117 7714 1183 7717
rect 560 7712 1183 7714
rect 560 7656 1122 7712
rect 1178 7656 1183 7712
rect 560 7654 1183 7656
rect 560 7624 960 7654
rect 1117 7651 1183 7654
rect 27429 7714 27495 7717
rect 28020 7714 28420 7744
rect 27429 7712 28420 7714
rect 27429 7656 27434 7712
rect 27490 7656 28420 7712
rect 27429 7654 28420 7656
rect 27429 7651 27495 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 28020 7624 28420 7654
rect 4870 7583 5186 7584
rect 6453 7578 6519 7581
rect 26233 7578 26299 7581
rect 6453 7576 26299 7578
rect 6453 7520 6458 7576
rect 6514 7520 26238 7576
rect 26294 7520 26299 7576
rect 6453 7518 26299 7520
rect 6453 7515 6519 7518
rect 26233 7515 26299 7518
rect 560 7442 960 7472
rect 1853 7442 1919 7445
rect 560 7440 1919 7442
rect 560 7384 1858 7440
rect 1914 7384 1919 7440
rect 560 7382 1919 7384
rect 560 7352 960 7382
rect 1853 7379 1919 7382
rect 2589 7442 2655 7445
rect 16573 7442 16639 7445
rect 2589 7440 16639 7442
rect 2589 7384 2594 7440
rect 2650 7384 16578 7440
rect 16634 7384 16639 7440
rect 2589 7382 16639 7384
rect 2589 7379 2655 7382
rect 16573 7379 16639 7382
rect 26693 7442 26759 7445
rect 28020 7442 28420 7472
rect 26693 7440 28420 7442
rect 26693 7384 26698 7440
rect 26754 7384 28420 7440
rect 26693 7382 28420 7384
rect 26693 7379 26759 7382
rect 28020 7352 28420 7382
rect 3325 7306 3391 7309
rect 7557 7306 7623 7309
rect 9397 7306 9463 7309
rect 3325 7304 9463 7306
rect 3325 7248 3330 7304
rect 3386 7248 7562 7304
rect 7618 7248 9402 7304
rect 9458 7248 9463 7304
rect 3325 7246 9463 7248
rect 3325 7243 3391 7246
rect 7557 7243 7623 7246
rect 9397 7243 9463 7246
rect 11421 7306 11487 7309
rect 25405 7306 25471 7309
rect 11421 7304 25471 7306
rect 11421 7248 11426 7304
rect 11482 7248 25410 7304
rect 25466 7248 25471 7304
rect 11421 7246 25471 7248
rect 11421 7243 11487 7246
rect 25405 7243 25471 7246
rect 560 7170 960 7200
rect 1485 7170 1551 7173
rect 560 7168 1551 7170
rect 560 7112 1490 7168
rect 1546 7112 1551 7168
rect 560 7110 1551 7112
rect 560 7080 960 7110
rect 1485 7107 1551 7110
rect 5901 7170 5967 7173
rect 21817 7170 21883 7173
rect 5901 7168 21883 7170
rect 5901 7112 5906 7168
rect 5962 7112 21822 7168
rect 21878 7112 21883 7168
rect 5901 7110 21883 7112
rect 5901 7107 5967 7110
rect 21817 7107 21883 7110
rect 27521 7170 27587 7173
rect 28020 7170 28420 7200
rect 27521 7168 28420 7170
rect 27521 7112 27526 7168
rect 27582 7112 28420 7168
rect 27521 7110 28420 7112
rect 27521 7107 27587 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 28020 7080 28420 7110
rect 4210 7039 4526 7040
rect 12065 7034 12131 7037
rect 14181 7034 14247 7037
rect 15469 7034 15535 7037
rect 12065 7032 15535 7034
rect 12065 6976 12070 7032
rect 12126 6976 14186 7032
rect 14242 6976 15474 7032
rect 15530 6976 15535 7032
rect 12065 6974 15535 6976
rect 12065 6971 12131 6974
rect 14181 6971 14247 6974
rect 15469 6971 15535 6974
rect 16665 7034 16731 7037
rect 27245 7034 27311 7037
rect 16665 7032 27311 7034
rect 16665 6976 16670 7032
rect 16726 6976 27250 7032
rect 27306 6976 27311 7032
rect 16665 6974 27311 6976
rect 16665 6971 16731 6974
rect 27245 6971 27311 6974
rect 560 6898 960 6928
rect 2405 6898 2471 6901
rect 560 6896 2471 6898
rect 560 6840 2410 6896
rect 2466 6840 2471 6896
rect 560 6838 2471 6840
rect 560 6808 960 6838
rect 2405 6835 2471 6838
rect 2681 6898 2747 6901
rect 16389 6898 16455 6901
rect 2681 6896 16455 6898
rect 2681 6840 2686 6896
rect 2742 6840 16394 6896
rect 16450 6840 16455 6896
rect 2681 6838 16455 6840
rect 2681 6835 2747 6838
rect 16389 6835 16455 6838
rect 17861 6898 17927 6901
rect 22369 6898 22435 6901
rect 17861 6896 22435 6898
rect 17861 6840 17866 6896
rect 17922 6840 22374 6896
rect 22430 6840 22435 6896
rect 17861 6838 22435 6840
rect 17861 6835 17927 6838
rect 22369 6835 22435 6838
rect 27061 6898 27127 6901
rect 28020 6898 28420 6928
rect 27061 6896 28420 6898
rect 27061 6840 27066 6896
rect 27122 6840 28420 6896
rect 27061 6838 28420 6840
rect 27061 6835 27127 6838
rect 28020 6808 28420 6838
rect 2405 6762 2471 6765
rect 12617 6762 12683 6765
rect 2405 6760 12683 6762
rect 2405 6704 2410 6760
rect 2466 6704 12622 6760
rect 12678 6704 12683 6760
rect 2405 6702 12683 6704
rect 2405 6699 2471 6702
rect 12617 6699 12683 6702
rect 12801 6762 12867 6765
rect 15561 6762 15627 6765
rect 12801 6760 15627 6762
rect 12801 6704 12806 6760
rect 12862 6704 15566 6760
rect 15622 6704 15627 6760
rect 12801 6702 15627 6704
rect 12801 6699 12867 6702
rect 15561 6699 15627 6702
rect 15745 6762 15811 6765
rect 18689 6762 18755 6765
rect 15745 6760 18755 6762
rect 15745 6704 15750 6760
rect 15806 6704 18694 6760
rect 18750 6704 18755 6760
rect 15745 6702 18755 6704
rect 15745 6699 15811 6702
rect 18689 6699 18755 6702
rect 560 6626 960 6656
rect 1301 6626 1367 6629
rect 560 6624 1367 6626
rect 560 6568 1306 6624
rect 1362 6568 1367 6624
rect 560 6566 1367 6568
rect 560 6536 960 6566
rect 1301 6563 1367 6566
rect 10777 6626 10843 6629
rect 18781 6626 18847 6629
rect 20989 6626 21055 6629
rect 10777 6624 21055 6626
rect 10777 6568 10782 6624
rect 10838 6568 18786 6624
rect 18842 6568 20994 6624
rect 21050 6568 21055 6624
rect 10777 6566 21055 6568
rect 10777 6563 10843 6566
rect 18781 6563 18847 6566
rect 20989 6563 21055 6566
rect 27429 6626 27495 6629
rect 28020 6626 28420 6656
rect 27429 6624 28420 6626
rect 27429 6568 27434 6624
rect 27490 6568 28420 6624
rect 27429 6566 28420 6568
rect 27429 6563 27495 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 28020 6536 28420 6566
rect 4870 6495 5186 6496
rect 6545 6490 6611 6493
rect 13905 6490 13971 6493
rect 6545 6488 13971 6490
rect 6545 6432 6550 6488
rect 6606 6432 13910 6488
rect 13966 6432 13971 6488
rect 6545 6430 13971 6432
rect 6545 6427 6611 6430
rect 13905 6427 13971 6430
rect 17769 6490 17835 6493
rect 19977 6490 20043 6493
rect 25681 6490 25747 6493
rect 26509 6490 26575 6493
rect 17769 6488 26575 6490
rect 17769 6432 17774 6488
rect 17830 6432 19982 6488
rect 20038 6432 25686 6488
rect 25742 6432 26514 6488
rect 26570 6432 26575 6488
rect 17769 6430 26575 6432
rect 17769 6427 17835 6430
rect 19977 6427 20043 6430
rect 25681 6427 25747 6430
rect 26509 6427 26575 6430
rect 560 6354 960 6384
rect 1209 6354 1275 6357
rect 560 6352 1275 6354
rect 560 6296 1214 6352
rect 1270 6296 1275 6352
rect 560 6294 1275 6296
rect 560 6264 960 6294
rect 1209 6291 1275 6294
rect 3417 6354 3483 6357
rect 3693 6354 3759 6357
rect 5809 6354 5875 6357
rect 3417 6352 5875 6354
rect 3417 6296 3422 6352
rect 3478 6296 3698 6352
rect 3754 6296 5814 6352
rect 5870 6296 5875 6352
rect 3417 6294 5875 6296
rect 3417 6291 3483 6294
rect 3693 6291 3759 6294
rect 5809 6291 5875 6294
rect 9305 6354 9371 6357
rect 14273 6354 14339 6357
rect 14733 6354 14799 6357
rect 26141 6354 26207 6357
rect 9305 6352 26207 6354
rect 9305 6296 9310 6352
rect 9366 6296 14278 6352
rect 14334 6296 14738 6352
rect 14794 6296 26146 6352
rect 26202 6296 26207 6352
rect 9305 6294 26207 6296
rect 9305 6291 9371 6294
rect 14273 6291 14339 6294
rect 14733 6291 14799 6294
rect 26141 6291 26207 6294
rect 27429 6354 27495 6357
rect 28020 6354 28420 6384
rect 27429 6352 28420 6354
rect 27429 6296 27434 6352
rect 27490 6296 28420 6352
rect 27429 6294 28420 6296
rect 27429 6291 27495 6294
rect 28020 6264 28420 6294
rect 5717 6218 5783 6221
rect 14089 6218 14155 6221
rect 20897 6218 20963 6221
rect 5717 6216 20963 6218
rect 5717 6160 5722 6216
rect 5778 6160 14094 6216
rect 14150 6160 20902 6216
rect 20958 6160 20963 6216
rect 5717 6158 20963 6160
rect 5717 6155 5783 6158
rect 14089 6155 14155 6158
rect 20897 6155 20963 6158
rect 560 6082 960 6112
rect 1233 6082 1299 6085
rect 560 6080 1299 6082
rect 560 6024 1238 6080
rect 1294 6024 1299 6080
rect 560 6022 1299 6024
rect 560 5992 960 6022
rect 1233 6019 1299 6022
rect 6637 6082 6703 6085
rect 9581 6082 9647 6085
rect 6637 6080 9647 6082
rect 6637 6024 6642 6080
rect 6698 6024 9586 6080
rect 9642 6024 9647 6080
rect 6637 6022 9647 6024
rect 6637 6019 6703 6022
rect 9581 6019 9647 6022
rect 12801 6082 12867 6085
rect 13261 6082 13327 6085
rect 12801 6080 13327 6082
rect 12801 6024 12806 6080
rect 12862 6024 13266 6080
rect 13322 6024 13327 6080
rect 12801 6022 13327 6024
rect 12801 6019 12867 6022
rect 13261 6019 13327 6022
rect 21173 6082 21239 6085
rect 23841 6082 23907 6085
rect 21173 6080 23907 6082
rect 21173 6024 21178 6080
rect 21234 6024 23846 6080
rect 23902 6024 23907 6080
rect 21173 6022 23907 6024
rect 21173 6019 21239 6022
rect 23841 6019 23907 6022
rect 26693 6082 26759 6085
rect 28020 6082 28420 6112
rect 26693 6080 28420 6082
rect 26693 6024 26698 6080
rect 26754 6024 28420 6080
rect 26693 6022 28420 6024
rect 26693 6019 26759 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 28020 5992 28420 6022
rect 4210 5951 4526 5952
rect 9305 5946 9371 5949
rect 8158 5944 9371 5946
rect 8158 5888 9310 5944
rect 9366 5888 9371 5944
rect 8158 5886 9371 5888
rect 560 5810 960 5840
rect 1165 5810 1231 5813
rect 560 5808 1231 5810
rect 560 5752 1170 5808
rect 1226 5752 1231 5808
rect 560 5750 1231 5752
rect 560 5720 960 5750
rect 1165 5747 1231 5750
rect 2037 5810 2103 5813
rect 8158 5810 8218 5886
rect 9305 5883 9371 5886
rect 12433 5946 12499 5949
rect 13537 5946 13603 5949
rect 27245 5946 27311 5949
rect 12433 5944 27311 5946
rect 12433 5888 12438 5944
rect 12494 5888 13542 5944
rect 13598 5888 27250 5944
rect 27306 5888 27311 5944
rect 12433 5886 27311 5888
rect 12433 5883 12499 5886
rect 13537 5883 13603 5886
rect 27245 5883 27311 5886
rect 2037 5808 8218 5810
rect 2037 5752 2042 5808
rect 2098 5752 8218 5808
rect 2037 5750 8218 5752
rect 8385 5810 8451 5813
rect 17585 5810 17651 5813
rect 19333 5810 19399 5813
rect 8385 5808 16590 5810
rect 8385 5752 8390 5808
rect 8446 5752 16590 5808
rect 8385 5750 16590 5752
rect 2037 5747 2103 5750
rect 8385 5747 8451 5750
rect 1669 5674 1735 5677
rect 8937 5674 9003 5677
rect 1669 5672 9003 5674
rect 1669 5616 1674 5672
rect 1730 5616 8942 5672
rect 8998 5616 9003 5672
rect 1669 5614 9003 5616
rect 16530 5674 16590 5750
rect 17585 5808 19399 5810
rect 17585 5752 17590 5808
rect 17646 5752 19338 5808
rect 19394 5752 19399 5808
rect 17585 5750 19399 5752
rect 17585 5747 17651 5750
rect 19333 5747 19399 5750
rect 19609 5810 19675 5813
rect 22093 5810 22159 5813
rect 19609 5808 22159 5810
rect 19609 5752 19614 5808
rect 19670 5752 22098 5808
rect 22154 5752 22159 5808
rect 19609 5750 22159 5752
rect 19609 5747 19675 5750
rect 22093 5747 22159 5750
rect 27061 5810 27127 5813
rect 28020 5810 28420 5840
rect 27061 5808 28420 5810
rect 27061 5752 27066 5808
rect 27122 5752 28420 5808
rect 27061 5750 28420 5752
rect 27061 5747 27127 5750
rect 28020 5720 28420 5750
rect 18505 5674 18571 5677
rect 20345 5674 20411 5677
rect 16530 5672 20411 5674
rect 16530 5616 18510 5672
rect 18566 5616 20350 5672
rect 20406 5616 20411 5672
rect 16530 5614 20411 5616
rect 1669 5611 1735 5614
rect 8937 5611 9003 5614
rect 18505 5611 18571 5614
rect 20345 5611 20411 5614
rect 20805 5674 20871 5677
rect 21449 5674 21515 5677
rect 24117 5674 24183 5677
rect 20805 5672 24183 5674
rect 20805 5616 20810 5672
rect 20866 5616 21454 5672
rect 21510 5616 24122 5672
rect 24178 5616 24183 5672
rect 20805 5614 24183 5616
rect 20805 5611 20871 5614
rect 21449 5611 21515 5614
rect 24117 5611 24183 5614
rect 560 5538 960 5568
rect 1853 5538 1919 5541
rect 560 5536 1919 5538
rect 560 5480 1858 5536
rect 1914 5480 1919 5536
rect 560 5478 1919 5480
rect 560 5448 960 5478
rect 1853 5475 1919 5478
rect 7373 5538 7439 5541
rect 8385 5538 8451 5541
rect 7373 5536 8451 5538
rect 7373 5480 7378 5536
rect 7434 5480 8390 5536
rect 8446 5480 8451 5536
rect 7373 5478 8451 5480
rect 7373 5475 7439 5478
rect 8385 5475 8451 5478
rect 14917 5538 14983 5541
rect 15745 5538 15811 5541
rect 14917 5536 15811 5538
rect 14917 5480 14922 5536
rect 14978 5480 15750 5536
rect 15806 5480 15811 5536
rect 14917 5478 15811 5480
rect 14917 5475 14983 5478
rect 15745 5475 15811 5478
rect 17033 5538 17099 5541
rect 17861 5538 17927 5541
rect 19425 5540 19491 5541
rect 19374 5538 19380 5540
rect 17033 5536 17927 5538
rect 17033 5480 17038 5536
rect 17094 5480 17866 5536
rect 17922 5480 17927 5536
rect 17033 5478 17927 5480
rect 19334 5478 19380 5538
rect 19444 5536 19491 5540
rect 19486 5480 19491 5536
rect 17033 5475 17099 5478
rect 17861 5475 17927 5478
rect 19374 5476 19380 5478
rect 19444 5476 19491 5480
rect 19425 5475 19491 5476
rect 27429 5538 27495 5541
rect 28020 5538 28420 5568
rect 27429 5536 28420 5538
rect 27429 5480 27434 5536
rect 27490 5480 28420 5536
rect 27429 5478 28420 5480
rect 27429 5475 27495 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 28020 5448 28420 5478
rect 4870 5407 5186 5408
rect 4429 5402 4495 5405
rect 4654 5402 4660 5404
rect 4429 5400 4660 5402
rect 4429 5344 4434 5400
rect 4490 5344 4660 5400
rect 4429 5342 4660 5344
rect 4429 5339 4495 5342
rect 4654 5340 4660 5342
rect 4724 5340 4730 5404
rect 13629 5402 13695 5405
rect 18873 5402 18939 5405
rect 13629 5400 18939 5402
rect 13629 5344 13634 5400
rect 13690 5344 18878 5400
rect 18934 5344 18939 5400
rect 13629 5342 18939 5344
rect 13629 5339 13695 5342
rect 18873 5339 18939 5342
rect 19057 5402 19123 5405
rect 26877 5402 26943 5405
rect 19057 5400 26943 5402
rect 19057 5344 19062 5400
rect 19118 5344 26882 5400
rect 26938 5344 26943 5400
rect 19057 5342 26943 5344
rect 19057 5339 19123 5342
rect 26877 5339 26943 5342
rect 560 5266 960 5296
rect 1149 5266 1215 5269
rect 560 5264 1215 5266
rect 560 5208 1154 5264
rect 1210 5208 1215 5264
rect 560 5206 1215 5208
rect 560 5176 960 5206
rect 1149 5203 1215 5206
rect 2221 5266 2287 5269
rect 7557 5266 7623 5269
rect 2221 5264 7623 5266
rect 2221 5208 2226 5264
rect 2282 5208 7562 5264
rect 7618 5208 7623 5264
rect 2221 5206 7623 5208
rect 2221 5203 2287 5206
rect 7557 5203 7623 5206
rect 7741 5266 7807 5269
rect 8293 5266 8359 5269
rect 7741 5264 8359 5266
rect 7741 5208 7746 5264
rect 7802 5208 8298 5264
rect 8354 5208 8359 5264
rect 7741 5206 8359 5208
rect 7741 5203 7807 5206
rect 8293 5203 8359 5206
rect 9121 5266 9187 5269
rect 9489 5266 9555 5269
rect 9765 5266 9831 5269
rect 9121 5264 9831 5266
rect 9121 5208 9126 5264
rect 9182 5208 9494 5264
rect 9550 5208 9770 5264
rect 9826 5208 9831 5264
rect 9121 5206 9831 5208
rect 9121 5203 9187 5206
rect 9489 5203 9555 5206
rect 9765 5203 9831 5206
rect 10777 5266 10843 5269
rect 16205 5266 16271 5269
rect 20989 5266 21055 5269
rect 10777 5264 21055 5266
rect 10777 5208 10782 5264
rect 10838 5208 16210 5264
rect 16266 5208 20994 5264
rect 21050 5208 21055 5264
rect 10777 5206 21055 5208
rect 10777 5203 10843 5206
rect 16205 5203 16271 5206
rect 20989 5203 21055 5206
rect 26693 5266 26759 5269
rect 28020 5266 28420 5296
rect 26693 5264 28420 5266
rect 26693 5208 26698 5264
rect 26754 5208 28420 5264
rect 26693 5206 28420 5208
rect 26693 5203 26759 5206
rect 28020 5176 28420 5206
rect 1761 5130 1827 5133
rect 15653 5130 15719 5133
rect 1761 5128 15719 5130
rect 1761 5072 1766 5128
rect 1822 5072 15658 5128
rect 15714 5072 15719 5128
rect 1761 5070 15719 5072
rect 1761 5067 1827 5070
rect 15653 5067 15719 5070
rect 21081 5130 21147 5133
rect 24669 5130 24735 5133
rect 21081 5128 24735 5130
rect 21081 5072 21086 5128
rect 21142 5072 24674 5128
rect 24730 5072 24735 5128
rect 21081 5070 24735 5072
rect 21081 5067 21147 5070
rect 24669 5067 24735 5070
rect 560 4994 960 5024
rect 1143 4994 1209 4997
rect 560 4992 1209 4994
rect 560 4936 1148 4992
rect 1204 4936 1209 4992
rect 560 4934 1209 4936
rect 560 4904 960 4934
rect 1143 4931 1209 4934
rect 4889 4994 4955 4997
rect 7465 4994 7531 4997
rect 4889 4992 7531 4994
rect 4889 4936 4894 4992
rect 4950 4936 7470 4992
rect 7526 4936 7531 4992
rect 4889 4934 7531 4936
rect 4889 4931 4955 4934
rect 7465 4931 7531 4934
rect 15745 4994 15811 4997
rect 22553 4994 22619 4997
rect 15745 4992 22619 4994
rect 15745 4936 15750 4992
rect 15806 4936 22558 4992
rect 22614 4936 22619 4992
rect 15745 4934 22619 4936
rect 15745 4931 15811 4934
rect 22553 4931 22619 4934
rect 27429 4994 27495 4997
rect 28020 4994 28420 5024
rect 27429 4992 28420 4994
rect 27429 4936 27434 4992
rect 27490 4936 28420 4992
rect 27429 4934 28420 4936
rect 27429 4931 27495 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 28020 4904 28420 4934
rect 4210 4863 4526 4864
rect 9949 4858 10015 4861
rect 12801 4858 12867 4861
rect 9949 4856 12867 4858
rect 9949 4800 9954 4856
rect 10010 4800 12806 4856
rect 12862 4800 12867 4856
rect 9949 4798 12867 4800
rect 9949 4795 10015 4798
rect 12801 4795 12867 4798
rect 13077 4858 13143 4861
rect 21173 4858 21239 4861
rect 13077 4856 21239 4858
rect 13077 4800 13082 4856
rect 13138 4800 21178 4856
rect 21234 4800 21239 4856
rect 13077 4798 21239 4800
rect 13077 4795 13143 4798
rect 21173 4795 21239 4798
rect 560 4722 960 4752
rect 1117 4722 1183 4725
rect 560 4720 1183 4722
rect 560 4664 1122 4720
rect 1178 4664 1183 4720
rect 560 4662 1183 4664
rect 560 4632 960 4662
rect 1117 4659 1183 4662
rect 1669 4722 1735 4725
rect 15837 4722 15903 4725
rect 1669 4720 15903 4722
rect 1669 4664 1674 4720
rect 1730 4664 15842 4720
rect 15898 4664 15903 4720
rect 1669 4662 15903 4664
rect 1669 4659 1735 4662
rect 15837 4659 15903 4662
rect 17033 4722 17099 4725
rect 21081 4722 21147 4725
rect 17033 4720 21147 4722
rect 17033 4664 17038 4720
rect 17094 4664 21086 4720
rect 21142 4664 21147 4720
rect 17033 4662 21147 4664
rect 17033 4659 17099 4662
rect 21081 4659 21147 4662
rect 22921 4722 22987 4725
rect 23381 4722 23447 4725
rect 24301 4722 24367 4725
rect 22921 4720 24367 4722
rect 22921 4664 22926 4720
rect 22982 4664 23386 4720
rect 23442 4664 24306 4720
rect 24362 4664 24367 4720
rect 22921 4662 24367 4664
rect 22921 4659 22987 4662
rect 23381 4659 23447 4662
rect 24301 4659 24367 4662
rect 26693 4722 26759 4725
rect 28020 4722 28420 4752
rect 26693 4720 28420 4722
rect 26693 4664 26698 4720
rect 26754 4664 28420 4720
rect 26693 4662 28420 4664
rect 26693 4659 26759 4662
rect 28020 4632 28420 4662
rect 1945 4586 2011 4589
rect 16757 4586 16823 4589
rect 1945 4584 16823 4586
rect 1945 4528 1950 4584
rect 2006 4528 16762 4584
rect 16818 4528 16823 4584
rect 1945 4526 16823 4528
rect 1945 4523 2011 4526
rect 16757 4523 16823 4526
rect 17125 4586 17191 4589
rect 18597 4586 18663 4589
rect 17125 4584 18663 4586
rect 17125 4528 17130 4584
rect 17186 4528 18602 4584
rect 18658 4528 18663 4584
rect 17125 4526 18663 4528
rect 17125 4523 17191 4526
rect 18597 4523 18663 4526
rect 18965 4586 19031 4589
rect 19149 4586 19215 4589
rect 18965 4584 19215 4586
rect 18965 4528 18970 4584
rect 19026 4528 19154 4584
rect 19210 4528 19215 4584
rect 18965 4526 19215 4528
rect 18965 4523 19031 4526
rect 19149 4523 19215 4526
rect 19701 4586 19767 4589
rect 21265 4586 21331 4589
rect 19701 4584 21331 4586
rect 19701 4528 19706 4584
rect 19762 4528 21270 4584
rect 21326 4528 21331 4584
rect 19701 4526 21331 4528
rect 19701 4523 19767 4526
rect 21265 4523 21331 4526
rect 560 4450 960 4480
rect 1485 4450 1551 4453
rect 560 4448 1551 4450
rect 560 4392 1490 4448
rect 1546 4392 1551 4448
rect 560 4390 1551 4392
rect 560 4360 960 4390
rect 1485 4387 1551 4390
rect 7925 4450 7991 4453
rect 8702 4450 8708 4452
rect 7925 4448 8708 4450
rect 7925 4392 7930 4448
rect 7986 4392 8708 4448
rect 7925 4390 8708 4392
rect 7925 4387 7991 4390
rect 8702 4388 8708 4390
rect 8772 4388 8778 4452
rect 16205 4450 16271 4453
rect 26509 4450 26575 4453
rect 16205 4448 26575 4450
rect 16205 4392 16210 4448
rect 16266 4392 26514 4448
rect 26570 4392 26575 4448
rect 16205 4390 26575 4392
rect 16205 4387 16271 4390
rect 26509 4387 26575 4390
rect 27061 4450 27127 4453
rect 28020 4450 28420 4480
rect 27061 4448 28420 4450
rect 27061 4392 27066 4448
rect 27122 4392 28420 4448
rect 27061 4390 28420 4392
rect 27061 4387 27127 4390
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 28020 4360 28420 4390
rect 4870 4319 5186 4320
rect 5441 4314 5507 4317
rect 5398 4312 5507 4314
rect 5398 4256 5446 4312
rect 5502 4256 5507 4312
rect 5398 4251 5507 4256
rect 8385 4314 8451 4317
rect 9673 4314 9739 4317
rect 13721 4314 13787 4317
rect 17769 4314 17835 4317
rect 8385 4312 17835 4314
rect 8385 4256 8390 4312
rect 8446 4256 9678 4312
rect 9734 4256 13726 4312
rect 13782 4256 17774 4312
rect 17830 4256 17835 4312
rect 8385 4254 17835 4256
rect 8385 4251 8451 4254
rect 9673 4251 9739 4254
rect 13721 4251 13787 4254
rect 17769 4251 17835 4254
rect 17953 4314 18019 4317
rect 18873 4314 18939 4317
rect 17953 4312 18939 4314
rect 17953 4256 17958 4312
rect 18014 4256 18878 4312
rect 18934 4256 18939 4312
rect 17953 4254 18939 4256
rect 17953 4251 18019 4254
rect 18873 4251 18939 4254
rect 20253 4314 20319 4317
rect 21173 4314 21239 4317
rect 20253 4312 21239 4314
rect 20253 4256 20258 4312
rect 20314 4256 21178 4312
rect 21234 4256 21239 4312
rect 20253 4254 21239 4256
rect 20253 4251 20319 4254
rect 21173 4251 21239 4254
rect 560 4178 960 4208
rect 1853 4178 1919 4181
rect 560 4176 1919 4178
rect 560 4120 1858 4176
rect 1914 4120 1919 4176
rect 560 4118 1919 4120
rect 560 4088 960 4118
rect 1853 4115 1919 4118
rect 5073 4178 5139 4181
rect 5398 4178 5458 4251
rect 16481 4178 16547 4181
rect 5073 4176 5458 4178
rect 5073 4120 5078 4176
rect 5134 4120 5458 4176
rect 5073 4118 5458 4120
rect 6870 4176 16547 4178
rect 6870 4120 16486 4176
rect 16542 4120 16547 4176
rect 6870 4118 16547 4120
rect 5073 4115 5139 4118
rect 1669 4042 1735 4045
rect 6870 4042 6930 4118
rect 16481 4115 16547 4118
rect 16941 4178 17007 4181
rect 20253 4178 20319 4181
rect 24025 4178 24091 4181
rect 24669 4178 24735 4181
rect 24853 4178 24919 4181
rect 16941 4176 24919 4178
rect 16941 4120 16946 4176
rect 17002 4120 20258 4176
rect 20314 4120 24030 4176
rect 24086 4120 24674 4176
rect 24730 4120 24858 4176
rect 24914 4120 24919 4176
rect 16941 4118 24919 4120
rect 16941 4115 17007 4118
rect 20253 4115 20319 4118
rect 24025 4115 24091 4118
rect 24669 4115 24735 4118
rect 24853 4115 24919 4118
rect 27429 4178 27495 4181
rect 28020 4178 28420 4208
rect 27429 4176 28420 4178
rect 27429 4120 27434 4176
rect 27490 4120 28420 4176
rect 27429 4118 28420 4120
rect 27429 4115 27495 4118
rect 28020 4088 28420 4118
rect 1669 4040 6930 4042
rect 1669 3984 1674 4040
rect 1730 3984 6930 4040
rect 1669 3982 6930 3984
rect 7373 4042 7439 4045
rect 8845 4042 8911 4045
rect 7373 4040 8911 4042
rect 7373 3984 7378 4040
rect 7434 3984 8850 4040
rect 8906 3984 8911 4040
rect 7373 3982 8911 3984
rect 1669 3979 1735 3982
rect 7373 3979 7439 3982
rect 8845 3979 8911 3982
rect 9673 4042 9739 4045
rect 10317 4042 10383 4045
rect 20529 4042 20595 4045
rect 9673 4040 20595 4042
rect 9673 3984 9678 4040
rect 9734 3984 10322 4040
rect 10378 3984 20534 4040
rect 20590 3984 20595 4040
rect 9673 3982 20595 3984
rect 9673 3979 9739 3982
rect 10317 3979 10383 3982
rect 20529 3979 20595 3982
rect 20897 4042 20963 4045
rect 24025 4042 24091 4045
rect 20897 4040 24091 4042
rect 20897 3984 20902 4040
rect 20958 3984 24030 4040
rect 24086 3984 24091 4040
rect 20897 3982 24091 3984
rect 20897 3979 20963 3982
rect 24025 3979 24091 3982
rect 560 3906 960 3936
rect 1301 3906 1367 3909
rect 560 3904 1367 3906
rect 560 3848 1306 3904
rect 1362 3848 1367 3904
rect 560 3846 1367 3848
rect 560 3816 960 3846
rect 1301 3843 1367 3846
rect 5165 3906 5231 3909
rect 6361 3906 6427 3909
rect 7189 3906 7255 3909
rect 8385 3906 8451 3909
rect 5165 3904 8451 3906
rect 5165 3848 5170 3904
rect 5226 3848 6366 3904
rect 6422 3848 7194 3904
rect 7250 3848 8390 3904
rect 8446 3848 8451 3904
rect 5165 3846 8451 3848
rect 5165 3843 5231 3846
rect 6361 3843 6427 3846
rect 7189 3843 7255 3846
rect 8385 3843 8451 3846
rect 9213 3906 9279 3909
rect 11789 3906 11855 3909
rect 14917 3906 14983 3909
rect 9213 3904 14983 3906
rect 9213 3848 9218 3904
rect 9274 3848 11794 3904
rect 11850 3848 14922 3904
rect 14978 3848 14983 3904
rect 9213 3846 14983 3848
rect 9213 3843 9279 3846
rect 11789 3843 11855 3846
rect 14917 3843 14983 3846
rect 15745 3906 15811 3909
rect 26509 3906 26575 3909
rect 15745 3904 26575 3906
rect 15745 3848 15750 3904
rect 15806 3848 26514 3904
rect 26570 3848 26575 3904
rect 15745 3846 26575 3848
rect 15745 3843 15811 3846
rect 26509 3843 26575 3846
rect 27429 3906 27495 3909
rect 28020 3906 28420 3936
rect 27429 3904 28420 3906
rect 27429 3848 27434 3904
rect 27490 3848 28420 3904
rect 27429 3846 28420 3848
rect 27429 3843 27495 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 28020 3816 28420 3846
rect 4210 3775 4526 3776
rect 3233 3770 3299 3773
rect 3601 3770 3667 3773
rect 3233 3768 3667 3770
rect 3233 3712 3238 3768
rect 3294 3712 3606 3768
rect 3662 3712 3667 3768
rect 3233 3710 3667 3712
rect 3233 3707 3299 3710
rect 3601 3707 3667 3710
rect 4797 3770 4863 3773
rect 7281 3770 7347 3773
rect 4797 3768 7347 3770
rect 4797 3712 4802 3768
rect 4858 3712 7286 3768
rect 7342 3712 7347 3768
rect 4797 3710 7347 3712
rect 4797 3707 4863 3710
rect 7281 3707 7347 3710
rect 8385 3770 8451 3773
rect 9857 3770 9923 3773
rect 10225 3770 10291 3773
rect 8385 3768 10291 3770
rect 8385 3712 8390 3768
rect 8446 3712 9862 3768
rect 9918 3712 10230 3768
rect 10286 3712 10291 3768
rect 8385 3710 10291 3712
rect 8385 3707 8451 3710
rect 9857 3707 9923 3710
rect 10225 3707 10291 3710
rect 17401 3770 17467 3773
rect 18413 3770 18479 3773
rect 17401 3768 18479 3770
rect 17401 3712 17406 3768
rect 17462 3712 18418 3768
rect 18474 3712 18479 3768
rect 17401 3710 18479 3712
rect 17401 3707 17467 3710
rect 18413 3707 18479 3710
rect 18597 3770 18663 3773
rect 24853 3770 24919 3773
rect 18597 3768 24919 3770
rect 18597 3712 18602 3768
rect 18658 3712 24858 3768
rect 24914 3712 24919 3768
rect 18597 3710 24919 3712
rect 18597 3707 18663 3710
rect 24853 3707 24919 3710
rect 560 3634 960 3664
rect 1209 3634 1275 3637
rect 560 3632 1275 3634
rect 560 3576 1214 3632
rect 1270 3576 1275 3632
rect 560 3574 1275 3576
rect 560 3544 960 3574
rect 1209 3571 1275 3574
rect 4654 3572 4660 3636
rect 4724 3634 4730 3636
rect 5349 3634 5415 3637
rect 4724 3632 5415 3634
rect 4724 3576 5354 3632
rect 5410 3576 5415 3632
rect 4724 3574 5415 3576
rect 4724 3572 4730 3574
rect 5349 3571 5415 3574
rect 7557 3634 7623 3637
rect 18873 3634 18939 3637
rect 7557 3632 18939 3634
rect 7557 3576 7562 3632
rect 7618 3576 18878 3632
rect 18934 3576 18939 3632
rect 7557 3574 18939 3576
rect 7557 3571 7623 3574
rect 18873 3571 18939 3574
rect 26693 3634 26759 3637
rect 28020 3634 28420 3664
rect 26693 3632 28420 3634
rect 26693 3576 26698 3632
rect 26754 3576 28420 3632
rect 26693 3574 28420 3576
rect 26693 3571 26759 3574
rect 28020 3544 28420 3574
rect 4245 3498 4311 3501
rect 5073 3498 5139 3501
rect 4245 3496 5139 3498
rect 4245 3440 4250 3496
rect 4306 3440 5078 3496
rect 5134 3440 5139 3496
rect 4245 3438 5139 3440
rect 4245 3435 4311 3438
rect 5073 3435 5139 3438
rect 5441 3498 5507 3501
rect 8109 3498 8175 3501
rect 5441 3496 8175 3498
rect 5441 3440 5446 3496
rect 5502 3440 8114 3496
rect 8170 3440 8175 3496
rect 5441 3438 8175 3440
rect 5441 3435 5507 3438
rect 8109 3435 8175 3438
rect 8702 3436 8708 3500
rect 8772 3498 8778 3500
rect 8845 3498 8911 3501
rect 8772 3496 8911 3498
rect 8772 3440 8850 3496
rect 8906 3440 8911 3496
rect 8772 3438 8911 3440
rect 8772 3436 8778 3438
rect 8845 3435 8911 3438
rect 12709 3498 12775 3501
rect 13261 3498 13327 3501
rect 12709 3496 13327 3498
rect 12709 3440 12714 3496
rect 12770 3440 13266 3496
rect 13322 3440 13327 3496
rect 12709 3438 13327 3440
rect 12709 3435 12775 3438
rect 13261 3435 13327 3438
rect 14641 3498 14707 3501
rect 26877 3498 26943 3501
rect 14641 3496 26943 3498
rect 14641 3440 14646 3496
rect 14702 3440 26882 3496
rect 26938 3440 26943 3496
rect 14641 3438 26943 3440
rect 14641 3435 14707 3438
rect 26877 3435 26943 3438
rect 560 3362 960 3392
rect 1301 3362 1367 3365
rect 560 3360 1367 3362
rect 560 3304 1306 3360
rect 1362 3304 1367 3360
rect 560 3302 1367 3304
rect 560 3272 960 3302
rect 1301 3299 1367 3302
rect 5717 3362 5783 3365
rect 12985 3362 13051 3365
rect 19609 3362 19675 3365
rect 5717 3360 10058 3362
rect 5717 3304 5722 3360
rect 5778 3304 10058 3360
rect 5717 3302 10058 3304
rect 5717 3299 5783 3302
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 5993 3226 6059 3229
rect 6453 3226 6519 3229
rect 7649 3226 7715 3229
rect 9305 3226 9371 3229
rect 5993 3224 9371 3226
rect 5993 3168 5998 3224
rect 6054 3168 6458 3224
rect 6514 3168 7654 3224
rect 7710 3168 9310 3224
rect 9366 3168 9371 3224
rect 5993 3166 9371 3168
rect 9998 3226 10058 3302
rect 12985 3360 19675 3362
rect 12985 3304 12990 3360
rect 13046 3304 19614 3360
rect 19670 3304 19675 3360
rect 12985 3302 19675 3304
rect 12985 3299 13051 3302
rect 19609 3299 19675 3302
rect 24853 3362 24919 3365
rect 26325 3362 26391 3365
rect 24853 3360 26391 3362
rect 24853 3304 24858 3360
rect 24914 3304 26330 3360
rect 26386 3304 26391 3360
rect 24853 3302 26391 3304
rect 24853 3299 24919 3302
rect 26325 3299 26391 3302
rect 27061 3362 27127 3365
rect 28020 3362 28420 3392
rect 27061 3360 28420 3362
rect 27061 3304 27066 3360
rect 27122 3304 28420 3360
rect 27061 3302 28420 3304
rect 27061 3299 27127 3302
rect 28020 3272 28420 3302
rect 10869 3226 10935 3229
rect 12709 3226 12775 3229
rect 9998 3224 12775 3226
rect 9998 3168 10874 3224
rect 10930 3168 12714 3224
rect 12770 3168 12775 3224
rect 9998 3166 12775 3168
rect 5993 3163 6059 3166
rect 6453 3163 6519 3166
rect 7649 3163 7715 3166
rect 9305 3163 9371 3166
rect 10869 3163 10935 3166
rect 12709 3163 12775 3166
rect 14917 3226 14983 3229
rect 19149 3226 19215 3229
rect 14917 3224 19215 3226
rect 14917 3168 14922 3224
rect 14978 3168 19154 3224
rect 19210 3168 19215 3224
rect 14917 3166 19215 3168
rect 14917 3163 14983 3166
rect 19149 3163 19215 3166
rect 19333 3228 19399 3229
rect 19333 3224 19380 3228
rect 19444 3226 19450 3228
rect 20437 3226 20503 3229
rect 23933 3226 23999 3229
rect 19333 3168 19338 3224
rect 19333 3164 19380 3168
rect 19444 3166 19490 3226
rect 20437 3224 23999 3226
rect 20437 3168 20442 3224
rect 20498 3168 23938 3224
rect 23994 3168 23999 3224
rect 20437 3166 23999 3168
rect 19444 3164 19450 3166
rect 19333 3163 19399 3164
rect 20437 3163 20503 3166
rect 23933 3163 23999 3166
rect 24117 3226 24183 3229
rect 26969 3226 27035 3229
rect 24117 3224 27035 3226
rect 24117 3168 24122 3224
rect 24178 3168 26974 3224
rect 27030 3168 27035 3224
rect 24117 3166 27035 3168
rect 24117 3163 24183 3166
rect 26969 3163 27035 3166
rect 560 3090 960 3120
rect 1485 3090 1551 3093
rect 560 3088 1551 3090
rect 560 3032 1490 3088
rect 1546 3032 1551 3088
rect 560 3030 1551 3032
rect 560 3000 960 3030
rect 1485 3027 1551 3030
rect 1945 3090 2011 3093
rect 12341 3090 12407 3093
rect 1945 3088 12407 3090
rect 1945 3032 1950 3088
rect 2006 3032 12346 3088
rect 12402 3032 12407 3088
rect 1945 3030 12407 3032
rect 1945 3027 2011 3030
rect 12341 3027 12407 3030
rect 14825 3090 14891 3093
rect 27245 3090 27311 3093
rect 14825 3088 27311 3090
rect 14825 3032 14830 3088
rect 14886 3032 27250 3088
rect 27306 3032 27311 3088
rect 14825 3030 27311 3032
rect 14825 3027 14891 3030
rect 27245 3027 27311 3030
rect 27429 3090 27495 3093
rect 28020 3090 28420 3120
rect 27429 3088 28420 3090
rect 27429 3032 27434 3088
rect 27490 3032 28420 3088
rect 27429 3030 28420 3032
rect 27429 3027 27495 3030
rect 28020 3000 28420 3030
rect 4245 2954 4311 2957
rect 4889 2954 4955 2957
rect 10409 2954 10475 2957
rect 11881 2954 11947 2957
rect 21449 2954 21515 2957
rect 25221 2954 25287 2957
rect 4245 2952 25287 2954
rect 4245 2896 4250 2952
rect 4306 2896 4894 2952
rect 4950 2896 10414 2952
rect 10470 2896 11886 2952
rect 11942 2896 21454 2952
rect 21510 2896 25226 2952
rect 25282 2896 25287 2952
rect 4245 2894 25287 2896
rect 4245 2891 4311 2894
rect 4889 2891 4955 2894
rect 10409 2891 10475 2894
rect 11881 2891 11947 2894
rect 21449 2891 21515 2894
rect 25221 2891 25287 2894
rect 560 2818 960 2848
rect 1853 2818 1919 2821
rect 560 2816 1919 2818
rect 560 2760 1858 2816
rect 1914 2760 1919 2816
rect 560 2758 1919 2760
rect 560 2728 960 2758
rect 1853 2755 1919 2758
rect 4981 2818 5047 2821
rect 13261 2818 13327 2821
rect 19149 2818 19215 2821
rect 4981 2816 19215 2818
rect 4981 2760 4986 2816
rect 5042 2760 13266 2816
rect 13322 2760 19154 2816
rect 19210 2760 19215 2816
rect 4981 2758 19215 2760
rect 4981 2755 5047 2758
rect 13261 2755 13327 2758
rect 19149 2755 19215 2758
rect 20805 2818 20871 2821
rect 22921 2818 22987 2821
rect 20805 2816 22987 2818
rect 20805 2760 20810 2816
rect 20866 2760 22926 2816
rect 22982 2760 22987 2816
rect 20805 2758 22987 2760
rect 20805 2755 20871 2758
rect 22921 2755 22987 2758
rect 25957 2818 26023 2821
rect 26693 2818 26759 2821
rect 28020 2818 28420 2848
rect 25957 2816 26066 2818
rect 25957 2760 25962 2816
rect 26018 2760 26066 2816
rect 25957 2755 26066 2760
rect 26693 2816 28420 2818
rect 26693 2760 26698 2816
rect 26754 2760 28420 2816
rect 26693 2758 28420 2760
rect 26693 2755 26759 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 21909 2682 21975 2685
rect 7606 2680 21975 2682
rect 7606 2624 21914 2680
rect 21970 2624 21975 2680
rect 7606 2622 21975 2624
rect 560 2546 960 2576
rect 1025 2546 1091 2549
rect 560 2544 1091 2546
rect 560 2488 1030 2544
rect 1086 2488 1091 2544
rect 560 2486 1091 2488
rect 560 2456 960 2486
rect 1025 2483 1091 2486
rect 2313 2546 2379 2549
rect 7606 2546 7666 2622
rect 21909 2619 21975 2622
rect 22553 2682 22619 2685
rect 24945 2682 25011 2685
rect 22553 2680 25011 2682
rect 22553 2624 22558 2680
rect 22614 2624 24950 2680
rect 25006 2624 25011 2680
rect 22553 2622 25011 2624
rect 22553 2619 22619 2622
rect 24945 2619 25011 2622
rect 24669 2546 24735 2549
rect 2313 2544 7666 2546
rect 2313 2488 2318 2544
rect 2374 2488 7666 2544
rect 2313 2486 7666 2488
rect 8526 2544 24735 2546
rect 8526 2488 24674 2544
rect 24730 2488 24735 2544
rect 8526 2486 24735 2488
rect 2313 2483 2379 2486
rect 5073 2410 5139 2413
rect 8526 2410 8586 2486
rect 24669 2483 24735 2486
rect 5073 2408 8586 2410
rect 5073 2352 5078 2408
rect 5134 2352 8586 2408
rect 5073 2350 8586 2352
rect 8661 2410 8727 2413
rect 25773 2410 25839 2413
rect 8661 2408 25839 2410
rect 8661 2352 8666 2408
rect 8722 2352 25778 2408
rect 25834 2352 25839 2408
rect 8661 2350 25839 2352
rect 5073 2347 5139 2350
rect 8661 2347 8727 2350
rect 25773 2347 25839 2350
rect 560 2274 960 2304
rect 1301 2274 1367 2277
rect 560 2272 1367 2274
rect 560 2216 1306 2272
rect 1362 2216 1367 2272
rect 560 2214 1367 2216
rect 560 2184 960 2214
rect 1301 2211 1367 2214
rect 9213 2274 9279 2277
rect 10041 2274 10107 2277
rect 23933 2274 23999 2277
rect 9213 2272 10107 2274
rect 9213 2216 9218 2272
rect 9274 2216 10046 2272
rect 10102 2216 10107 2272
rect 9213 2214 10107 2216
rect 9213 2211 9279 2214
rect 10041 2211 10107 2214
rect 17174 2272 23999 2274
rect 17174 2216 23938 2272
rect 23994 2216 23999 2272
rect 17174 2214 23999 2216
rect 26006 2274 26066 2755
rect 28020 2728 28420 2758
rect 26141 2546 26207 2549
rect 28020 2546 28420 2576
rect 26141 2544 28420 2546
rect 26141 2488 26146 2544
rect 26202 2488 28420 2544
rect 26141 2486 28420 2488
rect 26141 2483 26207 2486
rect 28020 2456 28420 2486
rect 28020 2274 28420 2304
rect 26006 2214 28420 2274
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 8201 2138 8267 2141
rect 17174 2138 17234 2214
rect 23933 2211 23999 2214
rect 28020 2184 28420 2214
rect 8201 2136 17234 2138
rect 8201 2080 8206 2136
rect 8262 2080 17234 2136
rect 8201 2078 17234 2080
rect 8201 2075 8267 2078
rect 560 2002 960 2032
rect 3969 2002 4035 2005
rect 560 2000 4035 2002
rect 560 1944 3974 2000
rect 4030 1944 4035 2000
rect 560 1942 4035 1944
rect 560 1912 960 1942
rect 3969 1939 4035 1942
rect 8109 2002 8175 2005
rect 25589 2002 25655 2005
rect 8109 2000 25655 2002
rect 8109 1944 8114 2000
rect 8170 1944 25594 2000
rect 25650 1944 25655 2000
rect 8109 1942 25655 1944
rect 8109 1939 8175 1942
rect 25589 1939 25655 1942
rect 25957 2002 26023 2005
rect 28020 2002 28420 2032
rect 25957 2000 28420 2002
rect 25957 1944 25962 2000
rect 26018 1944 28420 2000
rect 25957 1942 28420 1944
rect 25957 1939 26023 1942
rect 28020 1912 28420 1942
<< via3 >>
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 19380 5536 19444 5540
rect 19380 5480 19430 5536
rect 19430 5480 19444 5536
rect 19380 5476 19444 5480
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4660 5340 4724 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 8708 4388 8772 4452
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4660 3572 4724 3636
rect 8708 3436 8772 3500
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 19380 3224 19444 3228
rect 19380 3168 19394 3224
rect 19394 3168 19444 3224
rect 19380 3164 19444 3168
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 7104 4528 7664
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4868 7648 5188 7664
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 19379 5540 19445 5541
rect 19379 5476 19380 5540
rect 19444 5476 19445 5540
rect 19379 5475 19445 5476
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4659 5404 4725 5405
rect 4659 5340 4660 5404
rect 4724 5340 4725 5404
rect 4659 5339 4725 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4662 3637 4722 5339
rect 4868 4384 5188 5408
rect 8707 4452 8773 4453
rect 8707 4388 8708 4452
rect 8772 4388 8773 4452
rect 8707 4387 8773 4388
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4659 3636 4725 3637
rect 4659 3572 4660 3636
rect 4724 3572 4725 3636
rect 4659 3571 4725 3572
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 3296 5188 4320
rect 8710 3501 8770 4387
rect 8707 3500 8773 3501
rect 8707 3436 8708 3500
rect 8772 3436 8773 3500
rect 8707 3435 8773 3436
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 19382 3229 19442 5475
rect 19379 3228 19445 3229
rect 19379 3164 19380 3228
rect 19444 3164 19445 3228
rect 19379 3163 19445 3164
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1710522493
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1710522493
transform -1 0 23092 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1710522493
transform -1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1710522493
transform -1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1710522493
transform -1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1710522493
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1710522493
transform -1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1710522493
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1710522493
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1710522493
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1710522493
transform -1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1710522493
transform -1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1710522493
transform -1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1710522493
transform -1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1710522493
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1710522493
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__1
timestamp 1710522493
transform 1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 3772 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1710522493
transform -1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _177_
timestamp 1710522493
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1710522493
transform -1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1710522493
transform 1 0 8924 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1710522493
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1710522493
transform 1 0 10764 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1710522493
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1710522493
transform -1 0 11224 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1710522493
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 12972 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 25208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 17572 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1710522493
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7636 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _192_
timestamp 1710522493
transform -1 0 6440 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5152 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7728 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 6256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _196_
timestamp 1710522493
transform 1 0 7176 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _197_
timestamp 1710522493
transform 1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 8096 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _200_
timestamp 1710522493
transform 1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1710522493
transform 1 0 9384 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _202_
timestamp 1710522493
transform -1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _203_
timestamp 1710522493
transform 1 0 12604 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _204_
timestamp 1710522493
transform 1 0 13432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _205_
timestamp 1710522493
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _206_
timestamp 1710522493
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 16376 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _208_
timestamp 1710522493
transform 1 0 14904 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 15364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _210_
timestamp 1710522493
transform -1 0 15548 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _211_
timestamp 1710522493
transform -1 0 17848 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _212_
timestamp 1710522493
transform 1 0 17756 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _213_
timestamp 1710522493
transform -1 0 16560 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _214_
timestamp 1710522493
transform -1 0 19136 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _215_
timestamp 1710522493
transform 1 0 19228 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _216_
timestamp 1710522493
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _217_
timestamp 1710522493
transform 1 0 21252 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _218_
timestamp 1710522493
transform 1 0 19688 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _219_
timestamp 1710522493
transform -1 0 21620 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 7544 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 5152 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _223_
timestamp 1710522493
transform -1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp 1710522493
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _225_
timestamp 1710522493
transform -1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 1710522493
transform 1 0 4876 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 5428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1710522493
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 6900 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _231_
timestamp 1710522493
transform -1 0 9476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp 1710522493
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 1710522493
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _234_
timestamp 1710522493
transform 1 0 8740 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7820 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _236_
timestamp 1710522493
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1710522493
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 1710522493
transform -1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _239_
timestamp 1710522493
transform 1 0 9476 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _240_
timestamp 1710522493
transform -1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _241_
timestamp 1710522493
transform 1 0 10672 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1710522493
transform -1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1710522493
transform 1 0 12788 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _244_
timestamp 1710522493
transform -1 0 13156 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _245_
timestamp 1710522493
transform -1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1710522493
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _247_
timestamp 1710522493
transform 1 0 13892 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _248_
timestamp 1710522493
transform 1 0 13248 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 1710522493
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _250_
timestamp 1710522493
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _251_
timestamp 1710522493
transform 1 0 18124 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _252_
timestamp 1710522493
transform -1 0 15732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1710522493
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1710522493
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _255_
timestamp 1710522493
transform 1 0 18400 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _256_
timestamp 1710522493
transform 1 0 17296 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 1710522493
transform -1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1710522493
transform -1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _259_
timestamp 1710522493
transform 1 0 20332 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _260_
timestamp 1710522493
transform 1 0 17940 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp 1710522493
transform -1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1710522493
transform -1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 4416 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 6072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _267_
timestamp 1710522493
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _268_
timestamp 1710522493
transform 1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _269_
timestamp 1710522493
transform -1 0 6900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1710522493
transform -1 0 8740 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _271_
timestamp 1710522493
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1710522493
transform -1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _273_
timestamp 1710522493
transform 1 0 9936 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1710522493
transform -1 0 13248 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _275_
timestamp 1710522493
transform -1 0 12788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1710522493
transform 1 0 6072 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _277_
timestamp 1710522493
transform 1 0 6256 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 1710522493
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 16652 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1710522493
transform 1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1710522493
transform -1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1710522493
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _283_
timestamp 1710522493
transform -1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _284_
timestamp 1710522493
transform -1 0 10580 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _286_
timestamp 1710522493
transform -1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1710522493
transform 1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 1710522493
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _289_
timestamp 1710522493
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _290_
timestamp 1710522493
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _291_
timestamp 1710522493
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _292_
timestamp 1710522493
transform -1 0 14996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _293_
timestamp 1710522493
transform -1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _294_
timestamp 1710522493
transform 1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 1710522493
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _296_
timestamp 1710522493
transform -1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp 1710522493
transform -1 0 24012 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1710522493
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _299_
timestamp 1710522493
transform -1 0 24380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1710522493
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _301_
timestamp 1710522493
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 17940 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _303_
timestamp 1710522493
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 20424 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 13064 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _306_
timestamp 1710522493
transform 1 0 12420 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _307_
timestamp 1710522493
transform 1 0 19228 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 23552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _309_
timestamp 1710522493
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 24564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _311_
timestamp 1710522493
transform 1 0 25576 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _312_
timestamp 1710522493
transform 1 0 23000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1710522493
transform -1 0 24656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 24196 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _315_
timestamp 1710522493
transform 1 0 26128 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 23000 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _317_
timestamp 1710522493
transform -1 0 25576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _318_
timestamp 1710522493
transform -1 0 22448 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _319_
timestamp 1710522493
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 20240 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _321_
timestamp 1710522493
transform -1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _322_
timestamp 1710522493
transform -1 0 23460 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _323_
timestamp 1710522493
transform -1 0 22816 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _324_
timestamp 1710522493
transform 1 0 20516 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _326_
timestamp 1710522493
transform 1 0 19228 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _327_
timestamp 1710522493
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 1710522493
transform 1 0 17848 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1710522493
transform 1 0 18308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 15732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 1710522493
transform 1 0 15272 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1710522493
transform -1 0 16192 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _334_
timestamp 1710522493
transform -1 0 9200 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _335_
timestamp 1710522493
transform 1 0 9200 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _336_
timestamp 1710522493
transform -1 0 9936 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1710522493
transform 1 0 9292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _338_
timestamp 1710522493
transform -1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _339_
timestamp 1710522493
transform 1 0 14260 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 1710522493
transform -1 0 14536 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1710522493
transform -1 0 14628 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _342_
timestamp 1710522493
transform -1 0 8372 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _343_
timestamp 1710522493
transform -1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _344_
timestamp 1710522493
transform 1 0 7176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _345_
timestamp 1710522493
transform -1 0 8372 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1710522493
transform 1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19872 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _348_
timestamp 1710522493
transform 1 0 22264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _349_
timestamp 1710522493
transform 1 0 3496 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1710522493
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1710522493
transform -1 0 24288 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _352_
timestamp 1710522493
transform 1 0 21068 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _353_
timestamp 1710522493
transform -1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _354_
timestamp 1710522493
transform -1 0 4876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _355_
timestamp 1710522493
transform -1 0 4416 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _356_
timestamp 1710522493
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _357_
timestamp 1710522493
transform 1 0 10028 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _358_
timestamp 1710522493
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _359_
timestamp 1710522493
transform 1 0 14076 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _360_
timestamp 1710522493
transform 1 0 15824 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _361_
timestamp 1710522493
transform 1 0 17848 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _362_
timestamp 1710522493
transform 1 0 22724 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 23920 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _364_
timestamp 1710522493
transform -1 0 12604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _365_
timestamp 1710522493
transform -1 0 12972 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _366_
timestamp 1710522493
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _367_
timestamp 1710522493
transform 1 0 10672 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1710522493
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _369_
timestamp 1710522493
transform 1 0 4048 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _370_
timestamp 1710522493
transform -1 0 3680 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _371_
timestamp 1710522493
transform 1 0 4600 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1710522493
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1710522493
transform 1 0 24932 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_1  _374_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 17296 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _376_
timestamp 1710522493
transform 1 0 12144 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1710522493
transform 1 0 12144 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _378_
timestamp 1710522493
transform 1 0 4876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _379_
timestamp 1710522493
transform 1 0 5244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _380_
timestamp 1710522493
transform 1 0 5428 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1710522493
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19872 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19780 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1710522493
transform 1 0 18032 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _385_
timestamp 1710522493
transform 1 0 16008 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _386_
timestamp 1710522493
transform 1 0 8924 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1710522493
transform -1 0 16008 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _388_
timestamp 1710522493
transform 1 0 6716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1710522493
transform 1 0 1840 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1710522493
transform 1 0 22356 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 20516 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _392_
timestamp 1710522493
transform 1 0 2116 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _393_
timestamp 1710522493
transform 1 0 2208 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _394_
timestamp 1710522493
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _395_
timestamp 1710522493
transform 1 0 10304 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _396_
timestamp 1710522493
transform 1 0 12144 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _397_
timestamp 1710522493
transform -1 0 16376 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _398_
timestamp 1710522493
transform 1 0 16652 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _399_
timestamp 1710522493
transform -1 0 21344 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1710522493
transform -1 0 23828 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1710522493
transform 1 0 22448 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1710522493
transform 1 0 24380 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1710522493
transform 1 0 23092 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp 1710522493
transform -1 0 26220 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _405_
timestamp 1710522493
transform -1 0 12052 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _406_
timestamp 1710522493
transform 1 0 2116 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp 1710522493
transform 1 0 24380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _408_
timestamp 1710522493
transform 1 0 11684 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _409_
timestamp 1710522493
transform 1 0 4140 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 14996 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1710522493
transform -1 0 6992 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1710522493
transform 1 0 10488 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1710522493
transform 1 0 19872 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1710522493
transform 1 0 19872 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 7912 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout89 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 1710522493
transform -1 0 24288 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 1710522493
transform -1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 1710522493
transform -1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout94
timestamp 1710522493
transform -1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 14076 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout96
timestamp 1710522493
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout97
timestamp 1710522493
transform 1 0 6440 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 1710522493
transform -1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 1710522493
transform -1 0 13984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 1710522493
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout101
timestamp 1710522493
transform -1 0 17940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp 1710522493
transform -1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout103
timestamp 1710522493
transform -1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout104
timestamp 1710522493
transform -1 0 26036 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout105
timestamp 1710522493
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout106
timestamp 1710522493
transform -1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 1710522493
transform -1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 1710522493
transform -1 0 22172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 1710522493
transform -1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 1710522493
transform 1 0 9016 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 1710522493
transform -1 0 10580 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 1710522493
transform -1 0 22356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 1710522493
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1710522493
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1710522493
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_90
timestamp 1710522493
transform 1 0 9384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1710522493
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_117 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_155
timestamp 1710522493
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1710522493
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1710522493
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_175
timestamp 1710522493
transform 1 0 17204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_189
timestamp 1710522493
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1710522493
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_228
timestamp 1710522493
transform 1 0 22080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_257
timestamp 1710522493
transform 1 0 24748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_271
timestamp 1710522493
transform 1 0 26036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_281
timestamp 1710522493
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_48
timestamp 1710522493
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1710522493
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_198
timestamp 1710522493
transform 1 0 19320 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_210
timestamp 1710522493
transform 1 0 20424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_274
timestamp 1710522493
transform 1 0 26312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1710522493
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_58
timestamp 1710522493
transform 1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_63
timestamp 1710522493
transform 1 0 6900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1710522493
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_135
timestamp 1710522493
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_148
timestamp 1710522493
transform 1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_156
timestamp 1710522493
transform 1 0 15456 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_164
timestamp 1710522493
transform 1 0 16192 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_170 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_182
timestamp 1710522493
transform 1 0 17848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1710522493
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1710522493
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_35
timestamp 1710522493
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1710522493
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_86
timestamp 1710522493
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1710522493
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_130
timestamp 1710522493
transform 1 0 13064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_146
timestamp 1710522493
transform 1 0 14536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1710522493
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_176
timestamp 1710522493
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_180
timestamp 1710522493
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_188
timestamp 1710522493
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1710522493
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_242
timestamp 1710522493
transform 1 0 23368 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_252
timestamp 1710522493
transform 1 0 24288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_274
timestamp 1710522493
transform 1 0 26312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_7
timestamp 1710522493
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_70
timestamp 1710522493
transform 1 0 7544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1710522493
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1710522493
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1710522493
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_157
timestamp 1710522493
transform 1 0 15548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_169
timestamp 1710522493
transform 1 0 16652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_190
timestamp 1710522493
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1710522493
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_226
timestamp 1710522493
transform 1 0 21896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_276
timestamp 1710522493
transform 1 0 26496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_14
timestamp 1710522493
transform 1 0 2392 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_22
timestamp 1710522493
transform 1 0 3128 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_31
timestamp 1710522493
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_42
timestamp 1710522493
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_70
timestamp 1710522493
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_77
timestamp 1710522493
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_82
timestamp 1710522493
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_103
timestamp 1710522493
transform 1 0 10580 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_160
timestamp 1710522493
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_172
timestamp 1710522493
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1710522493
transform 1 0 19596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1710522493
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_256
timestamp 1710522493
transform 1 0 24656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_270 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 25944 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_281
timestamp 1710522493
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_11
timestamp 1710522493
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_19
timestamp 1710522493
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1710522493
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_96
timestamp 1710522493
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_119
timestamp 1710522493
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1710522493
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1710522493
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_151
timestamp 1710522493
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_167
timestamp 1710522493
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_273
timestamp 1710522493
transform 1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_34
timestamp 1710522493
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1710522493
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1710522493
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_79
timestamp 1710522493
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_84
timestamp 1710522493
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1710522493
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1710522493
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1710522493
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_132
timestamp 1710522493
transform 1 0 13248 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_137
timestamp 1710522493
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_154
timestamp 1710522493
transform 1 0 15272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1710522493
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_183
timestamp 1710522493
transform 1 0 17940 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_268
timestamp 1710522493
transform 1 0 25760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_281
timestamp 1710522493
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_15
timestamp 1710522493
transform 1 0 2484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1710522493
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1710522493
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_114
timestamp 1710522493
transform 1 0 11592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1710522493
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_207
timestamp 1710522493
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_220
timestamp 1710522493
transform 1 0 21344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_243
timestamp 1710522493
transform 1 0 23460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_250
timestamp 1710522493
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_20
timestamp 1710522493
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_24
timestamp 1710522493
transform 1 0 3312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_44
timestamp 1710522493
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_94
timestamp 1710522493
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_103
timestamp 1710522493
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1710522493
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1710522493
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_125
timestamp 1710522493
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_139
timestamp 1710522493
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_146
timestamp 1710522493
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1710522493
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1710522493
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1710522493
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_193
timestamp 1710522493
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_201
timestamp 1710522493
transform 1 0 19596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_237
timestamp 1710522493
transform 1 0 22908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_242
timestamp 1710522493
transform 1 0 23368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_253
timestamp 1710522493
transform 1 0 24380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_274
timestamp 1710522493
transform 1 0 26312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1710522493
transform 1 0 21988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1710522493
transform -1 0 25208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1710522493
transform -1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1710522493
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1710522493
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1710522493
transform 1 0 26036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1710522493
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1710522493
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1710522493
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1710522493
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1710522493
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1710522493
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1710522493
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1710522493
transform -1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1710522493
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1710522493
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1710522493
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1710522493
transform -1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1710522493
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1710522493
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1710522493
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1710522493
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1710522493
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1710522493
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1710522493
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1710522493
transform 1 0 13340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1710522493
transform 1 0 15732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  output27
timestamp 1710522493
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1710522493
transform 1 0 27048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1710522493
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1710522493
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1710522493
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1710522493
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1710522493
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1710522493
transform -1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1710522493
transform -1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1710522493
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1710522493
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1710522493
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1710522493
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1710522493
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1710522493
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1710522493
transform -1 0 19044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1710522493
transform -1 0 21712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1710522493
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1710522493
transform 1 0 27232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1710522493
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1710522493
transform 1 0 27232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1710522493
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1710522493
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1710522493
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1710522493
transform 1 0 27232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1710522493
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1710522493
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1710522493
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1710522493
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1710522493
transform -1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1710522493
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1710522493
transform -1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1710522493
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1710522493
transform -1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1710522493
transform -1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1710522493
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1710522493
transform -1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1710522493
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1710522493
transform -1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1710522493
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1710522493
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1710522493
transform 1 0 25760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1710522493
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1710522493
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1710522493
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1710522493
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1710522493
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1710522493
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1710522493
transform 1 0 27232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1710522493
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1710522493
transform -1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1710522493
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1710522493
transform -1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1710522493
transform -1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1710522493
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1710522493
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1710522493
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1710522493
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1710522493
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1710522493
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1710522493
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 1710522493
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1710522493
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 1710522493
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1710522493
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 1710522493
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1710522493
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 1710522493
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1710522493
transform -1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 1710522493
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1710522493
transform -1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 1710522493
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1710522493
transform -1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 1710522493
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1710522493
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 1710522493
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1710522493
transform -1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 1710522493
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1710522493
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 1710522493
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1710522493
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1710522493
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22
timestamp 1710522493
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1710522493
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp 1710522493
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 1710522493
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 1710522493
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp 1710522493
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp 1710522493
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 1710522493
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 1710522493
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_31
timestamp 1710522493
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_32
timestamp 1710522493
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_33
timestamp 1710522493
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_34
timestamp 1710522493
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_35
timestamp 1710522493
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1710522493
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1710522493
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1710522493
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1710522493
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1710522493
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_41
timestamp 1710522493
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 1710522493
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_43
timestamp 1710522493
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_44
timestamp 1710522493
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_45
timestamp 1710522493
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_46
timestamp 1710522493
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_47
timestamp 1710522493
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_48
timestamp 1710522493
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_49
timestamp 1710522493
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_50
timestamp 1710522493
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_51
timestamp 1710522493
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp 1710522493
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp 1710522493
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 1710522493
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 1710522493
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 1710522493
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1710522493
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_58
timestamp 1710522493
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_59
timestamp 1710522493
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_60
timestamp 1710522493
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_61
timestamp 1710522493
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1710522493
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1710522493
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_64
timestamp 1710522493
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 1710522493
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_66
timestamp 1710522493
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_67
timestamp 1710522493
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_68
timestamp 1710522493
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_69
timestamp 1710522493
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_70
timestamp 1710522493
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_71
timestamp 1710522493
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_72
timestamp 1710522493
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_73
timestamp 1710522493
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_74
timestamp 1710522493
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp 1710522493
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_76
timestamp 1710522493
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_77
timestamp 1710522493
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_78
timestamp 1710522493
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_79
timestamp 1710522493
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 4208 2128 4528 7664 0 FreeSans 1920 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4868 2128 5188 7664 0 FreeSans 1920 90 0 0 VSS
port 1 nsew ground bidirectional
rlabel metal1 14490 7072 14490 7072 0 VDD
rlabel metal1 14490 7616 14490 7616 0 VSS
rlabel metal1 24610 5746 24610 5746 0 _000_
rlabel metal1 20240 5338 20240 5338 0 _001_
rlabel metal1 20332 6970 20332 6970 0 _002_
rlabel metal2 18354 6630 18354 6630 0 _003_
rlabel metal1 16238 6426 16238 6426 0 _004_
rlabel metal2 9338 6698 9338 6698 0 _005_
rlabel metal2 14582 6698 14582 6698 0 _006_
rlabel metal1 7123 6970 7123 6970 0 _007_
rlabel metal1 2983 4794 2983 4794 0 _008_
rlabel metal1 22402 2924 22402 2924 0 _009_
rlabel metal1 20930 3162 20930 3162 0 _010_
rlabel metal1 2438 3128 2438 3128 0 _011_
rlabel metal1 3174 4046 3174 4046 0 _012_
rlabel metal1 2162 3400 2162 3400 0 _013_
rlabel metal2 10626 3298 10626 3298 0 _014_
rlabel metal1 12098 2924 12098 2924 0 _015_
rlabel metal1 14996 2618 14996 2618 0 _016_
rlabel metal1 16698 2618 16698 2618 0 _017_
rlabel metal1 18446 2312 18446 2312 0 _018_
rlabel metal2 23322 4403 23322 4403 0 _019_
rlabel metal1 23828 3366 23828 3366 0 _020_
rlabel metal1 11592 5066 11592 5066 0 _021_
rlabel metal2 3818 6052 3818 6052 0 _022_
rlabel metal2 24978 6562 24978 6562 0 _023_
rlabel metal1 12098 6426 12098 6426 0 _024_
rlabel metal1 4554 6426 4554 6426 0 _025_
rlabel metal1 22448 6290 22448 6290 0 _026_
rlabel metal2 7406 4692 7406 4692 0 _027_
rlabel metal2 22310 5542 22310 5542 0 _028_
rlabel metal1 16514 5678 16514 5678 0 _029_
rlabel metal2 14950 5627 14950 5627 0 _030_
rlabel via1 14674 5202 14674 5202 0 _031_
rlabel metal2 6210 4148 6210 4148 0 _032_
rlabel metal2 9430 5916 9430 5916 0 _033_
rlabel metal2 9614 4250 9614 4250 0 _034_
rlabel metal1 12742 5746 12742 5746 0 _035_
rlabel metal1 7590 4148 7590 4148 0 _036_
rlabel metal2 17250 6732 17250 6732 0 _037_
rlabel metal1 8096 2414 8096 2414 0 _038_
rlabel metal1 18124 4590 18124 4590 0 _039_
rlabel metal1 9430 2992 9430 2992 0 _040_
rlabel metal1 16054 4692 16054 4692 0 _041_
rlabel metal1 26266 3570 26266 3570 0 _042_
rlabel metal1 3726 7378 3726 7378 0 _044_
rlabel metal1 6026 7378 6026 7378 0 _045_
rlabel metal1 8602 7378 8602 7378 0 _046_
rlabel metal2 10810 7140 10810 7140 0 _047_
rlabel metal1 11224 6426 11224 6426 0 _048_
rlabel metal1 13570 4794 13570 4794 0 _049_
rlabel metal1 25806 3026 25806 3026 0 _050_
rlabel metal2 9246 4539 9246 4539 0 _051_
rlabel metal2 13754 4199 13754 4199 0 _052_
rlabel metal1 13478 4658 13478 4658 0 _053_
rlabel metal1 5888 3706 5888 3706 0 _054_
rlabel metal1 5887 4114 5887 4114 0 _055_
rlabel metal1 5934 3468 5934 3468 0 _056_
rlabel metal1 7314 3536 7314 3536 0 _057_
rlabel metal1 8372 5202 8372 5202 0 _058_
rlabel metal2 9614 3332 9614 3332 0 _059_
rlabel metal2 11178 4420 11178 4420 0 _060_
rlabel metal1 13294 4250 13294 4250 0 _061_
rlabel metal2 14306 3026 14306 3026 0 _062_
rlabel metal1 15364 3978 15364 3978 0 _063_
rlabel metal1 14996 3706 14996 3706 0 _064_
rlabel metal1 14766 5134 14766 5134 0 _065_
rlabel metal1 17986 4046 17986 4046 0 _066_
rlabel metal1 16008 5134 16008 5134 0 _067_
rlabel metal2 19458 4284 19458 4284 0 _068_
rlabel metal2 21482 3842 21482 3842 0 _069_
rlabel metal1 22034 5644 22034 5644 0 _070_
rlabel metal1 16284 4590 16284 4590 0 _071_
rlabel metal1 5060 4794 5060 4794 0 _072_
rlabel metal1 5106 4182 5106 4182 0 _073_
rlabel metal1 6899 4114 6899 4114 0 _074_
rlabel metal1 5658 3536 5658 3536 0 _075_
rlabel metal1 6762 5134 6762 5134 0 _076_
rlabel metal2 8786 6086 8786 6086 0 _077_
rlabel metal2 8786 3298 8786 3298 0 _078_
rlabel metal2 7866 3536 7866 3536 0 _079_
rlabel metal2 10074 4148 10074 4148 0 _080_
rlabel viali 10074 4114 10074 4114 0 _081_
rlabel metal2 10902 4284 10902 4284 0 _082_
rlabel metal1 12512 5746 12512 5746 0 _083_
rlabel metal1 12558 5236 12558 5236 0 _084_
rlabel metal2 13938 5253 13938 5253 0 _085_
rlabel metal1 13478 4182 13478 4182 0 _086_
rlabel metal1 17572 5882 17572 5882 0 _087_
rlabel metal2 15594 5372 15594 5372 0 _088_
rlabel metal1 17342 5236 17342 5236 0 _089_
rlabel metal1 17296 4590 17296 4590 0 _090_
rlabel metal2 18998 4335 18998 4335 0 _091_
rlabel metal1 16974 4556 16974 4556 0 _092_
rlabel metal1 6026 4080 6026 4080 0 _093_
rlabel metal1 7038 4080 7038 4080 0 _094_
rlabel metal1 6440 5202 6440 5202 0 _095_
rlabel metal2 8694 3332 8694 3332 0 _096_
rlabel metal1 9890 4114 9890 4114 0 _097_
rlabel metal2 12374 5916 12374 5916 0 _098_
rlabel metal2 6118 6324 6118 6324 0 _099_
rlabel metal1 16514 6154 16514 6154 0 _100_
rlabel metal1 17572 5202 17572 5202 0 _101_
rlabel via1 19178 4114 19178 4114 0 _102_
rlabel metal1 7130 2482 7130 2482 0 _103_
rlabel metal1 18906 5746 18906 5746 0 _104_
rlabel metal1 25852 3910 25852 3910 0 _105_
rlabel metal2 25530 6426 25530 6426 0 _106_
rlabel metal1 18906 3434 18906 3434 0 _107_
rlabel metal1 23690 2482 23690 2482 0 _108_
rlabel metal1 19642 2958 19642 2958 0 _109_
rlabel metal1 19366 3502 19366 3502 0 _110_
rlabel via2 19642 3349 19642 3349 0 _111_
rlabel metal1 20240 3638 20240 3638 0 _112_
rlabel metal1 24656 3026 24656 3026 0 _113_
rlabel metal2 26588 2516 26588 2516 0 _114_
rlabel metal2 21850 6987 21850 6987 0 _115_
rlabel metal1 20470 5236 20470 5236 0 _116_
rlabel via2 14122 6205 14122 6205 0 _117_
rlabel metal1 22540 5338 22540 5338 0 _118_
rlabel metal2 22586 6460 22586 6460 0 _119_
rlabel metal2 21206 6630 21206 6630 0 _120_
rlabel metal2 19550 5950 19550 5950 0 _121_
rlabel metal1 19780 5882 19780 5882 0 _122_
rlabel metal1 19136 6834 19136 6834 0 _123_
rlabel metal1 18768 6834 18768 6834 0 _124_
rlabel metal1 16264 5712 16264 5712 0 _125_
rlabel metal1 15686 5882 15686 5882 0 _126_
rlabel metal1 15732 6426 15732 6426 0 _127_
rlabel metal1 9339 5236 9339 5236 0 _128_
rlabel metal2 9890 5780 9890 5780 0 _129_
rlabel metal2 9522 6052 9522 6052 0 _130_
rlabel metal1 15295 5610 15295 5610 0 _131_
rlabel metal1 14168 5882 14168 5882 0 _132_
rlabel metal1 14168 6426 14168 6426 0 _133_
rlabel metal1 7682 5542 7682 5542 0 _134_
rlabel metal2 7682 5440 7682 5440 0 _135_
rlabel metal1 7498 5882 7498 5882 0 _136_
rlabel metal1 7820 6426 7820 6426 0 _137_
rlabel metal2 20838 2907 20838 2907 0 _138_
rlabel metal2 21114 2108 21114 2108 0 _139_
rlabel metal1 4048 4590 4048 4590 0 _140_
rlabel metal1 24058 4454 24058 4454 0 _141_
rlabel metal1 12006 4046 12006 4046 0 _142_
rlabel metal2 12006 4284 12006 4284 0 _143_
rlabel metal1 11822 4250 11822 4250 0 _144_
rlabel metal1 11546 5134 11546 5134 0 _145_
rlabel metal1 4600 4998 4600 4998 0 _146_
rlabel metal1 4830 5644 4830 5644 0 _147_
rlabel metal1 4554 5746 4554 5746 0 _148_
rlabel metal1 15318 4080 15318 4080 0 _149_
rlabel metal1 14582 4046 14582 4046 0 _150_
rlabel metal1 12604 6426 12604 6426 0 _151_
rlabel metal1 5520 3162 5520 3162 0 _152_
rlabel metal1 5612 5882 5612 5882 0 _153_
rlabel metal1 5382 6222 5382 6222 0 _154_
rlabel metal2 23414 6494 23414 6494 0 _155_
rlabel metal1 24058 4250 24058 4250 0 _156_
rlabel metal1 15088 5270 15088 5270 0 clk
rlabel metal1 6946 4624 6946 4624 0 clknet_0_clk
rlabel metal2 2162 6562 2162 6562 0 clknet_2_0__leaf_clk
rlabel metal1 11454 6766 11454 6766 0 clknet_2_1__leaf_clk
rlabel metal1 16514 3026 16514 3026 0 clknet_2_2__leaf_clk
rlabel metal1 21666 6188 21666 6188 0 clknet_2_3__leaf_clk
rlabel metal2 2990 1350 2990 1350 0 comp_p
rlabel metal1 23000 3502 23000 3502 0 counter\[0\]
rlabel metal2 22034 5542 22034 5542 0 counter\[10\]
rlabel metal1 25392 2414 25392 2414 0 counter\[11\]
rlabel metal1 5106 2482 5106 2482 0 counter\[1\]
rlabel metal2 12742 3417 12742 3417 0 counter\[2\]
rlabel metal2 12650 2686 12650 2686 0 counter\[3\]
rlabel metal1 4646 3536 4646 3536 0 counter\[4\]
rlabel metal2 9062 2924 9062 2924 0 counter\[5\]
rlabel metal1 13754 2516 13754 2516 0 counter\[6\]
rlabel metal1 12604 3502 12604 3502 0 counter\[7\]
rlabel metal1 17434 2380 17434 2380 0 counter\[8\]
rlabel metal1 16146 2482 16146 2482 0 counter\[9\]
rlabel metal1 26036 5202 26036 5202 0 counter_sample
rlabel metal2 2070 2676 2070 2676 0 en_comp
rlabel metal1 26818 6800 26818 6800 0 en_offset_cal
rlabel metal2 27830 1350 27830 1350 0 en_offset_cal_o
rlabel metal1 25622 2890 25622 2890 0 en_vcm_sw_o
rlabel metal1 4002 4454 4002 4454 0 net1
rlabel metal1 8786 2550 8786 2550 0 net10
rlabel metal1 15134 5202 15134 5202 0 net100
rlabel metal1 16330 4148 16330 4148 0 net101
rlabel metal1 19366 5746 19366 5746 0 net102
rlabel metal1 25852 6358 25852 6358 0 net103
rlabel metal2 20010 6579 20010 6579 0 net104
rlabel metal1 17756 7242 17756 7242 0 net105
rlabel metal1 18538 7310 18538 7310 0 net106
rlabel metal2 18262 4301 18262 4301 0 net107
rlabel metal2 26818 1972 26818 1972 0 net108
rlabel metal2 7038 7582 7038 7582 0 net109
rlabel metal1 9617 2414 9617 2414 0 net11
rlabel viali 9899 2482 9899 2482 0 net110
rlabel metal1 11921 3502 11921 3502 0 net111
rlabel metal1 21390 7310 21390 7310 0 net112
rlabel metal1 17671 6698 17671 6698 0 net113
rlabel metal1 24840 3026 24840 3026 0 net114
rlabel metal1 24150 5236 24150 5236 0 net115
rlabel metal1 22724 4114 22724 4114 0 net116
rlabel viali 23690 3500 23690 3500 0 net117
rlabel metal2 21114 3196 21114 3196 0 net118
rlabel metal1 12512 2618 12512 2618 0 net12
rlabel metal1 13662 2516 13662 2516 0 net13
rlabel metal1 15364 3570 15364 3570 0 net14
rlabel metal1 18216 2482 18216 2482 0 net15
rlabel metal2 18906 3196 18906 3196 0 net16
rlabel metal2 22034 2788 22034 2788 0 net17
rlabel metal1 18170 7242 18170 7242 0 net18
rlabel metal2 17986 7480 17986 7480 0 net19
rlabel metal1 25392 2550 25392 2550 0 net2
rlabel metal1 3772 3502 3772 3502 0 net20
rlabel metal2 4738 7310 4738 7310 0 net21
rlabel metal1 5704 7446 5704 7446 0 net22
rlabel metal1 8280 7446 8280 7446 0 net23
rlabel metal1 11408 7378 11408 7378 0 net24
rlabel metal1 12972 7446 12972 7446 0 net25
rlabel metal1 13754 5882 13754 5882 0 net26
rlabel metal2 2346 3859 2346 3859 0 net27
rlabel metal1 26588 2346 26588 2346 0 net28
rlabel metal1 25990 2992 25990 2992 0 net29
rlabel metal2 27002 4284 27002 4284 0 net3
rlabel metal2 26542 2822 26542 2822 0 net30
rlabel metal3 8556 2448 8556 2448 0 net31
rlabel metal2 8418 5729 8418 5729 0 net32
rlabel metal1 3404 4998 3404 4998 0 net33
rlabel metal1 23874 2380 23874 2380 0 net34
rlabel metal2 6118 2244 6118 2244 0 net35
rlabel metal1 7222 2380 7222 2380 0 net36
rlabel metal2 10074 2329 10074 2329 0 net37
rlabel metal1 11546 2380 11546 2380 0 net38
rlabel metal1 13110 2448 13110 2448 0 net39
rlabel metal1 19044 7242 19044 7242 0 net4
rlabel metal1 15042 2448 15042 2448 0 net40
rlabel metal1 16744 3366 16744 3366 0 net41
rlabel metal1 19044 2822 19044 2822 0 net42
rlabel metal1 21666 2448 21666 2448 0 net43
rlabel metal2 27370 6290 27370 6290 0 net44
rlabel metal2 15778 4811 15778 4811 0 net45
rlabel metal1 6624 3706 6624 3706 0 net46
rlabel metal1 8832 4998 8832 4998 0 net47
rlabel metal2 9890 3553 9890 3553 0 net48
rlabel metal1 11362 5270 11362 5270 0 net49
rlabel metal1 25760 6426 25760 6426 0 net5
rlabel metal2 27278 5797 27278 5797 0 net50
rlabel metal1 16652 4590 16652 4590 0 net51
rlabel metal1 19044 4454 19044 4454 0 net52
rlabel via2 21114 4709 21114 4709 0 net53
rlabel metal2 26542 7582 26542 7582 0 net54
rlabel metal1 2070 5168 2070 5168 0 net55
rlabel metal2 9982 6256 9982 6256 0 net56
rlabel metal2 2714 4862 2714 4862 0 net57
rlabel metal1 2484 5678 2484 5678 0 net58
rlabel via2 1702 5661 1702 5661 0 net59
rlabel metal2 23966 6970 23966 6970 0 net6
rlabel metal2 2070 6035 2070 6035 0 net60
rlabel via2 2438 6749 2438 6749 0 net61
rlabel metal1 1840 6290 1840 6290 0 net62
rlabel via2 2622 7395 2622 7395 0 net63
rlabel metal1 1886 6834 1886 6834 0 net64
rlabel metal2 2254 6001 2254 6001 0 net65
rlabel metal3 17204 2176 17204 2176 0 net66
rlabel via2 16238 4437 16238 4437 0 net67
rlabel metal3 16882 1972 16882 1972 0 net68
rlabel metal2 8694 2329 8694 2329 0 net69
rlabel metal1 5566 2584 5566 2584 0 net7
rlabel metal2 9982 2278 9982 2278 0 net70
rlabel metal2 14858 3757 14858 3757 0 net71
rlabel metal2 14674 3417 14674 3417 0 net72
rlabel via2 15778 3893 15778 3893 0 net73
rlabel metal1 27278 3570 27278 3570 0 net74
rlabel metal1 27278 4080 27278 4080 0 net75
rlabel metal1 22494 4760 22494 4760 0 net76
rlabel metal1 4784 4998 4784 4998 0 net77
rlabel metal2 1702 4641 1702 4641 0 net78
rlabel metal1 3036 2414 3036 2414 0 net79
rlabel metal1 22494 5134 22494 5134 0 net8
rlabel metal2 2438 2142 2438 2142 0 net80
rlabel metal2 2346 2244 2346 2244 0 net81
rlabel metal2 1702 2210 1702 2210 0 net82
rlabel via2 1978 3043 1978 3043 0 net83
rlabel metal2 1702 3519 1702 3519 0 net84
rlabel metal2 1794 4301 1794 4301 0 net85
rlabel metal2 2254 2754 2254 2754 0 net86
rlabel metal2 1978 4335 1978 4335 0 net87
rlabel metal2 14490 3332 14490 3332 0 net88
rlabel metal1 8648 5542 8648 5542 0 net89
rlabel metal1 6762 2618 6762 2618 0 net9
rlabel metal1 18078 2312 18078 2312 0 net90
rlabel metal1 19642 5678 19642 5678 0 net91
rlabel metal2 18262 2142 18262 2142 0 net92
rlabel metal1 4922 2380 4922 2380 0 net93
rlabel metal2 20562 4573 20562 4573 0 net94
rlabel metal1 14352 4590 14352 4590 0 net95
rlabel metal1 4554 4590 4554 4590 0 net96
rlabel metal2 5474 5440 5474 5440 0 net97
rlabel metal1 6210 5202 6210 5202 0 net98
rlabel metal1 14076 3366 14076 3366 0 net99
rlabel metal1 26818 2822 26818 2822 0 offset_cal_cycle
rlabel metal1 3864 5134 3864 5134 0 result\[0\]
rlabel via2 21022 6613 21022 6613 0 result\[10\]
rlabel metal2 21206 5015 21206 5015 0 result\[11\]
rlabel metal2 8142 3638 8142 3638 0 result\[1\]
rlabel metal1 9200 5882 9200 5882 0 result\[2\]
rlabel metal1 9522 6630 9522 6630 0 result\[3\]
rlabel metal1 10672 6426 10672 6426 0 result\[4\]
rlabel metal1 13386 5814 13386 5814 0 result\[5\]
rlabel metal1 6394 5610 6394 5610 0 result\[6\]
rlabel metal1 6578 5542 6578 5542 0 result\[7\]
rlabel metal1 9338 7310 9338 7310 0 result\[8\]
rlabel metal1 19596 6426 19596 6426 0 result\[9\]
rlabel metal1 18354 7378 18354 7378 0 rst_z
rlabel metal2 1150 1418 1150 1418 0 sample_o
rlabel metal1 25760 7378 25760 7378 0 single_ended
rlabel via2 14766 6307 14766 6307 0 single_ended_reg
rlabel metal1 24242 7412 24242 7412 0 start
rlabel metal1 25070 6086 25070 6086 0 state\[0\]
rlabel metal1 23782 5236 23782 5236 0 state\[1\]
rlabel metal2 3910 1316 3910 1316 0 vcm_o[0]
rlabel metal2 7590 1316 7590 1316 0 vcm_o[2]
rlabel metal2 9430 1316 9430 1316 0 vcm_o[3]
rlabel metal2 11270 1316 11270 1316 0 vcm_o[4]
rlabel metal2 13110 1316 13110 1316 0 vcm_o[5]
rlabel metal2 14950 1316 14950 1316 0 vcm_o[6]
rlabel metal2 16790 1316 16790 1316 0 vcm_o[7]
rlabel metal2 18630 1316 18630 1316 0 vcm_o[8]
rlabel metal2 20470 1486 20470 1486 0 vcm_o[9]
rlabel metal1 23230 3400 23230 3400 0 vcm_o_i[10]
rlabel metal2 6670 1384 6670 1384 0 vcm_o_i[1]
rlabel metal1 8832 3570 8832 3570 0 vcm_o_i[2]
rlabel metal2 10350 1384 10350 1384 0 vcm_o_i[3]
rlabel metal2 12190 1384 12190 1384 0 vcm_o_i[4]
rlabel metal2 14030 1350 14030 1350 0 vcm_o_i[5]
rlabel metal2 15870 1384 15870 1384 0 vcm_o_i[6]
rlabel metal1 17940 2958 17940 2958 0 vcm_o_i[7]
rlabel metal1 19642 3026 19642 3026 0 vcm_o_i[8]
rlabel metal2 21390 1350 21390 1350 0 vcm_o_i[9]
rlabel metal3 774 7956 774 7956 0 vin_p_sw_on
rlabel metal2 27462 4879 27462 4879 0 vref_z_n_o[0]
rlabel metal2 27462 7599 27462 7599 0 vref_z_n_o[10]
rlabel metal3 27746 5236 27746 5236 0 vref_z_n_o[1]
rlabel metal2 27462 5423 27462 5423 0 vref_z_n_o[2]
rlabel metal3 27746 6052 27746 6052 0 vref_z_n_o[4]
rlabel metal2 27462 6103 27462 6103 0 vref_z_n_o[5]
rlabel metal2 27462 6511 27462 6511 0 vref_z_n_o[6]
rlabel metal1 27508 6630 27508 6630 0 vref_z_n_o[8]
rlabel metal3 27746 7412 27746 7412 0 vref_z_n_o[9]
rlabel metal3 636 4964 636 4964 0 vref_z_p_o[0]
rlabel metal1 1610 7514 1610 7514 0 vref_z_p_o[10]
rlabel metal3 1096 5508 1096 5508 0 vref_z_p_o[2]
rlabel metal3 636 6052 636 6052 0 vref_z_p_o[4]
rlabel metal1 1748 6630 1748 6630 0 vref_z_p_o[5]
rlabel metal1 1426 6426 1426 6426 0 vref_z_p_o[6]
rlabel metal3 1372 6868 1372 6868 0 vref_z_p_o[7]
rlabel metal2 1518 7055 1518 7055 0 vref_z_p_o[8]
rlabel metal2 1886 7191 1886 7191 0 vref_z_p_o[9]
rlabel metal3 27378 1972 27378 1972 0 vss_n_o[0]
rlabel metal3 27746 4692 27746 4692 0 vss_n_o[10]
rlabel metal3 27401 2244 27401 2244 0 vss_n_o[1]
rlabel metal3 27470 2516 27470 2516 0 vss_n_o[2]
rlabel metal3 27746 2788 27746 2788 0 vss_n_o[3]
rlabel metal3 27746 3604 27746 3604 0 vss_n_o[6]
rlabel metal2 27462 3791 27462 3791 0 vss_n_o[7]
rlabel metal2 4002 2125 4002 2125 0 vss_p_o[0]
rlabel metal3 820 2244 820 2244 0 vss_p_o[1]
rlabel metal3 682 2516 682 2516 0 vss_p_o[2]
rlabel metal2 1886 2703 1886 2703 0 vss_p_o[3]
rlabel metal2 1518 2839 1518 2839 0 vss_p_o[4]
rlabel metal1 1610 3162 1610 3162 0 vss_p_o[5]
rlabel metal1 1380 2890 1380 2890 0 vss_p_o[6]
rlabel metal1 1426 3706 1426 3706 0 vss_p_o[7]
rlabel metal3 1096 4148 1096 4148 0 vss_p_o[8]
rlabel metal2 1518 4199 1518 4199 0 vss_p_o[9]
flabel metal3 s 560 7896 960 8016 0 FreeSans 480 0 0 0 vin_p_sw_on
port 45 nsew signal input
flabel metal3 s 560 4904 960 5024 0 FreeSans 480 0 0 0 vref_z_p_o[0]
port 57 nsew signal output
flabel metal3 s 560 7624 960 7744 0 FreeSans 480 0 0 0 vref_z_p_o[10]
port 58 nsew signal output
flabel metal3 s 560 5176 960 5296 0 FreeSans 480 0 0 0 vref_z_p_o[1]
port 59 nsew signal output
flabel metal3 s 560 5448 960 5568 0 FreeSans 480 0 0 0 vref_z_p_o[2]
port 60 nsew signal output
flabel metal3 s 560 5720 960 5840 0 FreeSans 480 0 0 0 vref_z_p_o[3]
port 61 nsew signal output
flabel metal3 s 560 5992 960 6112 0 FreeSans 480 0 0 0 vref_z_p_o[4]
port 62 nsew signal output
flabel metal3 s 560 6264 960 6384 0 FreeSans 480 0 0 0 vref_z_p_o[5]
port 63 nsew signal output
flabel metal3 s 560 6536 960 6656 0 FreeSans 480 0 0 0 vref_z_p_o[6]
port 64 nsew signal output
flabel metal3 s 560 6808 960 6928 0 FreeSans 480 0 0 0 vref_z_p_o[7]
port 65 nsew signal output
flabel metal3 s 560 7080 960 7200 0 FreeSans 480 0 0 0 vref_z_p_o[8]
port 66 nsew signal output
flabel metal3 s 560 7352 960 7472 0 FreeSans 480 0 0 0 vref_z_p_o[9]
port 67 nsew signal output
flabel metal3 s 560 1912 960 2032 0 FreeSans 480 0 0 0 vss_p_o[0]
port 79 nsew signal output
flabel metal3 s 560 4632 960 4752 0 FreeSans 480 0 0 0 vss_p_o[10]
port 80 nsew signal output
flabel metal3 s 560 2184 960 2304 0 FreeSans 480 0 0 0 vss_p_o[1]
port 81 nsew signal output
flabel metal3 s 560 2456 960 2576 0 FreeSans 480 0 0 0 vss_p_o[2]
port 82 nsew signal output
flabel metal3 s 560 2728 960 2848 0 FreeSans 480 0 0 0 vss_p_o[3]
port 83 nsew signal output
flabel metal3 s 560 3000 960 3120 0 FreeSans 480 0 0 0 vss_p_o[4]
port 84 nsew signal output
flabel metal3 s 560 3272 960 3392 0 FreeSans 480 0 0 0 vss_p_o[5]
port 85 nsew signal output
flabel metal3 s 560 3544 960 3664 0 FreeSans 480 0 0 0 vss_p_o[6]
port 86 nsew signal output
flabel metal3 s 560 3816 960 3936 0 FreeSans 480 0 0 0 vss_p_o[7]
port 87 nsew signal output
flabel metal3 s 560 4088 960 4208 0 FreeSans 480 0 0 0 vss_p_o[8]
port 88 nsew signal output
flabel metal3 s 560 4360 960 4480 0 FreeSans 480 0 0 0 vss_p_o[9]
port 89 nsew signal output
rlabel metal3 28036 7956 28036 7956 0 vin_n_sw_on
rlabel metal3 27990 5780 27990 5780 0 vref_z_n_o[3]
rlabel metal3 27990 6868 27990 6868 0 vref_z_n_o[7]
rlabel metal3 28174 3060 28174 3060 0 vss_n_o[4]
rlabel metal3 27990 3332 27990 3332 0 vss_n_o[5]
rlabel metal3 28174 4148 28174 4148 0 vss_n_o[8]
rlabel metal3 27990 4420 27990 4420 0 vss_n_o[9]
flabel metal3 s 28020 4360 28420 4480 0 FreeSans 480 0 0 0 vss_n_o[9]
port 78 nsew signal output
flabel metal3 s 28020 4088 28420 4208 0 FreeSans 480 0 0 0 vss_n_o[8]
port 77 nsew signal output
flabel metal3 s 28020 3816 28420 3936 0 FreeSans 480 0 0 0 vss_n_o[7]
port 76 nsew signal output
flabel metal3 s 28020 3544 28420 3664 0 FreeSans 480 0 0 0 vss_n_o[6]
port 75 nsew signal output
flabel metal3 s 28020 3272 28420 3392 0 FreeSans 480 0 0 0 vss_n_o[5]
port 74 nsew signal output
flabel metal3 s 28020 3000 28420 3120 0 FreeSans 480 0 0 0 vss_n_o[4]
port 73 nsew signal output
flabel metal3 s 28020 2728 28420 2848 0 FreeSans 480 0 0 0 vss_n_o[3]
port 72 nsew signal output
flabel metal3 s 28020 2456 28420 2576 0 FreeSans 480 0 0 0 vss_n_o[2]
port 71 nsew signal output
flabel metal3 s 28020 2184 28420 2304 0 FreeSans 480 0 0 0 vss_n_o[1]
port 70 nsew signal output
flabel metal3 s 28020 4632 28420 4752 0 FreeSans 480 0 0 0 vss_n_o[10]
port 69 nsew signal output
flabel metal3 s 28020 1912 28420 2032 0 FreeSans 480 0 0 0 vss_n_o[0]
port 68 nsew signal output
flabel metal3 s 28020 7352 28420 7472 0 FreeSans 480 0 0 0 vref_z_n_o[9]
port 56 nsew signal output
flabel metal3 s 28020 7080 28420 7200 0 FreeSans 480 0 0 0 vref_z_n_o[8]
port 55 nsew signal output
flabel metal3 s 28020 6808 28420 6928 0 FreeSans 480 0 0 0 vref_z_n_o[7]
port 54 nsew signal output
flabel metal3 s 28020 6536 28420 6656 0 FreeSans 480 0 0 0 vref_z_n_o[6]
port 53 nsew signal output
flabel metal3 s 28020 6264 28420 6384 0 FreeSans 480 0 0 0 vref_z_n_o[5]
port 52 nsew signal output
flabel metal3 s 28020 5992 28420 6112 0 FreeSans 480 0 0 0 vref_z_n_o[4]
port 51 nsew signal output
flabel metal3 s 28020 5720 28420 5840 0 FreeSans 480 0 0 0 vref_z_n_o[3]
port 50 nsew signal output
flabel metal3 s 28020 5448 28420 5568 0 FreeSans 480 0 0 0 vref_z_n_o[2]
port 49 nsew signal output
flabel metal3 s 28020 5176 28420 5296 0 FreeSans 480 0 0 0 vref_z_n_o[1]
port 48 nsew signal output
flabel metal3 s 28020 7624 28420 7744 0 FreeSans 480 0 0 0 vref_z_n_o[10]
port 47 nsew signal output
flabel metal3 s 28020 4904 28420 5024 0 FreeSans 480 0 0 0 vref_z_n_o[0]
port 46 nsew signal output
flabel metal3 s 28020 7896 28420 8016 0 FreeSans 480 0 0 0 vin_n_sw_on
port 44 nsew signal input
rlabel metal2 22310 1612 22310 1612 0 vcm_o[10]
flabel metal2 s 22834 7710 22890 8110 0 FreeSans 224 90 0 0 start
port 20 nsew signal input
flabel metal2 s 25226 7710 25282 8110 0 FreeSans 224 90 0 0 single_ended
port 19 nsew signal input
flabel metal2 s 18050 7710 18106 8110 0 FreeSans 224 90 0 0 rst_z
port 17 nsew signal input
flabel metal2 s 27618 7710 27674 8110 0 FreeSans 224 90 0 0 en_offset_cal
port 12 nsew signal input
flabel metal2 s 15658 7710 15714 8110 0 FreeSans 224 90 0 0 data[5]
port 10 nsew signal output
flabel metal2 s 13266 7710 13322 8110 0 FreeSans 224 90 0 0 data[4]
port 9 nsew signal output
flabel metal2 s 10874 7710 10930 8110 0 FreeSans 224 90 0 0 data[3]
port 8 nsew signal output
flabel metal2 s 8482 7710 8538 8110 0 FreeSans 224 90 0 0 data[2]
port 7 nsew signal output
flabel metal2 s 6090 7710 6146 8110 0 FreeSans 224 90 0 0 data[1]
port 6 nsew signal output
flabel metal2 s 3698 7710 3754 8110 0 FreeSans 224 90 0 0 data[0]
port 5 nsew signal output
flabel metal2 s 1306 7710 1362 8110 0 FreeSans 224 90 0 0 clk_data
port 3 nsew signal output
flabel metal2 s 20442 7710 20498 8110 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 21362 1200 21418 1600 0 FreeSans 224 90 0 0 vcm_o_i[9]
port 43 nsew signal input
flabel metal2 s 19522 1200 19578 1600 0 FreeSans 224 90 0 0 vcm_o_i[8]
port 42 nsew signal input
flabel metal2 s 17682 1200 17738 1600 0 FreeSans 224 90 0 0 vcm_o_i[7]
port 41 nsew signal input
flabel metal2 s 15842 1200 15898 1600 0 FreeSans 224 90 0 0 vcm_o_i[6]
port 40 nsew signal input
flabel metal2 s 14002 1200 14058 1600 0 FreeSans 224 90 0 0 vcm_o_i[5]
port 39 nsew signal input
flabel metal2 s 12162 1200 12218 1600 0 FreeSans 224 90 0 0 vcm_o_i[4]
port 38 nsew signal input
flabel metal2 s 10322 1200 10378 1600 0 FreeSans 224 90 0 0 vcm_o_i[3]
port 37 nsew signal input
flabel metal2 s 8482 1200 8538 1600 0 FreeSans 224 90 0 0 vcm_o_i[2]
port 36 nsew signal input
flabel metal2 s 6642 1200 6698 1600 0 FreeSans 224 90 0 0 vcm_o_i[1]
port 35 nsew signal input
flabel metal2 s 23202 1200 23258 1600 0 FreeSans 224 90 0 0 vcm_o_i[10]
port 34 nsew signal input
flabel metal2 s 4802 1200 4858 1600 0 FreeSans 224 90 0 0 vcm_o_i[0]
port 33 nsew signal input
flabel metal2 s 20442 1200 20498 1600 0 FreeSans 224 90 0 0 vcm_o[9]
port 32 nsew signal output
flabel metal2 s 18602 1200 18658 1600 0 FreeSans 224 90 0 0 vcm_o[8]
port 31 nsew signal output
flabel metal2 s 16762 1200 16818 1600 0 FreeSans 224 90 0 0 vcm_o[7]
port 30 nsew signal output
flabel metal2 s 14922 1200 14978 1600 0 FreeSans 224 90 0 0 vcm_o[6]
port 29 nsew signal output
flabel metal2 s 13082 1200 13138 1600 0 FreeSans 224 90 0 0 vcm_o[5]
port 28 nsew signal output
flabel metal2 s 11242 1200 11298 1600 0 FreeSans 224 90 0 0 vcm_o[4]
port 27 nsew signal output
flabel metal2 s 9402 1200 9458 1600 0 FreeSans 224 90 0 0 vcm_o[3]
port 26 nsew signal output
flabel metal2 s 7562 1200 7618 1600 0 FreeSans 224 90 0 0 vcm_o[2]
port 25 nsew signal output
flabel metal2 s 5722 1200 5778 1600 0 FreeSans 224 90 0 0 vcm_o[1]
port 24 nsew signal output
flabel metal2 s 22282 1200 22338 1600 0 FreeSans 224 90 0 0 vcm_o[10]
port 23 nsew signal output
flabel metal2 s 3882 1200 3938 1600 0 FreeSans 224 90 0 0 vcm_o[0]
port 22 nsew signal output
flabel metal2 s 24122 1200 24178 1600 0 FreeSans 224 90 0 0 vcm_dummy_o
port 21 nsew signal output
flabel metal2 s 1122 1200 1178 1600 0 FreeSans 224 90 0 0 sample_o
port 18 nsew signal output
flabel metal2 s 26882 1200 26938 1600 0 FreeSans 224 90 0 0 offset_cal_cycle
port 16 nsew signal output
flabel metal2 s 25962 1200 26018 1600 0 FreeSans 224 90 0 0 en_vcm_sw_o_i
port 15 nsew signal input
flabel metal2 s 25042 1200 25098 1600 0 FreeSans 224 90 0 0 en_vcm_sw_o
port 14 nsew signal output
flabel metal2 s 27802 1200 27858 1600 0 FreeSans 224 90 0 0 en_offset_cal_o
port 13 nsew signal output
flabel metal2 s 2042 1200 2098 1600 0 FreeSans 224 90 0 0 en_comp
port 11 nsew signal output
flabel metal2 s 2962 1200 3018 1600 0 FreeSans 224 90 0 0 comp_p
port 4 nsew signal input
rlabel metal2 25990 1355 25990 1355 0 en_vcm_sw_o_i
rlabel metal2 24150 1355 24150 1355 0 vcm_dummy_o
rlabel metal2 4830 1474 4830 1474 0 vcm_o_i[0]
rlabel metal2 5750 1375 5750 1375 0 vcm_o[1]
rlabel metal2 1334 7968 1334 7968 0 clk_data
rlabel metal2 3726 7832 3726 7832 0 data[0]
rlabel metal2 6118 8002 6118 8002 0 data[1]
rlabel metal2 8510 8002 8510 8002 0 data[2]
rlabel metal2 10902 8002 10902 8002 0 data[3]
rlabel metal2 13294 8002 13294 8002 0 data[4]
rlabel metal2 15686 7965 15686 7965 0 data[5]
rlabel metal3 724 5236 724 5236 0 vref_z_p_o[1]
rlabel metal3 632 5780 632 5780 0 vref_z_p_o[3]
rlabel metal3 632 4692 632 4692 0 vss_p_o[10]
<< properties >>
string FIXED_BBOX 0 0 29000 10000
<< end >>
