magic
tech sky130A
magscale 1 2
timestamp 1710680845
<< nwell >>
rect -6283 -594 6283 594
<< pmos >>
rect -6087 -375 -3087 375
rect -3029 -375 -29 375
rect 29 -375 3029 375
rect 3087 -375 6087 375
<< pdiff >>
rect -6145 363 -6087 375
rect -6145 -363 -6133 363
rect -6099 -363 -6087 363
rect -6145 -375 -6087 -363
rect -3087 363 -3029 375
rect -3087 -363 -3075 363
rect -3041 -363 -3029 363
rect -3087 -375 -3029 -363
rect -29 363 29 375
rect -29 -363 -17 363
rect 17 -363 29 363
rect -29 -375 29 -363
rect 3029 363 3087 375
rect 3029 -363 3041 363
rect 3075 -363 3087 363
rect 3029 -375 3087 -363
rect 6087 363 6145 375
rect 6087 -363 6099 363
rect 6133 -363 6145 363
rect 6087 -375 6145 -363
<< pdiffc >>
rect -6133 -363 -6099 363
rect -3075 -363 -3041 363
rect -17 -363 17 363
rect 3041 -363 3075 363
rect 6099 -363 6133 363
<< nsubdiff >>
rect -6247 524 -6151 558
rect 6151 524 6247 558
rect -6247 462 -6213 524
rect 6213 462 6247 524
rect -6247 -524 -6213 -462
rect 6213 -524 6247 -462
rect -6247 -558 -6151 -524
rect 6151 -558 6247 -524
<< nsubdiffcont >>
rect -6151 524 6151 558
rect -6247 -462 -6213 462
rect 6213 -462 6247 462
rect -6151 -558 6151 -524
<< poly >>
rect -6087 456 -3087 472
rect -6087 422 -6071 456
rect -3103 422 -3087 456
rect -6087 375 -3087 422
rect -3029 456 -29 472
rect -3029 422 -3013 456
rect -45 422 -29 456
rect -3029 375 -29 422
rect 29 456 3029 472
rect 29 422 45 456
rect 3013 422 3029 456
rect 29 375 3029 422
rect 3087 456 6087 472
rect 3087 422 3103 456
rect 6071 422 6087 456
rect 3087 375 6087 422
rect -6087 -422 -3087 -375
rect -6087 -456 -6071 -422
rect -3103 -456 -3087 -422
rect -6087 -472 -3087 -456
rect -3029 -422 -29 -375
rect -3029 -456 -3013 -422
rect -45 -456 -29 -422
rect -3029 -472 -29 -456
rect 29 -422 3029 -375
rect 29 -456 45 -422
rect 3013 -456 3029 -422
rect 29 -472 3029 -456
rect 3087 -422 6087 -375
rect 3087 -456 3103 -422
rect 6071 -456 6087 -422
rect 3087 -472 6087 -456
<< polycont >>
rect -6071 422 -3103 456
rect -3013 422 -45 456
rect 45 422 3013 456
rect 3103 422 6071 456
rect -6071 -456 -3103 -422
rect -3013 -456 -45 -422
rect 45 -456 3013 -422
rect 3103 -456 6071 -422
<< locali >>
rect -6247 524 -6151 558
rect 6151 524 6247 558
rect -6247 462 -6213 524
rect 6213 462 6247 524
rect -6087 422 -6071 456
rect -3103 422 -3087 456
rect -3029 422 -3013 456
rect -45 422 -29 456
rect 29 422 45 456
rect 3013 422 3029 456
rect 3087 422 3103 456
rect 6071 422 6087 456
rect -6133 363 -6099 379
rect -6133 -379 -6099 -363
rect -3075 363 -3041 379
rect -3075 -379 -3041 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 3041 363 3075 379
rect 3041 -379 3075 -363
rect 6099 363 6133 379
rect 6099 -379 6133 -363
rect -6087 -456 -6071 -422
rect -3103 -456 -3087 -422
rect -3029 -456 -3013 -422
rect -45 -456 -29 -422
rect 29 -456 45 -422
rect 3013 -456 3029 -422
rect 3087 -456 3103 -422
rect 6071 -456 6087 -422
rect -6247 -524 -6213 -462
rect 6213 -524 6247 -462
rect -6247 -558 -6151 -524
rect 6151 -558 6247 -524
<< viali >>
rect -6071 422 -3103 456
rect -3013 422 -45 456
rect 45 422 3013 456
rect 3103 422 6071 456
rect -6133 -363 -6099 363
rect -3075 -363 -3041 363
rect -17 -363 17 363
rect 3041 -363 3075 363
rect 6099 -363 6133 363
rect -6071 -456 -3103 -422
rect -3013 -456 -45 -422
rect 45 -456 3013 -422
rect 3103 -456 6071 -422
<< metal1 >>
rect -6083 456 -3091 462
rect -6083 422 -6071 456
rect -3103 422 -3091 456
rect -6083 416 -3091 422
rect -3025 456 -33 462
rect -3025 422 -3013 456
rect -45 422 -33 456
rect -3025 416 -33 422
rect 33 456 3025 462
rect 33 422 45 456
rect 3013 422 3025 456
rect 33 416 3025 422
rect 3091 456 6083 462
rect 3091 422 3103 456
rect 6071 422 6083 456
rect 3091 416 6083 422
rect -6139 363 -6093 375
rect -6139 -363 -6133 363
rect -6099 -363 -6093 363
rect -6139 -375 -6093 -363
rect -3081 363 -3035 375
rect -3081 -363 -3075 363
rect -3041 -363 -3035 363
rect -3081 -375 -3035 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 3035 363 3081 375
rect 3035 -363 3041 363
rect 3075 -363 3081 363
rect 3035 -375 3081 -363
rect 6093 363 6139 375
rect 6093 -363 6099 363
rect 6133 -363 6139 363
rect 6093 -375 6139 -363
rect -6083 -422 -3091 -416
rect -6083 -456 -6071 -422
rect -3103 -456 -3091 -422
rect -6083 -462 -3091 -456
rect -3025 -422 -33 -416
rect -3025 -456 -3013 -422
rect -45 -456 -33 -422
rect -3025 -462 -33 -456
rect 33 -422 3025 -416
rect 33 -456 45 -422
rect 3013 -456 3025 -422
rect 33 -462 3025 -456
rect 3091 -422 6083 -416
rect 3091 -456 3103 -422
rect 6071 -456 6083 -422
rect 3091 -462 6083 -456
<< properties >>
string FIXED_BBOX -6230 -541 6230 541
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.75 l 15.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
