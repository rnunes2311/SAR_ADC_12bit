magic
tech sky130A
magscale 1 2
timestamp 1711813427
<< error_p >>
rect -659 272 -601 278
rect -239 272 -181 278
rect 181 272 239 278
rect 601 272 659 278
rect -659 238 -647 272
rect -239 238 -227 272
rect 181 238 193 272
rect 601 238 613 272
rect -659 232 -601 238
rect -239 232 -181 238
rect 181 232 239 238
rect 601 232 659 238
rect -869 -238 -811 -232
rect -449 -238 -391 -232
rect -29 -238 29 -232
rect 391 -238 449 -232
rect 811 -238 869 -232
rect -869 -272 -857 -238
rect -449 -272 -437 -238
rect -29 -272 -17 -238
rect 391 -272 403 -238
rect 811 -272 823 -238
rect -869 -278 -811 -272
rect -449 -278 -391 -272
rect -29 -278 29 -272
rect 391 -278 449 -272
rect 811 -278 869 -272
<< nmoslvt >>
rect -855 -200 -825 200
rect -645 -200 -615 200
rect -435 -200 -405 200
rect -225 -200 -195 200
rect -15 -200 15 200
rect 195 -200 225 200
rect 405 -200 435 200
rect 615 -200 645 200
rect 825 -200 855 200
<< ndiff >>
rect -917 188 -855 200
rect -917 -188 -905 188
rect -871 -188 -855 188
rect -917 -200 -855 -188
rect -825 188 -763 200
rect -825 -188 -809 188
rect -775 -188 -763 188
rect -825 -200 -763 -188
rect -707 188 -645 200
rect -707 -188 -695 188
rect -661 -188 -645 188
rect -707 -200 -645 -188
rect -615 188 -553 200
rect -615 -188 -599 188
rect -565 -188 -553 188
rect -615 -200 -553 -188
rect -497 188 -435 200
rect -497 -188 -485 188
rect -451 -188 -435 188
rect -497 -200 -435 -188
rect -405 188 -343 200
rect -405 -188 -389 188
rect -355 -188 -343 188
rect -405 -200 -343 -188
rect -287 188 -225 200
rect -287 -188 -275 188
rect -241 -188 -225 188
rect -287 -200 -225 -188
rect -195 188 -133 200
rect -195 -188 -179 188
rect -145 -188 -133 188
rect -195 -200 -133 -188
rect -77 188 -15 200
rect -77 -188 -65 188
rect -31 -188 -15 188
rect -77 -200 -15 -188
rect 15 188 77 200
rect 15 -188 31 188
rect 65 -188 77 188
rect 15 -200 77 -188
rect 133 188 195 200
rect 133 -188 145 188
rect 179 -188 195 188
rect 133 -200 195 -188
rect 225 188 287 200
rect 225 -188 241 188
rect 275 -188 287 188
rect 225 -200 287 -188
rect 343 188 405 200
rect 343 -188 355 188
rect 389 -188 405 188
rect 343 -200 405 -188
rect 435 188 497 200
rect 435 -188 451 188
rect 485 -188 497 188
rect 435 -200 497 -188
rect 553 188 615 200
rect 553 -188 565 188
rect 599 -188 615 188
rect 553 -200 615 -188
rect 645 188 707 200
rect 645 -188 661 188
rect 695 -188 707 188
rect 645 -200 707 -188
rect 763 188 825 200
rect 763 -188 775 188
rect 809 -188 825 188
rect 763 -200 825 -188
rect 855 188 917 200
rect 855 -188 871 188
rect 905 -188 917 188
rect 855 -200 917 -188
<< ndiffc >>
rect -905 -188 -871 188
rect -809 -188 -775 188
rect -695 -188 -661 188
rect -599 -188 -565 188
rect -485 -188 -451 188
rect -389 -188 -355 188
rect -275 -188 -241 188
rect -179 -188 -145 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 145 -188 179 188
rect 241 -188 275 188
rect 355 -188 389 188
rect 451 -188 485 188
rect 565 -188 599 188
rect 661 -188 695 188
rect 775 -188 809 188
rect 871 -188 905 188
<< poly >>
rect -663 272 -597 288
rect -663 238 -647 272
rect -613 238 -597 272
rect -855 200 -825 226
rect -663 222 -597 238
rect -243 272 -177 288
rect -243 238 -227 272
rect -193 238 -177 272
rect -645 200 -615 222
rect -435 200 -405 226
rect -243 222 -177 238
rect 177 272 243 288
rect 177 238 193 272
rect 227 238 243 272
rect -225 200 -195 222
rect -15 200 15 226
rect 177 222 243 238
rect 597 272 663 288
rect 597 238 613 272
rect 647 238 663 272
rect 195 200 225 222
rect 405 200 435 226
rect 597 222 663 238
rect 615 200 645 222
rect 825 200 855 226
rect -855 -222 -825 -200
rect -873 -238 -807 -222
rect -645 -226 -615 -200
rect -435 -222 -405 -200
rect -873 -272 -857 -238
rect -823 -272 -807 -238
rect -873 -288 -807 -272
rect -453 -238 -387 -222
rect -225 -226 -195 -200
rect -15 -222 15 -200
rect -453 -272 -437 -238
rect -403 -272 -387 -238
rect -453 -288 -387 -272
rect -33 -238 33 -222
rect 195 -226 225 -200
rect 405 -222 435 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 387 -238 453 -222
rect 615 -226 645 -200
rect 825 -222 855 -200
rect 387 -272 403 -238
rect 437 -272 453 -238
rect 387 -288 453 -272
rect 807 -238 873 -222
rect 807 -272 823 -238
rect 857 -272 873 -238
rect 807 -288 873 -272
<< polycont >>
rect -647 238 -613 272
rect -227 238 -193 272
rect 193 238 227 272
rect 613 238 647 272
rect -857 -272 -823 -238
rect -437 -272 -403 -238
rect -17 -272 17 -238
rect 403 -272 437 -238
rect 823 -272 857 -238
<< locali >>
rect -663 238 -647 272
rect -613 238 -597 272
rect -243 238 -227 272
rect -193 238 -177 272
rect 177 238 193 272
rect 227 238 243 272
rect 597 238 613 272
rect 647 238 663 272
rect -905 188 -871 204
rect -905 -204 -871 -188
rect -809 188 -775 204
rect -809 -204 -775 -188
rect -695 188 -661 204
rect -695 -204 -661 -188
rect -599 188 -565 204
rect -599 -204 -565 -188
rect -485 188 -451 204
rect -485 -204 -451 -188
rect -389 188 -355 204
rect -389 -204 -355 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -179 188 -145 204
rect -179 -204 -145 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 145 188 179 204
rect 145 -204 179 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 355 188 389 204
rect 355 -204 389 -188
rect 451 188 485 204
rect 451 -204 485 -188
rect 565 188 599 204
rect 565 -204 599 -188
rect 661 188 695 204
rect 661 -204 695 -188
rect 775 188 809 204
rect 775 -204 809 -188
rect 871 188 905 204
rect 871 -204 905 -188
rect -873 -272 -857 -238
rect -823 -272 -807 -238
rect -453 -272 -437 -238
rect -403 -272 -387 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 387 -272 403 -238
rect 437 -272 453 -238
rect 807 -272 823 -238
rect 857 -272 873 -238
<< viali >>
rect -647 238 -613 272
rect -227 238 -193 272
rect 193 238 227 272
rect 613 238 647 272
rect -905 -188 -871 188
rect -809 -188 -775 188
rect -695 -188 -661 188
rect -599 -188 -565 188
rect -485 -188 -451 188
rect -389 -188 -355 188
rect -275 -188 -241 188
rect -179 -188 -145 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 145 -188 179 188
rect 241 -188 275 188
rect 355 -188 389 188
rect 451 -188 485 188
rect 565 -188 599 188
rect 661 -188 695 188
rect 775 -188 809 188
rect 871 -188 905 188
rect -857 -272 -823 -238
rect -437 -272 -403 -238
rect -17 -272 17 -238
rect 403 -272 437 -238
rect 823 -272 857 -238
<< metal1 >>
rect -659 272 -601 278
rect -659 238 -647 272
rect -613 238 -601 272
rect -659 232 -601 238
rect -239 272 -181 278
rect -239 238 -227 272
rect -193 238 -181 272
rect -239 232 -181 238
rect 181 272 239 278
rect 181 238 193 272
rect 227 238 239 272
rect 181 232 239 238
rect 601 272 659 278
rect 601 238 613 272
rect 647 238 659 272
rect 601 232 659 238
rect -911 188 -865 200
rect -911 -188 -905 188
rect -871 -188 -865 188
rect -911 -200 -865 -188
rect -815 188 -769 200
rect -815 -188 -809 188
rect -775 -188 -769 188
rect -815 -200 -769 -188
rect -701 188 -655 200
rect -701 -188 -695 188
rect -661 -188 -655 188
rect -701 -200 -655 -188
rect -605 188 -559 200
rect -605 -188 -599 188
rect -565 -188 -559 188
rect -605 -200 -559 -188
rect -491 188 -445 200
rect -491 -188 -485 188
rect -451 -188 -445 188
rect -491 -200 -445 -188
rect -395 188 -349 200
rect -395 -188 -389 188
rect -355 -188 -349 188
rect -395 -200 -349 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -185 188 -139 200
rect -185 -188 -179 188
rect -145 -188 -139 188
rect -185 -200 -139 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 139 188 185 200
rect 139 -188 145 188
rect 179 -188 185 188
rect 139 -200 185 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 349 188 395 200
rect 349 -188 355 188
rect 389 -188 395 188
rect 349 -200 395 -188
rect 445 188 491 200
rect 445 -188 451 188
rect 485 -188 491 188
rect 445 -200 491 -188
rect 559 188 605 200
rect 559 -188 565 188
rect 599 -188 605 188
rect 559 -200 605 -188
rect 655 188 701 200
rect 655 -188 661 188
rect 695 -188 701 188
rect 655 -200 701 -188
rect 769 188 815 200
rect 769 -188 775 188
rect 809 -188 815 188
rect 769 -200 815 -188
rect 865 188 911 200
rect 865 -188 871 188
rect 905 -188 911 188
rect 865 -200 911 -188
rect -869 -238 -811 -232
rect -869 -272 -857 -238
rect -823 -272 -811 -238
rect -869 -278 -811 -272
rect -449 -238 -391 -232
rect -449 -272 -437 -238
rect -403 -272 -391 -238
rect -449 -278 -391 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 391 -238 449 -232
rect 391 -272 403 -238
rect 437 -272 449 -238
rect 391 -278 449 -272
rect 811 -238 869 -232
rect 811 -272 823 -238
rect 857 -272 869 -238
rect 811 -278 869 -272
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 9 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
