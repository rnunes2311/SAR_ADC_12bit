magic
tech sky130A
magscale 1 2
timestamp 1711883348
<< error_p >>
rect -221 172 -163 178
rect -29 172 29 178
rect 163 172 221 178
rect -221 138 -209 172
rect -29 138 -17 172
rect 163 138 175 172
rect -221 132 -163 138
rect -29 132 29 138
rect 163 132 221 138
rect -317 -138 -259 -132
rect -125 -138 -67 -132
rect 67 -138 125 -132
rect 259 -138 317 -132
rect -317 -172 -305 -138
rect -125 -172 -113 -138
rect 67 -172 79 -138
rect 259 -172 271 -138
rect -317 -178 -259 -172
rect -125 -178 -67 -172
rect 67 -178 125 -172
rect 259 -178 317 -172
<< pwell >>
rect -503 -310 503 310
<< nmos >>
rect -303 -100 -273 100
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
rect 273 -100 303 100
<< ndiff >>
rect -365 88 -303 100
rect -365 -88 -353 88
rect -319 -88 -303 88
rect -365 -100 -303 -88
rect -273 88 -207 100
rect -273 -88 -257 88
rect -223 -88 -207 88
rect -273 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 273 100
rect 207 -88 223 88
rect 257 -88 273 88
rect 207 -100 273 -88
rect 303 88 365 100
rect 303 -88 319 88
rect 353 -88 365 88
rect 303 -100 365 -88
<< ndiffc >>
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
<< psubdiff >>
rect -467 240 -371 274
rect 371 240 467 274
rect -467 178 -433 240
rect 433 178 467 240
rect -467 -240 -433 -178
rect 433 -240 467 -178
rect -467 -274 -371 -240
rect 371 -274 467 -240
<< psubdiffcont >>
rect -371 240 371 274
rect -467 -178 -433 178
rect 433 -178 467 178
rect -371 -274 371 -240
<< poly >>
rect -225 172 -159 188
rect -225 138 -209 172
rect -175 138 -159 172
rect -303 100 -273 126
rect -225 122 -159 138
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -207 100 -177 122
rect -111 100 -81 126
rect -33 122 33 138
rect 159 172 225 188
rect 159 138 175 172
rect 209 138 225 172
rect -15 100 15 122
rect 81 100 111 126
rect 159 122 225 138
rect 177 100 207 122
rect 273 100 303 126
rect -303 -122 -273 -100
rect -321 -138 -255 -122
rect -207 -126 -177 -100
rect -111 -122 -81 -100
rect -321 -172 -305 -138
rect -271 -172 -255 -138
rect -321 -188 -255 -172
rect -129 -138 -63 -122
rect -15 -126 15 -100
rect 81 -122 111 -100
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect -129 -188 -63 -172
rect 63 -138 129 -122
rect 177 -126 207 -100
rect 273 -122 303 -100
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 63 -188 129 -172
rect 255 -138 321 -122
rect 255 -172 271 -138
rect 305 -172 321 -138
rect 255 -188 321 -172
<< polycont >>
rect -209 138 -175 172
rect -17 138 17 172
rect 175 138 209 172
rect -305 -172 -271 -138
rect -113 -172 -79 -138
rect 79 -172 113 -138
rect 271 -172 305 -138
<< locali >>
rect -467 240 -371 274
rect 371 240 467 274
rect -467 178 -433 240
rect 433 178 467 240
rect -225 138 -209 172
rect -175 138 -159 172
rect -33 138 -17 172
rect 17 138 33 172
rect 159 138 175 172
rect 209 138 225 172
rect -353 88 -319 104
rect -353 -104 -319 -88
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect 319 88 353 104
rect 319 -104 353 -88
rect -321 -172 -305 -138
rect -271 -172 -255 -138
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 255 -172 271 -138
rect 305 -172 321 -138
rect -467 -240 -433 -178
rect 433 -240 467 -178
rect -467 -274 -371 -240
rect 371 -274 467 -240
<< viali >>
rect -209 138 -175 172
rect -17 138 17 172
rect 175 138 209 172
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect -305 -172 -271 -138
rect -113 -172 -79 -138
rect 79 -172 113 -138
rect 271 -172 305 -138
<< metal1 >>
rect -221 172 -163 178
rect -221 138 -209 172
rect -175 138 -163 172
rect -221 132 -163 138
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect 163 172 221 178
rect 163 138 175 172
rect 209 138 221 172
rect 163 132 221 138
rect -359 88 -313 100
rect -359 -88 -353 88
rect -319 -88 -313 88
rect -359 -100 -313 -88
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect 313 88 359 100
rect 313 -88 319 88
rect 353 -88 359 88
rect 313 -100 359 -88
rect -317 -138 -259 -132
rect -317 -172 -305 -138
rect -271 -172 -259 -138
rect -317 -178 -259 -172
rect -125 -138 -67 -132
rect -125 -172 -113 -138
rect -79 -172 -67 -138
rect -125 -178 -67 -172
rect 67 -138 125 -132
rect 67 -172 79 -138
rect 113 -172 125 -138
rect 67 -178 125 -172
rect 259 -138 317 -132
rect 259 -172 271 -138
rect 305 -172 317 -138
rect 259 -178 317 -172
<< properties >>
string FIXED_BBOX -450 -257 450 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
