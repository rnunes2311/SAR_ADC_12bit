magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -555 272 -497 278
rect -344 272 -286 278
rect -134 272 -76 278
rect 76 272 134 278
rect 285 276 343 282
rect -555 238 -543 272
rect -344 238 -332 272
rect -134 238 -122 272
rect 76 238 88 272
rect 285 242 297 276
rect 496 272 554 278
rect -555 232 -497 238
rect -344 232 -286 238
rect -134 232 -76 238
rect 76 232 134 238
rect 285 236 343 242
rect 496 238 508 272
rect 496 232 554 238
rect -602 -200 -540 200
rect -510 -200 -448 200
rect -392 -200 -330 200
rect -300 -200 -238 200
rect -182 -200 -120 200
rect -90 -200 -28 200
rect 28 -200 90 200
rect 120 -200 182 200
rect 238 -200 300 200
rect 330 -200 392 200
rect 448 -200 510 200
rect 540 -200 602 200
<< pwell >>
rect -559 222 -493 288
rect -138 222 -72 288
rect 281 226 347 292
<< nmoslvt >>
rect -540 -200 -510 200
rect -330 -200 -300 200
rect -120 -200 -90 200
rect 90 -200 120 200
rect 300 -200 330 200
rect 510 -200 540 200
<< ndiff >>
rect -602 188 -540 200
rect -602 -188 -590 188
rect -556 -188 -540 188
rect -602 -200 -540 -188
rect -510 188 -448 200
rect -510 -188 -494 188
rect -460 -188 -448 188
rect -510 -200 -448 -188
rect -392 188 -330 200
rect -392 -188 -380 188
rect -346 -188 -330 188
rect -392 -200 -330 -188
rect -300 188 -238 200
rect -300 -188 -284 188
rect -250 -188 -238 188
rect -300 -200 -238 -188
rect -182 188 -120 200
rect -182 -188 -170 188
rect -136 -188 -120 188
rect -182 -200 -120 -188
rect -90 188 -28 200
rect -90 -188 -74 188
rect -40 -188 -28 188
rect -90 -200 -28 -188
rect 28 188 90 200
rect 28 -188 40 188
rect 74 -188 90 188
rect 28 -200 90 -188
rect 120 188 182 200
rect 120 -188 136 188
rect 170 -188 182 188
rect 120 -200 182 -188
rect 238 188 300 200
rect 238 -188 250 188
rect 284 -188 300 188
rect 238 -200 300 -188
rect 330 188 392 200
rect 330 -188 346 188
rect 380 -188 392 188
rect 330 -200 392 -188
rect 448 188 510 200
rect 448 -188 460 188
rect 494 -188 510 188
rect 448 -200 510 -188
rect 540 188 602 200
rect 540 -188 556 188
rect 590 -188 602 188
rect 540 -200 602 -188
<< ndiffc >>
rect -590 -188 -556 188
rect -494 -188 -460 188
rect -380 -188 -346 188
rect -284 -188 -250 188
rect -170 -188 -136 188
rect -74 -188 -40 188
rect 40 -188 74 188
rect 136 -188 170 188
rect 250 -188 284 188
rect 346 -188 380 188
rect 460 -188 494 188
rect 556 -188 590 188
<< poly >>
rect -559 272 -493 288
rect -559 238 -543 272
rect -509 238 -493 272
rect -559 222 -493 238
rect -348 272 -282 288
rect -348 238 -332 272
rect -298 238 -282 272
rect -348 222 -282 238
rect -138 272 -72 288
rect -138 238 -122 272
rect -88 238 -72 272
rect -138 222 -72 238
rect 72 272 138 288
rect 72 238 88 272
rect 122 238 138 272
rect 72 222 138 238
rect 281 276 347 292
rect 281 242 297 276
rect 331 242 347 276
rect 281 226 347 242
rect 492 272 558 288
rect 492 238 508 272
rect 542 238 558 272
rect -540 200 -510 222
rect -330 200 -300 222
rect -120 200 -90 222
rect 90 200 120 222
rect 300 200 330 226
rect 492 222 558 238
rect 510 200 540 222
rect -540 -226 -510 -200
rect -330 -226 -300 -200
rect -120 -226 -90 -200
rect 90 -226 120 -200
rect 300 -226 330 -200
rect 510 -226 540 -200
<< polycont >>
rect -543 238 -509 272
rect -332 238 -298 272
rect -122 238 -88 272
rect 88 238 122 272
rect 297 242 331 276
rect 508 238 542 272
<< locali >>
rect -559 238 -543 272
rect -509 238 -493 272
rect -348 238 -332 272
rect -298 238 -282 272
rect -138 238 -122 272
rect -88 238 -72 272
rect 72 238 88 272
rect 122 238 138 272
rect 281 242 297 276
rect 331 242 347 276
rect 492 238 508 272
rect 542 238 558 272
rect -590 188 -556 204
rect -590 -204 -556 -188
rect -494 188 -460 204
rect -494 -204 -460 -188
rect -380 188 -346 204
rect -380 -204 -346 -188
rect -284 188 -250 204
rect -284 -204 -250 -188
rect -170 188 -136 204
rect -170 -204 -136 -188
rect -74 188 -40 204
rect -74 -204 -40 -188
rect 40 188 74 204
rect 40 -204 74 -188
rect 136 188 170 204
rect 136 -204 170 -188
rect 250 188 284 204
rect 250 -204 284 -188
rect 346 188 380 204
rect 346 -204 380 -188
rect 460 188 494 204
rect 460 -204 494 -188
rect 556 188 590 204
rect 556 -204 590 -188
<< viali >>
rect -543 238 -509 272
rect -332 238 -298 272
rect -122 238 -88 272
rect 88 238 122 272
rect 297 242 331 276
rect 508 238 542 272
rect -590 -188 -556 188
rect -494 -188 -460 188
rect -380 -188 -346 188
rect -284 -188 -250 188
rect -170 -188 -136 188
rect -74 -188 -40 188
rect 40 -188 74 188
rect 136 -188 170 188
rect 250 -188 284 188
rect 346 -188 380 188
rect 460 -188 494 188
rect 556 -188 590 188
<< metal1 >>
rect -555 272 -497 278
rect -555 238 -543 272
rect -509 238 -497 272
rect -555 232 -497 238
rect -344 272 -286 278
rect -344 238 -332 272
rect -298 238 -286 272
rect -344 232 -286 238
rect -134 272 -76 278
rect -134 238 -122 272
rect -88 238 -76 272
rect -134 232 -76 238
rect 76 272 134 278
rect 76 238 88 272
rect 122 238 134 272
rect 76 232 134 238
rect 285 276 343 282
rect 285 242 297 276
rect 331 242 343 276
rect 285 236 343 242
rect 496 272 554 278
rect 496 238 508 272
rect 542 238 554 272
rect 496 232 554 238
rect -596 188 -550 200
rect -596 -188 -590 188
rect -556 -188 -550 188
rect -596 -200 -550 -188
rect -500 188 -454 200
rect -500 -188 -494 188
rect -460 -188 -454 188
rect -500 -200 -454 -188
rect -386 188 -340 200
rect -386 -188 -380 188
rect -346 -188 -340 188
rect -386 -200 -340 -188
rect -290 188 -244 200
rect -290 -188 -284 188
rect -250 -188 -244 188
rect -290 -200 -244 -188
rect -176 188 -130 200
rect -176 -188 -170 188
rect -136 -188 -130 188
rect -176 -200 -130 -188
rect -80 188 -34 200
rect -80 -188 -74 188
rect -40 -188 -34 188
rect -80 -200 -34 -188
rect 34 188 80 200
rect 34 -188 40 188
rect 74 -188 80 188
rect 34 -200 80 -188
rect 130 188 176 200
rect 130 -188 136 188
rect 170 -188 176 188
rect 130 -200 176 -188
rect 244 188 290 200
rect 244 -188 250 188
rect 284 -188 290 188
rect 244 -200 290 -188
rect 340 188 386 200
rect 340 -188 346 188
rect 380 -188 386 188
rect 340 -200 386 -188
rect 454 188 500 200
rect 454 -188 460 188
rect 494 -188 500 188
rect 454 -200 500 -188
rect 550 188 596 200
rect 550 -188 556 188
rect 590 -188 596 188
rect 550 -200 596 -188
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
