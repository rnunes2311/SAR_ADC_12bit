magic
tech sky130A
magscale 1 2
timestamp 1711831168
<< nwell >>
rect -3225 -1087 3225 1087
<< pmos >>
rect -3029 118 -29 868
rect 29 118 3029 868
rect -3029 -868 -29 -118
rect 29 -868 3029 -118
<< pdiff >>
rect -3087 856 -3029 868
rect -3087 130 -3075 856
rect -3041 130 -3029 856
rect -3087 118 -3029 130
rect -29 856 29 868
rect -29 130 -17 856
rect 17 130 29 856
rect -29 118 29 130
rect 3029 856 3087 868
rect 3029 130 3041 856
rect 3075 130 3087 856
rect 3029 118 3087 130
rect -3087 -130 -3029 -118
rect -3087 -856 -3075 -130
rect -3041 -856 -3029 -130
rect -3087 -868 -3029 -856
rect -29 -130 29 -118
rect -29 -856 -17 -130
rect 17 -856 29 -130
rect -29 -868 29 -856
rect 3029 -130 3087 -118
rect 3029 -856 3041 -130
rect 3075 -856 3087 -130
rect 3029 -868 3087 -856
<< pdiffc >>
rect -3075 130 -3041 856
rect -17 130 17 856
rect 3041 130 3075 856
rect -3075 -856 -3041 -130
rect -17 -856 17 -130
rect 3041 -856 3075 -130
<< nsubdiff >>
rect -3189 1017 -3093 1051
rect 3093 1017 3189 1051
rect -3189 955 -3155 1017
rect 3155 955 3189 1017
rect -3189 -1017 -3155 -955
rect 3155 -1017 3189 -955
rect -3189 -1051 -3093 -1017
rect 3093 -1051 3189 -1017
<< nsubdiffcont >>
rect -3093 1017 3093 1051
rect -3189 -955 -3155 955
rect 3155 -955 3189 955
rect -3093 -1051 3093 -1017
<< poly >>
rect -3029 949 -29 965
rect -3029 915 -3013 949
rect -45 915 -29 949
rect -3029 868 -29 915
rect 29 949 3029 965
rect 29 915 45 949
rect 3013 915 3029 949
rect 29 868 3029 915
rect -3029 71 -29 118
rect -3029 37 -3013 71
rect -45 37 -29 71
rect -3029 21 -29 37
rect 29 71 3029 118
rect 29 37 45 71
rect 3013 37 3029 71
rect 29 21 3029 37
rect -3029 -37 -29 -21
rect -3029 -71 -3013 -37
rect -45 -71 -29 -37
rect -3029 -118 -29 -71
rect 29 -37 3029 -21
rect 29 -71 45 -37
rect 3013 -71 3029 -37
rect 29 -118 3029 -71
rect -3029 -915 -29 -868
rect -3029 -949 -3013 -915
rect -45 -949 -29 -915
rect -3029 -965 -29 -949
rect 29 -915 3029 -868
rect 29 -949 45 -915
rect 3013 -949 3029 -915
rect 29 -965 3029 -949
<< polycont >>
rect -3013 915 -45 949
rect 45 915 3013 949
rect -3013 37 -45 71
rect 45 37 3013 71
rect -3013 -71 -45 -37
rect 45 -71 3013 -37
rect -3013 -949 -45 -915
rect 45 -949 3013 -915
<< locali >>
rect -3189 1017 -3093 1051
rect 3093 1017 3189 1051
rect -3189 955 -3155 1017
rect 3155 955 3189 1017
rect -3029 915 -3013 949
rect -45 915 -29 949
rect 29 915 45 949
rect 3013 915 3029 949
rect -3075 856 -3041 872
rect -3075 114 -3041 130
rect -17 856 17 872
rect -17 114 17 130
rect 3041 856 3075 872
rect 3041 114 3075 130
rect -3029 37 -3013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 3013 37 3029 71
rect -3029 -71 -3013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 3013 -71 3029 -37
rect -3075 -130 -3041 -114
rect -3075 -872 -3041 -856
rect -17 -130 17 -114
rect -17 -872 17 -856
rect 3041 -130 3075 -114
rect 3041 -872 3075 -856
rect -3029 -949 -3013 -915
rect -45 -949 -29 -915
rect 29 -949 45 -915
rect 3013 -949 3029 -915
rect -3189 -1017 -3155 -955
rect 3155 -1017 3189 -955
rect -3189 -1051 -3093 -1017
rect 3093 -1051 3189 -1017
<< viali >>
rect -3013 915 -45 949
rect 45 915 3013 949
rect -3075 130 -3041 856
rect -17 130 17 856
rect 3041 130 3075 856
rect -3013 37 -45 71
rect 45 37 3013 71
rect -3013 -71 -45 -37
rect 45 -71 3013 -37
rect -3075 -856 -3041 -130
rect -17 -856 17 -130
rect 3041 -856 3075 -130
rect -3013 -949 -45 -915
rect 45 -949 3013 -915
<< metal1 >>
rect -3025 949 -33 955
rect -3025 915 -3013 949
rect -45 915 -33 949
rect -3025 909 -33 915
rect 33 949 3025 955
rect 33 915 45 949
rect 3013 915 3025 949
rect 33 909 3025 915
rect -3081 856 -3035 868
rect -3081 130 -3075 856
rect -3041 130 -3035 856
rect -3081 118 -3035 130
rect -23 856 23 868
rect -23 130 -17 856
rect 17 130 23 856
rect -23 118 23 130
rect 3035 856 3081 868
rect 3035 130 3041 856
rect 3075 130 3081 856
rect 3035 118 3081 130
rect -3025 71 -33 77
rect -3025 37 -3013 71
rect -45 37 -33 71
rect -3025 31 -33 37
rect 33 71 3025 77
rect 33 37 45 71
rect 3013 37 3025 71
rect 33 31 3025 37
rect -3025 -37 -33 -31
rect -3025 -71 -3013 -37
rect -45 -71 -33 -37
rect -3025 -77 -33 -71
rect 33 -37 3025 -31
rect 33 -71 45 -37
rect 3013 -71 3025 -37
rect 33 -77 3025 -71
rect -3081 -130 -3035 -118
rect -3081 -856 -3075 -130
rect -3041 -856 -3035 -130
rect -3081 -868 -3035 -856
rect -23 -130 23 -118
rect -23 -856 -17 -130
rect 17 -856 23 -130
rect -23 -868 23 -856
rect 3035 -130 3081 -118
rect 3035 -856 3041 -130
rect 3075 -856 3081 -130
rect 3035 -868 3081 -856
rect -3025 -915 -33 -909
rect -3025 -949 -3013 -915
rect -45 -949 -33 -915
rect -3025 -955 -33 -949
rect 33 -915 3025 -909
rect 33 -949 45 -915
rect 3013 -949 3025 -915
rect 33 -955 3025 -949
<< properties >>
string FIXED_BBOX -3172 -1034 3172 1034
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.75 l 15.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
