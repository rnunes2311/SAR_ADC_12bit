magic
tech sky130A
magscale 1 2
timestamp 1717081718
<< nwell >>
rect 15679 1323 15712 2118
rect 15638 1203 16023 1323
rect 15679 1140 15909 1203
rect 15679 714 15930 1140
rect 20064 964 20329 1107
rect 15690 610 15930 714
rect 20024 870 20329 964
rect 20024 696 20328 870
rect 15900 560 15930 610
<< pwell >>
rect 19509 1204 20003 1304
rect 19509 1022 19996 1204
rect 19468 135 19846 340
rect 19468 84 20279 135
rect 19531 83 20279 84
<< psubdiff >>
rect 19545 1234 19569 1268
rect 19975 1234 19999 1268
rect 19554 96 19583 130
rect 20169 96 20198 130
<< nsubdiff >>
rect 20104 910 20194 940
rect 20104 690 20194 781
<< psubdiffcont >>
rect 19569 1234 19975 1268
rect 19583 96 20169 130
<< nsubdiffcont >>
rect 20104 781 20194 910
<< poly >>
rect 16106 1129 16442 1200
<< locali >>
rect 19553 1234 19569 1268
rect 19975 1234 19991 1268
rect 19590 964 19624 1002
rect 19899 967 19937 1001
rect 20084 910 20213 931
rect 20084 781 20104 910
rect 20194 781 20213 910
rect 20084 698 20213 781
rect 19623 685 20213 698
rect 19623 664 20179 685
rect 19566 358 19604 392
rect 19718 352 19892 402
rect 20220 352 20254 390
rect 16830 120 16900 160
rect 17994 120 18204 160
rect 19404 154 19444 160
rect 19404 153 19569 154
rect 19404 130 19597 153
rect 19404 127 19583 130
rect 19404 122 19558 127
rect 19404 120 19583 122
rect 19531 119 19583 120
rect 19537 96 19583 119
rect 20169 96 20237 122
<< viali >>
rect 12499 2049 15466 2083
rect 16100 1272 16500 1306
rect 19590 1002 19624 1038
rect 8643 301 8677 980
rect 15626 315 15660 994
rect 16553 307 16587 986
rect 19863 967 19899 1001
rect 19937 967 19973 1001
rect 19590 928 19624 964
rect 19530 358 19566 392
rect 19604 358 19640 392
rect 20220 390 20254 426
rect 20220 316 20254 352
rect 12508 120 15475 154
rect 16110 120 16510 154
rect 16900 120 17994 160
rect 18204 120 19404 160
<< metal1 >>
rect 8607 2083 15690 2120
rect 8607 2049 12499 2083
rect 15466 2049 15690 2083
rect 8607 2023 15690 2049
rect 8607 1868 8704 2023
rect 9980 1918 9990 1988
rect 10050 1918 10080 1988
rect 10140 1918 10150 1988
rect 11770 1918 11780 1988
rect 11840 1918 11870 1988
rect 11930 1918 11940 1988
rect 12950 1918 12960 1988
rect 13020 1918 13050 1988
rect 13110 1918 13120 1988
rect 15220 1928 15230 1988
rect 15290 1928 15330 1988
rect 15390 1928 15400 1988
rect 15591 1868 15690 2023
rect 8607 1439 15690 1868
rect 8607 980 8704 1439
rect 15591 1322 15690 1439
rect 15591 1306 16624 1322
rect 15591 1272 16100 1306
rect 16500 1272 16624 1306
rect 15591 1266 16624 1272
rect 15591 1225 16157 1266
rect 16470 1225 16624 1266
rect 8798 1130 15496 1178
rect 8798 1078 9995 1130
rect 10056 1078 10089 1130
rect 10150 1078 11775 1130
rect 11836 1078 11869 1130
rect 11930 1078 12955 1130
rect 13016 1078 13049 1130
rect 13110 1078 15225 1130
rect 15286 1078 15319 1130
rect 15380 1078 15496 1130
rect 8798 1016 15496 1078
rect 15591 1140 16003 1225
rect 16230 1193 16291 1203
rect 16189 1144 16230 1190
rect 8607 301 8643 980
rect 8677 864 8704 980
rect 15591 994 15690 1140
rect 15829 1038 15839 1099
rect 15891 1038 15901 1099
rect 15840 1005 15890 1038
rect 15591 864 15626 994
rect 8677 435 15626 864
rect 8677 301 8704 435
rect 8607 185 8704 301
rect 15591 315 15626 435
rect 15660 652 15690 994
rect 15829 944 15839 1005
rect 15891 944 15901 1005
rect 15660 474 15688 652
rect 15660 326 15748 474
rect 15840 350 15890 944
rect 15930 560 16003 1140
rect 16324 1193 16385 1203
rect 16291 1144 16324 1190
rect 16230 1131 16291 1141
rect 16385 1144 16428 1190
rect 16324 1131 16385 1141
rect 16527 986 16624 1225
rect 16141 696 16151 757
rect 16203 696 16213 757
rect 16333 696 16343 757
rect 16395 696 16405 757
rect 16141 602 16151 663
rect 16203 602 16213 663
rect 16333 602 16343 663
rect 16395 602 16405 663
rect 15932 552 16003 560
rect 15932 551 16104 552
rect 15932 490 16047 551
rect 16099 490 16109 551
rect 16229 490 16239 551
rect 16291 490 16301 551
rect 16421 490 16431 551
rect 16483 490 16493 551
rect 15932 457 16104 490
rect 15932 396 16047 457
rect 16099 396 16109 457
rect 16229 396 16239 457
rect 16291 396 16301 457
rect 16421 396 16431 457
rect 16483 396 16493 457
rect 15660 315 15688 326
rect 9993 278 10054 288
rect 8806 226 9993 262
rect 10087 278 10148 288
rect 10054 226 10087 262
rect 11765 278 11826 288
rect 10148 226 11765 262
rect 11859 278 11920 288
rect 11826 226 11859 262
rect 12945 278 13006 288
rect 11920 226 12945 262
rect 13039 278 13100 288
rect 13006 226 13039 262
rect 15221 276 15282 286
rect 13100 226 15221 262
rect 8806 224 15221 226
rect 15315 276 15376 286
rect 15282 224 15315 262
rect 15376 224 15496 262
rect 8806 216 15496 224
rect 15221 214 15282 216
rect 15315 214 15376 216
rect 15591 185 15688 315
rect 15723 265 15784 275
rect 15723 203 15784 213
rect 15817 265 15878 275
rect 15817 203 15878 213
rect 8607 167 15688 185
rect 15932 185 16003 396
rect 16527 307 16553 986
rect 16587 307 16624 986
rect 16527 185 16624 307
rect 15932 167 16624 185
rect 8607 154 16624 167
rect 8607 120 12508 154
rect 15475 120 16110 154
rect 16510 120 16624 154
rect 8607 88 16624 120
rect 16790 1306 20014 1388
rect 16790 185 16868 1306
rect 16986 1243 17396 1264
rect 16986 1191 17116 1243
rect 17177 1191 17210 1243
rect 17271 1191 17396 1243
rect 16986 1168 17396 1191
rect 17155 992 17165 1053
rect 17217 992 17227 1053
rect 17155 898 17165 959
rect 17217 898 17227 959
rect 16917 664 16927 725
rect 16979 664 16989 725
rect 17393 664 17403 725
rect 17455 664 17465 725
rect 16917 570 16927 631
rect 16979 570 16989 631
rect 17393 570 17403 631
rect 17455 570 17465 631
rect 17526 185 17614 1306
rect 17655 1243 17974 1264
rect 17655 1191 17785 1243
rect 17846 1191 17879 1243
rect 17940 1191 17974 1243
rect 17655 1162 17974 1191
rect 18040 1234 20014 1306
rect 18040 1050 18198 1234
rect 18312 1184 18467 1194
rect 18373 1132 18406 1184
rect 18312 1122 18467 1132
rect 17665 666 17675 727
rect 17727 666 17737 727
rect 17665 572 17675 633
rect 17727 572 17737 633
rect 17903 468 17913 529
rect 17965 468 17975 529
rect 17903 374 17913 435
rect 17965 374 17975 435
rect 18040 366 18278 1050
rect 18343 992 18353 1053
rect 18405 992 18415 1053
rect 18558 1050 18622 1234
rect 18343 898 18353 959
rect 18405 898 18415 959
rect 18040 185 18198 366
rect 18476 364 18622 1050
rect 18981 1004 19043 1234
rect 19149 1184 19304 1194
rect 19210 1132 19243 1184
rect 19149 1122 19304 1132
rect 19370 1004 19459 1234
rect 19566 1024 19576 1085
rect 19628 1024 19638 1085
rect 18773 828 18783 889
rect 18835 828 18845 889
rect 18773 734 18783 795
rect 18835 734 18845 795
rect 18669 575 18679 636
rect 18731 575 18741 636
rect 18867 575 18877 636
rect 18929 575 18939 636
rect 18669 481 18679 542
rect 18731 481 18741 542
rect 18867 481 18877 542
rect 18929 481 18939 542
rect 18558 185 18622 364
rect 18981 357 19125 1004
rect 19183 818 19193 879
rect 19245 818 19255 879
rect 19183 724 19193 785
rect 19245 724 19255 785
rect 18727 256 18788 266
rect 18727 194 18788 204
rect 18821 256 18882 266
rect 18821 194 18882 204
rect 16790 166 18622 185
rect 18981 185 19043 357
rect 19321 351 19459 1004
rect 19584 1002 19590 1024
rect 19624 1002 19630 1024
rect 19860 1012 19921 1022
rect 19584 991 19630 1002
rect 19566 930 19576 991
rect 19628 930 19638 991
rect 19851 961 19860 1007
rect 19954 1012 20015 1022
rect 19921 1001 19954 1007
rect 19921 967 19937 1001
rect 19921 961 19954 967
rect 19860 950 19921 960
rect 19954 950 20015 960
rect 19584 928 19590 930
rect 19624 928 19630 930
rect 19584 916 19630 928
rect 19603 644 19613 718
rect 20188 644 20198 718
rect 20215 438 20225 459
rect 20214 426 20225 438
rect 19527 404 19588 414
rect 19518 352 19527 398
rect 19621 404 19682 414
rect 19588 392 19621 398
rect 19588 358 19604 392
rect 19588 352 19621 358
rect 19370 185 19459 351
rect 19527 342 19588 352
rect 19621 342 19682 352
rect 20214 390 20220 426
rect 20277 398 20287 459
rect 20254 390 20260 398
rect 20214 365 20260 390
rect 20214 352 20225 365
rect 20214 316 20220 352
rect 20214 304 20225 316
rect 20277 304 20287 365
rect 18981 166 19581 185
rect 16790 160 19581 166
rect 16790 159 16900 160
rect 17994 159 18204 160
rect 19404 159 19581 160
rect 16790 99 16833 159
rect 19424 120 19581 159
rect 19598 120 19608 158
rect 19424 99 19608 120
rect 16790 96 19608 99
rect 20204 96 20214 158
rect 16790 89 19628 96
<< via1 >>
rect 9990 1918 10050 1988
rect 10080 1918 10140 1988
rect 11780 1918 11840 1988
rect 11870 1918 11930 1988
rect 12960 1918 13020 1988
rect 13050 1918 13110 1988
rect 15230 1928 15290 1988
rect 15330 1928 15390 1988
rect 9995 1078 10056 1130
rect 10089 1078 10150 1130
rect 11775 1078 11836 1130
rect 11869 1078 11930 1130
rect 12955 1078 13016 1130
rect 13049 1078 13110 1130
rect 15225 1078 15286 1130
rect 15319 1078 15380 1130
rect 15839 1038 15891 1099
rect 15839 944 15891 1005
rect 16230 1141 16291 1193
rect 16324 1141 16385 1193
rect 16151 696 16203 757
rect 16343 696 16395 757
rect 16151 602 16203 663
rect 16343 602 16395 663
rect 16047 490 16099 551
rect 16239 490 16291 551
rect 16431 490 16483 551
rect 16047 396 16099 457
rect 16239 396 16291 457
rect 16431 396 16483 457
rect 9993 226 10054 278
rect 10087 226 10148 278
rect 11765 226 11826 278
rect 11859 226 11920 278
rect 12945 226 13006 278
rect 13039 226 13100 278
rect 15221 224 15282 276
rect 15315 224 15376 276
rect 15723 213 15784 265
rect 15817 213 15878 265
rect 17116 1191 17177 1243
rect 17210 1191 17271 1243
rect 17165 992 17217 1053
rect 17165 898 17217 959
rect 16927 664 16979 725
rect 17403 664 17455 725
rect 16927 570 16979 631
rect 17403 570 17455 631
rect 17785 1191 17846 1243
rect 17879 1191 17940 1243
rect 18312 1132 18373 1184
rect 18406 1132 18467 1184
rect 17675 666 17727 727
rect 17675 572 17727 633
rect 17913 468 17965 529
rect 17913 374 17965 435
rect 18353 992 18405 1053
rect 18353 898 18405 959
rect 19149 1132 19210 1184
rect 19243 1132 19304 1184
rect 19576 1038 19628 1085
rect 19576 1024 19590 1038
rect 19590 1024 19624 1038
rect 19624 1024 19628 1038
rect 18783 828 18835 889
rect 18783 734 18835 795
rect 18679 575 18731 636
rect 18877 575 18929 636
rect 18679 481 18731 542
rect 18877 481 18929 542
rect 19193 818 19245 879
rect 19193 724 19245 785
rect 18727 204 18788 256
rect 18821 204 18882 256
rect 19576 964 19628 991
rect 19576 930 19590 964
rect 19590 930 19624 964
rect 19624 930 19628 964
rect 19860 1001 19921 1012
rect 19954 1001 20015 1012
rect 19860 967 19863 1001
rect 19863 967 19899 1001
rect 19899 967 19921 1001
rect 19954 967 19973 1001
rect 19973 967 20015 1001
rect 19860 960 19921 967
rect 19954 960 20015 967
rect 19613 644 20188 718
rect 20225 426 20277 459
rect 19527 392 19588 404
rect 19621 392 19682 404
rect 19527 358 19530 392
rect 19530 358 19566 392
rect 19566 358 19588 392
rect 19621 358 19640 392
rect 19640 358 19682 392
rect 19527 352 19588 358
rect 19621 352 19682 358
rect 20225 398 20254 426
rect 20254 398 20277 426
rect 20225 352 20277 365
rect 20225 316 20254 352
rect 20254 316 20277 352
rect 20225 304 20277 316
rect 16833 120 16900 159
rect 16900 120 17994 159
rect 17994 120 18204 159
rect 18204 120 19404 159
rect 19404 120 19424 159
rect 16833 99 19424 120
rect 19608 96 20204 158
<< metal2 >>
rect 9990 1988 10050 1998
rect 10080 1988 10140 1998
rect 10050 1918 10080 1958
rect 9990 1908 10140 1918
rect 11780 1988 11840 1998
rect 11870 1988 11930 1998
rect 11840 1918 11870 1958
rect 11780 1908 11930 1918
rect 12960 1988 13020 1998
rect 13050 1988 13110 1998
rect 13020 1918 13050 1968
rect 15230 1988 15390 1998
rect 15290 1928 15330 1988
rect 15230 1918 15390 1928
rect 12960 1908 13110 1918
rect 10020 1130 10120 1908
rect 11780 1130 11880 1908
rect 12970 1130 13070 1908
rect 15240 1130 15340 1918
rect 15618 1265 20198 1388
rect 15618 1212 16157 1265
rect 16470 1243 20198 1265
rect 16470 1212 17116 1243
rect 9985 1078 9995 1130
rect 10056 1078 10089 1130
rect 10150 1078 10160 1130
rect 11765 1078 11775 1130
rect 11836 1078 11869 1130
rect 11930 1078 11940 1130
rect 12945 1078 12955 1130
rect 13016 1078 13049 1130
rect 13110 1078 13120 1130
rect 15215 1078 15225 1130
rect 15286 1078 15319 1130
rect 15380 1078 15390 1130
rect 15850 1109 15880 1212
rect 16194 1141 16230 1193
rect 16291 1141 16324 1193
rect 16385 1170 16395 1193
rect 17106 1191 17116 1212
rect 17177 1191 17210 1243
rect 17271 1212 17785 1243
rect 17271 1191 17281 1212
rect 17775 1191 17785 1212
rect 17846 1191 17879 1243
rect 17940 1212 20198 1243
rect 17940 1191 17950 1212
rect 19798 1187 19998 1212
rect 16385 1141 16946 1170
rect 16194 1133 16946 1141
rect 18264 1133 18312 1184
rect 16194 1132 18312 1133
rect 18373 1132 18406 1184
rect 18467 1170 18477 1184
rect 19139 1170 19149 1184
rect 18467 1132 19149 1170
rect 19210 1132 19243 1184
rect 19304 1170 19314 1184
rect 19304 1132 19614 1170
rect 16194 1130 19614 1132
rect 15839 1099 15891 1109
rect 10020 278 10120 1078
rect 11780 278 11880 1078
rect 12970 278 13070 1078
rect 15240 850 15340 1078
rect 16897 1093 18312 1130
rect 19584 1095 19614 1130
rect 19576 1085 19628 1095
rect 15839 1005 15891 1038
rect 15839 934 15891 944
rect 17165 1053 17217 1063
rect 18353 1053 18405 1063
rect 17217 992 18353 1004
rect 17165 959 18405 992
rect 17217 956 18353 959
rect 17165 888 17217 898
rect 19576 991 19628 1024
rect 19576 920 19628 930
rect 19849 1012 20049 1078
rect 19849 960 19860 1012
rect 19921 960 19954 1012
rect 20015 960 20049 1012
rect 18353 888 18405 898
rect 18783 889 18835 899
rect 15240 828 18783 850
rect 19193 879 19245 889
rect 18835 828 19193 850
rect 15240 818 19193 828
rect 19849 878 20049 960
rect 15240 800 19245 818
rect 9983 226 9993 278
rect 10054 226 10087 278
rect 10148 226 10158 278
rect 11755 226 11765 278
rect 11826 226 11859 278
rect 11920 226 11930 278
rect 12935 226 12945 278
rect 13006 226 13039 278
rect 13100 226 13110 278
rect 15240 276 15340 800
rect 18783 795 18835 800
rect 16151 757 16203 767
rect 16343 757 16395 767
rect 16203 696 16343 700
rect 16840 725 17040 740
rect 16840 700 16927 725
rect 16395 696 16927 700
rect 16151 686 16927 696
rect 15936 664 16927 686
rect 16979 700 17040 725
rect 17403 725 17455 735
rect 16979 664 17403 700
rect 17675 727 17727 737
rect 17455 666 17675 700
rect 18783 724 18835 734
rect 19193 785 19245 800
rect 20106 728 20197 1212
rect 19193 714 19245 724
rect 19613 718 20197 728
rect 17455 664 17727 666
rect 15936 663 17727 664
rect 15936 654 16151 663
rect 15211 224 15221 276
rect 15282 224 15315 276
rect 15376 224 15386 276
rect 15713 213 15723 265
rect 15784 213 15817 265
rect 15878 257 15888 265
rect 15936 257 15968 654
rect 16203 648 16343 663
rect 16151 592 16203 602
rect 16395 648 17727 663
rect 16343 592 16395 602
rect 16840 631 17040 648
rect 16840 570 16927 631
rect 16979 570 17040 631
rect 16047 551 16099 561
rect 16239 551 16291 561
rect 16099 490 16239 494
rect 16431 551 16483 561
rect 16291 490 16431 494
rect 16840 540 17040 570
rect 17403 631 17455 648
rect 17403 560 17455 570
rect 17675 633 17727 648
rect 18708 646 18908 660
rect 17675 562 17727 572
rect 18679 636 18929 646
rect 18731 575 18877 636
rect 20188 644 20197 718
rect 19613 634 20197 644
rect 18679 542 18929 575
rect 16047 457 16483 490
rect 16099 442 16239 457
rect 16047 386 16099 396
rect 16291 442 16431 457
rect 16239 386 16291 396
rect 16431 386 16483 396
rect 17913 529 17965 539
rect 18731 481 18877 542
rect 18679 471 18929 481
rect 17913 435 17965 468
rect 18708 460 18908 471
rect 20143 459 20343 479
rect 17965 374 19527 404
rect 17913 364 19527 374
rect 17914 352 19527 364
rect 19588 352 19621 404
rect 19682 352 19692 404
rect 20143 398 20225 459
rect 20277 398 20343 459
rect 20143 365 20343 398
rect 15878 256 18717 257
rect 15878 225 18727 256
rect 15878 213 15888 225
rect 18717 204 18727 225
rect 18788 204 18821 256
rect 18882 204 18892 256
rect 19831 170 20031 347
rect 20143 304 20225 365
rect 20277 304 20343 365
rect 20143 279 20343 304
rect 16787 159 20290 170
rect 16787 99 16833 159
rect 19424 158 20290 159
rect 19424 99 19608 158
rect 16787 96 19608 99
rect 20204 96 20290 158
rect 16787 77 20290 96
use sky130_fd_pr__pfet_01v8_CMU2ES  sky130_fd_pr__pfet_01v8_CMU2ES_0
timestamp 1717081077
transform 1 0 12151 0 1 1101
box -3545 -1017 3545 1017
use sky130_fd_pr__pfet_01v8_XG6TDL  sky130_fd_pr__pfet_01v8_XG6TDL_0
timestamp 1710675123
transform 1 0 16265 0 1 703
box -359 -619 359 619
use sky130_fd_sc_hd__inv_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 20014 0 -1 1225
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19554 0 1 137
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x3
timestamp 1710522493
transform 1 0 19830 0 1 137
box -38 -48 498 592
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1710675955
transform 1 0 15801 0 1 403
box -211 -319 211 319
use sky130_fd_pr__nfet_05v0_nvt_F93ZEE  XM3
timestamp 1715417500
transform 1 0 17191 0 1 730
box -437 -658 441 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM4
timestamp 1710677421
transform 1 0 18383 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_01v8_6EHS5V  XM5
timestamp 1710677421
transform 1 0 19223 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_05v0_nvt_JFFQEL  XM7
timestamp 1710675123
transform 1 0 17820 0 1 730
box -318 -658 318 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM8
timestamp 1710677421
transform 1 0 18803 0 -1 694
box -263 -610 263 610
<< labels >>
flabel metal2 16840 540 17040 740 0 FreeSans 256 0 0 0 VGATE
port 5 nsew
flabel metal2 17806 968 17830 982 0 FreeSans 800 0 0 0 Vd
flabel metal2 18620 360 18650 390 0 FreeSans 800 0 0 0 VGATE_1V8
flabel metal2 18978 810 19010 829 0 FreeSans 800 0 0 0 Vbottom
flabel metal2 19071 1141 19097 1157 0 FreeSans 800 0 0 0 EN_Z
flabel metal2 18708 460 18908 660 0 FreeSans 256 0 0 0 VIN
port 2 nsew
flabel metal2 19849 878 20049 1078 0 FreeSans 256 0 0 0 EN
port 4 nsew
flabel metal2 20143 279 20343 479 0 FreeSans 256 0 0 0 SW_ON
port 3 nsew
flabel metal2 19831 147 20031 347 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal2 19798 1187 19998 1387 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 11069 1604 11129 1664 0 FreeSans 800 0 0 0 Vtop
flabel metal2 16238 666 16278 688 0 FreeSans 800 0 0 0 Vgate
flabel metal1 11070 600 11130 660 0 FreeSans 800 0 0 0 Vtop
flabel metal2 15707 1286 15763 1337 0 FreeSans 800 0 0 0 VDD
<< end >>
