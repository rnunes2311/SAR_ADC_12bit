* SPICE3 file created from CDAC_mim_12bit_flat.ext - technology: sky130A
* Empty netlist for LVS

.subckt CDAC_12bit C0_dummy C0 C1 C2 C3 C4 C5 C6 C7 C8 C9 C10 Ctop VSS
.ends
