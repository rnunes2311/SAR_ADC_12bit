magic
tech sky130A
magscale 1 2
timestamp 1711964565
<< nwell >>
rect -1742 -1019 1742 1019
<< pmos >>
rect -1546 -800 -1446 800
rect -1274 -800 -1174 800
rect -1002 -800 -902 800
rect -730 -800 -630 800
rect -458 -800 -358 800
rect -186 -800 -86 800
rect 86 -800 186 800
rect 358 -800 458 800
rect 630 -800 730 800
rect 902 -800 1002 800
rect 1174 -800 1274 800
rect 1446 -800 1546 800
<< pdiff >>
rect -1604 788 -1546 800
rect -1604 -788 -1592 788
rect -1558 -788 -1546 788
rect -1604 -800 -1546 -788
rect -1446 788 -1388 800
rect -1446 -788 -1434 788
rect -1400 -788 -1388 788
rect -1446 -800 -1388 -788
rect -1332 788 -1274 800
rect -1332 -788 -1320 788
rect -1286 -788 -1274 788
rect -1332 -800 -1274 -788
rect -1174 788 -1116 800
rect -1174 -788 -1162 788
rect -1128 -788 -1116 788
rect -1174 -800 -1116 -788
rect -1060 788 -1002 800
rect -1060 -788 -1048 788
rect -1014 -788 -1002 788
rect -1060 -800 -1002 -788
rect -902 788 -844 800
rect -902 -788 -890 788
rect -856 -788 -844 788
rect -902 -800 -844 -788
rect -788 788 -730 800
rect -788 -788 -776 788
rect -742 -788 -730 788
rect -788 -800 -730 -788
rect -630 788 -572 800
rect -630 -788 -618 788
rect -584 -788 -572 788
rect -630 -800 -572 -788
rect -516 788 -458 800
rect -516 -788 -504 788
rect -470 -788 -458 788
rect -516 -800 -458 -788
rect -358 788 -300 800
rect -358 -788 -346 788
rect -312 -788 -300 788
rect -358 -800 -300 -788
rect -244 788 -186 800
rect -244 -788 -232 788
rect -198 -788 -186 788
rect -244 -800 -186 -788
rect -86 788 -28 800
rect -86 -788 -74 788
rect -40 -788 -28 788
rect -86 -800 -28 -788
rect 28 788 86 800
rect 28 -788 40 788
rect 74 -788 86 788
rect 28 -800 86 -788
rect 186 788 244 800
rect 186 -788 198 788
rect 232 -788 244 788
rect 186 -800 244 -788
rect 300 788 358 800
rect 300 -788 312 788
rect 346 -788 358 788
rect 300 -800 358 -788
rect 458 788 516 800
rect 458 -788 470 788
rect 504 -788 516 788
rect 458 -800 516 -788
rect 572 788 630 800
rect 572 -788 584 788
rect 618 -788 630 788
rect 572 -800 630 -788
rect 730 788 788 800
rect 730 -788 742 788
rect 776 -788 788 788
rect 730 -800 788 -788
rect 844 788 902 800
rect 844 -788 856 788
rect 890 -788 902 788
rect 844 -800 902 -788
rect 1002 788 1060 800
rect 1002 -788 1014 788
rect 1048 -788 1060 788
rect 1002 -800 1060 -788
rect 1116 788 1174 800
rect 1116 -788 1128 788
rect 1162 -788 1174 788
rect 1116 -800 1174 -788
rect 1274 788 1332 800
rect 1274 -788 1286 788
rect 1320 -788 1332 788
rect 1274 -800 1332 -788
rect 1388 788 1446 800
rect 1388 -788 1400 788
rect 1434 -788 1446 788
rect 1388 -800 1446 -788
rect 1546 788 1604 800
rect 1546 -788 1558 788
rect 1592 -788 1604 788
rect 1546 -800 1604 -788
<< pdiffc >>
rect -1592 -788 -1558 788
rect -1434 -788 -1400 788
rect -1320 -788 -1286 788
rect -1162 -788 -1128 788
rect -1048 -788 -1014 788
rect -890 -788 -856 788
rect -776 -788 -742 788
rect -618 -788 -584 788
rect -504 -788 -470 788
rect -346 -788 -312 788
rect -232 -788 -198 788
rect -74 -788 -40 788
rect 40 -788 74 788
rect 198 -788 232 788
rect 312 -788 346 788
rect 470 -788 504 788
rect 584 -788 618 788
rect 742 -788 776 788
rect 856 -788 890 788
rect 1014 -788 1048 788
rect 1128 -788 1162 788
rect 1286 -788 1320 788
rect 1400 -788 1434 788
rect 1558 -788 1592 788
<< nsubdiff >>
rect -1706 949 -1610 983
rect 1610 949 1706 983
rect -1706 887 -1672 949
rect 1672 887 1706 949
rect -1706 -949 -1672 -887
rect 1672 -949 1706 -887
rect -1706 -983 -1610 -949
rect 1610 -983 1706 -949
<< nsubdiffcont >>
rect -1610 949 1610 983
rect -1706 -887 -1672 887
rect 1672 -887 1706 887
rect -1610 -983 1610 -949
<< poly >>
rect -1546 881 -1446 897
rect -1546 847 -1530 881
rect -1462 847 -1446 881
rect -1546 800 -1446 847
rect -1274 881 -1174 897
rect -1274 847 -1258 881
rect -1190 847 -1174 881
rect -1274 800 -1174 847
rect -1002 881 -902 897
rect -1002 847 -986 881
rect -918 847 -902 881
rect -1002 800 -902 847
rect -730 881 -630 897
rect -730 847 -714 881
rect -646 847 -630 881
rect -730 800 -630 847
rect -458 881 -358 897
rect -458 847 -442 881
rect -374 847 -358 881
rect -458 800 -358 847
rect -186 881 -86 897
rect -186 847 -170 881
rect -102 847 -86 881
rect -186 800 -86 847
rect 86 881 186 897
rect 86 847 102 881
rect 170 847 186 881
rect 86 800 186 847
rect 358 881 458 897
rect 358 847 374 881
rect 442 847 458 881
rect 358 800 458 847
rect 630 881 730 897
rect 630 847 646 881
rect 714 847 730 881
rect 630 800 730 847
rect 902 881 1002 897
rect 902 847 918 881
rect 986 847 1002 881
rect 902 800 1002 847
rect 1174 881 1274 897
rect 1174 847 1190 881
rect 1258 847 1274 881
rect 1174 800 1274 847
rect 1446 881 1546 897
rect 1446 847 1462 881
rect 1530 847 1546 881
rect 1446 800 1546 847
rect -1546 -847 -1446 -800
rect -1546 -881 -1530 -847
rect -1462 -881 -1446 -847
rect -1546 -897 -1446 -881
rect -1274 -847 -1174 -800
rect -1274 -881 -1258 -847
rect -1190 -881 -1174 -847
rect -1274 -897 -1174 -881
rect -1002 -847 -902 -800
rect -1002 -881 -986 -847
rect -918 -881 -902 -847
rect -1002 -897 -902 -881
rect -730 -847 -630 -800
rect -730 -881 -714 -847
rect -646 -881 -630 -847
rect -730 -897 -630 -881
rect -458 -847 -358 -800
rect -458 -881 -442 -847
rect -374 -881 -358 -847
rect -458 -897 -358 -881
rect -186 -847 -86 -800
rect -186 -881 -170 -847
rect -102 -881 -86 -847
rect -186 -897 -86 -881
rect 86 -847 186 -800
rect 86 -881 102 -847
rect 170 -881 186 -847
rect 86 -897 186 -881
rect 358 -847 458 -800
rect 358 -881 374 -847
rect 442 -881 458 -847
rect 358 -897 458 -881
rect 630 -847 730 -800
rect 630 -881 646 -847
rect 714 -881 730 -847
rect 630 -897 730 -881
rect 902 -847 1002 -800
rect 902 -881 918 -847
rect 986 -881 1002 -847
rect 902 -897 1002 -881
rect 1174 -847 1274 -800
rect 1174 -881 1190 -847
rect 1258 -881 1274 -847
rect 1174 -897 1274 -881
rect 1446 -847 1546 -800
rect 1446 -881 1462 -847
rect 1530 -881 1546 -847
rect 1446 -897 1546 -881
<< polycont >>
rect -1530 847 -1462 881
rect -1258 847 -1190 881
rect -986 847 -918 881
rect -714 847 -646 881
rect -442 847 -374 881
rect -170 847 -102 881
rect 102 847 170 881
rect 374 847 442 881
rect 646 847 714 881
rect 918 847 986 881
rect 1190 847 1258 881
rect 1462 847 1530 881
rect -1530 -881 -1462 -847
rect -1258 -881 -1190 -847
rect -986 -881 -918 -847
rect -714 -881 -646 -847
rect -442 -881 -374 -847
rect -170 -881 -102 -847
rect 102 -881 170 -847
rect 374 -881 442 -847
rect 646 -881 714 -847
rect 918 -881 986 -847
rect 1190 -881 1258 -847
rect 1462 -881 1530 -847
<< locali >>
rect -1706 949 -1610 983
rect 1610 949 1706 983
rect -1706 887 -1672 949
rect 1672 887 1706 949
rect -1546 847 -1530 881
rect -1462 847 -1446 881
rect -1274 847 -1258 881
rect -1190 847 -1174 881
rect -1002 847 -986 881
rect -918 847 -902 881
rect -730 847 -714 881
rect -646 847 -630 881
rect -458 847 -442 881
rect -374 847 -358 881
rect -186 847 -170 881
rect -102 847 -86 881
rect 86 847 102 881
rect 170 847 186 881
rect 358 847 374 881
rect 442 847 458 881
rect 630 847 646 881
rect 714 847 730 881
rect 902 847 918 881
rect 986 847 1002 881
rect 1174 847 1190 881
rect 1258 847 1274 881
rect 1446 847 1462 881
rect 1530 847 1546 881
rect -1592 788 -1558 804
rect -1592 -804 -1558 -788
rect -1434 788 -1400 804
rect -1434 -804 -1400 -788
rect -1320 788 -1286 804
rect -1320 -804 -1286 -788
rect -1162 788 -1128 804
rect -1162 -804 -1128 -788
rect -1048 788 -1014 804
rect -1048 -804 -1014 -788
rect -890 788 -856 804
rect -890 -804 -856 -788
rect -776 788 -742 804
rect -776 -804 -742 -788
rect -618 788 -584 804
rect -618 -804 -584 -788
rect -504 788 -470 804
rect -504 -804 -470 -788
rect -346 788 -312 804
rect -346 -804 -312 -788
rect -232 788 -198 804
rect -232 -804 -198 -788
rect -74 788 -40 804
rect -74 -804 -40 -788
rect 40 788 74 804
rect 40 -804 74 -788
rect 198 788 232 804
rect 198 -804 232 -788
rect 312 788 346 804
rect 312 -804 346 -788
rect 470 788 504 804
rect 470 -804 504 -788
rect 584 788 618 804
rect 584 -804 618 -788
rect 742 788 776 804
rect 742 -804 776 -788
rect 856 788 890 804
rect 856 -804 890 -788
rect 1014 788 1048 804
rect 1014 -804 1048 -788
rect 1128 788 1162 804
rect 1128 -804 1162 -788
rect 1286 788 1320 804
rect 1286 -804 1320 -788
rect 1400 788 1434 804
rect 1400 -804 1434 -788
rect 1558 788 1592 804
rect 1558 -804 1592 -788
rect -1546 -881 -1530 -847
rect -1462 -881 -1446 -847
rect -1274 -881 -1258 -847
rect -1190 -881 -1174 -847
rect -1002 -881 -986 -847
rect -918 -881 -902 -847
rect -730 -881 -714 -847
rect -646 -881 -630 -847
rect -458 -881 -442 -847
rect -374 -881 -358 -847
rect -186 -881 -170 -847
rect -102 -881 -86 -847
rect 86 -881 102 -847
rect 170 -881 186 -847
rect 358 -881 374 -847
rect 442 -881 458 -847
rect 630 -881 646 -847
rect 714 -881 730 -847
rect 902 -881 918 -847
rect 986 -881 1002 -847
rect 1174 -881 1190 -847
rect 1258 -881 1274 -847
rect 1446 -881 1462 -847
rect 1530 -881 1546 -847
rect -1706 -949 -1672 -887
rect 1672 -949 1706 -887
rect -1706 -983 -1610 -949
rect 1610 -983 1706 -949
<< viali >>
rect -1530 847 -1462 881
rect -1258 847 -1190 881
rect -986 847 -918 881
rect -714 847 -646 881
rect -442 847 -374 881
rect -170 847 -102 881
rect 102 847 170 881
rect 374 847 442 881
rect 646 847 714 881
rect 918 847 986 881
rect 1190 847 1258 881
rect 1462 847 1530 881
rect -1592 -788 -1558 788
rect -1434 -788 -1400 788
rect -1320 -788 -1286 788
rect -1162 -788 -1128 788
rect -1048 -788 -1014 788
rect -890 -788 -856 788
rect -776 -788 -742 788
rect -618 -788 -584 788
rect -504 -788 -470 788
rect -346 -788 -312 788
rect -232 -788 -198 788
rect -74 -788 -40 788
rect 40 -788 74 788
rect 198 -788 232 788
rect 312 -788 346 788
rect 470 -788 504 788
rect 584 -788 618 788
rect 742 -788 776 788
rect 856 -788 890 788
rect 1014 -788 1048 788
rect 1128 -788 1162 788
rect 1286 -788 1320 788
rect 1400 -788 1434 788
rect 1558 -788 1592 788
rect -1530 -881 -1462 -847
rect -1258 -881 -1190 -847
rect -986 -881 -918 -847
rect -714 -881 -646 -847
rect -442 -881 -374 -847
rect -170 -881 -102 -847
rect 102 -881 170 -847
rect 374 -881 442 -847
rect 646 -881 714 -847
rect 918 -881 986 -847
rect 1190 -881 1258 -847
rect 1462 -881 1530 -847
<< metal1 >>
rect -1542 881 -1450 887
rect -1542 847 -1530 881
rect -1462 847 -1450 881
rect -1542 841 -1450 847
rect -1270 881 -1178 887
rect -1270 847 -1258 881
rect -1190 847 -1178 881
rect -1270 841 -1178 847
rect -998 881 -906 887
rect -998 847 -986 881
rect -918 847 -906 881
rect -998 841 -906 847
rect -726 881 -634 887
rect -726 847 -714 881
rect -646 847 -634 881
rect -726 841 -634 847
rect -454 881 -362 887
rect -454 847 -442 881
rect -374 847 -362 881
rect -454 841 -362 847
rect -182 881 -90 887
rect -182 847 -170 881
rect -102 847 -90 881
rect -182 841 -90 847
rect 90 881 182 887
rect 90 847 102 881
rect 170 847 182 881
rect 90 841 182 847
rect 362 881 454 887
rect 362 847 374 881
rect 442 847 454 881
rect 362 841 454 847
rect 634 881 726 887
rect 634 847 646 881
rect 714 847 726 881
rect 634 841 726 847
rect 906 881 998 887
rect 906 847 918 881
rect 986 847 998 881
rect 906 841 998 847
rect 1178 881 1270 887
rect 1178 847 1190 881
rect 1258 847 1270 881
rect 1178 841 1270 847
rect 1450 881 1542 887
rect 1450 847 1462 881
rect 1530 847 1542 881
rect 1450 841 1542 847
rect -1598 788 -1552 800
rect -1598 -788 -1592 788
rect -1558 -788 -1552 788
rect -1598 -800 -1552 -788
rect -1440 788 -1394 800
rect -1440 -788 -1434 788
rect -1400 -788 -1394 788
rect -1440 -800 -1394 -788
rect -1326 788 -1280 800
rect -1326 -788 -1320 788
rect -1286 -788 -1280 788
rect -1326 -800 -1280 -788
rect -1168 788 -1122 800
rect -1168 -788 -1162 788
rect -1128 -788 -1122 788
rect -1168 -800 -1122 -788
rect -1054 788 -1008 800
rect -1054 -788 -1048 788
rect -1014 -788 -1008 788
rect -1054 -800 -1008 -788
rect -896 788 -850 800
rect -896 -788 -890 788
rect -856 -788 -850 788
rect -896 -800 -850 -788
rect -782 788 -736 800
rect -782 -788 -776 788
rect -742 -788 -736 788
rect -782 -800 -736 -788
rect -624 788 -578 800
rect -624 -788 -618 788
rect -584 -788 -578 788
rect -624 -800 -578 -788
rect -510 788 -464 800
rect -510 -788 -504 788
rect -470 -788 -464 788
rect -510 -800 -464 -788
rect -352 788 -306 800
rect -352 -788 -346 788
rect -312 -788 -306 788
rect -352 -800 -306 -788
rect -238 788 -192 800
rect -238 -788 -232 788
rect -198 -788 -192 788
rect -238 -800 -192 -788
rect -80 788 -34 800
rect -80 -788 -74 788
rect -40 -788 -34 788
rect -80 -800 -34 -788
rect 34 788 80 800
rect 34 -788 40 788
rect 74 -788 80 788
rect 34 -800 80 -788
rect 192 788 238 800
rect 192 -788 198 788
rect 232 -788 238 788
rect 192 -800 238 -788
rect 306 788 352 800
rect 306 -788 312 788
rect 346 -788 352 788
rect 306 -800 352 -788
rect 464 788 510 800
rect 464 -788 470 788
rect 504 -788 510 788
rect 464 -800 510 -788
rect 578 788 624 800
rect 578 -788 584 788
rect 618 -788 624 788
rect 578 -800 624 -788
rect 736 788 782 800
rect 736 -788 742 788
rect 776 -788 782 788
rect 736 -800 782 -788
rect 850 788 896 800
rect 850 -788 856 788
rect 890 -788 896 788
rect 850 -800 896 -788
rect 1008 788 1054 800
rect 1008 -788 1014 788
rect 1048 -788 1054 788
rect 1008 -800 1054 -788
rect 1122 788 1168 800
rect 1122 -788 1128 788
rect 1162 -788 1168 788
rect 1122 -800 1168 -788
rect 1280 788 1326 800
rect 1280 -788 1286 788
rect 1320 -788 1326 788
rect 1280 -800 1326 -788
rect 1394 788 1440 800
rect 1394 -788 1400 788
rect 1434 -788 1440 788
rect 1394 -800 1440 -788
rect 1552 788 1598 800
rect 1552 -788 1558 788
rect 1592 -788 1598 788
rect 1552 -800 1598 -788
rect -1542 -847 -1450 -841
rect -1542 -881 -1530 -847
rect -1462 -881 -1450 -847
rect -1542 -887 -1450 -881
rect -1270 -847 -1178 -841
rect -1270 -881 -1258 -847
rect -1190 -881 -1178 -847
rect -1270 -887 -1178 -881
rect -998 -847 -906 -841
rect -998 -881 -986 -847
rect -918 -881 -906 -847
rect -998 -887 -906 -881
rect -726 -847 -634 -841
rect -726 -881 -714 -847
rect -646 -881 -634 -847
rect -726 -887 -634 -881
rect -454 -847 -362 -841
rect -454 -881 -442 -847
rect -374 -881 -362 -847
rect -454 -887 -362 -881
rect -182 -847 -90 -841
rect -182 -881 -170 -847
rect -102 -881 -90 -847
rect -182 -887 -90 -881
rect 90 -847 182 -841
rect 90 -881 102 -847
rect 170 -881 182 -847
rect 90 -887 182 -881
rect 362 -847 454 -841
rect 362 -881 374 -847
rect 442 -881 454 -847
rect 362 -887 454 -881
rect 634 -847 726 -841
rect 634 -881 646 -847
rect 714 -881 726 -847
rect 634 -887 726 -881
rect 906 -847 998 -841
rect 906 -881 918 -847
rect 986 -881 998 -847
rect 906 -887 998 -881
rect 1178 -847 1270 -841
rect 1178 -881 1190 -847
rect 1258 -881 1270 -847
rect 1178 -887 1270 -881
rect 1450 -847 1542 -841
rect 1450 -881 1462 -847
rect 1530 -881 1542 -847
rect 1450 -887 1542 -881
<< properties >>
string FIXED_BBOX -1689 -966 1689 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
