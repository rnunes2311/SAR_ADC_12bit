magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< error_p >>
rect -29 881 29 887
rect -29 847 -17 881
rect -29 841 29 847
rect -29 -847 29 -841
rect -29 -881 -17 -847
rect -29 -887 29 -881
<< nwell >>
rect -211 -1019 211 1019
<< pmoshvt >>
rect -15 -800 15 800
<< pdiff >>
rect -73 788 -15 800
rect -73 -788 -61 788
rect -27 -788 -15 788
rect -73 -800 -15 -788
rect 15 788 73 800
rect 15 -788 27 788
rect 61 -788 73 788
rect 15 -800 73 -788
<< pdiffc >>
rect -61 -788 -27 788
rect 27 -788 61 788
<< nsubdiff >>
rect -175 949 -79 983
rect 79 949 175 983
rect -175 887 -141 949
rect 141 887 175 949
rect -175 -949 -141 -887
rect 141 -949 175 -887
rect -175 -983 -79 -949
rect 79 -983 175 -949
<< nsubdiffcont >>
rect -79 949 79 983
rect -175 -887 -141 887
rect 141 -887 175 887
rect -79 -983 79 -949
<< poly >>
rect -33 881 33 897
rect -33 847 -17 881
rect 17 847 33 881
rect -33 831 33 847
rect -15 800 15 831
rect -15 -831 15 -800
rect -33 -847 33 -831
rect -33 -881 -17 -847
rect 17 -881 33 -847
rect -33 -897 33 -881
<< polycont >>
rect -17 847 17 881
rect -17 -881 17 -847
<< locali >>
rect -175 949 -79 983
rect 79 949 175 983
rect -175 887 -141 949
rect 141 887 175 949
rect -33 847 -17 881
rect 17 847 33 881
rect -61 788 -27 804
rect -61 -804 -27 -788
rect 27 788 61 804
rect 27 -804 61 -788
rect -33 -881 -17 -847
rect 17 -881 33 -847
rect -175 -949 -141 -887
rect 141 -949 175 -887
rect -175 -983 -79 -949
rect 79 -983 175 -949
<< viali >>
rect -17 847 17 881
rect -61 -788 -27 788
rect 27 -788 61 788
rect -17 -881 17 -847
<< metal1 >>
rect -29 881 29 887
rect -29 847 -17 881
rect 17 847 29 881
rect -29 841 29 847
rect -67 788 -21 800
rect -67 -788 -61 788
rect -27 -788 -21 788
rect -67 -800 -21 -788
rect 21 788 67 800
rect 21 -788 27 788
rect 61 -788 67 788
rect 21 -800 67 -788
rect -29 -847 29 -841
rect -29 -881 -17 -847
rect 17 -881 29 -847
rect -29 -887 29 -881
<< properties >>
string FIXED_BBOX -158 -966 158 966
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 8.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
