magic
tech sky130A
magscale 1 2
timestamp 1715417773
<< metal1 >>
rect -645 27755 -615 30892
rect -585 27845 -555 30892
rect -525 27935 -495 30892
rect -465 28025 -435 30892
rect -405 28115 -375 30892
rect -345 28205 -315 30892
rect -285 28295 -255 30892
rect -225 28475 -195 30892
rect -165 28565 -135 30892
rect -105 28655 -75 30892
rect -45 28745 -15 30892
rect 15 28835 45 30892
rect 75 28925 105 30892
rect 135 29015 165 30892
rect 195 29105 225 30892
rect 255 29195 285 30892
rect 315 29285 345 30892
rect 375 29375 405 30892
rect 435 29465 465 30892
rect 495 29555 525 30892
rect 555 29645 585 30892
rect 615 29760 645 30892
rect 705 30810 735 30892
rect 680 30750 690 30810
rect 750 30750 760 30810
rect 2585 30165 2900 30195
rect 615 29750 675 29760
rect 615 29690 620 29750
rect 615 29680 675 29690
rect 2345 29660 2405 29670
rect 555 29615 2345 29645
rect 2345 29590 2405 29600
rect 3350 29555 3360 29570
rect 495 29525 3360 29555
rect 3350 29510 3360 29525
rect 3420 29510 3430 29570
rect 3870 29465 3880 29480
rect 435 29435 3880 29465
rect 3870 29420 3880 29435
rect 3940 29420 3950 29480
rect 4120 29375 4130 29390
rect 375 29345 4130 29375
rect 4120 29330 4130 29345
rect 4190 29330 4200 29390
rect 4360 29285 4370 29300
rect 315 29255 4370 29285
rect 4360 29240 4370 29255
rect 4430 29240 4440 29300
rect 4610 29195 4620 29210
rect 255 29165 4620 29195
rect 4610 29150 4620 29165
rect 4680 29150 4690 29210
rect 4850 29105 4860 29120
rect 195 29075 4860 29105
rect 4850 29060 4860 29075
rect 4920 29060 4930 29120
rect 5090 29015 5100 29030
rect 135 28985 5100 29015
rect 5090 28970 5100 28985
rect 5160 28970 5170 29030
rect 5340 28925 5350 28940
rect 75 28895 5350 28925
rect 5340 28880 5350 28895
rect 5410 28880 5420 28940
rect 5570 28835 5580 28850
rect 15 28805 5580 28835
rect 5570 28790 5580 28805
rect 5640 28790 5650 28850
rect 8090 28790 8100 28850
rect 8160 28835 8170 28850
rect 8160 28805 15040 28835
rect 8160 28790 8170 28805
rect 6120 28745 6130 28760
rect -45 28715 6130 28745
rect 6120 28700 6130 28715
rect 6190 28700 6200 28760
rect 8860 28700 8870 28760
rect 8930 28745 8940 28760
rect 8930 28715 15040 28745
rect 8930 28700 8940 28715
rect 6890 28655 6900 28670
rect -105 28625 6900 28655
rect 6890 28610 6900 28625
rect 6960 28610 6970 28670
rect 9630 28610 9640 28670
rect 9700 28655 9710 28670
rect 9700 28625 15040 28655
rect 9700 28610 9710 28625
rect 7280 28565 7290 28580
rect -165 28535 7290 28565
rect 7280 28520 7290 28535
rect 7350 28520 7360 28580
rect 10010 28520 10020 28580
rect 10080 28565 10090 28580
rect 10080 28535 15040 28565
rect 10080 28520 10090 28535
rect 7450 28475 7460 28490
rect -225 28445 7460 28475
rect 7450 28430 7460 28445
rect 7520 28430 7530 28490
rect 10200 28430 10210 28490
rect 10270 28475 10280 28490
rect 10270 28445 15040 28475
rect 10270 28430 10280 28445
rect 5834 28340 5844 28400
rect 5904 28385 5914 28400
rect 7670 28385 7680 28400
rect 5904 28355 7680 28385
rect 5904 28340 5914 28355
rect 7670 28340 7680 28355
rect 7740 28340 7750 28400
rect 11690 28340 11700 28400
rect 11760 28385 11770 28400
rect 11760 28355 15040 28385
rect 11760 28340 11770 28355
rect 10410 28295 10420 28310
rect -285 28265 10420 28295
rect 10410 28250 10420 28265
rect 10480 28250 10490 28310
rect 11850 28250 11860 28310
rect 11920 28295 11930 28310
rect 11920 28265 15040 28295
rect 11920 28250 11930 28265
rect 10600 28205 10610 28220
rect -345 28175 10610 28205
rect 10600 28160 10610 28175
rect 10670 28160 10680 28220
rect 12010 28160 12020 28220
rect 12080 28205 12090 28220
rect 12080 28175 15040 28205
rect 12080 28160 12090 28175
rect 10720 28115 10730 28130
rect -405 28085 10730 28115
rect 10720 28070 10730 28085
rect 10790 28070 10800 28130
rect 12170 28070 12180 28130
rect 12240 28115 12250 28130
rect 12240 28085 15040 28115
rect 12240 28070 12250 28085
rect 10930 28025 10940 28040
rect -465 27995 10940 28025
rect 10930 27980 10940 27995
rect 11000 27980 11010 28040
rect 11770 27980 11780 28040
rect 11840 28025 11850 28040
rect 11840 27995 15040 28025
rect 11840 27980 11850 27995
rect 11140 27935 11150 27950
rect -525 27905 11150 27935
rect 11140 27890 11150 27905
rect 11210 27890 11220 27950
rect 11930 27890 11940 27950
rect 12000 27935 12010 27950
rect 12000 27905 15040 27935
rect 12000 27890 12010 27905
rect 11350 27845 11360 27860
rect -585 27815 11360 27845
rect 11350 27800 11360 27815
rect 11420 27800 11430 27860
rect 12090 27800 12100 27860
rect 12160 27845 12170 27860
rect 12160 27815 15040 27845
rect 12160 27800 12170 27815
rect 11560 27755 11570 27770
rect -645 27725 11570 27755
rect 11560 27710 11570 27725
rect 11630 27710 11640 27770
rect 12250 27710 12260 27770
rect 12320 27755 12330 27770
rect 12320 27725 15040 27755
rect 12320 27710 12330 27725
rect 6210 25660 6220 25720
rect 6790 25660 6800 25720
rect 8940 25660 8950 25720
rect 9520 25660 9530 25720
rect 13620 25565 13630 25580
rect 13600 25535 13630 25565
rect 13620 25520 13630 25535
rect 13690 25520 13700 25580
rect 13710 25475 13720 25490
rect 13600 25445 13720 25475
rect 13710 25430 13720 25445
rect 13780 25430 13790 25490
rect 13800 25385 13810 25400
rect 13600 25355 13810 25385
rect 13800 25340 13810 25355
rect 13870 25340 13880 25400
rect 13890 25295 13900 25310
rect 13600 25265 13900 25295
rect 13890 25250 13900 25265
rect 13960 25250 13970 25310
rect 13980 25205 13990 25220
rect 13600 25175 13990 25205
rect 13980 25160 13990 25175
rect 14050 25160 14060 25220
rect 14070 25115 14080 25130
rect 13600 25085 14080 25115
rect 14070 25070 14080 25085
rect 14140 25070 14150 25130
rect 14160 25025 14170 25040
rect 13600 24995 14170 25025
rect 14160 24980 14170 24995
rect 14230 24980 14240 25040
rect 14610 24935 14620 24950
rect 13600 24905 14620 24935
rect 14610 24890 14620 24905
rect 14680 24890 14690 24950
rect 14250 24845 14260 24860
rect 13600 24815 14260 24845
rect 14250 24800 14260 24815
rect 14320 24800 14330 24860
rect 14520 24755 14530 24770
rect 13600 24725 14530 24755
rect 14520 24710 14530 24725
rect 14590 24710 14600 24770
rect 14430 24665 14440 24680
rect 13600 24635 14440 24665
rect 14430 24620 14440 24635
rect 14500 24620 14510 24680
rect 14340 24575 14350 24590
rect 13600 24545 14350 24575
rect 14340 24530 14350 24545
rect 14410 24530 14420 24590
rect 14608 13160 14692 13166
rect 14608 13150 14620 13160
rect 13600 13110 14620 13150
rect 14608 13100 14620 13110
rect 14680 13100 14692 13160
rect 14608 13094 14692 13100
rect 14518 12790 14602 12796
rect 14518 12780 14530 12790
rect 13600 12740 14530 12780
rect 14518 12730 14530 12740
rect 14590 12730 14602 12790
rect 14518 12724 14602 12730
rect 14428 12420 14512 12426
rect 14428 12410 14440 12420
rect 13600 12370 14440 12410
rect 14428 12360 14440 12370
rect 14500 12360 14512 12420
rect 14428 12354 14512 12360
rect 14338 12050 14422 12056
rect 14338 12040 14350 12050
rect 13600 12000 14350 12040
rect 14338 11990 14350 12000
rect 14410 11990 14422 12050
rect 14338 11984 14422 11990
rect 14248 11680 14332 11686
rect 14248 11670 14260 11680
rect 13600 11630 14260 11670
rect 14248 11620 14260 11630
rect 14320 11620 14332 11680
rect 14248 11614 14332 11620
rect 14158 11310 14242 11316
rect 14158 11300 14170 11310
rect 13600 11260 14170 11300
rect 14158 11250 14170 11260
rect 14230 11250 14242 11310
rect 14158 11244 14242 11250
rect 14068 10570 14152 10576
rect 14068 10560 14080 10570
rect 13600 10520 14080 10560
rect 14068 10510 14080 10520
rect 14140 10510 14152 10570
rect 14068 10504 14152 10510
rect 13978 10200 14062 10206
rect 13978 10190 13990 10200
rect 13600 10150 13990 10190
rect 13978 10140 13990 10150
rect 14050 10140 14062 10200
rect 13978 10134 14062 10140
rect 13888 9460 13972 9466
rect 13888 9450 13900 9460
rect 13600 9410 13900 9450
rect 13888 9400 13900 9410
rect 13960 9400 13972 9460
rect 13888 9394 13972 9400
rect 13798 8350 13882 8356
rect 13798 8340 13810 8350
rect 13600 8300 13810 8340
rect 13798 8290 13810 8300
rect 13870 8290 13882 8350
rect 13798 8284 13882 8290
rect 13708 6500 13792 6506
rect 13708 6490 13720 6500
rect 13600 6450 13720 6490
rect 13708 6440 13720 6450
rect 13780 6440 13792 6500
rect 13708 6434 13792 6440
rect 13628 4280 13712 4286
rect 13628 4220 13640 4280
rect 13700 4220 13712 4280
rect 13628 4214 13712 4220
<< via1 >>
rect 690 30750 750 30810
rect 620 29690 675 29750
rect 2345 29600 2405 29660
rect 3360 29510 3420 29570
rect 3880 29420 3940 29480
rect 4130 29330 4190 29390
rect 4370 29240 4430 29300
rect 4620 29150 4680 29210
rect 4860 29060 4920 29120
rect 5100 28970 5160 29030
rect 5350 28880 5410 28940
rect 5580 28790 5640 28850
rect 8100 28790 8160 28850
rect 6130 28700 6190 28760
rect 8870 28700 8930 28760
rect 6900 28610 6960 28670
rect 9640 28610 9700 28670
rect 7290 28520 7350 28580
rect 10020 28520 10080 28580
rect 7460 28430 7520 28490
rect 10210 28430 10270 28490
rect 5844 28340 5904 28400
rect 7680 28340 7740 28400
rect 11700 28340 11760 28400
rect 10420 28250 10480 28310
rect 11860 28250 11920 28310
rect 10610 28160 10670 28220
rect 12020 28160 12080 28220
rect 10730 28070 10790 28130
rect 12180 28070 12240 28130
rect 10940 27980 11000 28040
rect 11780 27980 11840 28040
rect 11150 27890 11210 27950
rect 11940 27890 12000 27950
rect 11360 27800 11420 27860
rect 12100 27800 12160 27860
rect 11570 27710 11630 27770
rect 12260 27710 12320 27770
rect 6220 25660 6790 25720
rect 8950 25660 9520 25720
rect 13630 25520 13690 25580
rect 13720 25430 13780 25490
rect 13810 25340 13870 25400
rect 13900 25250 13960 25310
rect 13990 25160 14050 25220
rect 14080 25070 14140 25130
rect 14170 24980 14230 25040
rect 14620 24890 14680 24950
rect 14260 24800 14320 24860
rect 14530 24710 14590 24770
rect 14440 24620 14500 24680
rect 14350 24530 14410 24590
rect 14620 13100 14680 13160
rect 14530 12730 14590 12790
rect 14440 12360 14500 12420
rect 14350 11990 14410 12050
rect 14260 11620 14320 11680
rect 14170 11250 14230 11310
rect 14080 10510 14140 10570
rect 13990 10140 14050 10200
rect 13900 9400 13960 9460
rect 13810 8290 13870 8350
rect 13720 6440 13780 6500
rect 13640 4220 13700 4280
<< metal2 >>
rect 690 30810 750 30820
rect 750 30800 765 30810
rect 750 30760 2588 30800
rect 750 30750 765 30760
rect 690 30740 750 30750
rect -710 30630 -650 30640
rect -650 30580 3998 30620
rect -710 30560 -650 30570
rect 5844 30560 5904 30570
rect 5844 30490 5904 30500
rect -320 29990 -250 30000
rect -260 29956 -250 29990
rect -260 29930 2941 29956
rect -320 29900 2941 29930
rect -260 29840 2941 29900
rect -320 29810 2941 29840
rect -260 29780 2941 29810
rect -260 29750 -250 29780
rect -320 29740 -250 29750
rect 605 29740 620 29750
rect 300 29700 620 29740
rect 300 27620 340 29700
rect 605 29690 620 29700
rect 675 29690 685 29750
rect 5844 29690 5904 29700
rect 2345 29660 2405 29670
rect 5844 29620 5904 29630
rect 2345 29590 2405 29600
rect 2345 27670 2385 29590
rect 3360 29570 3420 29580
rect 3360 29500 3420 29510
rect 3370 27660 3410 29500
rect 3880 29480 3940 29490
rect 3880 29410 3940 29420
rect 3890 27680 3930 29410
rect 4130 29390 4190 29400
rect 4130 29320 4190 29330
rect 4140 27660 4180 29320
rect 4370 29300 4430 29310
rect 4370 29230 4430 29240
rect 4380 27660 4420 29230
rect 4620 29210 4680 29220
rect 4620 29140 4680 29150
rect 4630 27660 4670 29140
rect 4860 29120 4920 29130
rect 4860 29050 4920 29060
rect 4870 27660 4910 29050
rect 5100 29030 5160 29040
rect 5100 28960 5160 28970
rect 5110 27680 5150 28960
rect 5350 28940 5410 28950
rect 5350 28870 5410 28880
rect 5360 27700 5400 28870
rect 5580 28850 5640 28860
rect 5580 28780 5640 28790
rect 5590 27680 5630 28780
rect 5854 28410 5894 29620
rect 8100 28850 8160 28860
rect 8100 28780 8160 28790
rect 6130 28760 6190 28770
rect 6130 28690 6190 28700
rect 5844 28400 5904 28410
rect 5844 28330 5904 28340
rect 6140 27670 6180 28690
rect 6900 28670 6960 28680
rect 6900 28600 6960 28610
rect 6910 27660 6950 28600
rect 7290 28580 7350 28590
rect 7290 28510 7350 28520
rect 7300 27670 7340 28510
rect 7460 28490 7520 28500
rect 7460 28420 7520 28430
rect 7470 27640 7510 28420
rect 7680 28400 7740 28410
rect 7680 28330 7740 28340
rect 7690 27670 7730 28330
rect 8110 27700 8150 28780
rect 8870 28760 8930 28770
rect 8870 28690 8930 28700
rect 8880 27710 8920 28690
rect 9640 28670 9700 28680
rect 9640 28600 9700 28610
rect 9650 27700 9690 28600
rect 10020 28580 10080 28590
rect 10020 28510 10080 28520
rect 10030 27700 10070 28510
rect 10210 28490 10270 28500
rect 10210 28420 10270 28430
rect 10220 27700 10260 28420
rect 11700 28400 11760 28410
rect 11700 28330 11760 28340
rect 10420 28310 10480 28320
rect 10420 28240 10480 28250
rect 10430 27680 10470 28240
rect 10610 28220 10670 28230
rect 10610 28150 10670 28160
rect 10620 27680 10660 28150
rect 10730 28130 10790 28140
rect 10730 28060 10790 28070
rect 10740 27680 10780 28060
rect 10940 28040 11000 28050
rect 10940 27970 11000 27980
rect 10950 27660 10990 27970
rect 11150 27950 11210 27960
rect 11150 27880 11210 27890
rect 11160 27680 11200 27880
rect 11360 27860 11420 27870
rect 11360 27790 11420 27800
rect 11370 27670 11410 27790
rect 11570 27770 11630 27780
rect 11570 27700 11630 27710
rect 11710 27700 11750 28330
rect 11860 28310 11920 28320
rect 11860 28240 11920 28250
rect 11780 28040 11840 28050
rect 11780 27970 11840 27980
rect 11790 27700 11830 27970
rect 11870 27700 11910 28240
rect 12020 28220 12080 28230
rect 12020 28150 12080 28160
rect 11940 27950 12000 27960
rect 11940 27880 12000 27890
rect 11950 27700 11990 27880
rect 12030 27700 12070 28150
rect 12180 28130 12240 28140
rect 12180 28060 12240 28070
rect 12100 27860 12160 27870
rect 12100 27790 12160 27800
rect 12110 27700 12150 27790
rect 12190 27700 12230 28060
rect 12260 27770 12320 27780
rect 12260 27700 12320 27710
rect -190 27360 -130 27370
rect -130 27315 90 27355
rect -190 27290 -130 27300
rect -320 27060 -260 27070
rect -260 27015 90 27055
rect -320 26990 -260 27000
rect -450 26750 -390 26760
rect -390 26705 90 26745
rect -450 26680 -390 26690
rect -580 26340 -520 26350
rect -520 26295 90 26335
rect -580 26270 -520 26280
rect -710 26210 -650 26220
rect -650 26165 90 26205
rect -710 26140 -650 26150
rect 6220 25720 6790 25730
rect 6220 25650 6790 25660
rect 8950 25720 9520 25730
rect 8950 25650 9520 25660
rect 13630 25580 13690 25590
rect 13630 25510 13690 25520
rect 13640 4290 13680 25510
rect 13720 25490 13780 25500
rect 13720 25420 13780 25430
rect 13730 6510 13770 25420
rect 13810 25400 13870 25410
rect 13810 25330 13870 25340
rect 13820 8360 13860 25330
rect 13900 25310 13960 25320
rect 13900 25240 13960 25250
rect 13910 9470 13950 25240
rect 13990 25220 14050 25230
rect 13990 25150 14050 25160
rect 14000 10210 14040 25150
rect 14080 25130 14140 25140
rect 14080 25060 14140 25070
rect 14090 10580 14130 25060
rect 14170 25040 14230 25050
rect 14170 24970 14230 24980
rect 14180 11320 14220 24970
rect 14620 24950 14680 24960
rect 14620 24880 14680 24890
rect 14260 24860 14320 24870
rect 14260 24790 14320 24800
rect 14270 11690 14310 24790
rect 14530 24770 14590 24780
rect 14530 24700 14590 24710
rect 14440 24680 14500 24690
rect 14440 24610 14500 24620
rect 14350 24590 14410 24600
rect 14350 24520 14410 24530
rect 14360 12060 14400 24520
rect 14450 12430 14490 24610
rect 14540 12800 14580 24700
rect 14630 13170 14670 24880
rect 14620 13160 14680 13170
rect 14620 13090 14680 13100
rect 14530 12790 14590 12800
rect 14530 12720 14590 12730
rect 14440 12420 14500 12430
rect 14440 12350 14500 12360
rect 14350 12050 14410 12060
rect 14350 11980 14410 11990
rect 14260 11680 14320 11690
rect 14260 11610 14320 11620
rect 14170 11310 14230 11320
rect 14170 11240 14230 11250
rect 14080 10570 14140 10580
rect 14080 10500 14140 10510
rect 13990 10200 14050 10210
rect 13990 10130 14050 10140
rect 13900 9460 13960 9470
rect 13900 9390 13960 9400
rect 13810 8350 13870 8360
rect 13810 8280 13870 8290
rect 13720 6500 13780 6510
rect 13720 6430 13780 6440
rect 13640 4280 13700 4290
rect 13640 4210 13700 4220
<< via2 >>
rect -710 30570 -650 30630
rect 5844 30500 5904 30560
rect -320 29930 -260 29990
rect -320 29840 -260 29900
rect -320 29750 -260 29810
rect 5844 29630 5904 29690
rect -190 27300 -130 27360
rect -320 27000 -260 27060
rect -450 26690 -390 26750
rect -580 26280 -520 26340
rect -710 26150 -650 26210
rect 6220 25660 6790 25720
rect 8950 25660 9520 25720
<< metal3 >>
rect -720 30630 -640 30635
rect -720 30570 -710 30630
rect -650 30570 -640 30630
rect -720 30565 -640 30570
rect -710 26215 -650 30565
rect 5834 30560 5914 30570
rect 5834 30500 5844 30560
rect 5904 30500 5914 30560
rect 5834 30490 5914 30500
rect -330 29990 -250 29995
rect -330 29930 -320 29990
rect -260 29930 -250 29990
rect -330 29900 -250 29930
rect -330 29840 -320 29900
rect -260 29840 -250 29900
rect -330 29810 -250 29840
rect -330 29750 -320 29810
rect -260 29750 -250 29810
rect -330 29745 -250 29750
rect -320 27065 -260 29745
rect 5844 29700 5904 30490
rect 5834 29690 5914 29700
rect 5834 29630 5844 29690
rect 5904 29630 5914 29690
rect 5834 29620 5914 29630
rect -190 27365 -130 27400
rect -200 27360 -120 27365
rect -200 27300 -190 27360
rect -130 27300 -120 27360
rect -200 27295 -120 27300
rect -190 27260 -130 27295
rect -330 27060 -250 27065
rect -330 27000 -320 27060
rect -260 27000 -250 27060
rect -330 26995 -250 27000
rect -450 26755 -390 26790
rect -460 26750 -380 26755
rect -460 26690 -450 26750
rect -390 26690 -380 26750
rect -460 26685 -380 26690
rect -450 26650 -390 26685
rect -580 26345 -520 26380
rect -590 26340 -510 26345
rect -590 26280 -580 26340
rect -520 26280 -510 26340
rect -590 26275 -510 26280
rect -580 26240 -520 26275
rect -720 26210 -640 26215
rect -720 26150 -710 26210
rect -650 26150 -640 26210
rect -720 26145 -640 26150
rect 6210 25720 6800 25725
rect 6210 25660 6220 25720
rect 6790 25660 6800 25720
rect 6210 25655 6800 25660
rect 8940 25720 9530 25725
rect 8940 25660 8950 25720
rect 9520 25660 9530 25720
rect 8940 25655 9530 25660
use bootstrap  bootstrap_0 ~/Desktop/SAR_ADC_12bit/layout/subcells/bootstrap
timestamp 1715417500
transform -1 0 22799 0 -1 31168
box 9245 72 20313 2258
use CDAC_mim_12bit  CDAC_mim_12bit_1 ~/Desktop/SAR_ADC_12bit/layout/subcells/CDAC
timestamp 1715383943
transform 1 0 400 0 1 370
box -400 -380 13390 24190
use switches  switches_0 ~/Desktop/SAR_ADC_12bit/layout/subcells/switches
timestamp 1714328045
transform 1 0 220 0 1 23665
box -200 855 13477 4090
<< end >>
