magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< nwell >>
rect -246 -1019 246 1019
<< pmos >>
rect -50 -800 50 800
<< pdiff >>
rect -108 788 -50 800
rect -108 -788 -96 788
rect -62 -788 -50 788
rect -108 -800 -50 -788
rect 50 788 108 800
rect 50 -788 62 788
rect 96 -788 108 788
rect 50 -800 108 -788
<< pdiffc >>
rect -96 -788 -62 788
rect 62 -788 96 788
<< nsubdiff >>
rect -210 949 -114 983
rect 114 949 210 983
rect -210 887 -176 949
rect 176 887 210 949
rect -210 -949 -176 -887
rect 176 -949 210 -887
rect -210 -983 -114 -949
rect 114 -983 210 -949
<< nsubdiffcont >>
rect -114 949 114 983
rect -210 -887 -176 887
rect 176 -887 210 887
rect -114 -983 114 -949
<< poly >>
rect -50 881 50 897
rect -50 847 -34 881
rect 34 847 50 881
rect -50 800 50 847
rect -50 -847 50 -800
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect -50 -897 50 -881
<< polycont >>
rect -34 847 34 881
rect -34 -881 34 -847
<< locali >>
rect -210 949 -114 983
rect 114 949 210 983
rect -210 887 -176 949
rect 176 887 210 949
rect -50 847 -34 881
rect 34 847 50 881
rect -96 788 -62 804
rect -96 -804 -62 -788
rect 62 788 96 804
rect 62 -804 96 -788
rect -50 -881 -34 -847
rect 34 -881 50 -847
rect -210 -949 -176 -887
rect 176 -949 210 -887
rect -210 -983 -114 -949
rect 114 -983 210 -949
<< viali >>
rect -34 847 34 881
rect -96 -788 -62 788
rect 62 -788 96 788
rect -34 -881 34 -847
<< metal1 >>
rect -46 881 46 887
rect -46 847 -34 881
rect 34 847 46 881
rect -46 841 46 847
rect -102 788 -56 800
rect -102 -788 -96 788
rect -62 -788 -56 788
rect -102 -800 -56 -788
rect 56 788 102 800
rect 56 -788 62 788
rect 96 -788 102 788
rect 56 -800 102 -788
rect -46 -847 46 -841
rect -46 -881 -34 -847
rect 34 -881 46 -847
rect -46 -887 46 -881
<< properties >>
string FIXED_BBOX -193 -966 193 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
