** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/break_before_make/break_before_make.sch

.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt break_before_make EN_VSS_I[10] EN_VSS_I[9] EN_VSS_I[8] EN_VSS_I[7] EN_VSS_I[6] EN_VSS_I[5] EN_VSS_I[4] EN_VSS_I[3]
+ EN_VSS_I[2] EN_VSS_I[1] EN_VSS_I[0] VDD VSS EN_VSS_O[10] EN_VSS_O[9] EN_VSS_O[8] EN_VSS_O[7] EN_VSS_O[6] EN_VSS_O[5] EN_VSS_O[4] EN_VSS_O[3]
+ EN_VSS_O[2] EN_VSS_O[1] EN_VSS_O[0] EN_VREF_Z_O[10] EN_VREF_Z_O[9] EN_VREF_Z_O[8] EN_VREF_Z_O[7] EN_VREF_Z_O[6] EN_VREF_Z_O[5] EN_VREF_Z_O[4]
+ EN_VREF_Z_O[3] EN_VREF_Z_O[2] EN_VREF_Z_O[1] EN_VREF_Z_O[0] EN_VREF_Z_I[10] EN_VREF_Z_I[9] EN_VREF_Z_I[8] EN_VREF_Z_I[7] EN_VREF_Z_I[6]
+ EN_VREF_Z_I[5] EN_VREF_Z_I[4] EN_VREF_Z_I[3] EN_VREF_Z_I[2] EN_VREF_Z_I[1] EN_VREF_Z_I[0]
*.PININFO EN_VSS_I[10:0]:I EN_VREF_Z_I[10:0]:I VDD:I VSS:I EN_VSS_O[10:0]:O EN_VREF_Z_O[10:0]:O
x1[10] EN_VSS_I[10] EN_VREF_Z_O[10] VSS VSS VDD VDD EN_VSS_O[10] sky130_fd_sc_hd__and2_4
x1[9] EN_VSS_I[9] EN_VREF_Z_O[9] VSS VSS VDD VDD EN_VSS_O[9] sky130_fd_sc_hd__and2_4
x1[8] EN_VSS_I[8] EN_VREF_Z_O[8] VSS VSS VDD VDD EN_VSS_O[8] sky130_fd_sc_hd__and2_4
x1[7] EN_VSS_I[7] EN_VREF_Z_O[7] VSS VSS VDD VDD EN_VSS_O[7] sky130_fd_sc_hd__and2_4
x1[6] EN_VSS_I[6] EN_VREF_Z_O[6] VSS VSS VDD VDD EN_VSS_O[6] sky130_fd_sc_hd__and2_4
x1[5] EN_VSS_I[5] EN_VREF_Z_O[5] VSS VSS VDD VDD EN_VSS_O[5] sky130_fd_sc_hd__and2_4
x1[4] EN_VSS_I[4] EN_VREF_Z_O[4] VSS VSS VDD VDD EN_VSS_O[4] sky130_fd_sc_hd__and2_4
x1[3] EN_VSS_I[3] EN_VREF_Z_O[3] VSS VSS VDD VDD EN_VSS_O[3] sky130_fd_sc_hd__and2_4
x1[2] EN_VSS_I[2] EN_VREF_Z_O[2] VSS VSS VDD VDD EN_VSS_O[2] sky130_fd_sc_hd__and2_4
x1[1] EN_VSS_I[1] EN_VREF_Z_O[1] VSS VSS VDD VDD EN_VSS_O[1] sky130_fd_sc_hd__and2_4
x1[0] EN_VSS_I[0] EN_VREF_Z_O[0] VSS VSS VDD VDD EN_VSS_O[0] sky130_fd_sc_hd__and2_4
x2[10] EN_VSS_O[10] EN_VREF_Z_I[10] VSS VSS VDD VDD EN_VREF_Z_O[10] sky130_fd_sc_hd__or2_4
x2[9] EN_VSS_O[9] EN_VREF_Z_I[9] VSS VSS VDD VDD EN_VREF_Z_O[9] sky130_fd_sc_hd__or2_4
x2[8] EN_VSS_O[8] EN_VREF_Z_I[8] VSS VSS VDD VDD EN_VREF_Z_O[8] sky130_fd_sc_hd__or2_4
x2[7] EN_VSS_O[7] EN_VREF_Z_I[7] VSS VSS VDD VDD EN_VREF_Z_O[7] sky130_fd_sc_hd__or2_4
x2[6] EN_VSS_O[6] EN_VREF_Z_I[6] VSS VSS VDD VDD EN_VREF_Z_O[6] sky130_fd_sc_hd__or2_4
x2[5] EN_VSS_O[5] EN_VREF_Z_I[5] VSS VSS VDD VDD EN_VREF_Z_O[5] sky130_fd_sc_hd__or2_4
x2[4] EN_VSS_O[4] EN_VREF_Z_I[4] VSS VSS VDD VDD EN_VREF_Z_O[4] sky130_fd_sc_hd__or2_4
x2[3] EN_VSS_O[3] EN_VREF_Z_I[3] VSS VSS VDD VDD EN_VREF_Z_O[3] sky130_fd_sc_hd__or2_4
x2[2] EN_VSS_O[2] EN_VREF_Z_I[2] VSS VSS VDD VDD EN_VREF_Z_O[2] sky130_fd_sc_hd__or2_4
x2[1] EN_VSS_O[1] EN_VREF_Z_I[1] VSS VSS VDD VDD EN_VREF_Z_O[1] sky130_fd_sc_hd__or2_4
x2[0] EN_VSS_O[0] EN_VREF_Z_I[0] VSS VSS VDD VDD EN_VREF_Z_O[0] sky130_fd_sc_hd__or2_4
.ends
.end
