** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/SAR_ADC_12bit.sch

.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/subcells/state_machine/state_machine_openlane_generated.spice

.subckt CDAC_12bit C0_dummy_btm C0_btm C1_btm C2_btm C3_btm C4_btm C5_btm C6_btm C7_btm C8_btm C9_btm C10_btm VDAC VSS
.ends

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START
+ EN_OFFSET_CAL CLK VREF_GND SINGLE_ENDED
*.PININFO VIN_P:I VDD:I VREF:I VCM:I VSS:I VIN_N:I RST_Z:I START:I CLK_DATA:O DATA[5:0]:O EN_OFFSET_CAL:I CLK:I VREF_GND:I
*+ SINGLE_ENDED:I
x1 C0_dummy_N_btm C0_N_btm C1_N_btm C2_N_btm C3_N_btm C4_N_btm C5_N_btm C6_N_btm C7_N_btm C8_N_btm C9_N_btm C10_N_btm VDAC_N VSS
+ CDAC_12bit
x2 C0_dummy_P_btm C0_P_btm C1_P_btm C2_P_btm C3_P_btm C4_P_btm C5_P_btm C6_P_btm C7_P_btm C8_P_btm C9_P_btm C10_P_btm VDAC_P VSS
+ CDAC_12bit
x3 VCM VREF_GND VREF VIN_P EN_VIN_BSTR_P EN_REF_Z_P[10] EN_REF_Z_P[9] EN_REF_Z_P[8] EN_REF_Z_P[7] EN_REF_Z_P[6] EN_REF_Z_P[5]
+ EN_REF_Z_P[4] EN_REF_Z_P[3] EN_REF_Z_P[2] EN_REF_Z_P[1] EN_REF_Z_P[0] EN_VSS_P[10] EN_VSS_P[9] EN_VSS_P[8] EN_VSS_P[7] EN_VSS_P[6] EN_VSS_P[5]
+ EN_VSS_P[4] EN_VSS_P[3] EN_VSS_P[2] EN_VSS_P[1] EN_VSS_P[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3]
+ EN_VCM[2] EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY C8_P_btm C7_P_btm C0_P_btm C6_P_btm C5_P_btm C0_dummy_P_btm C4_P_btm C3_P_btm VDAC_P
+ C10_P_btm C9_P_btm C2_P_btm C1_P_btm VDD VSS switches
x4 VCM VREF_GND VREF VIN_N EN_VIN_BSTR_N EN_REF_Z_N[10] EN_REF_Z_N[9] EN_REF_Z_N[8] EN_REF_Z_N[7] EN_REF_Z_N[6] EN_REF_Z_N[5]
+ EN_REF_Z_N[4] EN_REF_Z_N[3] EN_REF_Z_N[2] EN_REF_Z_N[1] EN_REF_Z_N[0] EN_VSS_N[10] EN_VSS_N[9] EN_VSS_N[8] EN_VSS_N[7] EN_VSS_N[6] EN_VSS_N[5]
+ EN_VSS_N[4] EN_VSS_N[3] EN_VSS_N[2] EN_VSS_N[1] EN_VSS_N[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3]
+ EN_VCM[2] EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY C8_N_btm C7_N_btm C0_N_btm C6_N_btm C5_N_btm C0_dummy_N_btm C4_N_btm C3_N_btm VDAC_N
+ C10_N_btm C9_N_btm C2_N_btm C1_N_btm VDD VSS switches
x5 VDAC_N VDAC_P VDD RST_Z VDAC_Pi VDAC_Ni VSS CAL_P CAL_N preamplifier
x6 VDD VDAC_Pi VDAC_Ni EN_COMP COMP_P COMP_N VSS latched_comparator
x7 VDD COMP_P EN_COMP CAL_P CAL_N EN_VOS_CAL VSS OFFSET_CAL_CYCLE offset_calibration
x8 VDD VSS RST_Z START COMP_P SMPL EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2]
+ EN_VCM[1] EN_VCM[0] EN_COMP SMPL_ON_P SMPL_ON_N EN_VCM_DUMMY EN_VCM_SW EN_OFFSET_CAL OFFSET_CAL_CYCLE EN_VOS_CAL CLK_DATA DATA[5] DATA[4]
+ DATA[3] DATA[2] DATA[1] DATA[0] EN_VSS_N[10] EN_VSS_N[9] EN_VSS_N[8] EN_VSS_N[7] EN_VSS_N[6] EN_VSS_N[5] EN_VSS_N[4] EN_VSS_N[3]
+ EN_VSS_N[2] EN_VSS_N[1] EN_VSS_N[0] EN_REF_Z_N[10] EN_REF_Z_N[9] EN_REF_Z_N[8] EN_REF_Z_N[7] EN_REF_Z_N[6] EN_REF_Z_N[5] EN_REF_Z_N[4]
+ EN_REF_Z_N[3] EN_REF_Z_N[2] EN_REF_Z_N[1] EN_REF_Z_N[0] EN_VSS_P_BBM[10] EN_VSS_P_BBM[9] EN_VSS_P_BBM[8] EN_VSS_P_BBM[7] EN_VSS_P_BBM[6]
+ EN_VSS_P_BBM[5] EN_VSS_P_BBM[4] EN_VSS_P_BBM[3] EN_VSS_P_BBM[2] EN_VSS_P_BBM[1] EN_VSS_P_BBM[0] EN_REF_Z_P_BBM[10] EN_REF_Z_P_BBM[9]
+ EN_REF_Z_P_BBM[8] EN_REF_Z_P_BBM[7] EN_REF_Z_P_BBM[6] EN_REF_Z_P_BBM[5] EN_REF_Z_P_BBM[4] EN_REF_Z_P_BBM[3] EN_REF_Z_P_BBM[2] EN_REF_Z_P_BBM[1]
+ EN_REF_Z_P_BBM[0] CLK EN_VCM_SW EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2] EN_VCM[1] EN_VCM[0]
+ SINGLE_ENDED state_machine
x11 VDD VSS VIN_P SMPL_ON_P SMPL EN_VIN_BSTR_P bootstrap
x12 VDD VSS VIN_N SMPL_ON_N SMPL EN_VIN_BSTR_N bootstrap
x9 EN_VSS_P_BBM[10] EN_VSS_P_BBM[9] EN_VSS_P_BBM[8] EN_VSS_P_BBM[7] EN_VSS_P_BBM[6] EN_VSS_P_BBM[5] EN_VSS_P_BBM[4]
+ EN_VSS_P_BBM[3] EN_VSS_P_BBM[2] EN_VSS_P_BBM[1] EN_VSS_P_BBM[0] VDD VSS EN_VSS_P[10] EN_VSS_P[9] EN_VSS_P[8] EN_VSS_P[7] EN_VSS_P[6] EN_VSS_P[5]
+ EN_VSS_P[4] EN_VSS_P[3] EN_VSS_P[2] EN_VSS_P[1] EN_VSS_P[0] EN_REF_Z_P[10] EN_REF_Z_P[9] EN_REF_Z_P[8] EN_REF_Z_P[7] EN_REF_Z_P[6]
+ EN_REF_Z_P[5] EN_REF_Z_P[4] EN_REF_Z_P[3] EN_REF_Z_P[2] EN_REF_Z_P[1] EN_REF_Z_P[0] EN_REF_Z_P_BBM[10] EN_REF_Z_P_BBM[9] EN_REF_Z_P_BBM[8]
+ EN_REF_Z_P_BBM[7] EN_REF_Z_P_BBM[6] EN_REF_Z_P_BBM[5] EN_REF_Z_P_BBM[4] EN_REF_Z_P_BBM[3] EN_REF_Z_P_BBM[2] EN_REF_Z_P_BBM[1] EN_REF_Z_P_BBM[0]
+ break_before_make
.ends

* expanding   symbol:  subcells/switches/switches.sym # of pins=25
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/switches/switches.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/switches/switches.sch
.subckt switches VCM VREF_GND VREF VIN EN_VIN EN_VREF_Z[10] EN_VREF_Z[9] EN_VREF_Z[8] EN_VREF_Z[7] EN_VREF_Z[6] EN_VREF_Z[5]
+ EN_VREF_Z[4] EN_VREF_Z[3] EN_VREF_Z[2] EN_VREF_Z[1] EN_VREF_Z[0] EN_VSS[10] EN_VSS[9] EN_VSS[8] EN_VSS[7] EN_VSS[6] EN_VSS[5] EN_VSS[4]
+ EN_VSS[3] EN_VSS[2] EN_VSS[1] EN_VSS[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2]
+ EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY Cbtm_8 Cbtm_7 Cbtm_0 Cbtm_6 Cbtm_5 Cbtm_0_dummy Cbtm_4 Cbtm_3 VDAC Cbtm_10 Cbtm_9 Cbtm_2 Cbtm_1
+ VDD VSS
*.PININFO VCM:I VREF_GND:I VREF:I VIN:I VDD:I Cbtm_0_dummy:O Cbtm_0:O Cbtm_1:O Cbtm_2:O Cbtm_3:O Cbtm_4:O Cbtm_5:O Cbtm_6:O
*+ Cbtm_7:O Cbtm_8:O Cbtm_9:O Cbtm_10:O VDAC:O EN_VIN:I EN_VREF_Z[10:0]:I EN_VSS[10:0]:I EN_VCM[10:0]:I EN_VCM_DUMMY:I EN_VCM_SW:I VSS:I
x1 VCM EN_VCM_SW VDAC VDD VSS switch_VCM
x2 VCM VREF_GND VIN VREF EN_VCM[10] EN_VREF_Z[10] Cbtm_10 VDD EN_VSS[10] EN_VIN VSS switch_C10
x3 VCM VREF_GND VIN VREF EN_VCM[9] EN_VREF_Z[9] Cbtm_9 VDD EN_VSS[9] EN_VIN VSS switch_C9
x4 VCM VREF_GND VIN VREF EN_VCM[8] EN_VREF_Z[8] Cbtm_8 VDD EN_VSS[8] EN_VIN VSS switch_C8
x5 VCM VREF_GND VIN VREF EN_VCM[7] EN_VREF_Z[7] Cbtm_7 VDD EN_VSS[7] EN_VIN VSS switch_C7
x6 VCM VREF_GND VIN VREF EN_VCM[6] EN_VREF_Z[6] Cbtm_6 VDD EN_VSS[6] EN_VIN VSS switch_C6
x7 VCM VREF_GND VIN VREF EN_VCM[5] EN_VREF_Z[5] Cbtm_5 VDD EN_VSS[5] EN_VIN VSS switch_C5
x8 VCM VREF_GND VIN VREF EN_VCM[4] EN_VREF_Z[4] Cbtm_4 VDD EN_VSS[4] EN_VIN VSS switch_C5
x9 VCM VREF_GND VIN VREF EN_VCM[3] EN_VREF_Z[3] Cbtm_3 VDD EN_VSS[3] EN_VIN VSS switch_C5
x10 VCM VREF_GND VIN VREF EN_VCM[2] EN_VREF_Z[2] Cbtm_2 VDD EN_VSS[2] EN_VIN VSS switch_C5
x11 VCM VREF_GND VIN VREF EN_VCM[1] EN_VREF_Z[1] Cbtm_1 VDD EN_VSS[1] EN_VIN VSS switch_C5
x12 VCM VREF_GND VIN VREF EN_VCM[0] EN_VREF_Z[0] Cbtm_0 VDD EN_VSS[0] EN_VIN VSS switch_C5
x13 VCM VIN EN_VCM_DUMMY Cbtm_0_dummy EN_VIN VSS switch_C0_dummy
.ends


* expanding   symbol:  subcells/preamplifier/preamplifier.sym # of pins=9
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/preamplifier/preamplifier.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/preamplifier/preamplifier.sch
.subckt preamplifier IN_N IN_P VDD EN OUT_P OUT_N VSS CAL_P CAL_N
*.PININFO VDD:I VSS:I IN_P:I IN_N:I OUT_P:O OUT_N:O EN:I CAL_P:I CAL_N:I
XM4 net1 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 m=6
XM5 net5 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 m=1
XM7 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM12 OUT_N net5 net9 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=4
XM14 OUT_P net5 net10 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=4
XM8 net9 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 m=1
XM6 net10 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 m=1
XM16 net8 EN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=1
XM17 net3 EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM18 net5 EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
x1 EN VSS VSS VDD VDD EN_Z sky130_fd_sc_hd__inv_1
XM20 net6 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=2
XM19 VDD OUT_N net6 VSS sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.5 nf=1 m=1
XM21 VDD OUT_P net6 VSS sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.5 nf=1 m=1
XM1 net12 IN_P net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=24 nf=4 m=4
XM2 net7 IN_N net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=24 nf=4 m=4
XM15 net9 CAL_P net11 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM22 net10 CAL_N net11 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM3 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 m=1
XR6 net2 net3 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM23 net11 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 m=3
XR3 net8 net2 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[3] rn[0] OUT_N VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[2] rn[1] rn[0] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[1] rn[2] rn[1] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[0] common rn[2] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR5 net4 net5 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM9 OUT_P VSS net7 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=8 nf=1 m=1
XM10 OUT_N VSS net12 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=8 nf=1 m=1
XR1[3] rp[0] OUT_P VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[2] rp[1] rp[0] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[1] rp[2] rp[1] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[0] common rp[2] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM11 VDD net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 m=2
XM13 VSS net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=2
XM24 net10 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 m=1
XM25 net9 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 m=1
.ends


* expanding   symbol:  subcells/latched_comparator/latched_comparator.sym # of pins=7
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/latched_comparator/latched_comparator.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/latched_comparator/latched_comparator.sch
.subckt latched_comparator VDD VIN_P VIN_N EN OUT_P OUT_N VSS
*.PININFO VIN_P:I VIN_N:I VDD:I VSS:I EN:I OUT_N:O OUT_P:O
x1 EN VSS VSS VDD VDD ENi sky130_fd_sc_hd__buf_4
XM10 net2 ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 OUT_Ni ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 OUT_Ni OUT_Pi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
XM9 OUT_Pi OUT_Ni VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 m=1
XM3 OUT_Ni OUT_Pi net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 OUT_Pi OUT_Ni net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM18 net1 ENi VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=2
XM16 net3 VIN_N net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM1 net2 VIN_P net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM11 OUT_Pi ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 net3 ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
x4 OUT_Pi VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x5 OUT_Ni VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x6 net5 VSS VSS VDD VDD OUT_N sky130_fd_sc_hd__inv_4
x7 net4 VSS VSS VDD VDD OUT_P sky130_fd_sc_hd__inv_4
XM2 net1 net1 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=2
.ends


* expanding   symbol:  subcells/offset_calibration/offset_calibration.sym # of pins=8
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/offset_calibration/offset_calibration.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/offset_calibration/offset_calibration.sch
.subckt offset_calibration VDD CAL_RESULT EN_COMP CAL_P CAL_N EN VSS CAL_CYCLE
*.PININFO EN_COMP:I CAL_N:O CAL_P:O VDD:I VSS:I EN:I CAL_RESULT:I CAL_CYCLE:I
XM26 net2 EN_COMPi net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM27 net1 CAL_RESULTi VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM28 net2 EN_COMP_Z net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM29 net3 CAL_RESULTi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM30 net2 LOAD_CALi CAL_P VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM31 net2 LOAD_CAL_Z CAL_P VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
x22 EN net8 net7 VSS VSS VDD VDD LOAD_CAL_Z sky130_fd_sc_hd__nand3_1
x3 LOAD_CAL_Z VSS VSS VDD VDD LOAD_CALi sky130_fd_sc_hd__inv_1
XM32 net5 LOAD_CAL_Z CAL_N VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM33 net5 LOAD_CALi CAL_N VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM34 net5 EN_COMP_Z net6 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM35 net6 CAL_RESULT_Z VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM36 net5 EN_COMPi net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM37 net4 CAL_RESULT_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM24 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=10 nf=1 m=3
XM25 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=10 nf=1 m=3
XM1 CAL_N EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 CAL_P EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
x1 CAL_RESULT CAL_CYCLE VSS VSS VDD VDD CAL_RESULT_Z sky130_fd_sc_hd__nand2_1
x4 CAL_RESULT_Z VSS VSS VDD VDD CAL_RESULTi sky130_fd_sc_hd__inv_1
x2 EN_COMP CAL_CYCLE VSS VSS VDD VDD EN_COMP_Z sky130_fd_sc_hd__nand2_1
x5 EN_COMP_Z VSS VSS VDD VDD EN_COMPi sky130_fd_sc_hd__inv_1
x6 EN_COMPi VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_1
x7 CAL_CYCLE VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  subcells/bootstrap/bootstrap.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/bootstrap/bootstrap.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/bootstrap/bootstrap.sch
.subckt bootstrap VDD VSS VIN SW_ON EN VGATE
*.PININFO VDD:I VSS:I VIN:I VGATE:O EN:I SW_ON:O
XM1 VDD VGATE Vtop Vtop sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 VGATE EN_Z_LVL_SHFT Vtop Vtop sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=4 m=1
XM3 VGATE VDD Vd VSS sky130_fd_pr__nfet_05v0_nvt L=0.9 W=8 nf=2 m=1
XM4 Vd EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 m=1
XM5 Vbottom EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 m=1
XM6 Vtop Vbottom Vtop Vtop sky130_fd_pr__pfet_01v8 L=16.6 W=13.6 nf=4 m=1
x1 EN VSS VSS VDD VDD EN_Z sky130_fd_sc_hd__inv_4
XM8 VIN VGATE Vbottom VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 m=1
XM7 VGATE VDD VGATE_1V8 VSS sky130_fd_pr__nfet_05v0_nvt L=0.9 W=4 nf=1 m=1
x2 VGATE_1V8 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_2
x3 net1 VSS VSS VDD VDD SW_ON sky130_fd_sc_hd__inv_4
XM9 EN_Z_LVL_SHFT EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 EN_Z_LVL_SHFT EN Vbottom VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM11 EN_Z_LVL_SHFT VGATE Vbottom VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=2 m=1
.ends


* expanding   symbol:  subcells/break_before_make/break_before_make.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/break_before_make/break_before_make.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/break_before_make/break_before_make.sch
.subckt break_before_make EN_VSS_I[10] EN_VSS_I[9] EN_VSS_I[8] EN_VSS_I[7] EN_VSS_I[6] EN_VSS_I[5] EN_VSS_I[4] EN_VSS_I[3]
+ EN_VSS_I[2] EN_VSS_I[1] EN_VSS_I[0] VDD VSS EN_VSS_O[10] EN_VSS_O[9] EN_VSS_O[8] EN_VSS_O[7] EN_VSS_O[6] EN_VSS_O[5] EN_VSS_O[4] EN_VSS_O[3]
+ EN_VSS_O[2] EN_VSS_O[1] EN_VSS_O[0] EN_VREF_Z_O[10] EN_VREF_Z_O[9] EN_VREF_Z_O[8] EN_VREF_Z_O[7] EN_VREF_Z_O[6] EN_VREF_Z_O[5] EN_VREF_Z_O[4]
+ EN_VREF_Z_O[3] EN_VREF_Z_O[2] EN_VREF_Z_O[1] EN_VREF_Z_O[0] EN_VREF_Z_I[10] EN_VREF_Z_I[9] EN_VREF_Z_I[8] EN_VREF_Z_I[7] EN_VREF_Z_I[6]
+ EN_VREF_Z_I[5] EN_VREF_Z_I[4] EN_VREF_Z_I[3] EN_VREF_Z_I[2] EN_VREF_Z_I[1] EN_VREF_Z_I[0]
*.PININFO EN_VSS_I[10:0]:I EN_VREF_Z_I[10:0]:I VDD:I VSS:I EN_VSS_O[10:0]:O EN_VREF_Z_O[10:0]:O
x1[10] EN_VSS_I[10] EN_VREF_Z_O[10] VSS VSS VDD VDD EN_VSS_O[10] sky130_fd_sc_hd__and2_4
x1[9] EN_VSS_I[9] EN_VREF_Z_O[9] VSS VSS VDD VDD EN_VSS_O[9] sky130_fd_sc_hd__and2_4
x1[8] EN_VSS_I[8] EN_VREF_Z_O[8] VSS VSS VDD VDD EN_VSS_O[8] sky130_fd_sc_hd__and2_4
x1[7] EN_VSS_I[7] EN_VREF_Z_O[7] VSS VSS VDD VDD EN_VSS_O[7] sky130_fd_sc_hd__and2_4
x1[6] EN_VSS_I[6] EN_VREF_Z_O[6] VSS VSS VDD VDD EN_VSS_O[6] sky130_fd_sc_hd__and2_4
x1[5] EN_VSS_I[5] EN_VREF_Z_O[5] VSS VSS VDD VDD EN_VSS_O[5] sky130_fd_sc_hd__and2_4
x1[4] EN_VSS_I[4] EN_VREF_Z_O[4] VSS VSS VDD VDD EN_VSS_O[4] sky130_fd_sc_hd__and2_4
x1[3] EN_VSS_I[3] EN_VREF_Z_O[3] VSS VSS VDD VDD EN_VSS_O[3] sky130_fd_sc_hd__and2_4
x1[2] EN_VSS_I[2] EN_VREF_Z_O[2] VSS VSS VDD VDD EN_VSS_O[2] sky130_fd_sc_hd__and2_4
x1[1] EN_VSS_I[1] EN_VREF_Z_O[1] VSS VSS VDD VDD EN_VSS_O[1] sky130_fd_sc_hd__and2_4
x1[0] EN_VSS_I[0] EN_VREF_Z_O[0] VSS VSS VDD VDD EN_VSS_O[0] sky130_fd_sc_hd__and2_4
x2[10] EN_VSS_O[10] EN_VREF_Z_I[10] VSS VSS VDD VDD EN_VREF_Z_O[10] sky130_fd_sc_hd__or2_4
x2[9] EN_VSS_O[9] EN_VREF_Z_I[9] VSS VSS VDD VDD EN_VREF_Z_O[9] sky130_fd_sc_hd__or2_4
x2[8] EN_VSS_O[8] EN_VREF_Z_I[8] VSS VSS VDD VDD EN_VREF_Z_O[8] sky130_fd_sc_hd__or2_4
x2[7] EN_VSS_O[7] EN_VREF_Z_I[7] VSS VSS VDD VDD EN_VREF_Z_O[7] sky130_fd_sc_hd__or2_4
x2[6] EN_VSS_O[6] EN_VREF_Z_I[6] VSS VSS VDD VDD EN_VREF_Z_O[6] sky130_fd_sc_hd__or2_4
x2[5] EN_VSS_O[5] EN_VREF_Z_I[5] VSS VSS VDD VDD EN_VREF_Z_O[5] sky130_fd_sc_hd__or2_4
x2[4] EN_VSS_O[4] EN_VREF_Z_I[4] VSS VSS VDD VDD EN_VREF_Z_O[4] sky130_fd_sc_hd__or2_4
x2[3] EN_VSS_O[3] EN_VREF_Z_I[3] VSS VSS VDD VDD EN_VREF_Z_O[3] sky130_fd_sc_hd__or2_4
x2[2] EN_VSS_O[2] EN_VREF_Z_I[2] VSS VSS VDD VDD EN_VREF_Z_O[2] sky130_fd_sc_hd__or2_4
x2[1] EN_VSS_O[1] EN_VREF_Z_I[1] VSS VSS VDD VDD EN_VREF_Z_O[1] sky130_fd_sc_hd__or2_4
x2[0] EN_VSS_O[0] EN_VREF_Z_I[0] VSS VSS VDD VDD EN_VREF_Z_O[0] sky130_fd_sc_hd__or2_4
x1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_12
x2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
.ends


* expanding   symbol:  subcells/individual_switches/switch_VCM.sym # of pins=5
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_VCM.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_VCM.sch
.subckt switch_VCM VCM EN_VCM Cbtm VDD VSS
*.PININFO VCM:I EN_VCM:I Cbtm:O VSS:I VDD:I
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=64 nf=8 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C10.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C10.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C10.sch
.subckt switch_C10 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=2 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=64 nf=8 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=128 nf=16 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=64 nf=8 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C9.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C9.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C9.sch
.subckt switch_C9 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=32 nf=4 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=64 nf=8 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=32 nf=4 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C8.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C8.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C8.sch
.subckt switch_C8 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=2 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=32 nf=4 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=16 nf=2 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C7.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C7.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C7.sch
.subckt switch_C7 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=2 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C6.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C6.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C6.sch
.subckt switch_C6 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=8 nf=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C5.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C5.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C5.sch
.subckt switch_C5 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VREF_GND:I VREF:I VCM:I EN_VCM:I Cbtm:O VDD:I EN_VSS:I EN_VREF_Z:I VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C0_dummy.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C0_dummy.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C0_dummy.sch
.subckt switch_C0_dummy VCM VIN EN_VCM Cbtm EN_VIN VSS
*.PININFO VIN:I EN_VIN:I VCM:I EN_VCM:I Cbtm:O VSS:I
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
.ends

.end
