magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< error_p >>
rect -29 262 29 268
rect -29 228 -17 262
rect -29 222 29 228
rect -29 -228 29 -222
rect -29 -262 -17 -228
rect -29 -268 29 -262
<< pwell >>
rect -211 -400 211 400
<< nmoslvt >>
rect -15 -190 15 190
<< ndiff >>
rect -73 178 -15 190
rect -73 -178 -61 178
rect -27 -178 -15 178
rect -73 -190 -15 -178
rect 15 178 73 190
rect 15 -178 27 178
rect 61 -178 73 178
rect 15 -190 73 -178
<< ndiffc >>
rect -61 -178 -27 178
rect 27 -178 61 178
<< psubdiff >>
rect -175 330 -79 364
rect 79 330 175 364
rect -175 268 -141 330
rect 141 268 175 330
rect -175 -330 -141 -268
rect 141 -330 175 -268
rect -175 -364 -79 -330
rect 79 -364 175 -330
<< psubdiffcont >>
rect -79 330 79 364
rect -175 -268 -141 268
rect 141 -268 175 268
rect -79 -364 79 -330
<< poly >>
rect -33 262 33 278
rect -33 228 -17 262
rect 17 228 33 262
rect -33 212 33 228
rect -15 190 15 212
rect -15 -212 15 -190
rect -33 -228 33 -212
rect -33 -262 -17 -228
rect 17 -262 33 -228
rect -33 -278 33 -262
<< polycont >>
rect -17 228 17 262
rect -17 -262 17 -228
<< locali >>
rect -175 330 -79 364
rect 79 330 175 364
rect -175 268 -141 330
rect 141 268 175 330
rect -33 228 -17 262
rect 17 228 33 262
rect -61 178 -27 194
rect -61 -194 -27 -178
rect 27 178 61 194
rect 27 -194 61 -178
rect -33 -262 -17 -228
rect 17 -262 33 -228
rect -175 -330 -141 -268
rect 141 -330 175 -268
rect -175 -364 -79 -330
rect 79 -364 175 -330
<< viali >>
rect -17 228 17 262
rect -61 -178 -27 178
rect 27 -178 61 178
rect -17 -262 17 -228
<< metal1 >>
rect -29 262 29 268
rect -29 228 -17 262
rect 17 228 29 262
rect -29 222 29 228
rect -67 178 -21 190
rect -67 -178 -61 178
rect -27 -178 -21 178
rect -67 -190 -21 -178
rect 21 178 67 190
rect 21 -178 27 178
rect 61 -178 67 178
rect 21 -190 67 -178
rect -29 -228 29 -222
rect -29 -262 -17 -228
rect 17 -262 29 -228
rect -29 -268 29 -262
<< properties >>
string FIXED_BBOX -158 -347 158 347
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.9 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
