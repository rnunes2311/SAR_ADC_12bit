magic
tech sky130A
magscale 1 2
timestamp 1711310191
<< metal3 >>
rect -1086 1122 1086 1150
rect -1086 -1122 1002 1122
rect 1066 -1122 1086 1122
rect -1086 -1150 1086 -1122
<< via3 >>
rect 1002 -1122 1066 1122
<< mimcap >>
rect -1046 1070 754 1110
rect -1046 -1070 -1006 1070
rect 714 -1070 754 1070
rect -1046 -1110 754 -1070
<< mimcapcontact >>
rect -1006 -1070 714 1070
<< metal4 >>
rect 986 1122 1082 1138
rect -1007 1070 715 1071
rect -1007 -1070 -1006 1070
rect 714 -1070 715 1070
rect -1007 -1071 715 -1070
rect 986 -1122 1002 1122
rect 1066 -1122 1082 1122
rect 986 -1138 1082 -1122
<< properties >>
string FIXED_BBOX -1086 -1150 794 1150
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 9 l 11.1 val 207.438 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
