magic
tech sky130A
magscale 1 2
timestamp 1711995413
<< error_p >>
rect -77 123 -19 129
rect 115 123 173 129
rect -77 89 -65 123
rect 115 89 127 123
rect -77 83 -19 89
rect 115 83 173 89
rect -173 -89 -115 -83
rect 19 -89 77 -83
rect -173 -123 -161 -89
rect 19 -123 31 -89
rect -173 -129 -115 -123
rect 19 -129 77 -123
<< nwell >>
rect -359 -261 359 261
<< pmos >>
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
<< pdiff >>
rect -221 30 -159 42
rect -221 -30 -209 30
rect -175 -30 -159 30
rect -221 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 221 42
rect 159 -30 175 30
rect 209 -30 221 30
rect 159 -42 221 -30
<< pdiffc >>
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
<< nsubdiff >>
rect -323 191 -227 225
rect 227 191 323 225
rect -323 -191 -289 191
rect 289 129 323 191
rect 289 -191 323 -129
rect -323 -225 -227 -191
rect 227 -225 323 -191
<< nsubdiffcont >>
rect -227 191 227 225
rect 289 -129 323 129
rect -227 -225 227 -191
<< poly >>
rect -81 123 -15 139
rect -81 89 -65 123
rect -31 89 -15 123
rect -81 73 -15 89
rect 111 123 177 139
rect 111 89 127 123
rect 161 89 177 123
rect 111 73 177 89
rect -159 42 -129 68
rect -63 42 -33 73
rect 33 42 63 68
rect 129 42 159 73
rect -159 -73 -129 -42
rect -63 -68 -33 -42
rect 33 -73 63 -42
rect 129 -68 159 -42
rect -177 -89 -111 -73
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect -177 -139 -111 -123
rect 15 -89 81 -73
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 15 -139 81 -123
<< polycont >>
rect -65 89 -31 123
rect 127 89 161 123
rect -161 -123 -127 -89
rect 31 -123 65 -89
<< locali >>
rect -323 191 -227 225
rect 227 191 323 225
rect -323 -191 -289 191
rect 289 129 323 191
rect -81 89 -65 123
rect -31 89 -15 123
rect 111 89 127 123
rect 161 89 177 123
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect -177 -123 -161 -89
rect -127 -123 -111 -89
rect 15 -123 31 -89
rect 65 -123 81 -89
rect 289 -191 323 -129
rect -323 -225 -227 -191
rect 227 -225 323 -191
<< viali >>
rect -65 89 -31 123
rect 127 89 161 123
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect -161 -123 -127 -89
rect 31 -123 65 -89
<< metal1 >>
rect -77 123 -19 129
rect -77 89 -65 123
rect -31 89 -19 123
rect -77 83 -19 89
rect 115 123 173 129
rect 115 89 127 123
rect 161 89 173 123
rect 115 83 173 89
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect -173 -89 -115 -83
rect -173 -123 -161 -89
rect -127 -123 -115 -89
rect -173 -129 -115 -123
rect 19 -89 77 -83
rect 19 -123 31 -89
rect 65 -123 77 -89
rect 19 -129 77 -123
<< properties >>
string FIXED_BBOX -306 -208 306 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
