magic
tech sky130A
magscale 1 2
timestamp 1711801860
<< error_p >>
rect -749 872 -691 878
rect -557 872 -499 878
rect -365 872 -307 878
rect -173 872 -115 878
rect 19 872 77 878
rect 211 872 269 878
rect 403 872 461 878
rect 595 872 653 878
rect 787 872 845 878
rect -749 838 -737 872
rect -557 838 -545 872
rect -365 838 -353 872
rect -173 838 -161 872
rect 19 838 31 872
rect 211 838 223 872
rect 403 838 415 872
rect 595 838 607 872
rect 787 838 799 872
rect -749 832 -691 838
rect -557 832 -499 838
rect -365 832 -307 838
rect -173 832 -115 838
rect 19 832 77 838
rect 211 832 269 838
rect 403 832 461 838
rect 595 832 653 838
rect 787 832 845 838
rect -845 -838 -787 -832
rect -653 -838 -595 -832
rect -461 -838 -403 -832
rect -269 -838 -211 -832
rect -77 -838 -19 -832
rect 115 -838 173 -832
rect 307 -838 365 -832
rect 499 -838 557 -832
rect 691 -838 749 -832
rect -845 -872 -833 -838
rect -653 -872 -641 -838
rect -461 -872 -449 -838
rect -269 -872 -257 -838
rect -77 -872 -65 -838
rect 115 -872 127 -838
rect 307 -872 319 -838
rect 499 -872 511 -838
rect 691 -872 703 -838
rect -845 -878 -787 -872
rect -653 -878 -595 -872
rect -461 -878 -403 -872
rect -269 -878 -211 -872
rect -77 -878 -19 -872
rect 115 -878 173 -872
rect 307 -878 365 -872
rect 499 -878 557 -872
rect 691 -878 749 -872
<< pwell >>
rect -1031 -1010 5371 1010
<< nmos >>
rect -831 -800 -801 800
rect -735 -800 -705 800
rect -639 -800 -609 800
rect -543 -800 -513 800
rect -447 -800 -417 800
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
rect 417 -800 447 800
rect 513 -800 543 800
rect 609 -800 639 800
rect 705 -800 735 800
rect 801 -800 831 800
<< ndiff >>
rect -893 788 -831 800
rect -893 -788 -881 788
rect -847 -788 -831 788
rect -893 -800 -831 -788
rect -801 788 -735 800
rect -801 -788 -785 788
rect -751 -788 -735 788
rect -801 -800 -735 -788
rect -705 788 -639 800
rect -705 -788 -689 788
rect -655 -788 -639 788
rect -705 -800 -639 -788
rect -609 788 -543 800
rect -609 -788 -593 788
rect -559 -788 -543 788
rect -609 -800 -543 -788
rect -513 788 -447 800
rect -513 -788 -497 788
rect -463 -788 -447 788
rect -513 -800 -447 -788
rect -417 788 -351 800
rect -417 -788 -401 788
rect -367 -788 -351 788
rect -417 -800 -351 -788
rect -321 788 -255 800
rect -321 -788 -305 788
rect -271 -788 -255 788
rect -321 -800 -255 -788
rect -225 788 -159 800
rect -225 -788 -209 788
rect -175 -788 -159 788
rect -225 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 225 800
rect 159 -788 175 788
rect 209 -788 225 788
rect 159 -800 225 -788
rect 255 788 321 800
rect 255 -788 271 788
rect 305 -788 321 788
rect 255 -800 321 -788
rect 351 788 417 800
rect 351 -788 367 788
rect 401 -788 417 788
rect 351 -800 417 -788
rect 447 788 513 800
rect 447 -788 463 788
rect 497 -788 513 788
rect 447 -800 513 -788
rect 543 788 609 800
rect 543 -788 559 788
rect 593 -788 609 788
rect 543 -800 609 -788
rect 639 788 705 800
rect 639 -788 655 788
rect 689 -788 705 788
rect 639 -800 705 -788
rect 735 788 801 800
rect 735 -788 751 788
rect 785 -788 801 788
rect 735 -800 801 -788
rect 831 788 893 800
rect 831 -788 847 788
rect 881 -788 893 788
rect 831 -800 893 -788
<< ndiffc >>
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
<< psubdiff >>
rect -995 940 -899 974
rect 899 940 5335 974
rect -995 878 -961 940
rect 5301 878 5335 940
rect -995 -940 -961 -878
rect 5301 -940 5335 -878
rect -995 -974 -899 -940
rect 899 -974 5335 -940
<< psubdiffcont >>
rect -899 940 899 974
rect -995 -878 -961 878
rect 5301 -878 5335 878
rect -899 -974 899 -940
<< poly >>
rect -753 872 -687 888
rect -831 800 -801 857
rect -753 838 -737 872
rect -703 838 -687 872
rect -561 872 -495 888
rect -753 822 -687 838
rect -735 800 -705 822
rect -639 800 -609 858
rect -561 838 -545 872
rect -511 838 -495 872
rect -369 872 -303 888
rect -561 822 -495 838
rect -543 800 -513 822
rect -447 800 -417 856
rect -369 838 -353 872
rect -319 838 -303 872
rect -177 872 -111 888
rect -369 822 -303 838
rect -351 800 -321 822
rect -255 800 -225 857
rect -177 838 -161 872
rect -127 838 -111 872
rect 15 872 81 888
rect -177 822 -111 838
rect -159 800 -129 822
rect -63 800 -33 857
rect 15 838 31 872
rect 65 838 81 872
rect 207 872 273 888
rect 15 822 81 838
rect 33 800 63 822
rect 129 800 159 854
rect 207 838 223 872
rect 257 838 273 872
rect 399 872 465 888
rect 207 822 273 838
rect 225 800 255 822
rect 321 800 351 856
rect 399 838 415 872
rect 449 838 465 872
rect 591 872 657 888
rect 399 822 465 838
rect 417 800 447 822
rect 513 800 543 856
rect 591 838 607 872
rect 641 838 657 872
rect 783 872 849 888
rect 591 822 657 838
rect 609 800 639 822
rect 705 800 735 856
rect 783 838 799 872
rect 833 838 849 872
rect 783 822 849 838
rect 801 800 831 822
rect -831 -822 -801 -800
rect -849 -838 -783 -822
rect -735 -826 -705 -800
rect -639 -822 -609 -800
rect -849 -872 -833 -838
rect -799 -872 -783 -838
rect -849 -888 -783 -872
rect -657 -838 -591 -822
rect -543 -826 -513 -800
rect -447 -822 -417 -800
rect -657 -872 -641 -838
rect -607 -872 -591 -838
rect -657 -888 -591 -872
rect -465 -838 -399 -822
rect -351 -826 -321 -800
rect -255 -822 -225 -800
rect -465 -872 -449 -838
rect -415 -872 -399 -838
rect -465 -888 -399 -872
rect -273 -838 -207 -822
rect -159 -826 -129 -800
rect -63 -822 -33 -800
rect -273 -872 -257 -838
rect -223 -872 -207 -838
rect -273 -888 -207 -872
rect -81 -838 -15 -822
rect 33 -826 63 -800
rect 129 -822 159 -800
rect -81 -872 -65 -838
rect -31 -872 -15 -838
rect -81 -888 -15 -872
rect 111 -838 177 -822
rect 225 -826 255 -800
rect 321 -822 351 -800
rect 111 -872 127 -838
rect 161 -872 177 -838
rect 111 -888 177 -872
rect 303 -838 369 -822
rect 417 -826 447 -800
rect 513 -822 543 -800
rect 303 -872 319 -838
rect 353 -872 369 -838
rect 303 -888 369 -872
rect 495 -838 561 -822
rect 609 -826 639 -800
rect 705 -822 735 -800
rect 495 -872 511 -838
rect 545 -872 561 -838
rect 495 -888 561 -872
rect 687 -838 753 -822
rect 801 -826 831 -800
rect 687 -872 703 -838
rect 737 -872 753 -838
rect 687 -888 753 -872
<< polycont >>
rect -737 838 -703 872
rect -545 838 -511 872
rect -353 838 -319 872
rect -161 838 -127 872
rect 31 838 65 872
rect 223 838 257 872
rect 415 838 449 872
rect 607 838 641 872
rect 799 838 833 872
rect -833 -872 -799 -838
rect -641 -872 -607 -838
rect -449 -872 -415 -838
rect -257 -872 -223 -838
rect -65 -872 -31 -838
rect 127 -872 161 -838
rect 319 -872 353 -838
rect 511 -872 545 -838
rect 703 -872 737 -838
<< locali >>
rect -995 940 -899 974
rect 899 940 5335 974
rect -995 878 -961 940
rect 5301 878 5335 940
rect -753 838 -737 872
rect -703 838 -687 872
rect -561 838 -545 872
rect -511 838 -495 872
rect -369 838 -353 872
rect -319 838 -303 872
rect -177 838 -161 872
rect -127 838 -111 872
rect 15 838 31 872
rect 65 838 81 872
rect 207 838 223 872
rect 257 838 273 872
rect 399 838 415 872
rect 449 838 465 872
rect 591 838 607 872
rect 641 838 657 872
rect 783 838 799 872
rect 833 838 849 872
rect -881 788 -847 804
rect -881 -804 -847 -788
rect -785 788 -751 804
rect -785 -804 -751 -788
rect -689 788 -655 804
rect -689 -804 -655 -788
rect -593 788 -559 804
rect -593 -804 -559 -788
rect -497 788 -463 804
rect -497 -804 -463 -788
rect -401 788 -367 804
rect -401 -804 -367 -788
rect -305 788 -271 804
rect -305 -804 -271 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 271 788 305 804
rect 271 -804 305 -788
rect 367 788 401 804
rect 367 -804 401 -788
rect 463 788 497 804
rect 463 -804 497 -788
rect 559 788 593 804
rect 559 -804 593 -788
rect 655 788 689 804
rect 655 -804 689 -788
rect 751 788 785 804
rect 751 -804 785 -788
rect 847 788 881 804
rect 847 -804 881 -788
rect -849 -872 -833 -838
rect -799 -872 -783 -838
rect -657 -872 -641 -838
rect -607 -872 -591 -838
rect -465 -872 -449 -838
rect -415 -872 -399 -838
rect -273 -872 -257 -838
rect -223 -872 -207 -838
rect -81 -872 -65 -838
rect -31 -872 -15 -838
rect 111 -872 127 -838
rect 161 -872 177 -838
rect 303 -872 319 -838
rect 353 -872 369 -838
rect 495 -872 511 -838
rect 545 -872 561 -838
rect 687 -872 703 -838
rect 737 -872 753 -838
rect -995 -940 -961 -878
rect 5301 -940 5335 -878
rect -995 -974 -899 -940
rect 899 -974 5335 -940
<< viali >>
rect -737 838 -703 872
rect -545 838 -511 872
rect -353 838 -319 872
rect -161 838 -127 872
rect 31 838 65 872
rect 223 838 257 872
rect 415 838 449 872
rect 607 838 641 872
rect 799 838 833 872
rect -881 -788 -847 788
rect -785 -788 -751 788
rect -689 -788 -655 788
rect -593 -788 -559 788
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect 559 -788 593 788
rect 655 -788 689 788
rect 751 -788 785 788
rect 847 -788 881 788
rect -833 -872 -799 -838
rect -641 -872 -607 -838
rect -449 -872 -415 -838
rect -257 -872 -223 -838
rect -65 -872 -31 -838
rect 127 -872 161 -838
rect 319 -872 353 -838
rect 511 -872 545 -838
rect 703 -872 737 -838
<< metal1 >>
rect -749 872 -691 878
rect -749 838 -737 872
rect -703 838 -691 872
rect -749 832 -691 838
rect -557 872 -499 878
rect -557 838 -545 872
rect -511 838 -499 872
rect -557 832 -499 838
rect -365 872 -307 878
rect -365 838 -353 872
rect -319 838 -307 872
rect -365 832 -307 838
rect -173 872 -115 878
rect -173 838 -161 872
rect -127 838 -115 872
rect -173 832 -115 838
rect 19 872 77 878
rect 19 838 31 872
rect 65 838 77 872
rect 19 832 77 838
rect 211 872 269 878
rect 211 838 223 872
rect 257 838 269 872
rect 211 832 269 838
rect 403 872 461 878
rect 403 838 415 872
rect 449 838 461 872
rect 403 832 461 838
rect 595 872 653 878
rect 595 838 607 872
rect 641 838 653 872
rect 595 832 653 838
rect 787 872 845 878
rect 787 838 799 872
rect 833 838 845 872
rect 787 832 845 838
rect -887 788 -841 800
rect -887 -788 -881 788
rect -847 -788 -841 788
rect -887 -800 -841 -788
rect -791 788 -745 800
rect -791 -788 -785 788
rect -751 -788 -745 788
rect -791 -800 -745 -788
rect -695 788 -649 800
rect -695 -788 -689 788
rect -655 -788 -649 788
rect -695 -800 -649 -788
rect -599 788 -553 800
rect -599 -788 -593 788
rect -559 -788 -553 788
rect -599 -800 -553 -788
rect -503 788 -457 800
rect -503 -788 -497 788
rect -463 -788 -457 788
rect -503 -800 -457 -788
rect -407 788 -361 800
rect -407 -788 -401 788
rect -367 -788 -361 788
rect -407 -800 -361 -788
rect -311 788 -265 800
rect -311 -788 -305 788
rect -271 -788 -265 788
rect -311 -800 -265 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 265 788 311 800
rect 265 -788 271 788
rect 305 -788 311 788
rect 265 -800 311 -788
rect 361 788 407 800
rect 361 -788 367 788
rect 401 -788 407 788
rect 361 -800 407 -788
rect 457 788 503 800
rect 457 -788 463 788
rect 497 -788 503 788
rect 457 -800 503 -788
rect 553 788 599 800
rect 553 -788 559 788
rect 593 -788 599 788
rect 553 -800 599 -788
rect 649 788 695 800
rect 649 -788 655 788
rect 689 -788 695 788
rect 649 -800 695 -788
rect 745 788 791 800
rect 745 -788 751 788
rect 785 -788 791 788
rect 745 -800 791 -788
rect 841 788 887 800
rect 841 -788 847 788
rect 881 -788 887 788
rect 841 -800 887 -788
rect -845 -838 -787 -832
rect -845 -872 -833 -838
rect -799 -872 -787 -838
rect -845 -878 -787 -872
rect -653 -838 -595 -832
rect -653 -872 -641 -838
rect -607 -872 -595 -838
rect -653 -878 -595 -872
rect -461 -838 -403 -832
rect -461 -872 -449 -838
rect -415 -872 -403 -838
rect -461 -878 -403 -872
rect -269 -838 -211 -832
rect -269 -872 -257 -838
rect -223 -872 -211 -838
rect -269 -878 -211 -872
rect -77 -838 -19 -832
rect -77 -872 -65 -838
rect -31 -872 -19 -838
rect -77 -878 -19 -872
rect 115 -838 173 -832
rect 115 -872 127 -838
rect 161 -872 173 -838
rect 115 -878 173 -872
rect 307 -838 365 -832
rect 307 -872 319 -838
rect 353 -872 365 -838
rect 307 -878 365 -872
rect 499 -838 557 -832
rect 499 -872 511 -838
rect 545 -872 557 -838
rect 499 -878 557 -872
rect 691 -838 749 -832
rect 691 -872 703 -838
rect 737 -872 749 -838
rect 691 -878 749 -872
<< properties >>
string FIXED_BBOX -978 -957 978 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.150 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
