magic
tech sky130A
magscale 1 2
timestamp 1715417500
<< nwell >>
rect 15679 1323 15712 2253
rect 15638 1203 16023 1323
rect 15679 1140 15909 1203
rect 15679 714 15930 1140
rect 20034 964 20299 1107
rect 15690 610 15930 714
rect 19994 870 20299 964
rect 19994 696 20298 870
rect 15900 560 15930 610
<< pwell >>
rect 19479 1204 19973 1304
rect 19479 1022 19966 1204
rect 19468 135 19816 340
rect 19468 84 20249 135
rect 19501 83 20249 84
<< psubdiff >>
rect 19515 1234 19539 1268
rect 19945 1234 19969 1268
rect 19524 96 19553 130
rect 20139 96 20168 130
<< nsubdiff >>
rect 20074 910 20164 940
rect 20074 690 20164 781
<< psubdiffcont >>
rect 19539 1234 19945 1268
rect 19553 96 20139 130
<< nsubdiffcont >>
rect 20074 781 20164 910
<< poly >>
rect 16106 1129 16442 1200
<< locali >>
rect 19523 1234 19539 1268
rect 19945 1234 19961 1268
rect 19560 964 19594 1002
rect 19869 967 19907 1001
rect 20054 910 20183 931
rect 20054 781 20074 910
rect 20164 781 20183 910
rect 20054 698 20183 781
rect 19593 685 20183 698
rect 19593 664 20149 685
rect 19536 358 19574 392
rect 19688 352 19862 402
rect 20190 352 20224 390
rect 16830 120 16900 160
rect 17994 120 18204 160
rect 19404 154 19444 160
rect 19404 153 19539 154
rect 19404 130 19567 153
rect 19404 127 19553 130
rect 19404 122 19528 127
rect 19404 120 19553 122
rect 19501 119 19553 120
rect 19507 96 19553 119
rect 20139 96 20207 122
<< viali >>
rect 12499 2183 15466 2217
rect 16100 1272 16500 1306
rect 19560 1002 19594 1038
rect 9281 301 9315 980
rect 15626 315 15660 994
rect 16553 307 16587 986
rect 19833 967 19869 1001
rect 19907 967 19943 1001
rect 19560 928 19594 964
rect 19500 358 19536 392
rect 19574 358 19610 392
rect 20190 390 20224 426
rect 20190 316 20224 352
rect 12508 120 15475 154
rect 16110 120 16510 154
rect 16900 120 17994 160
rect 18204 120 19404 160
<< metal1 >>
rect 9245 2217 15690 2254
rect 9245 2183 12499 2217
rect 15466 2183 15690 2217
rect 9245 2157 15690 2183
rect 9245 1868 9342 2157
rect 9980 2050 9990 2120
rect 10050 2050 10080 2120
rect 10140 2050 10150 2120
rect 11770 2050 11780 2120
rect 11840 2050 11870 2120
rect 11930 2050 11940 2120
rect 12950 2050 12960 2120
rect 13020 2050 13050 2120
rect 13110 2050 13120 2120
rect 15220 2060 15230 2120
rect 15290 2060 15330 2120
rect 15390 2060 15400 2120
rect 15591 1868 15690 2157
rect 9245 1439 15690 1868
rect 9245 980 9342 1439
rect 15591 1322 15690 1439
rect 15591 1306 16624 1322
rect 15591 1272 16100 1306
rect 16500 1272 16624 1306
rect 15591 1266 16624 1272
rect 9464 1140 12425 1226
rect 12533 1140 15494 1229
rect 15591 1225 16157 1266
rect 16470 1225 16624 1266
rect 15591 1140 16003 1225
rect 16230 1193 16291 1203
rect 16189 1144 16230 1190
rect 9445 1130 15496 1140
rect 9445 1094 9995 1130
rect 10056 1094 10089 1130
rect 9995 1068 10056 1078
rect 10150 1094 11775 1130
rect 10089 1068 10150 1078
rect 11836 1094 11869 1130
rect 11775 1068 11836 1078
rect 11930 1094 12955 1130
rect 11869 1068 11930 1078
rect 13016 1094 13049 1130
rect 12955 1068 13016 1078
rect 13110 1094 15225 1130
rect 13049 1068 13110 1078
rect 15286 1094 15319 1130
rect 15225 1068 15286 1078
rect 15380 1094 15496 1130
rect 15319 1068 15380 1078
rect 9245 301 9281 980
rect 9315 864 9342 980
rect 15591 994 15690 1140
rect 15829 1038 15839 1099
rect 15891 1038 15901 1099
rect 15840 1005 15890 1038
rect 15591 864 15626 994
rect 9315 435 15626 864
rect 9315 301 9342 435
rect 9245 185 9342 301
rect 15591 315 15626 435
rect 15660 652 15690 994
rect 15829 944 15839 1005
rect 15891 944 15901 1005
rect 15660 474 15688 652
rect 15660 326 15748 474
rect 15840 350 15890 944
rect 15930 560 16003 1140
rect 16324 1193 16385 1203
rect 16291 1144 16324 1190
rect 16230 1131 16291 1141
rect 16385 1144 16428 1190
rect 16324 1131 16385 1141
rect 16527 986 16624 1225
rect 16141 696 16151 757
rect 16203 696 16213 757
rect 16333 696 16343 757
rect 16395 696 16405 757
rect 16141 602 16151 663
rect 16203 602 16213 663
rect 16333 602 16343 663
rect 16395 602 16405 663
rect 15932 552 16003 560
rect 15932 551 16104 552
rect 15932 490 16047 551
rect 16099 490 16109 551
rect 16229 490 16239 551
rect 16291 490 16301 551
rect 16421 490 16431 551
rect 16483 490 16493 551
rect 15932 457 16104 490
rect 15932 396 16047 457
rect 16099 396 16109 457
rect 16229 396 16239 457
rect 16291 396 16301 457
rect 16421 396 16431 457
rect 16483 396 16493 457
rect 15660 315 15688 326
rect 9993 278 10054 288
rect 9445 226 9993 262
rect 10087 278 10148 288
rect 10054 226 10087 262
rect 11765 278 11826 288
rect 10148 226 11765 262
rect 11859 278 11920 288
rect 11826 226 11859 262
rect 12945 278 13006 288
rect 11920 226 12945 262
rect 13039 278 13100 288
rect 13006 226 13039 262
rect 15221 276 15282 286
rect 13100 226 15221 262
rect 9445 224 15221 226
rect 15315 276 15376 286
rect 15282 224 15315 262
rect 15376 224 15496 262
rect 9445 216 15496 224
rect 15221 214 15282 216
rect 15315 214 15376 216
rect 15591 185 15688 315
rect 15723 265 15784 275
rect 15723 203 15784 213
rect 15817 265 15878 275
rect 15817 203 15878 213
rect 9245 167 15688 185
rect 15932 185 16003 396
rect 16527 307 16553 986
rect 16587 307 16624 986
rect 16527 185 16624 307
rect 15932 167 16624 185
rect 9245 154 16624 167
rect 9245 120 12508 154
rect 15475 120 16110 154
rect 16510 120 16624 154
rect 9245 88 16624 120
rect 16790 1306 19984 1388
rect 16790 185 16868 1306
rect 16986 1243 17396 1264
rect 16986 1191 17116 1243
rect 17177 1191 17210 1243
rect 17271 1191 17396 1243
rect 16986 1168 17396 1191
rect 17155 992 17165 1053
rect 17217 992 17227 1053
rect 17155 898 17165 959
rect 17217 898 17227 959
rect 16917 664 16927 725
rect 16979 664 16989 725
rect 17393 664 17403 725
rect 17455 664 17465 725
rect 16917 570 16927 631
rect 16979 570 16989 631
rect 17393 570 17403 631
rect 17455 570 17465 631
rect 17526 185 17614 1306
rect 17655 1243 17974 1264
rect 17655 1191 17785 1243
rect 17846 1191 17879 1243
rect 17940 1191 17974 1243
rect 17655 1162 17974 1191
rect 18040 1234 19984 1306
rect 18040 1050 18198 1234
rect 18312 1184 18467 1194
rect 18373 1132 18406 1184
rect 18312 1122 18467 1132
rect 17665 666 17675 727
rect 17727 666 17737 727
rect 17665 572 17675 633
rect 17727 572 17737 633
rect 17903 468 17913 529
rect 17965 468 17975 529
rect 17903 374 17913 435
rect 17965 374 17975 435
rect 18040 366 18278 1050
rect 18343 992 18353 1053
rect 18405 992 18415 1053
rect 18558 1050 18622 1234
rect 18343 898 18353 959
rect 18405 898 18415 959
rect 18040 185 18198 366
rect 18476 364 18622 1050
rect 18981 1004 19043 1234
rect 19149 1184 19304 1194
rect 19210 1132 19243 1184
rect 19149 1122 19304 1132
rect 19370 1004 19459 1234
rect 19536 1024 19546 1085
rect 19598 1024 19608 1085
rect 18773 828 18783 889
rect 18835 828 18845 889
rect 18773 734 18783 795
rect 18835 734 18845 795
rect 18669 575 18679 636
rect 18731 575 18741 636
rect 18867 575 18877 636
rect 18929 575 18939 636
rect 18669 481 18679 542
rect 18731 481 18741 542
rect 18867 481 18877 542
rect 18929 481 18939 542
rect 18558 185 18622 364
rect 18981 357 19125 1004
rect 19183 818 19193 879
rect 19245 818 19255 879
rect 19183 724 19193 785
rect 19245 724 19255 785
rect 18727 256 18788 266
rect 18727 194 18788 204
rect 18821 256 18882 266
rect 18821 194 18882 204
rect 16790 166 18622 185
rect 18981 185 19043 357
rect 19321 351 19459 1004
rect 19554 1002 19560 1024
rect 19594 1002 19600 1024
rect 19830 1012 19891 1022
rect 19554 991 19600 1002
rect 19536 930 19546 991
rect 19598 930 19608 991
rect 19821 961 19830 1007
rect 19924 1012 19985 1022
rect 19891 1001 19924 1007
rect 19891 967 19907 1001
rect 19891 961 19924 967
rect 19830 950 19891 960
rect 19924 950 19985 960
rect 19554 928 19560 930
rect 19594 928 19600 930
rect 19554 916 19600 928
rect 19573 644 19583 718
rect 20158 644 20168 718
rect 20185 438 20195 459
rect 20184 426 20195 438
rect 19497 404 19558 414
rect 19488 352 19497 398
rect 19591 404 19652 414
rect 19558 392 19591 398
rect 19558 358 19574 392
rect 19558 352 19591 358
rect 19370 185 19459 351
rect 19497 342 19558 352
rect 19591 342 19652 352
rect 20184 390 20190 426
rect 20247 398 20257 459
rect 20224 390 20230 398
rect 20184 365 20230 390
rect 20184 352 20195 365
rect 20184 316 20190 352
rect 20184 304 20195 316
rect 20247 304 20257 365
rect 18981 166 19551 185
rect 16790 160 19551 166
rect 16790 159 16900 160
rect 17994 159 18204 160
rect 19404 159 19551 160
rect 16790 99 16833 159
rect 19424 120 19551 159
rect 19568 120 19578 158
rect 19424 99 19578 120
rect 16790 96 19578 99
rect 20174 96 20184 158
rect 16790 89 19598 96
<< via1 >>
rect 9990 2050 10050 2120
rect 10080 2050 10140 2120
rect 11780 2050 11840 2120
rect 11870 2050 11930 2120
rect 12960 2050 13020 2120
rect 13050 2050 13110 2120
rect 15230 2060 15290 2120
rect 15330 2060 15390 2120
rect 9995 1078 10056 1130
rect 10089 1078 10150 1130
rect 11775 1078 11836 1130
rect 11869 1078 11930 1130
rect 12955 1078 13016 1130
rect 13049 1078 13110 1130
rect 15225 1078 15286 1130
rect 15319 1078 15380 1130
rect 15839 1038 15891 1099
rect 15839 944 15891 1005
rect 16230 1141 16291 1193
rect 16324 1141 16385 1193
rect 16151 696 16203 757
rect 16343 696 16395 757
rect 16151 602 16203 663
rect 16343 602 16395 663
rect 16047 490 16099 551
rect 16239 490 16291 551
rect 16431 490 16483 551
rect 16047 396 16099 457
rect 16239 396 16291 457
rect 16431 396 16483 457
rect 9993 226 10054 278
rect 10087 226 10148 278
rect 11765 226 11826 278
rect 11859 226 11920 278
rect 12945 226 13006 278
rect 13039 226 13100 278
rect 15221 224 15282 276
rect 15315 224 15376 276
rect 15723 213 15784 265
rect 15817 213 15878 265
rect 17116 1191 17177 1243
rect 17210 1191 17271 1243
rect 17165 992 17217 1053
rect 17165 898 17217 959
rect 16927 664 16979 725
rect 17403 664 17455 725
rect 16927 570 16979 631
rect 17403 570 17455 631
rect 17785 1191 17846 1243
rect 17879 1191 17940 1243
rect 18312 1132 18373 1184
rect 18406 1132 18467 1184
rect 17675 666 17727 727
rect 17675 572 17727 633
rect 17913 468 17965 529
rect 17913 374 17965 435
rect 18353 992 18405 1053
rect 18353 898 18405 959
rect 19149 1132 19210 1184
rect 19243 1132 19304 1184
rect 19546 1038 19598 1085
rect 19546 1024 19560 1038
rect 19560 1024 19594 1038
rect 19594 1024 19598 1038
rect 18783 828 18835 889
rect 18783 734 18835 795
rect 18679 575 18731 636
rect 18877 575 18929 636
rect 18679 481 18731 542
rect 18877 481 18929 542
rect 19193 818 19245 879
rect 19193 724 19245 785
rect 18727 204 18788 256
rect 18821 204 18882 256
rect 19546 964 19598 991
rect 19546 930 19560 964
rect 19560 930 19594 964
rect 19594 930 19598 964
rect 19830 1001 19891 1012
rect 19924 1001 19985 1012
rect 19830 967 19833 1001
rect 19833 967 19869 1001
rect 19869 967 19891 1001
rect 19924 967 19943 1001
rect 19943 967 19985 1001
rect 19830 960 19891 967
rect 19924 960 19985 967
rect 19583 644 20158 718
rect 20195 426 20247 459
rect 19497 392 19558 404
rect 19591 392 19652 404
rect 19497 358 19500 392
rect 19500 358 19536 392
rect 19536 358 19558 392
rect 19591 358 19610 392
rect 19610 358 19652 392
rect 19497 352 19558 358
rect 19591 352 19652 358
rect 20195 398 20224 426
rect 20224 398 20247 426
rect 20195 352 20247 365
rect 20195 316 20224 352
rect 20224 316 20247 352
rect 20195 304 20247 316
rect 16833 120 16900 159
rect 16900 120 17994 159
rect 17994 120 18204 159
rect 18204 120 19404 159
rect 19404 120 19424 159
rect 16833 99 19424 120
rect 19578 96 20174 158
<< metal2 >>
rect 9990 2120 10050 2130
rect 10080 2120 10140 2130
rect 10050 2050 10080 2090
rect 9990 2040 10140 2050
rect 11780 2120 11840 2130
rect 11870 2120 11930 2130
rect 11840 2050 11870 2090
rect 11780 2040 11930 2050
rect 12960 2120 13020 2130
rect 13050 2120 13110 2130
rect 13020 2050 13050 2100
rect 15230 2120 15390 2130
rect 15290 2060 15330 2120
rect 15230 2050 15390 2060
rect 12960 2040 13110 2050
rect 10020 1130 10120 2040
rect 11780 1130 11880 2040
rect 12970 1130 13070 2040
rect 15240 1130 15340 2050
rect 15618 1265 20168 1388
rect 15618 1212 16157 1265
rect 16470 1243 20168 1265
rect 16470 1212 17116 1243
rect 9985 1078 9995 1130
rect 10056 1078 10089 1130
rect 10150 1078 10160 1130
rect 11765 1078 11775 1130
rect 11836 1078 11869 1130
rect 11930 1078 11940 1130
rect 12945 1078 12955 1130
rect 13016 1078 13049 1130
rect 13110 1078 13120 1130
rect 15215 1078 15225 1130
rect 15286 1078 15319 1130
rect 15380 1078 15390 1130
rect 15850 1109 15880 1212
rect 16194 1141 16230 1193
rect 16291 1141 16324 1193
rect 16385 1170 16395 1193
rect 17106 1191 17116 1212
rect 17177 1191 17210 1243
rect 17271 1212 17785 1243
rect 17271 1191 17281 1212
rect 17775 1191 17785 1212
rect 17846 1191 17879 1243
rect 17940 1212 20168 1243
rect 17940 1191 17950 1212
rect 19768 1187 19968 1212
rect 16385 1141 16946 1170
rect 16194 1133 16946 1141
rect 18264 1133 18312 1184
rect 16194 1132 18312 1133
rect 18373 1132 18406 1184
rect 18467 1170 18477 1184
rect 19139 1170 19149 1184
rect 18467 1132 19149 1170
rect 19210 1132 19243 1184
rect 19304 1170 19314 1184
rect 19304 1132 19584 1170
rect 16194 1130 19584 1132
rect 15839 1099 15891 1109
rect 10020 278 10120 1078
rect 11780 278 11880 1078
rect 12970 278 13070 1078
rect 15240 850 15340 1078
rect 16897 1093 18312 1130
rect 19554 1095 19584 1130
rect 19546 1085 19598 1095
rect 15839 1005 15891 1038
rect 15839 934 15891 944
rect 17165 1053 17217 1063
rect 18353 1053 18405 1063
rect 17217 992 18353 1004
rect 17165 959 18405 992
rect 17217 956 18353 959
rect 17165 888 17217 898
rect 19546 991 19598 1024
rect 19546 920 19598 930
rect 19819 1012 20019 1078
rect 19819 960 19830 1012
rect 19891 960 19924 1012
rect 19985 960 20019 1012
rect 18353 888 18405 898
rect 18783 889 18835 899
rect 15240 828 18783 850
rect 19193 879 19245 889
rect 18835 828 19193 850
rect 15240 818 19193 828
rect 19819 878 20019 960
rect 15240 800 19245 818
rect 9983 226 9993 278
rect 10054 226 10087 278
rect 10148 226 10158 278
rect 11755 226 11765 278
rect 11826 226 11859 278
rect 11920 226 11930 278
rect 12935 226 12945 278
rect 13006 226 13039 278
rect 13100 226 13110 278
rect 15240 276 15340 800
rect 18783 795 18835 800
rect 16151 757 16203 767
rect 16343 757 16395 767
rect 16203 696 16343 700
rect 16840 725 17040 740
rect 16840 700 16927 725
rect 16395 696 16927 700
rect 16151 686 16927 696
rect 15936 664 16927 686
rect 16979 700 17040 725
rect 17403 725 17455 735
rect 16979 664 17403 700
rect 17675 727 17727 737
rect 17455 666 17675 700
rect 18783 724 18835 734
rect 19193 785 19245 800
rect 20076 728 20167 1212
rect 19193 714 19245 724
rect 19583 718 20167 728
rect 17455 664 17727 666
rect 15936 663 17727 664
rect 15936 654 16151 663
rect 15211 224 15221 276
rect 15282 224 15315 276
rect 15376 224 15386 276
rect 15713 213 15723 265
rect 15784 213 15817 265
rect 15878 257 15888 265
rect 15936 257 15968 654
rect 16203 648 16343 663
rect 16151 592 16203 602
rect 16395 648 17727 663
rect 16343 592 16395 602
rect 16840 631 17040 648
rect 16840 570 16927 631
rect 16979 570 17040 631
rect 16047 551 16099 561
rect 16239 551 16291 561
rect 16099 490 16239 494
rect 16431 551 16483 561
rect 16291 490 16431 494
rect 16840 540 17040 570
rect 17403 631 17455 648
rect 17403 560 17455 570
rect 17675 633 17727 648
rect 18708 646 18908 660
rect 17675 562 17727 572
rect 18679 636 18929 646
rect 18731 575 18877 636
rect 20158 644 20167 718
rect 19583 634 20167 644
rect 18679 542 18929 575
rect 16047 457 16483 490
rect 16099 442 16239 457
rect 16047 386 16099 396
rect 16291 442 16431 457
rect 16239 386 16291 396
rect 16431 386 16483 396
rect 17913 529 17965 539
rect 18731 481 18877 542
rect 18679 471 18929 481
rect 17913 435 17965 468
rect 18708 460 18908 471
rect 20113 459 20313 479
rect 17965 374 19497 404
rect 17913 364 19497 374
rect 17914 352 19497 364
rect 19558 352 19591 404
rect 19652 352 19662 404
rect 20113 398 20195 459
rect 20247 398 20313 459
rect 20113 365 20313 398
rect 15878 256 18717 257
rect 15878 225 18727 256
rect 15878 213 15888 225
rect 18717 204 18727 225
rect 18788 204 18821 256
rect 18882 204 18892 256
rect 19801 170 20001 347
rect 20113 304 20195 365
rect 20247 304 20313 365
rect 20113 279 20313 304
rect 16787 159 20260 170
rect 16787 99 16833 159
rect 19424 158 20260 159
rect 19424 99 19578 158
rect 16787 96 19578 99
rect 20174 96 20260 158
rect 16787 77 20260 96
use sky130_fd_pr__pfet_01v8_7FRQHJ  sky130_fd_pr__pfet_01v8_7FRQHJ_0
timestamp 1711831168
transform 1 0 12471 0 1 1171
box -3225 -1087 3225 1087
use sky130_fd_pr__pfet_01v8_XG6TDL  sky130_fd_pr__pfet_01v8_XG6TDL_0
timestamp 1710675123
transform 1 0 16265 0 1 703
box -359 -619 359 619
use sky130_fd_sc_hd__inv_4  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 19984 0 -1 1225
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19524 0 1 137
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x3
timestamp 1710522493
transform 1 0 19800 0 1 137
box -38 -48 498 592
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1710675955
transform 1 0 15801 0 1 403
box -211 -319 211 319
use sky130_fd_pr__nfet_05v0_nvt_F93ZEE  XM3
timestamp 1715417500
transform 1 0 17191 0 1 730
box -437 -658 441 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM4
timestamp 1710677421
transform 1 0 18383 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_01v8_6EHS5V  XM5
timestamp 1710677421
transform 1 0 19223 0 1 694
box -263 -610 263 610
use sky130_fd_pr__nfet_05v0_nvt_JFFQEL  XM7
timestamp 1710675123
transform 1 0 17820 0 1 730
box -318 -658 318 658
use sky130_fd_pr__nfet_01v8_6EHS5V  XM8
timestamp 1710677421
transform 1 0 18803 0 -1 694
box -263 -610 263 610
<< labels >>
flabel metal2 15707 1286 15763 1337 0 FreeSans 800 0 0 0 VDD
flabel metal1 11070 600 11130 660 0 FreeSans 800 0 0 0 Vtop
flabel metal2 16238 666 16278 688 0 FreeSans 800 0 0 0 Vgate
flabel metal1 11069 1604 11129 1664 0 FreeSans 800 0 0 0 Vtop
flabel metal2 16840 540 17040 740 0 FreeSans 256 0 0 0 VGATE
port 5 nsew
flabel metal2 17806 968 17830 982 0 FreeSans 800 0 0 0 Vd
flabel metal2 18620 360 18650 390 0 FreeSans 800 0 0 0 VGATE_1V8
flabel metal2 18978 810 19010 829 0 FreeSans 800 0 0 0 Vbottom
flabel metal2 19071 1141 19097 1157 0 FreeSans 800 0 0 0 EN_Z
flabel metal2 19819 878 20019 1078 0 FreeSans 256 0 0 0 EN
port 4 nsew
flabel metal2 20113 279 20313 479 0 FreeSans 256 0 0 0 SW_ON
port 3 nsew
flabel metal2 18708 460 18908 660 0 FreeSans 256 0 0 0 VIN
port 2 nsew
flabel metal2 19801 147 20001 347 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal2 19768 1187 19968 1387 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
