magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< pwell >>
rect -437 -658 441 658
<< mvnnmos >>
rect -209 -400 -29 400
rect 29 -400 209 400
<< mvndiff >>
rect -267 388 -209 400
rect -267 -388 -255 388
rect -221 -388 -209 388
rect -267 -400 -209 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 209 388 267 400
rect 209 -388 221 388
rect 255 -388 267 388
rect 209 -400 267 -388
<< mvndiffc >>
rect -255 -388 -221 388
rect -17 -388 17 388
rect 221 -388 255 388
<< mvpsubdiff >>
rect -401 610 405 622
rect -401 576 -293 610
rect 293 576 405 610
rect -401 564 405 576
rect -401 514 -343 564
rect -401 -514 -389 514
rect -355 -514 -343 514
rect 347 514 405 564
rect -401 -564 -343 -514
rect 347 -514 359 514
rect 393 -514 405 514
rect 347 -564 405 -514
rect -401 -576 405 -564
rect -401 -610 -293 -576
rect 293 -610 405 -576
rect -401 -622 405 -610
<< mvpsubdiffcont >>
rect -293 576 293 610
rect -389 -514 -355 514
rect 359 -514 393 514
rect -293 -610 293 -576
<< poly >>
rect -209 472 -29 488
rect -209 438 -193 472
rect -45 438 -29 472
rect -209 400 -29 438
rect 29 472 209 488
rect 29 438 45 472
rect 193 438 209 472
rect 29 400 209 438
rect -209 -438 -29 -400
rect -209 -472 -193 -438
rect -45 -472 -29 -438
rect -209 -488 -29 -472
rect 29 -438 209 -400
rect 29 -472 45 -438
rect 193 -472 209 -438
rect 29 -488 209 -472
<< polycont >>
rect -193 438 -45 472
rect 45 438 193 472
rect -193 -472 -45 -438
rect 45 -472 193 -438
<< locali >>
rect -389 576 -293 610
rect 293 576 393 610
rect -389 514 -355 576
rect 359 514 393 576
rect -209 438 -193 472
rect -45 438 -29 472
rect 29 438 45 472
rect 193 438 209 472
rect -255 388 -221 404
rect -255 -404 -221 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 221 388 255 404
rect 221 -404 255 -388
rect -209 -472 -193 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 193 -472 209 -438
rect -389 -576 -355 -514
rect 359 -576 393 -514
rect -389 -610 -293 -576
rect 293 -610 393 -576
<< viali >>
rect -193 438 -45 472
rect 45 438 193 472
rect -255 -388 -221 388
rect -17 -388 17 388
rect 221 -388 255 388
rect -193 -472 -45 -438
rect 45 -472 193 -438
<< metal1 >>
rect -205 472 -33 478
rect -205 438 -193 472
rect -45 438 -33 472
rect -205 432 -33 438
rect 33 472 205 478
rect 33 438 45 472
rect 193 438 205 472
rect 33 432 205 438
rect -261 388 -215 400
rect -261 -388 -255 388
rect -221 -388 -215 388
rect -261 -400 -215 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 215 388 261 400
rect 215 -388 221 388
rect 255 -388 261 388
rect 215 -400 261 -388
rect -205 -438 -33 -432
rect -205 -472 -193 -438
rect -45 -472 -33 -438
rect -205 -478 -33 -472
rect 33 -438 205 -432
rect 33 -472 45 -438
rect 193 -472 205 -438
rect 33 -478 205 -472
<< properties >>
string FIXED_BBOX -372 -593 372 593
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 4.0 l 0.9 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
