magic
tech sky130A
magscale 1 2
timestamp 1711996804
<< nwell >>
rect -3254 -3455 3254 3455
<< pmoslvt >>
rect -3058 1236 -1058 3236
rect -1000 1236 1000 3236
rect 1058 1236 3058 3236
rect -3058 -1000 -1058 1000
rect -1000 -1000 1000 1000
rect 1058 -1000 3058 1000
rect -3058 -3236 -1058 -1236
rect -1000 -3236 1000 -1236
rect 1058 -3236 3058 -1236
<< pdiff >>
rect -3116 3224 -3058 3236
rect -3116 1248 -3104 3224
rect -3070 1248 -3058 3224
rect -3116 1236 -3058 1248
rect -1058 3224 -1000 3236
rect -1058 1248 -1046 3224
rect -1012 1248 -1000 3224
rect -1058 1236 -1000 1248
rect 1000 3224 1058 3236
rect 1000 1248 1012 3224
rect 1046 1248 1058 3224
rect 1000 1236 1058 1248
rect 3058 3224 3116 3236
rect 3058 1248 3070 3224
rect 3104 1248 3116 3224
rect 3058 1236 3116 1248
rect -3116 988 -3058 1000
rect -3116 -988 -3104 988
rect -3070 -988 -3058 988
rect -3116 -1000 -3058 -988
rect -1058 988 -1000 1000
rect -1058 -988 -1046 988
rect -1012 -988 -1000 988
rect -1058 -1000 -1000 -988
rect 1000 988 1058 1000
rect 1000 -988 1012 988
rect 1046 -988 1058 988
rect 1000 -1000 1058 -988
rect 3058 988 3116 1000
rect 3058 -988 3070 988
rect 3104 -988 3116 988
rect 3058 -1000 3116 -988
rect -3116 -1248 -3058 -1236
rect -3116 -3224 -3104 -1248
rect -3070 -3224 -3058 -1248
rect -3116 -3236 -3058 -3224
rect -1058 -1248 -1000 -1236
rect -1058 -3224 -1046 -1248
rect -1012 -3224 -1000 -1248
rect -1058 -3236 -1000 -3224
rect 1000 -1248 1058 -1236
rect 1000 -3224 1012 -1248
rect 1046 -3224 1058 -1248
rect 1000 -3236 1058 -3224
rect 3058 -1248 3116 -1236
rect 3058 -3224 3070 -1248
rect 3104 -3224 3116 -1248
rect 3058 -3236 3116 -3224
<< pdiffc >>
rect -3104 1248 -3070 3224
rect -1046 1248 -1012 3224
rect 1012 1248 1046 3224
rect 3070 1248 3104 3224
rect -3104 -988 -3070 988
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect 3070 -988 3104 988
rect -3104 -3224 -3070 -1248
rect -1046 -3224 -1012 -1248
rect 1012 -3224 1046 -1248
rect 3070 -3224 3104 -1248
<< nsubdiff >>
rect -3218 3385 -3122 3419
rect 3122 3385 3218 3419
rect -3218 3323 -3184 3385
rect 3184 3323 3218 3385
rect -3218 -3385 -3184 -3323
rect 3184 -3385 3218 -3323
rect -3218 -3419 -3122 -3385
rect 3122 -3419 3218 -3385
<< nsubdiffcont >>
rect -3122 3385 3122 3419
rect -3218 -3323 -3184 3323
rect 3184 -3323 3218 3323
rect -3122 -3419 3122 -3385
<< poly >>
rect -3058 3317 -1058 3333
rect -3058 3283 -3042 3317
rect -1074 3283 -1058 3317
rect -3058 3236 -1058 3283
rect -1000 3317 1000 3333
rect -1000 3283 -984 3317
rect 984 3283 1000 3317
rect -1000 3236 1000 3283
rect 1058 3317 3058 3333
rect 1058 3283 1074 3317
rect 3042 3283 3058 3317
rect 1058 3236 3058 3283
rect -3058 1189 -1058 1236
rect -3058 1155 -3042 1189
rect -1074 1155 -1058 1189
rect -3058 1139 -1058 1155
rect -1000 1189 1000 1236
rect -1000 1155 -984 1189
rect 984 1155 1000 1189
rect -1000 1139 1000 1155
rect 1058 1189 3058 1236
rect 1058 1155 1074 1189
rect 3042 1155 3058 1189
rect 1058 1139 3058 1155
rect -3058 1081 -1058 1097
rect -3058 1047 -3042 1081
rect -1074 1047 -1058 1081
rect -3058 1000 -1058 1047
rect -1000 1081 1000 1097
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1000 1000 1000 1047
rect 1058 1081 3058 1097
rect 1058 1047 1074 1081
rect 3042 1047 3058 1081
rect 1058 1000 3058 1047
rect -3058 -1047 -1058 -1000
rect -3058 -1081 -3042 -1047
rect -1074 -1081 -1058 -1047
rect -3058 -1097 -1058 -1081
rect -1000 -1047 1000 -1000
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1000 -1097 1000 -1081
rect 1058 -1047 3058 -1000
rect 1058 -1081 1074 -1047
rect 3042 -1081 3058 -1047
rect 1058 -1097 3058 -1081
rect -3058 -1155 -1058 -1139
rect -3058 -1189 -3042 -1155
rect -1074 -1189 -1058 -1155
rect -3058 -1236 -1058 -1189
rect -1000 -1155 1000 -1139
rect -1000 -1189 -984 -1155
rect 984 -1189 1000 -1155
rect -1000 -1236 1000 -1189
rect 1058 -1155 3058 -1139
rect 1058 -1189 1074 -1155
rect 3042 -1189 3058 -1155
rect 1058 -1236 3058 -1189
rect -3058 -3283 -1058 -3236
rect -3058 -3317 -3042 -3283
rect -1074 -3317 -1058 -3283
rect -3058 -3333 -1058 -3317
rect -1000 -3283 1000 -3236
rect -1000 -3317 -984 -3283
rect 984 -3317 1000 -3283
rect -1000 -3333 1000 -3317
rect 1058 -3283 3058 -3236
rect 1058 -3317 1074 -3283
rect 3042 -3317 3058 -3283
rect 1058 -3333 3058 -3317
<< polycont >>
rect -3042 3283 -1074 3317
rect -984 3283 984 3317
rect 1074 3283 3042 3317
rect -3042 1155 -1074 1189
rect -984 1155 984 1189
rect 1074 1155 3042 1189
rect -3042 1047 -1074 1081
rect -984 1047 984 1081
rect 1074 1047 3042 1081
rect -3042 -1081 -1074 -1047
rect -984 -1081 984 -1047
rect 1074 -1081 3042 -1047
rect -3042 -1189 -1074 -1155
rect -984 -1189 984 -1155
rect 1074 -1189 3042 -1155
rect -3042 -3317 -1074 -3283
rect -984 -3317 984 -3283
rect 1074 -3317 3042 -3283
<< locali >>
rect -3218 3385 -3122 3419
rect 3122 3385 3218 3419
rect -3218 3323 -3184 3385
rect 3184 3323 3218 3385
rect -3058 3283 -3042 3317
rect -1074 3283 -1058 3317
rect -1000 3283 -984 3317
rect 984 3283 1000 3317
rect 1058 3283 1074 3317
rect 3042 3283 3058 3317
rect -3104 3224 -3070 3240
rect -3104 1232 -3070 1248
rect -1046 3224 -1012 3240
rect -1046 1232 -1012 1248
rect 1012 3224 1046 3240
rect 1012 1232 1046 1248
rect 3070 3224 3104 3240
rect 3070 1232 3104 1248
rect -3058 1155 -3042 1189
rect -1074 1155 -1058 1189
rect -1000 1155 -984 1189
rect 984 1155 1000 1189
rect 1058 1155 1074 1189
rect 3042 1155 3058 1189
rect -3058 1047 -3042 1081
rect -1074 1047 -1058 1081
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect 1058 1047 1074 1081
rect 3042 1047 3058 1081
rect -3104 988 -3070 1004
rect -3104 -1004 -3070 -988
rect -1046 988 -1012 1004
rect -1046 -1004 -1012 -988
rect 1012 988 1046 1004
rect 1012 -1004 1046 -988
rect 3070 988 3104 1004
rect 3070 -1004 3104 -988
rect -3058 -1081 -3042 -1047
rect -1074 -1081 -1058 -1047
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect 1058 -1081 1074 -1047
rect 3042 -1081 3058 -1047
rect -3058 -1189 -3042 -1155
rect -1074 -1189 -1058 -1155
rect -1000 -1189 -984 -1155
rect 984 -1189 1000 -1155
rect 1058 -1189 1074 -1155
rect 3042 -1189 3058 -1155
rect -3104 -1248 -3070 -1232
rect -3104 -3240 -3070 -3224
rect -1046 -1248 -1012 -1232
rect -1046 -3240 -1012 -3224
rect 1012 -1248 1046 -1232
rect 1012 -3240 1046 -3224
rect 3070 -1248 3104 -1232
rect 3070 -3240 3104 -3224
rect -3058 -3317 -3042 -3283
rect -1074 -3317 -1058 -3283
rect -1000 -3317 -984 -3283
rect 984 -3317 1000 -3283
rect 1058 -3317 1074 -3283
rect 3042 -3317 3058 -3283
rect -3218 -3385 -3184 -3323
rect 3184 -3385 3218 -3323
rect -3218 -3419 -3122 -3385
rect 3122 -3419 3218 -3385
<< viali >>
rect -3042 3283 -1074 3317
rect -984 3283 984 3317
rect 1074 3283 3042 3317
rect -3104 1248 -3070 3224
rect -1046 1248 -1012 3224
rect 1012 1248 1046 3224
rect 3070 1248 3104 3224
rect -3042 1155 -1074 1189
rect -984 1155 984 1189
rect 1074 1155 3042 1189
rect -3042 1047 -1074 1081
rect -984 1047 984 1081
rect 1074 1047 3042 1081
rect -3104 -988 -3070 988
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect 3070 -988 3104 988
rect -3042 -1081 -1074 -1047
rect -984 -1081 984 -1047
rect 1074 -1081 3042 -1047
rect -3042 -1189 -1074 -1155
rect -984 -1189 984 -1155
rect 1074 -1189 3042 -1155
rect -3104 -3224 -3070 -1248
rect -1046 -3224 -1012 -1248
rect 1012 -3224 1046 -1248
rect 3070 -3224 3104 -1248
rect -3042 -3317 -1074 -3283
rect -984 -3317 984 -3283
rect 1074 -3317 3042 -3283
<< metal1 >>
rect -3054 3317 -1062 3323
rect -3054 3283 -3042 3317
rect -1074 3283 -1062 3317
rect -3054 3277 -1062 3283
rect -996 3317 996 3323
rect -996 3283 -984 3317
rect 984 3283 996 3317
rect -996 3277 996 3283
rect 1062 3317 3054 3323
rect 1062 3283 1074 3317
rect 3042 3283 3054 3317
rect 1062 3277 3054 3283
rect -3110 3224 -3064 3236
rect -3110 1248 -3104 3224
rect -3070 1248 -3064 3224
rect -3110 1236 -3064 1248
rect -1052 3224 -1006 3236
rect -1052 1248 -1046 3224
rect -1012 1248 -1006 3224
rect -1052 1236 -1006 1248
rect 1006 3224 1052 3236
rect 1006 1248 1012 3224
rect 1046 1248 1052 3224
rect 1006 1236 1052 1248
rect 3064 3224 3110 3236
rect 3064 1248 3070 3224
rect 3104 1248 3110 3224
rect 3064 1236 3110 1248
rect -3054 1189 -1062 1195
rect -3054 1155 -3042 1189
rect -1074 1155 -1062 1189
rect -3054 1149 -1062 1155
rect -996 1189 996 1195
rect -996 1155 -984 1189
rect 984 1155 996 1189
rect -996 1149 996 1155
rect 1062 1189 3054 1195
rect 1062 1155 1074 1189
rect 3042 1155 3054 1189
rect 1062 1149 3054 1155
rect -3054 1081 -1062 1087
rect -3054 1047 -3042 1081
rect -1074 1047 -1062 1081
rect -3054 1041 -1062 1047
rect -996 1081 996 1087
rect -996 1047 -984 1081
rect 984 1047 996 1081
rect -996 1041 996 1047
rect 1062 1081 3054 1087
rect 1062 1047 1074 1081
rect 3042 1047 3054 1081
rect 1062 1041 3054 1047
rect -3110 988 -3064 1000
rect -3110 -988 -3104 988
rect -3070 -988 -3064 988
rect -3110 -1000 -3064 -988
rect -1052 988 -1006 1000
rect -1052 -988 -1046 988
rect -1012 -988 -1006 988
rect -1052 -1000 -1006 -988
rect 1006 988 1052 1000
rect 1006 -988 1012 988
rect 1046 -988 1052 988
rect 1006 -1000 1052 -988
rect 3064 988 3110 1000
rect 3064 -988 3070 988
rect 3104 -988 3110 988
rect 3064 -1000 3110 -988
rect -3054 -1047 -1062 -1041
rect -3054 -1081 -3042 -1047
rect -1074 -1081 -1062 -1047
rect -3054 -1087 -1062 -1081
rect -996 -1047 996 -1041
rect -996 -1081 -984 -1047
rect 984 -1081 996 -1047
rect -996 -1087 996 -1081
rect 1062 -1047 3054 -1041
rect 1062 -1081 1074 -1047
rect 3042 -1081 3054 -1047
rect 1062 -1087 3054 -1081
rect -3054 -1155 -1062 -1149
rect -3054 -1189 -3042 -1155
rect -1074 -1189 -1062 -1155
rect -3054 -1195 -1062 -1189
rect -996 -1155 996 -1149
rect -996 -1189 -984 -1155
rect 984 -1189 996 -1155
rect -996 -1195 996 -1189
rect 1062 -1155 3054 -1149
rect 1062 -1189 1074 -1155
rect 3042 -1189 3054 -1155
rect 1062 -1195 3054 -1189
rect -3110 -1248 -3064 -1236
rect -3110 -3224 -3104 -1248
rect -3070 -3224 -3064 -1248
rect -3110 -3236 -3064 -3224
rect -1052 -1248 -1006 -1236
rect -1052 -3224 -1046 -1248
rect -1012 -3224 -1006 -1248
rect -1052 -3236 -1006 -3224
rect 1006 -1248 1052 -1236
rect 1006 -3224 1012 -1248
rect 1046 -3224 1052 -1248
rect 1006 -3236 1052 -3224
rect 3064 -1248 3110 -1236
rect 3064 -3224 3070 -1248
rect 3104 -3224 3110 -1248
rect 3064 -3236 3110 -3224
rect -3054 -3283 -1062 -3277
rect -3054 -3317 -3042 -3283
rect -1074 -3317 -1062 -3283
rect -3054 -3323 -1062 -3317
rect -996 -3283 996 -3277
rect -996 -3317 -984 -3283
rect 984 -3317 996 -3283
rect -996 -3323 996 -3317
rect 1062 -3283 3054 -3277
rect 1062 -3317 1074 -3283
rect 3042 -3317 3054 -3283
rect 1062 -3323 3054 -3317
<< properties >>
string FIXED_BBOX -3201 -3402 3201 3402
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 10.0 m 3 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
