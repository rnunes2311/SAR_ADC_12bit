magic
tech sky130A
magscale 1 2
timestamp 1711982102
<< nwell >>
rect 2362 9826 2784 9828
rect -3416 9260 2784 9826
rect -3416 7796 2362 9260
rect -3418 7788 2362 7796
rect -3418 7475 -3066 7788
rect -2092 7326 -1242 7788
rect 232 6752 2362 7788
rect 4856 6752 6186 7590
<< pwell >>
rect 2784 9224 7548 9828
rect -3338 7235 -3152 7417
rect -3338 7231 -3317 7235
rect -3351 7197 -3317 7231
rect -1064 6944 206 7764
rect 2362 7766 7548 9224
rect 2362 7306 2784 7766
rect 2362 6752 3486 7306
rect 3810 6752 4528 7552
rect 6218 6752 7548 7572
<< nmos >>
rect -864 7154 -834 7554
rect -654 7154 -624 7554
rect -444 7154 -414 7554
rect -234 7154 -204 7554
rect -24 7154 6 7554
rect 2558 8814 2588 9014
rect 2558 6962 2588 8562
rect 6418 6962 6448 7362
rect 6514 6962 6544 7362
rect 6610 6962 6640 7362
rect 6706 6962 6736 7362
rect 7030 6962 7060 7362
rect 7126 6962 7156 7362
rect 7222 6962 7252 7362
rect 7318 6962 7348 7362
<< scnmos >>
rect -3260 7261 -3230 7391
<< pmos >>
rect -3220 8007 -3120 9607
rect -2948 8007 -2848 9607
rect -2676 8007 -2576 9607
rect -2404 8007 -2304 9607
rect -2132 8007 -2032 9607
rect -1860 8007 -1760 9607
rect -1588 8007 -1488 9607
rect -1316 8007 -1216 9607
rect -1044 8007 -944 9607
rect -772 8007 -672 9607
rect -500 8007 -400 9607
rect -228 8007 -128 9607
rect 44 8007 144 9607
rect 428 8407 468 9607
rect 526 8407 566 9607
rect 624 8407 664 9607
rect 722 8407 762 9607
rect 820 8407 860 9607
rect 918 8407 958 9607
rect 1016 8407 1056 9607
rect 1114 8407 1154 9607
rect 428 6971 468 8171
rect 526 6971 566 8171
rect 624 6971 664 8171
rect 722 6971 762 8171
rect 820 6971 860 8171
rect 918 6971 958 8171
rect 1016 6971 1056 8171
rect 1114 6971 1154 8171
rect 1440 8407 1480 9607
rect 1538 8407 1578 9607
rect 1636 8407 1676 9607
rect 1734 8407 1774 9607
rect 1832 8407 1872 9607
rect 1930 8407 1970 9607
rect 2028 8407 2068 9607
rect 2126 8407 2166 9607
rect 1440 6971 1480 8171
rect 1538 6971 1578 8171
rect 1636 6971 1676 8171
rect 1734 6971 1774 8171
rect 1832 6971 1872 8171
rect 1930 6971 1970 8171
rect 2028 6971 2068 8171
rect 2126 6971 2166 8171
rect 2558 9480 2588 9680
<< scpmoshvt >>
rect -3260 7511 -3230 7711
<< nnmos >>
rect 3000 7010 3100 7110
rect 3158 7010 3258 7110
<< pmoslvt >>
rect -1896 7546 -1696 7746
rect -1638 7546 -1438 7746
<< pmoshvt >>
rect 5056 6971 5086 7371
rect 5152 6971 5182 7371
rect 5248 6971 5278 7371
rect 5344 6971 5374 7371
rect 5668 6971 5698 7371
rect 5764 6971 5794 7371
rect 5860 6971 5890 7371
rect 5956 6971 5986 7371
<< nmoslvt >>
rect 4010 6962 4040 7342
rect 4106 6962 4136 7342
rect 4202 6962 4232 7342
rect 4298 6962 4328 7342
<< ndiff >>
rect -3312 7379 -3260 7391
rect -3312 7345 -3304 7379
rect -3270 7345 -3260 7379
rect -3312 7311 -3260 7345
rect -3312 7277 -3304 7311
rect -3270 7277 -3260 7311
rect -3312 7261 -3260 7277
rect -3230 7379 -3178 7391
rect -3230 7345 -3220 7379
rect -3186 7345 -3178 7379
rect -3230 7311 -3178 7345
rect -3230 7277 -3220 7311
rect -3186 7277 -3178 7311
rect -3230 7261 -3178 7277
rect -926 7542 -864 7554
rect -926 7166 -914 7542
rect -880 7166 -864 7542
rect -926 7154 -864 7166
rect -834 7542 -772 7554
rect -834 7166 -818 7542
rect -784 7166 -772 7542
rect -834 7154 -772 7166
rect -716 7542 -654 7554
rect -716 7166 -704 7542
rect -670 7166 -654 7542
rect -716 7154 -654 7166
rect -624 7542 -562 7554
rect -624 7166 -608 7542
rect -574 7166 -562 7542
rect -624 7154 -562 7166
rect -506 7542 -444 7554
rect -506 7166 -494 7542
rect -460 7166 -444 7542
rect -506 7154 -444 7166
rect -414 7542 -352 7554
rect -414 7166 -398 7542
rect -364 7166 -352 7542
rect -414 7154 -352 7166
rect -296 7542 -234 7554
rect -296 7166 -284 7542
rect -250 7166 -234 7542
rect -296 7154 -234 7166
rect -204 7542 -142 7554
rect -204 7166 -188 7542
rect -154 7166 -142 7542
rect -204 7154 -142 7166
rect -86 7542 -24 7554
rect -86 7166 -74 7542
rect -40 7166 -24 7542
rect -86 7154 -24 7166
rect 6 7542 68 7554
rect 6 7166 22 7542
rect 56 7166 68 7542
rect 6 7154 68 7166
rect 2500 9002 2558 9014
rect 2500 8826 2512 9002
rect 2546 8826 2558 9002
rect 2500 8814 2558 8826
rect 2588 9002 2646 9014
rect 2588 8826 2600 9002
rect 2634 8826 2646 9002
rect 2588 8814 2646 8826
rect 2500 8550 2558 8562
rect 2500 6974 2512 8550
rect 2546 6974 2558 8550
rect 2500 6962 2558 6974
rect 2588 8550 2646 8562
rect 2588 6974 2600 8550
rect 2634 6974 2646 8550
rect 2588 6962 2646 6974
rect 3948 7330 4010 7342
rect 3948 6974 3960 7330
rect 3994 6974 4010 7330
rect 3948 6962 4010 6974
rect 4040 7330 4106 7342
rect 4040 6974 4056 7330
rect 4090 6974 4106 7330
rect 4040 6962 4106 6974
rect 4136 7330 4202 7342
rect 4136 6974 4152 7330
rect 4186 6974 4202 7330
rect 4136 6962 4202 6974
rect 4232 7330 4298 7342
rect 4232 6974 4248 7330
rect 4282 6974 4298 7330
rect 4232 6962 4298 6974
rect 4328 7330 4390 7342
rect 4328 6974 4344 7330
rect 4378 6974 4390 7330
rect 4328 6962 4390 6974
rect 6356 7350 6418 7362
rect 6356 6974 6368 7350
rect 6402 6974 6418 7350
rect 6356 6962 6418 6974
rect 6448 7350 6514 7362
rect 6448 6974 6464 7350
rect 6498 6974 6514 7350
rect 6448 6962 6514 6974
rect 6544 7350 6610 7362
rect 6544 6974 6560 7350
rect 6594 6974 6610 7350
rect 6544 6962 6610 6974
rect 6640 7350 6706 7362
rect 6640 6974 6656 7350
rect 6690 6974 6706 7350
rect 6640 6962 6706 6974
rect 6736 7350 6798 7362
rect 6736 6974 6752 7350
rect 6786 6974 6798 7350
rect 6736 6962 6798 6974
rect 6968 7350 7030 7362
rect 6968 6974 6980 7350
rect 7014 6974 7030 7350
rect 6968 6962 7030 6974
rect 7060 7350 7126 7362
rect 7060 6974 7076 7350
rect 7110 6974 7126 7350
rect 7060 6962 7126 6974
rect 7156 7350 7222 7362
rect 7156 6974 7172 7350
rect 7206 6974 7222 7350
rect 7156 6962 7222 6974
rect 7252 7350 7318 7362
rect 7252 6974 7268 7350
rect 7302 6974 7318 7350
rect 7252 6962 7318 6974
rect 7348 7350 7410 7362
rect 7348 6974 7364 7350
rect 7398 6974 7410 7350
rect 7348 6962 7410 6974
<< pdiff >>
rect -3278 9595 -3220 9607
rect -3278 8019 -3266 9595
rect -3232 8019 -3220 9595
rect -3278 8007 -3220 8019
rect -3120 9595 -3062 9607
rect -3120 8019 -3108 9595
rect -3074 8019 -3062 9595
rect -3120 8007 -3062 8019
rect -3006 9595 -2948 9607
rect -3006 8019 -2994 9595
rect -2960 8019 -2948 9595
rect -3006 8007 -2948 8019
rect -2848 9595 -2790 9607
rect -2848 8019 -2836 9595
rect -2802 8019 -2790 9595
rect -2848 8007 -2790 8019
rect -2734 9595 -2676 9607
rect -2734 8019 -2722 9595
rect -2688 8019 -2676 9595
rect -2734 8007 -2676 8019
rect -2576 9595 -2518 9607
rect -2576 8019 -2564 9595
rect -2530 8019 -2518 9595
rect -2576 8007 -2518 8019
rect -2462 9595 -2404 9607
rect -2462 8019 -2450 9595
rect -2416 8019 -2404 9595
rect -2462 8007 -2404 8019
rect -2304 9595 -2246 9607
rect -2304 8019 -2292 9595
rect -2258 8019 -2246 9595
rect -2304 8007 -2246 8019
rect -2190 9595 -2132 9607
rect -2190 8019 -2178 9595
rect -2144 8019 -2132 9595
rect -2190 8007 -2132 8019
rect -2032 9595 -1974 9607
rect -2032 8019 -2020 9595
rect -1986 8019 -1974 9595
rect -2032 8007 -1974 8019
rect -1918 9595 -1860 9607
rect -1918 8019 -1906 9595
rect -1872 8019 -1860 9595
rect -1918 8007 -1860 8019
rect -1760 9595 -1702 9607
rect -1760 8019 -1748 9595
rect -1714 8019 -1702 9595
rect -1760 8007 -1702 8019
rect -1646 9595 -1588 9607
rect -1646 8019 -1634 9595
rect -1600 8019 -1588 9595
rect -1646 8007 -1588 8019
rect -1488 9595 -1430 9607
rect -1488 8019 -1476 9595
rect -1442 8019 -1430 9595
rect -1488 8007 -1430 8019
rect -1374 9595 -1316 9607
rect -1374 8019 -1362 9595
rect -1328 8019 -1316 9595
rect -1374 8007 -1316 8019
rect -1216 9595 -1158 9607
rect -1216 8019 -1204 9595
rect -1170 8019 -1158 9595
rect -1216 8007 -1158 8019
rect -1102 9595 -1044 9607
rect -1102 8019 -1090 9595
rect -1056 8019 -1044 9595
rect -1102 8007 -1044 8019
rect -944 9595 -886 9607
rect -944 8019 -932 9595
rect -898 8019 -886 9595
rect -944 8007 -886 8019
rect -830 9595 -772 9607
rect -830 8019 -818 9595
rect -784 8019 -772 9595
rect -830 8007 -772 8019
rect -672 9595 -614 9607
rect -672 8019 -660 9595
rect -626 8019 -614 9595
rect -672 8007 -614 8019
rect -558 9595 -500 9607
rect -558 8019 -546 9595
rect -512 8019 -500 9595
rect -558 8007 -500 8019
rect -400 9595 -342 9607
rect -400 8019 -388 9595
rect -354 8019 -342 9595
rect -400 8007 -342 8019
rect -286 9595 -228 9607
rect -286 8019 -274 9595
rect -240 8019 -228 9595
rect -286 8007 -228 8019
rect -128 9595 -70 9607
rect -128 8019 -116 9595
rect -82 8019 -70 9595
rect -128 8007 -70 8019
rect -14 9595 44 9607
rect -14 8019 -2 9595
rect 32 8019 44 9595
rect -14 8007 44 8019
rect 144 9595 202 9607
rect 144 8019 156 9595
rect 190 8019 202 9595
rect 144 8007 202 8019
rect 370 9595 428 9607
rect 370 8419 382 9595
rect 416 8419 428 9595
rect 370 8407 428 8419
rect 468 9595 526 9607
rect 468 8419 480 9595
rect 514 8419 526 9595
rect 468 8407 526 8419
rect 566 9595 624 9607
rect 566 8419 578 9595
rect 612 8419 624 9595
rect 566 8407 624 8419
rect 664 9595 722 9607
rect 664 8419 676 9595
rect 710 8419 722 9595
rect 664 8407 722 8419
rect 762 9595 820 9607
rect 762 8419 774 9595
rect 808 8419 820 9595
rect 762 8407 820 8419
rect 860 9595 918 9607
rect 860 8419 872 9595
rect 906 8419 918 9595
rect 860 8407 918 8419
rect 958 9595 1016 9607
rect 958 8419 970 9595
rect 1004 8419 1016 9595
rect 958 8407 1016 8419
rect 1056 9595 1114 9607
rect 1056 8419 1068 9595
rect 1102 8419 1114 9595
rect 1056 8407 1114 8419
rect 1154 9595 1212 9607
rect 1154 8419 1166 9595
rect 1200 8419 1212 9595
rect 1154 8407 1212 8419
rect 370 8159 428 8171
rect -3312 7699 -3260 7711
rect -3312 7665 -3304 7699
rect -3270 7665 -3260 7699
rect -3312 7631 -3260 7665
rect -3312 7597 -3304 7631
rect -3270 7597 -3260 7631
rect -3312 7563 -3260 7597
rect -3312 7529 -3304 7563
rect -3270 7529 -3260 7563
rect -3312 7511 -3260 7529
rect -3230 7699 -3178 7711
rect -3230 7665 -3220 7699
rect -3186 7665 -3178 7699
rect -3230 7631 -3178 7665
rect -3230 7597 -3220 7631
rect -3186 7597 -3178 7631
rect -3230 7563 -3178 7597
rect -3230 7529 -3220 7563
rect -3186 7529 -3178 7563
rect -3230 7511 -3178 7529
rect -1954 7734 -1896 7746
rect -1954 7558 -1942 7734
rect -1908 7558 -1896 7734
rect -1954 7546 -1896 7558
rect -1696 7734 -1638 7746
rect -1696 7558 -1684 7734
rect -1650 7558 -1638 7734
rect -1696 7546 -1638 7558
rect -1438 7734 -1380 7746
rect -1438 7558 -1426 7734
rect -1392 7558 -1380 7734
rect -1438 7546 -1380 7558
rect 370 6983 382 8159
rect 416 6983 428 8159
rect 370 6971 428 6983
rect 468 8159 526 8171
rect 468 6983 480 8159
rect 514 6983 526 8159
rect 468 6971 526 6983
rect 566 8159 624 8171
rect 566 6983 578 8159
rect 612 6983 624 8159
rect 566 6971 624 6983
rect 664 8159 722 8171
rect 664 6983 676 8159
rect 710 6983 722 8159
rect 664 6971 722 6983
rect 762 8159 820 8171
rect 762 6983 774 8159
rect 808 6983 820 8159
rect 762 6971 820 6983
rect 860 8159 918 8171
rect 860 6983 872 8159
rect 906 6983 918 8159
rect 860 6971 918 6983
rect 958 8159 1016 8171
rect 958 6983 970 8159
rect 1004 6983 1016 8159
rect 958 6971 1016 6983
rect 1056 8159 1114 8171
rect 1056 6983 1068 8159
rect 1102 6983 1114 8159
rect 1056 6971 1114 6983
rect 1154 8159 1212 8171
rect 1154 6983 1166 8159
rect 1200 6983 1212 8159
rect 1154 6971 1212 6983
rect 1382 9595 1440 9607
rect 1382 8419 1394 9595
rect 1428 8419 1440 9595
rect 1382 8407 1440 8419
rect 1480 9595 1538 9607
rect 1480 8419 1492 9595
rect 1526 8419 1538 9595
rect 1480 8407 1538 8419
rect 1578 9595 1636 9607
rect 1578 8419 1590 9595
rect 1624 8419 1636 9595
rect 1578 8407 1636 8419
rect 1676 9595 1734 9607
rect 1676 8419 1688 9595
rect 1722 8419 1734 9595
rect 1676 8407 1734 8419
rect 1774 9595 1832 9607
rect 1774 8419 1786 9595
rect 1820 8419 1832 9595
rect 1774 8407 1832 8419
rect 1872 9595 1930 9607
rect 1872 8419 1884 9595
rect 1918 8419 1930 9595
rect 1872 8407 1930 8419
rect 1970 9595 2028 9607
rect 1970 8419 1982 9595
rect 2016 8419 2028 9595
rect 1970 8407 2028 8419
rect 2068 9595 2126 9607
rect 2068 8419 2080 9595
rect 2114 8419 2126 9595
rect 2068 8407 2126 8419
rect 2166 9595 2224 9607
rect 2166 8419 2178 9595
rect 2212 8419 2224 9595
rect 2166 8407 2224 8419
rect 1382 8159 1440 8171
rect 1382 6983 1394 8159
rect 1428 6983 1440 8159
rect 1382 6971 1440 6983
rect 1480 8159 1538 8171
rect 1480 6983 1492 8159
rect 1526 6983 1538 8159
rect 1480 6971 1538 6983
rect 1578 8159 1636 8171
rect 1578 6983 1590 8159
rect 1624 6983 1636 8159
rect 1578 6971 1636 6983
rect 1676 8159 1734 8171
rect 1676 6983 1688 8159
rect 1722 6983 1734 8159
rect 1676 6971 1734 6983
rect 1774 8159 1832 8171
rect 1774 6983 1786 8159
rect 1820 6983 1832 8159
rect 1774 6971 1832 6983
rect 1872 8159 1930 8171
rect 1872 6983 1884 8159
rect 1918 6983 1930 8159
rect 1872 6971 1930 6983
rect 1970 8159 2028 8171
rect 1970 6983 1982 8159
rect 2016 6983 2028 8159
rect 1970 6971 2028 6983
rect 2068 8159 2126 8171
rect 2068 6983 2080 8159
rect 2114 6983 2126 8159
rect 2068 6971 2126 6983
rect 2166 8159 2224 8171
rect 2166 6983 2178 8159
rect 2212 6983 2224 8159
rect 2166 6971 2224 6983
rect 2500 9668 2558 9680
rect 2500 9492 2512 9668
rect 2546 9492 2558 9668
rect 2500 9480 2558 9492
rect 2588 9668 2646 9680
rect 2588 9492 2600 9668
rect 2634 9492 2646 9668
rect 2588 9480 2646 9492
rect 4994 7359 5056 7371
rect 4994 6983 5006 7359
rect 5040 6983 5056 7359
rect 4994 6971 5056 6983
rect 5086 7359 5152 7371
rect 5086 6983 5102 7359
rect 5136 6983 5152 7359
rect 5086 6971 5152 6983
rect 5182 7359 5248 7371
rect 5182 6983 5198 7359
rect 5232 6983 5248 7359
rect 5182 6971 5248 6983
rect 5278 7359 5344 7371
rect 5278 6983 5294 7359
rect 5328 6983 5344 7359
rect 5278 6971 5344 6983
rect 5374 7359 5436 7371
rect 5374 6983 5390 7359
rect 5424 6983 5436 7359
rect 5374 6971 5436 6983
rect 5606 7359 5668 7371
rect 5606 6983 5618 7359
rect 5652 6983 5668 7359
rect 5606 6971 5668 6983
rect 5698 7359 5764 7371
rect 5698 6983 5714 7359
rect 5748 6983 5764 7359
rect 5698 6971 5764 6983
rect 5794 7359 5860 7371
rect 5794 6983 5810 7359
rect 5844 6983 5860 7359
rect 5794 6971 5860 6983
rect 5890 7359 5956 7371
rect 5890 6983 5906 7359
rect 5940 6983 5956 7359
rect 5890 6971 5956 6983
rect 5986 7359 6048 7371
rect 5986 6983 6002 7359
rect 6036 6983 6048 7359
rect 5986 6971 6048 6983
<< mvndiff >>
rect 2942 7098 3000 7110
rect 2942 7022 2954 7098
rect 2988 7022 3000 7098
rect 2942 7010 3000 7022
rect 3100 7098 3158 7110
rect 3100 7022 3112 7098
rect 3146 7022 3158 7098
rect 3100 7010 3158 7022
rect 3258 7098 3316 7110
rect 3258 7022 3270 7098
rect 3304 7022 3316 7098
rect 3258 7010 3316 7022
<< ndiffc >>
rect -3304 7345 -3270 7379
rect -3304 7277 -3270 7311
rect -3220 7345 -3186 7379
rect -3220 7277 -3186 7311
rect -914 7166 -880 7542
rect -818 7166 -784 7542
rect -704 7166 -670 7542
rect -608 7166 -574 7542
rect -494 7166 -460 7542
rect -398 7166 -364 7542
rect -284 7166 -250 7542
rect -188 7166 -154 7542
rect -74 7166 -40 7542
rect 22 7166 56 7542
rect 2512 8826 2546 9002
rect 2600 8826 2634 9002
rect 2512 6974 2546 8550
rect 2600 6974 2634 8550
rect 3960 6974 3994 7330
rect 4056 6974 4090 7330
rect 4152 6974 4186 7330
rect 4248 6974 4282 7330
rect 4344 6974 4378 7330
rect 6368 6974 6402 7350
rect 6464 6974 6498 7350
rect 6560 6974 6594 7350
rect 6656 6974 6690 7350
rect 6752 6974 6786 7350
rect 6980 6974 7014 7350
rect 7076 6974 7110 7350
rect 7172 6974 7206 7350
rect 7268 6974 7302 7350
rect 7364 6974 7398 7350
<< pdiffc >>
rect -3266 8019 -3232 9595
rect -3108 8019 -3074 9595
rect -2994 8019 -2960 9595
rect -2836 8019 -2802 9595
rect -2722 8019 -2688 9595
rect -2564 8019 -2530 9595
rect -2450 8019 -2416 9595
rect -2292 8019 -2258 9595
rect -2178 8019 -2144 9595
rect -2020 8019 -1986 9595
rect -1906 8019 -1872 9595
rect -1748 8019 -1714 9595
rect -1634 8019 -1600 9595
rect -1476 8019 -1442 9595
rect -1362 8019 -1328 9595
rect -1204 8019 -1170 9595
rect -1090 8019 -1056 9595
rect -932 8019 -898 9595
rect -818 8019 -784 9595
rect -660 8019 -626 9595
rect -546 8019 -512 9595
rect -388 8019 -354 9595
rect -274 8019 -240 9595
rect -116 8019 -82 9595
rect -2 8019 32 9595
rect 156 8019 190 9595
rect 382 8419 416 9595
rect 480 8419 514 9595
rect 578 8419 612 9595
rect 676 8419 710 9595
rect 774 8419 808 9595
rect 872 8419 906 9595
rect 970 8419 1004 9595
rect 1068 8419 1102 9595
rect 1166 8419 1200 9595
rect -3304 7665 -3270 7699
rect -3304 7597 -3270 7631
rect -3304 7529 -3270 7563
rect -3220 7665 -3186 7699
rect -3220 7597 -3186 7631
rect -3220 7529 -3186 7563
rect -1942 7558 -1908 7734
rect -1684 7558 -1650 7734
rect -1426 7558 -1392 7734
rect 382 6983 416 8159
rect 480 6983 514 8159
rect 578 6983 612 8159
rect 676 6983 710 8159
rect 774 6983 808 8159
rect 872 6983 906 8159
rect 970 6983 1004 8159
rect 1068 6983 1102 8159
rect 1166 6983 1200 8159
rect 1394 8419 1428 9595
rect 1492 8419 1526 9595
rect 1590 8419 1624 9595
rect 1688 8419 1722 9595
rect 1786 8419 1820 9595
rect 1884 8419 1918 9595
rect 1982 8419 2016 9595
rect 2080 8419 2114 9595
rect 2178 8419 2212 9595
rect 1394 6983 1428 8159
rect 1492 6983 1526 8159
rect 1590 6983 1624 8159
rect 1688 6983 1722 8159
rect 1786 6983 1820 8159
rect 1884 6983 1918 8159
rect 1982 6983 2016 8159
rect 2080 6983 2114 8159
rect 2178 6983 2212 8159
rect 2512 9492 2546 9668
rect 2600 9492 2634 9668
rect 5006 6983 5040 7359
rect 5102 6983 5136 7359
rect 5198 6983 5232 7359
rect 5294 6983 5328 7359
rect 5390 6983 5424 7359
rect 5618 6983 5652 7359
rect 5714 6983 5748 7359
rect 5810 6983 5844 7359
rect 5906 6983 5940 7359
rect 6002 6983 6036 7359
<< mvndiffc >>
rect 2954 7022 2988 7098
rect 3112 7022 3146 7098
rect 3270 7022 3304 7098
<< psubdiff >>
rect -1028 7694 -932 7728
rect 74 7694 170 7728
rect -1028 7632 -994 7694
rect 136 7632 170 7694
rect -1028 7014 -994 7076
rect 136 7014 170 7076
rect -1028 6980 -932 7014
rect 74 6980 170 7014
rect 2820 9758 2916 9792
rect 7416 9758 7512 9792
rect 2820 9696 2854 9758
rect 2398 9154 2494 9188
rect 2652 9154 2748 9188
rect 2398 9092 2432 9154
rect 2714 9092 2748 9154
rect 2398 8736 2432 8798
rect 2714 8736 2748 8798
rect 2398 8702 2494 8736
rect 2652 8702 2748 8736
rect 2398 8640 2432 8702
rect 2714 8640 2748 8702
rect 2398 6822 2432 6884
rect 7478 9696 7512 9758
rect 2820 7836 2854 7898
rect 7478 7836 7512 7898
rect 2820 7802 2916 7836
rect 7416 7802 7512 7836
rect 3846 7482 3942 7516
rect 4396 7482 4492 7516
rect 3846 7420 3880 7482
rect 2714 6822 2748 6884
rect 2398 6788 2494 6822
rect 2652 6788 2748 6822
rect 4458 7420 4492 7482
rect 3846 6822 3880 6884
rect 4458 6822 4492 6884
rect 3846 6788 3942 6822
rect 4396 6788 4492 6822
rect 6254 7502 6350 7536
rect 6804 7502 6962 7536
rect 7416 7502 7512 7536
rect 6254 7440 6288 7502
rect 6866 7440 6900 7502
rect 6254 6822 6288 6884
rect 7478 7440 7512 7502
rect 6866 6822 6900 6884
rect 7478 6822 7512 6884
rect 6254 6788 6350 6822
rect 6804 6788 6962 6822
rect 7416 6788 7512 6822
<< nsubdiff >>
rect -3380 9756 -3284 9790
rect 208 9756 364 9790
rect 1218 9756 1376 9790
rect 2230 9756 2326 9790
rect -3380 9694 -3346 9756
rect 268 9694 304 9756
rect -3380 7858 -3346 7920
rect 268 7920 270 9694
rect 1280 9694 1314 9756
rect 268 7858 304 7920
rect -3380 7824 -3284 7858
rect 208 7824 304 7858
rect -2056 7761 -2022 7824
rect -1312 7761 -1278 7824
rect -2056 7396 -2022 7459
rect -1312 7396 -1278 7459
rect -2056 7362 -1960 7396
rect -1374 7362 -1278 7396
rect 268 6822 302 7824
rect 2292 9694 2326 9756
rect 1280 6822 1314 6884
rect 2398 9758 2494 9792
rect 2652 9758 2748 9792
rect 2398 9695 2432 9758
rect 2714 9695 2748 9758
rect 2398 9330 2432 9393
rect 2714 9330 2748 9393
rect 2398 9296 2494 9330
rect 2652 9296 2748 9330
rect 2292 6822 2326 6884
rect 268 6788 364 6822
rect 1218 6788 1376 6822
rect 2230 6788 2326 6822
rect 4892 7520 4988 7554
rect 5442 7520 5600 7554
rect 6054 7520 6150 7554
rect 4892 7458 4926 7520
rect 5504 7458 5538 7520
rect 4892 6822 4926 6884
rect 6116 7458 6150 7520
rect 5504 6822 5538 6884
rect 6116 6822 6150 6884
rect 4892 6788 4988 6822
rect 5442 6788 5600 6822
rect 6054 6788 6150 6822
<< mvpsubdiff >>
rect 2808 7258 3450 7270
rect 2808 7224 2916 7258
rect 3342 7224 3450 7258
rect 2808 7212 3450 7224
rect 2808 7162 2866 7212
rect 2808 6896 2820 7162
rect 2854 6896 2866 7162
rect 3392 7162 3450 7212
rect 2808 6846 2866 6896
rect 3392 6896 3404 7162
rect 3438 6896 3450 7162
rect 3392 6846 3450 6896
rect 2808 6834 3450 6846
rect 2808 6800 2916 6834
rect 3342 6800 3450 6834
rect 2808 6788 3450 6800
<< psubdiffcont >>
rect -932 7694 74 7728
rect -1028 7076 -994 7632
rect 136 7076 170 7632
rect -932 6980 74 7014
rect 2916 9758 7416 9792
rect 2494 9154 2652 9188
rect 2398 8798 2432 9092
rect 2714 8798 2748 9092
rect 2494 8702 2652 8736
rect 2398 6884 2432 8640
rect 2714 6884 2748 8640
rect 2820 7898 2854 9696
rect 7478 7898 7512 9696
rect 2916 7802 7416 7836
rect 3942 7482 4396 7516
rect 2494 6788 2652 6822
rect 3846 6884 3880 7420
rect 4458 6884 4492 7420
rect 3942 6788 4396 6822
rect 6350 7502 6804 7536
rect 6962 7502 7416 7536
rect 6254 6884 6288 7440
rect 6866 6884 6900 7440
rect 7478 6884 7512 7440
rect 6350 6788 6804 6822
rect 6962 6788 7416 6822
<< nsubdiffcont >>
rect -3284 9756 208 9790
rect 364 9756 1218 9790
rect 1376 9756 2230 9790
rect -3380 7920 -3346 9694
rect 270 7920 304 9694
rect -3284 7824 208 7858
rect -2056 7459 -2022 7761
rect -1312 7459 -1278 7761
rect -1960 7362 -1374 7396
rect 1280 6884 1314 9694
rect 2292 6884 2326 9694
rect 2494 9758 2652 9792
rect 2398 9393 2432 9695
rect 2714 9393 2748 9695
rect 2494 9296 2652 9330
rect 364 6788 1218 6822
rect 1376 6788 2230 6822
rect 4988 7520 5442 7554
rect 5600 7520 6054 7554
rect 4892 6884 4926 7458
rect 5504 6884 5538 7458
rect 6116 6884 6150 7458
rect 4988 6788 5442 6822
rect 5600 6788 6054 6822
<< mvpsubdiffcont >>
rect 2916 7224 3342 7258
rect 2820 6896 2854 7162
rect 3404 6896 3438 7162
rect 2916 6800 3342 6834
<< poly >>
rect -3220 9688 -3120 9704
rect -3220 9654 -3204 9688
rect -3136 9654 -3120 9688
rect -3220 9607 -3120 9654
rect -2948 9688 -2848 9704
rect -2948 9654 -2932 9688
rect -2864 9654 -2848 9688
rect -2948 9607 -2848 9654
rect -2676 9688 -2576 9704
rect -2676 9654 -2660 9688
rect -2592 9654 -2576 9688
rect -2676 9607 -2576 9654
rect -2404 9688 -2304 9704
rect -2404 9654 -2388 9688
rect -2320 9654 -2304 9688
rect -2404 9607 -2304 9654
rect -2132 9688 -2032 9704
rect -2132 9654 -2116 9688
rect -2048 9654 -2032 9688
rect -2132 9607 -2032 9654
rect -1860 9688 -1760 9704
rect -1860 9654 -1844 9688
rect -1776 9654 -1760 9688
rect -1860 9607 -1760 9654
rect -1588 9688 -1488 9704
rect -1588 9654 -1572 9688
rect -1504 9654 -1488 9688
rect -1588 9607 -1488 9654
rect -1316 9688 -1216 9704
rect -1316 9654 -1300 9688
rect -1232 9654 -1216 9688
rect -1316 9607 -1216 9654
rect -1044 9688 -944 9704
rect -1044 9654 -1028 9688
rect -960 9654 -944 9688
rect -1044 9607 -944 9654
rect -772 9688 -672 9704
rect -772 9654 -756 9688
rect -688 9654 -672 9688
rect -772 9607 -672 9654
rect -500 9688 -400 9704
rect -500 9654 -484 9688
rect -416 9654 -400 9688
rect -500 9607 -400 9654
rect -228 9688 -128 9704
rect -228 9654 -212 9688
rect -144 9654 -128 9688
rect -228 9607 -128 9654
rect 44 9688 144 9704
rect 44 9654 60 9688
rect 128 9654 144 9688
rect 44 9607 144 9654
rect -3220 7960 -3120 8007
rect -3220 7926 -3204 7960
rect -3136 7926 -3120 7960
rect -3220 7910 -3120 7926
rect -2948 7960 -2848 8007
rect -2948 7926 -2932 7960
rect -2864 7926 -2848 7960
rect -2948 7910 -2848 7926
rect -2676 7960 -2576 8007
rect -2676 7926 -2660 7960
rect -2592 7926 -2576 7960
rect -2676 7910 -2576 7926
rect -2404 7960 -2304 8007
rect -2404 7926 -2388 7960
rect -2320 7926 -2304 7960
rect -2404 7910 -2304 7926
rect -2132 7960 -2032 8007
rect -2132 7926 -2116 7960
rect -2048 7926 -2032 7960
rect -2132 7910 -2032 7926
rect -1860 7960 -1760 8007
rect -1860 7926 -1844 7960
rect -1776 7926 -1760 7960
rect -1860 7910 -1760 7926
rect -1588 7960 -1488 8007
rect -1588 7926 -1572 7960
rect -1504 7926 -1488 7960
rect -1588 7910 -1488 7926
rect -1316 7960 -1216 8007
rect -1316 7926 -1300 7960
rect -1232 7926 -1216 7960
rect -1316 7910 -1216 7926
rect -1044 7960 -944 8007
rect -1044 7926 -1028 7960
rect -960 7926 -944 7960
rect -1044 7910 -944 7926
rect -772 7960 -672 8007
rect -772 7926 -756 7960
rect -688 7926 -672 7960
rect -772 7910 -672 7926
rect -500 7960 -400 8007
rect -500 7926 -484 7960
rect -416 7926 -400 7960
rect -500 7910 -400 7926
rect -228 7960 -128 8007
rect -228 7926 -212 7960
rect -144 7926 -128 7960
rect -228 7910 -128 7926
rect 44 7960 144 8007
rect 44 7926 60 7960
rect 128 7926 144 7960
rect 44 7910 144 7926
rect 415 9688 481 9704
rect 415 9654 431 9688
rect 465 9654 481 9688
rect 415 9638 481 9654
rect 611 9688 677 9704
rect 611 9654 627 9688
rect 661 9654 677 9688
rect 611 9638 677 9654
rect 807 9688 873 9704
rect 807 9654 823 9688
rect 857 9654 873 9688
rect 807 9638 873 9654
rect 1003 9688 1069 9704
rect 1003 9654 1019 9688
rect 1053 9654 1069 9688
rect 1003 9638 1069 9654
rect 428 9607 468 9638
rect 526 9607 566 9633
rect 624 9607 664 9638
rect 722 9607 762 9633
rect 820 9607 860 9638
rect 918 9607 958 9633
rect 1016 9607 1056 9638
rect 1114 9607 1154 9633
rect 428 8381 468 8407
rect 526 8376 566 8407
rect 624 8381 664 8407
rect 722 8376 762 8407
rect 820 8381 860 8407
rect 918 8376 958 8407
rect 1016 8381 1056 8407
rect 1114 8376 1154 8407
rect 513 8360 579 8376
rect 513 8326 529 8360
rect 563 8326 579 8360
rect 513 8310 579 8326
rect 709 8360 775 8376
rect 709 8326 725 8360
rect 759 8326 775 8360
rect 709 8310 775 8326
rect 905 8360 971 8376
rect 905 8326 921 8360
rect 955 8326 971 8360
rect 905 8310 971 8326
rect 1101 8360 1167 8376
rect 1101 8326 1117 8360
rect 1151 8326 1167 8360
rect 1101 8310 1167 8326
rect 513 8252 579 8268
rect 513 8218 529 8252
rect 563 8218 579 8252
rect 513 8202 579 8218
rect 709 8252 775 8268
rect 709 8218 725 8252
rect 759 8218 775 8252
rect 709 8202 775 8218
rect 905 8252 971 8268
rect 905 8218 921 8252
rect 955 8218 971 8252
rect 905 8202 971 8218
rect 1101 8252 1167 8268
rect 1101 8218 1117 8252
rect 1151 8218 1167 8252
rect 1101 8202 1167 8218
rect 428 8171 468 8197
rect 526 8171 566 8202
rect 624 8171 664 8197
rect 722 8171 762 8202
rect 820 8171 860 8197
rect 918 8171 958 8202
rect 1016 8171 1056 8197
rect 1114 8171 1154 8202
rect -3260 7711 -3230 7737
rect -3260 7479 -3230 7511
rect -3316 7463 -3230 7479
rect -3316 7429 -3300 7463
rect -3266 7429 -3230 7463
rect -3316 7413 -3230 7429
rect -3260 7391 -3230 7413
rect -1896 7746 -1696 7772
rect -1638 7746 -1438 7772
rect -1896 7499 -1696 7546
rect -1896 7465 -1880 7499
rect -1712 7465 -1696 7499
rect -1896 7449 -1696 7465
rect -1638 7499 -1438 7546
rect -1638 7465 -1622 7499
rect -1454 7465 -1438 7499
rect -1638 7449 -1438 7465
rect -3260 7235 -3230 7261
rect -672 7626 -606 7642
rect -672 7592 -656 7626
rect -622 7592 -606 7626
rect -864 7554 -834 7580
rect -672 7576 -606 7592
rect -252 7626 -186 7642
rect -252 7592 -236 7626
rect -202 7592 -186 7626
rect -654 7554 -624 7576
rect -444 7554 -414 7580
rect -252 7576 -186 7592
rect -234 7554 -204 7576
rect -24 7554 6 7580
rect -864 7132 -834 7154
rect -882 7116 -816 7132
rect -654 7128 -624 7154
rect -444 7132 -414 7154
rect -882 7082 -866 7116
rect -832 7082 -816 7116
rect -882 7066 -816 7082
rect -462 7116 -396 7132
rect -234 7128 -204 7154
rect -24 7132 6 7154
rect -462 7082 -446 7116
rect -412 7082 -396 7116
rect -462 7066 -396 7082
rect -42 7116 24 7132
rect -42 7082 -26 7116
rect 8 7082 24 7116
rect -42 7066 24 7082
rect 428 6940 468 6971
rect 526 6945 566 6971
rect 624 6940 664 6971
rect 722 6945 762 6971
rect 820 6940 860 6971
rect 918 6945 958 6971
rect 1016 6940 1056 6971
rect 1114 6945 1154 6971
rect 415 6924 481 6940
rect 415 6890 431 6924
rect 465 6890 481 6924
rect 415 6874 481 6890
rect 611 6924 677 6940
rect 611 6890 627 6924
rect 661 6890 677 6924
rect 611 6874 677 6890
rect 807 6924 873 6940
rect 807 6890 823 6924
rect 857 6890 873 6924
rect 807 6874 873 6890
rect 1003 6924 1069 6940
rect 1003 6890 1019 6924
rect 1053 6890 1069 6924
rect 1003 6874 1069 6890
rect 1427 9688 1493 9704
rect 1427 9654 1443 9688
rect 1477 9654 1493 9688
rect 1427 9638 1493 9654
rect 1623 9688 1689 9704
rect 1623 9654 1639 9688
rect 1673 9654 1689 9688
rect 1623 9638 1689 9654
rect 1819 9688 1885 9704
rect 1819 9654 1835 9688
rect 1869 9654 1885 9688
rect 1819 9638 1885 9654
rect 2015 9688 2081 9704
rect 2015 9654 2031 9688
rect 2065 9654 2081 9688
rect 2015 9638 2081 9654
rect 1440 9607 1480 9638
rect 1538 9607 1578 9633
rect 1636 9607 1676 9638
rect 1734 9607 1774 9633
rect 1832 9607 1872 9638
rect 1930 9607 1970 9633
rect 2028 9607 2068 9638
rect 2126 9607 2166 9633
rect 1440 8381 1480 8407
rect 1538 8376 1578 8407
rect 1636 8381 1676 8407
rect 1734 8376 1774 8407
rect 1832 8381 1872 8407
rect 1930 8376 1970 8407
rect 2028 8381 2068 8407
rect 2126 8376 2166 8407
rect 1525 8360 1591 8376
rect 1525 8326 1541 8360
rect 1575 8326 1591 8360
rect 1525 8310 1591 8326
rect 1721 8360 1787 8376
rect 1721 8326 1737 8360
rect 1771 8326 1787 8360
rect 1721 8310 1787 8326
rect 1917 8360 1983 8376
rect 1917 8326 1933 8360
rect 1967 8326 1983 8360
rect 1917 8310 1983 8326
rect 2113 8360 2179 8376
rect 2113 8326 2129 8360
rect 2163 8326 2179 8360
rect 2113 8310 2179 8326
rect 1525 8252 1591 8268
rect 1525 8218 1541 8252
rect 1575 8218 1591 8252
rect 1525 8202 1591 8218
rect 1721 8252 1787 8268
rect 1721 8218 1737 8252
rect 1771 8218 1787 8252
rect 1721 8202 1787 8218
rect 1917 8252 1983 8268
rect 1917 8218 1933 8252
rect 1967 8218 1983 8252
rect 1917 8202 1983 8218
rect 2113 8252 2179 8268
rect 2113 8218 2129 8252
rect 2163 8218 2179 8252
rect 2113 8202 2179 8218
rect 1440 8171 1480 8197
rect 1538 8171 1578 8202
rect 1636 8171 1676 8197
rect 1734 8171 1774 8202
rect 1832 8171 1872 8197
rect 1930 8171 1970 8202
rect 2028 8171 2068 8197
rect 2126 8171 2166 8202
rect 1440 6940 1480 6971
rect 1538 6945 1578 6971
rect 1636 6940 1676 6971
rect 1734 6945 1774 6971
rect 1832 6940 1872 6971
rect 1930 6945 1970 6971
rect 2028 6940 2068 6971
rect 2126 6945 2166 6971
rect 1427 6924 1493 6940
rect 1427 6890 1443 6924
rect 1477 6890 1493 6924
rect 1427 6874 1493 6890
rect 1623 6924 1689 6940
rect 1623 6890 1639 6924
rect 1673 6890 1689 6924
rect 1623 6874 1689 6890
rect 1819 6924 1885 6940
rect 1819 6890 1835 6924
rect 1869 6890 1885 6924
rect 1819 6874 1885 6890
rect 2015 6924 2081 6940
rect 2015 6890 2031 6924
rect 2065 6890 2081 6924
rect 2015 6874 2081 6890
rect 2558 9680 2588 9706
rect 2558 9449 2588 9480
rect 2540 9433 2606 9449
rect 2540 9399 2556 9433
rect 2590 9399 2606 9433
rect 2540 9383 2606 9399
rect 2540 9086 2606 9102
rect 2540 9052 2556 9086
rect 2590 9052 2606 9086
rect 2540 9036 2606 9052
rect 2558 9014 2588 9036
rect 2558 8788 2588 8814
rect 2540 8634 2606 8650
rect 2540 8600 2556 8634
rect 2590 8600 2606 8634
rect 2540 8584 2606 8600
rect 2558 8562 2588 8584
rect 2558 6940 2588 6962
rect 2540 6924 2606 6940
rect 2540 6890 2556 6924
rect 2590 6890 2606 6924
rect 2540 6874 2606 6890
rect 3000 7110 3100 7136
rect 3158 7110 3258 7136
rect 3000 6972 3100 7010
rect 3000 6938 3016 6972
rect 3084 6938 3100 6972
rect 3000 6922 3100 6938
rect 3158 6972 3258 7010
rect 3158 6938 3174 6972
rect 3242 6938 3258 6972
rect 3158 6922 3258 6938
rect 4088 7414 4154 7430
rect 4088 7380 4104 7414
rect 4138 7380 4154 7414
rect 4010 7342 4040 7368
rect 4088 7364 4154 7380
rect 4280 7414 4346 7430
rect 4280 7380 4296 7414
rect 4330 7380 4346 7414
rect 4106 7342 4136 7364
rect 4202 7342 4232 7368
rect 4280 7364 4346 7380
rect 4298 7342 4328 7364
rect 4010 6940 4040 6962
rect 3992 6924 4058 6940
rect 4106 6936 4136 6962
rect 4202 6940 4232 6962
rect 3992 6890 4008 6924
rect 4042 6890 4058 6924
rect 3992 6874 4058 6890
rect 4184 6924 4250 6940
rect 4298 6936 4328 6962
rect 4184 6890 4200 6924
rect 4234 6890 4250 6924
rect 4184 6874 4250 6890
rect 5134 7452 5200 7468
rect 5134 7418 5150 7452
rect 5184 7418 5200 7452
rect 5134 7402 5200 7418
rect 5326 7452 5392 7468
rect 5326 7418 5342 7452
rect 5376 7418 5392 7452
rect 5326 7402 5392 7418
rect 5056 7371 5086 7397
rect 5152 7371 5182 7402
rect 5248 7371 5278 7397
rect 5344 7371 5374 7402
rect 5056 6940 5086 6971
rect 5152 6945 5182 6971
rect 5248 6940 5278 6971
rect 5344 6945 5374 6971
rect 5038 6924 5104 6940
rect 5038 6890 5054 6924
rect 5088 6890 5104 6924
rect 5038 6874 5104 6890
rect 5230 6924 5296 6940
rect 5230 6890 5246 6924
rect 5280 6890 5296 6924
rect 5230 6874 5296 6890
rect 5746 7452 5812 7468
rect 5746 7418 5762 7452
rect 5796 7418 5812 7452
rect 5746 7402 5812 7418
rect 5938 7452 6004 7468
rect 5938 7418 5954 7452
rect 5988 7418 6004 7452
rect 5938 7402 6004 7418
rect 5668 7371 5698 7397
rect 5764 7371 5794 7402
rect 5860 7371 5890 7397
rect 5956 7371 5986 7402
rect 5668 6940 5698 6971
rect 5764 6945 5794 6971
rect 5860 6940 5890 6971
rect 5956 6945 5986 6971
rect 5650 6924 5716 6940
rect 5650 6890 5666 6924
rect 5700 6890 5716 6924
rect 5650 6874 5716 6890
rect 5842 6924 5908 6940
rect 5842 6890 5858 6924
rect 5892 6890 5908 6924
rect 5842 6874 5908 6890
rect 6496 7434 6562 7450
rect 6496 7400 6512 7434
rect 6546 7400 6562 7434
rect 6418 7362 6448 7388
rect 6496 7384 6562 7400
rect 6688 7434 6754 7450
rect 6688 7400 6704 7434
rect 6738 7400 6754 7434
rect 6514 7362 6544 7384
rect 6610 7362 6640 7388
rect 6688 7384 6754 7400
rect 6706 7362 6736 7384
rect 6418 6940 6448 6962
rect 6400 6924 6466 6940
rect 6514 6936 6544 6962
rect 6610 6940 6640 6962
rect 6400 6890 6416 6924
rect 6450 6890 6466 6924
rect 6400 6874 6466 6890
rect 6592 6924 6658 6940
rect 6706 6936 6736 6962
rect 6592 6890 6608 6924
rect 6642 6890 6658 6924
rect 6592 6874 6658 6890
rect 7108 7434 7174 7450
rect 7108 7400 7124 7434
rect 7158 7400 7174 7434
rect 7030 7362 7060 7388
rect 7108 7384 7174 7400
rect 7300 7434 7366 7450
rect 7300 7400 7316 7434
rect 7350 7400 7366 7434
rect 7126 7362 7156 7384
rect 7222 7362 7252 7388
rect 7300 7384 7366 7400
rect 7318 7362 7348 7384
rect 7030 6940 7060 6962
rect 7012 6924 7078 6940
rect 7126 6936 7156 6962
rect 7222 6940 7252 6962
rect 7012 6890 7028 6924
rect 7062 6890 7078 6924
rect 7012 6874 7078 6890
rect 7204 6924 7270 6940
rect 7318 6936 7348 6962
rect 7204 6890 7220 6924
rect 7254 6890 7270 6924
rect 7204 6874 7270 6890
<< polycont >>
rect -3204 9654 -3136 9688
rect -2932 9654 -2864 9688
rect -2660 9654 -2592 9688
rect -2388 9654 -2320 9688
rect -2116 9654 -2048 9688
rect -1844 9654 -1776 9688
rect -1572 9654 -1504 9688
rect -1300 9654 -1232 9688
rect -1028 9654 -960 9688
rect -756 9654 -688 9688
rect -484 9654 -416 9688
rect -212 9654 -144 9688
rect 60 9654 128 9688
rect -3204 7926 -3136 7960
rect -2932 7926 -2864 7960
rect -2660 7926 -2592 7960
rect -2388 7926 -2320 7960
rect -2116 7926 -2048 7960
rect -1844 7926 -1776 7960
rect -1572 7926 -1504 7960
rect -1300 7926 -1232 7960
rect -1028 7926 -960 7960
rect -756 7926 -688 7960
rect -484 7926 -416 7960
rect -212 7926 -144 7960
rect 60 7926 128 7960
rect 431 9654 465 9688
rect 627 9654 661 9688
rect 823 9654 857 9688
rect 1019 9654 1053 9688
rect 529 8326 563 8360
rect 725 8326 759 8360
rect 921 8326 955 8360
rect 1117 8326 1151 8360
rect 529 8218 563 8252
rect 725 8218 759 8252
rect 921 8218 955 8252
rect 1117 8218 1151 8252
rect -3300 7429 -3266 7463
rect -1880 7465 -1712 7499
rect -1622 7465 -1454 7499
rect -656 7592 -622 7626
rect -236 7592 -202 7626
rect -866 7082 -832 7116
rect -446 7082 -412 7116
rect -26 7082 8 7116
rect 431 6890 465 6924
rect 627 6890 661 6924
rect 823 6890 857 6924
rect 1019 6890 1053 6924
rect 1443 9654 1477 9688
rect 1639 9654 1673 9688
rect 1835 9654 1869 9688
rect 2031 9654 2065 9688
rect 1541 8326 1575 8360
rect 1737 8326 1771 8360
rect 1933 8326 1967 8360
rect 2129 8326 2163 8360
rect 1541 8218 1575 8252
rect 1737 8218 1771 8252
rect 1933 8218 1967 8252
rect 2129 8218 2163 8252
rect 1443 6890 1477 6924
rect 1639 6890 1673 6924
rect 1835 6890 1869 6924
rect 2031 6890 2065 6924
rect 2556 9399 2590 9433
rect 2556 9052 2590 9086
rect 2556 8600 2590 8634
rect 2556 6890 2590 6924
rect 3016 6938 3084 6972
rect 3174 6938 3242 6972
rect 4104 7380 4138 7414
rect 4296 7380 4330 7414
rect 4008 6890 4042 6924
rect 4200 6890 4234 6924
rect 5150 7418 5184 7452
rect 5342 7418 5376 7452
rect 5054 6890 5088 6924
rect 5246 6890 5280 6924
rect 5762 7418 5796 7452
rect 5954 7418 5988 7452
rect 5666 6890 5700 6924
rect 5858 6890 5892 6924
rect 6512 7400 6546 7434
rect 6704 7400 6738 7434
rect 6416 6890 6450 6924
rect 6608 6890 6642 6924
rect 7124 7400 7158 7434
rect 7316 7400 7350 7434
rect 7028 6890 7062 6924
rect 7220 6890 7254 6924
<< xpolycontact >>
rect 2950 9592 3382 9662
rect 6950 9592 7382 9662
rect 2950 9426 3382 9496
rect 6950 9426 7382 9496
rect 2950 9260 3382 9330
rect 6950 9260 7382 9330
rect 2950 9094 3382 9164
rect 6950 9094 7382 9164
rect 2950 8928 3382 8998
rect 6950 8928 7382 8998
rect 2950 8762 3382 8832
rect 6950 8762 7382 8832
rect 2950 8596 3382 8666
rect 6950 8596 7382 8666
rect 2950 8430 3382 8500
rect 6950 8430 7382 8500
rect 2950 8264 3382 8334
rect 6950 8264 7382 8334
rect 2950 8098 3382 8168
rect 6950 8098 7382 8168
rect 2950 7932 3382 8002
rect 6950 7932 7382 8002
<< ppolyres >>
rect 3382 9592 6950 9662
rect 3382 9426 6950 9496
rect 3382 9260 6950 9330
rect 3382 9094 6950 9164
rect 3382 8928 6950 8998
rect 3382 8762 6950 8832
rect 3382 8596 6950 8666
rect 3382 8430 6950 8500
rect 3382 8264 6950 8334
rect 3382 8098 6950 8168
rect 3382 7932 6950 8002
<< locali >>
rect -3490 9890 2730 9930
rect -3490 9850 -3390 9890
rect 2640 9850 2730 9890
rect -3490 9792 2730 9850
rect 2840 9890 7620 9930
rect 2840 9840 2880 9890
rect 7490 9840 7620 9890
rect 2840 9820 7620 9840
rect 2840 9792 7530 9820
rect -3490 9790 2494 9792
rect -3490 7810 -3460 9790
rect -3400 9756 -3284 9790
rect 208 9756 364 9790
rect 1218 9756 1376 9790
rect 2230 9770 2494 9790
rect 2230 9756 2326 9770
rect -3400 9694 -3346 9756
rect -3400 7920 -3380 9694
rect 268 9694 304 9756
rect -3220 9654 -3204 9688
rect -3136 9654 -3120 9688
rect -2948 9654 -2932 9688
rect -2864 9654 -2848 9688
rect -2676 9654 -2660 9688
rect -2592 9654 -2576 9688
rect -2404 9654 -2388 9688
rect -2320 9654 -2304 9688
rect -2132 9654 -2116 9688
rect -2048 9654 -2032 9688
rect -1860 9654 -1844 9688
rect -1776 9654 -1760 9688
rect -1588 9654 -1572 9688
rect -1504 9654 -1488 9688
rect -1316 9654 -1300 9688
rect -1232 9654 -1216 9688
rect -1044 9654 -1028 9688
rect -960 9654 -944 9688
rect -772 9654 -756 9688
rect -688 9654 -672 9688
rect -500 9654 -484 9688
rect -416 9654 -400 9688
rect -228 9654 -212 9688
rect -144 9654 -128 9688
rect 44 9654 60 9688
rect 128 9654 144 9688
rect -3266 9595 -3232 9611
rect -3266 8003 -3232 8019
rect -3108 9595 -3074 9611
rect -3108 8003 -3074 8019
rect -2994 9595 -2960 9611
rect -2994 8003 -2960 8019
rect -2836 9595 -2802 9611
rect -2836 8003 -2802 8019
rect -2722 9595 -2688 9611
rect -2722 8003 -2688 8019
rect -2564 9595 -2530 9611
rect -2564 8003 -2530 8019
rect -2450 9595 -2416 9611
rect -2450 8003 -2416 8019
rect -2292 9595 -2258 9611
rect -2292 8003 -2258 8019
rect -2178 9595 -2144 9611
rect -2178 8003 -2144 8019
rect -2020 9595 -1986 9611
rect -2020 8003 -1986 8019
rect -1906 9595 -1872 9611
rect -1906 8003 -1872 8019
rect -1748 9595 -1714 9611
rect -1748 8003 -1714 8019
rect -1634 9595 -1600 9611
rect -1634 8003 -1600 8019
rect -1476 9595 -1442 9611
rect -1476 8003 -1442 8019
rect -1362 9595 -1328 9611
rect -1362 8003 -1328 8019
rect -1204 9595 -1170 9611
rect -1204 8003 -1170 8019
rect -1090 9595 -1056 9611
rect -1090 8003 -1056 8019
rect -932 9595 -898 9611
rect -932 8003 -898 8019
rect -818 9595 -784 9611
rect -818 8003 -784 8019
rect -660 9595 -626 9611
rect -660 8003 -626 8019
rect -546 9595 -512 9611
rect -546 8003 -512 8019
rect -388 9595 -354 9611
rect -388 8003 -354 8019
rect -274 9595 -240 9611
rect -274 8003 -240 8019
rect -116 9595 -82 9611
rect -116 8003 -82 8019
rect -2 9595 32 9611
rect -2 8003 32 8019
rect 156 9595 190 9611
rect 156 8003 190 8019
rect -3220 7926 -3204 7960
rect -3136 7926 -3120 7960
rect -2948 7926 -2932 7960
rect -2864 7926 -2848 7960
rect -2676 7926 -2660 7960
rect -2592 7926 -2576 7960
rect -2404 7926 -2388 7960
rect -2320 7926 -2304 7960
rect -2132 7926 -2116 7960
rect -2048 7926 -2032 7960
rect -1860 7926 -1844 7960
rect -1776 7926 -1760 7960
rect -1588 7926 -1572 7960
rect -1504 7926 -1488 7960
rect -1316 7926 -1300 7960
rect -1232 7926 -1216 7960
rect -1044 7926 -1028 7960
rect -960 7926 -944 7960
rect -772 7926 -756 7960
rect -688 7926 -672 7960
rect -500 7926 -484 7960
rect -416 7926 -400 7960
rect -228 7926 -212 7960
rect -144 7926 -128 7960
rect 44 7926 60 7960
rect 128 7926 144 7960
rect -3400 7858 -3346 7920
rect 268 7920 270 9694
rect 1280 9694 1314 9756
rect 415 9654 431 9688
rect 465 9654 481 9688
rect 611 9654 627 9688
rect 661 9654 677 9688
rect 807 9654 823 9688
rect 857 9654 873 9688
rect 1003 9654 1019 9688
rect 1053 9654 1069 9688
rect 382 9595 416 9611
rect 382 8403 416 8419
rect 480 9595 514 9611
rect 480 8403 514 8419
rect 578 9595 612 9611
rect 578 8403 612 8419
rect 676 9595 710 9611
rect 676 8403 710 8419
rect 774 9595 808 9611
rect 774 8403 808 8419
rect 872 9595 906 9611
rect 872 8403 906 8419
rect 970 9595 1004 9611
rect 970 8403 1004 8419
rect 1068 9595 1102 9611
rect 1068 8403 1102 8419
rect 1166 9595 1200 9611
rect 1166 8403 1200 8419
rect 513 8326 529 8360
rect 563 8326 579 8360
rect 709 8326 725 8360
rect 759 8326 775 8360
rect 905 8326 921 8360
rect 955 8326 971 8360
rect 1101 8326 1117 8360
rect 1151 8326 1167 8360
rect 513 8218 529 8252
rect 563 8218 579 8252
rect 709 8218 725 8252
rect 759 8218 775 8252
rect 905 8218 921 8252
rect 955 8218 971 8252
rect 1101 8218 1117 8252
rect 1151 8218 1167 8252
rect 268 7858 304 7920
rect -3400 7824 -3284 7858
rect 208 7824 304 7858
rect 382 8159 416 8175
rect -3400 7820 -2022 7824
rect -3400 7810 -2600 7820
rect -3490 7775 -2600 7810
rect -3490 7741 -3351 7775
rect -3317 7741 -3259 7775
rect -3225 7741 -3167 7775
rect -3133 7760 -2600 7775
rect -2080 7761 -2022 7820
rect -2080 7760 -2056 7761
rect -3133 7741 -2056 7760
rect -3490 7710 -3360 7741
rect -3312 7699 -3270 7741
rect -3150 7740 -2056 7741
rect -3312 7665 -3304 7699
rect -3312 7631 -3270 7665
rect -3312 7597 -3304 7631
rect -3312 7563 -3270 7597
rect -3312 7529 -3304 7563
rect -3312 7513 -3270 7529
rect -3236 7699 -3170 7707
rect -3236 7665 -3220 7699
rect -3186 7665 -3170 7699
rect -3236 7631 -3170 7665
rect -3236 7597 -3220 7631
rect -3186 7597 -3170 7631
rect -3236 7570 -3170 7597
rect -3236 7520 -3230 7570
rect -3180 7520 -3170 7570
rect -3236 7511 -3170 7520
rect -3316 7429 -3314 7477
rect -3260 7429 -3250 7477
rect -3316 7379 -3270 7395
rect -3216 7391 -3170 7511
rect -3316 7345 -3304 7379
rect -3316 7311 -3270 7345
rect -3316 7277 -3304 7311
rect -3316 7231 -3270 7277
rect -3236 7379 -3170 7391
rect -3236 7345 -3220 7379
rect -3186 7345 -3170 7379
rect -1312 7761 -1278 7824
rect -1942 7734 -1908 7750
rect -1942 7542 -1908 7558
rect -1684 7734 -1650 7750
rect -1684 7542 -1650 7558
rect -1426 7734 -1392 7750
rect -1426 7542 -1392 7558
rect -1896 7465 -1880 7499
rect -1712 7465 -1696 7499
rect -1638 7465 -1622 7499
rect -1454 7465 -1438 7499
rect -2056 7396 -2022 7459
rect -1312 7396 -1278 7459
rect -2056 7362 -1960 7396
rect -1374 7362 -1278 7396
rect -1028 7694 -932 7728
rect 74 7694 170 7728
rect -1028 7632 -994 7694
rect -3236 7311 -3170 7345
rect -3236 7277 -3220 7311
rect -3186 7277 -3170 7311
rect -3236 7265 -3170 7277
rect -3380 7220 -3351 7231
rect -3490 7197 -3351 7220
rect -3317 7197 -3259 7231
rect -3225 7197 -3167 7231
rect -3133 7197 -3104 7231
rect -3490 6800 -3110 7197
rect 136 7632 170 7694
rect -672 7592 -656 7626
rect -622 7592 -606 7626
rect -252 7592 -236 7626
rect -202 7592 -186 7626
rect -914 7542 -880 7558
rect -914 7150 -880 7166
rect -818 7542 -784 7558
rect -818 7150 -784 7166
rect -704 7542 -670 7558
rect -704 7150 -670 7166
rect -608 7542 -574 7558
rect -608 7150 -574 7166
rect -494 7542 -460 7558
rect -494 7150 -460 7166
rect -398 7542 -364 7558
rect -398 7150 -364 7166
rect -284 7542 -250 7558
rect -284 7150 -250 7166
rect -188 7542 -154 7558
rect -188 7150 -154 7166
rect -74 7542 -40 7558
rect -74 7150 -40 7166
rect 22 7542 56 7558
rect 22 7150 56 7166
rect -882 7082 -866 7116
rect -832 7082 -816 7116
rect -462 7082 -446 7116
rect -412 7082 -396 7116
rect -42 7082 -26 7116
rect 8 7082 24 7116
rect -1028 7014 -994 7076
rect 136 7014 170 7076
rect -1028 6980 -932 7014
rect 74 6980 170 7014
rect -1020 6800 160 6980
rect -3490 6720 160 6800
rect 268 6822 302 7824
rect 382 6967 416 6983
rect 480 8159 514 8175
rect 480 6967 514 6983
rect 578 8159 612 8175
rect 578 6967 612 6983
rect 676 8159 710 8175
rect 676 6967 710 6983
rect 774 8159 808 8175
rect 774 6967 808 6983
rect 872 8159 906 8175
rect 872 6967 906 6983
rect 970 8159 1004 8175
rect 970 6967 1004 6983
rect 1068 8159 1102 8175
rect 1068 6967 1102 6983
rect 1166 8159 1200 8175
rect 1166 6967 1200 6983
rect 415 6890 431 6924
rect 465 6890 481 6924
rect 611 6890 627 6924
rect 661 6890 677 6924
rect 807 6890 823 6924
rect 857 6890 873 6924
rect 1003 6890 1019 6924
rect 1053 6890 1069 6924
rect 2292 9694 2326 9756
rect 1427 9654 1443 9688
rect 1477 9654 1493 9688
rect 1623 9654 1639 9688
rect 1673 9654 1689 9688
rect 1819 9654 1835 9688
rect 1869 9654 1885 9688
rect 2015 9654 2031 9688
rect 2065 9654 2081 9688
rect 1394 9595 1428 9611
rect 1394 8403 1428 8419
rect 1492 9595 1526 9611
rect 1492 8403 1526 8419
rect 1590 9595 1624 9611
rect 1590 8403 1624 8419
rect 1688 9595 1722 9611
rect 1688 8403 1722 8419
rect 1786 9595 1820 9611
rect 1786 8403 1820 8419
rect 1884 9595 1918 9611
rect 1884 8403 1918 8419
rect 1982 9595 2016 9611
rect 1982 8403 2016 8419
rect 2080 9595 2114 9611
rect 2080 8403 2114 8419
rect 2178 9595 2212 9611
rect 2178 8403 2212 8419
rect 1525 8326 1541 8360
rect 1575 8326 1591 8360
rect 1721 8326 1737 8360
rect 1771 8326 1787 8360
rect 1917 8326 1933 8360
rect 1967 8326 1983 8360
rect 2113 8326 2129 8360
rect 2163 8326 2179 8360
rect 1525 8218 1541 8252
rect 1575 8218 1591 8252
rect 1721 8218 1737 8252
rect 1771 8218 1787 8252
rect 1917 8218 1933 8252
rect 1967 8218 1983 8252
rect 2113 8218 2129 8252
rect 2163 8218 2179 8252
rect 1394 8159 1428 8175
rect 1394 6967 1428 6983
rect 1492 8159 1526 8175
rect 1492 6967 1526 6983
rect 1590 8159 1624 8175
rect 1590 6967 1624 6983
rect 1688 8159 1722 8175
rect 1688 6967 1722 6983
rect 1786 8159 1820 8175
rect 1786 6967 1820 6983
rect 1884 8159 1918 8175
rect 1884 6967 1918 6983
rect 1982 8159 2016 8175
rect 1982 6967 2016 6983
rect 2080 8159 2114 8175
rect 2080 6967 2114 6983
rect 2178 8159 2212 8175
rect 2178 6967 2212 6983
rect 1427 6890 1443 6924
rect 1477 6890 1493 6924
rect 1623 6890 1639 6924
rect 1673 6890 1689 6924
rect 1819 6890 1835 6924
rect 1869 6890 1885 6924
rect 2015 6890 2031 6924
rect 2065 6890 2081 6924
rect 1280 6822 1314 6884
rect 2398 9758 2494 9770
rect 2652 9758 2748 9792
rect 2398 9695 2432 9758
rect 2714 9695 2748 9758
rect 2512 9668 2546 9684
rect 2512 9476 2546 9492
rect 2600 9668 2634 9684
rect 2600 9476 2634 9492
rect 2540 9399 2556 9433
rect 2590 9399 2606 9433
rect 2398 9330 2432 9393
rect 2714 9330 2748 9393
rect 2398 9296 2494 9330
rect 2652 9296 2748 9330
rect 2820 9758 2916 9792
rect 7416 9758 7530 9792
rect 2820 9696 2854 9758
rect 2292 6822 2326 6884
rect 268 6788 364 6822
rect 1218 6788 1376 6822
rect 2230 6788 2326 6822
rect 2398 9154 2494 9188
rect 2652 9154 2748 9188
rect 2398 9092 2432 9154
rect 2714 9092 2748 9154
rect 2540 9052 2556 9086
rect 2590 9052 2606 9086
rect 2512 9002 2546 9018
rect 2512 8810 2546 8826
rect 2600 9002 2634 9018
rect 2600 8810 2634 8826
rect 2398 8736 2432 8798
rect 2714 8736 2748 8798
rect 2398 8702 2494 8736
rect 2652 8702 2748 8736
rect 2398 8640 2432 8702
rect 2714 8640 2748 8702
rect 2540 8600 2556 8634
rect 2590 8600 2606 8634
rect 2512 8550 2546 8566
rect 2432 6974 2512 7030
rect 2432 6970 2546 6974
rect 2432 6884 2460 6970
rect 2512 6958 2546 6970
rect 2600 8550 2634 8566
rect 2600 6958 2634 6974
rect 2540 6890 2556 6924
rect 2590 6890 2606 6924
rect 2398 6822 2460 6884
rect 7478 9696 7530 9758
rect 2820 7836 2854 7898
rect 7512 7898 7530 9696
rect 7478 7836 7530 7898
rect 2820 7802 2916 7836
rect 7416 7802 7530 7836
rect 4910 7610 6130 7640
rect 4910 7554 4940 7610
rect 6080 7554 6130 7610
rect 4892 7550 4940 7554
rect 6080 7550 6150 7554
rect 4892 7520 4988 7550
rect 5442 7520 5600 7550
rect 6054 7520 6150 7550
rect 7490 7536 7530 7802
rect 3846 7482 3942 7516
rect 4396 7482 4492 7516
rect 3846 7420 3880 7482
rect 2714 6822 2748 6884
rect 2398 6788 2494 6822
rect 2652 6800 2748 6822
rect 2820 7224 2916 7258
rect 3342 7224 3438 7258
rect 2820 7162 2854 7224
rect 3404 7162 3438 7224
rect 2954 7098 2988 7114
rect 2954 7006 2988 7022
rect 3112 7098 3146 7114
rect 3112 7006 3146 7022
rect 3270 7098 3304 7114
rect 3270 7006 3304 7022
rect 3000 6938 3016 6972
rect 3084 6938 3100 6972
rect 3158 6938 3174 6972
rect 3242 6938 3258 6972
rect 2820 6834 2854 6896
rect 3404 6834 3438 6896
rect 2820 6800 2916 6834
rect 3342 6800 3438 6834
rect 4458 7420 4492 7482
rect 4088 7380 4104 7414
rect 4138 7380 4154 7414
rect 4280 7380 4296 7414
rect 4330 7380 4346 7414
rect 3960 7330 3994 7346
rect 3960 6958 3994 6974
rect 4056 7330 4090 7346
rect 4056 6958 4090 6974
rect 4152 7330 4186 7346
rect 4152 6958 4186 6974
rect 4248 7330 4282 7346
rect 4248 6958 4282 6974
rect 4344 7330 4378 7346
rect 4344 6958 4378 6974
rect 3992 6890 4008 6924
rect 4042 6890 4058 6924
rect 4184 6890 4200 6924
rect 4234 6890 4250 6924
rect 3846 6822 3880 6884
rect 4458 6822 4492 6884
rect 3846 6800 3942 6822
rect 2652 6788 3942 6800
rect 4396 6788 4492 6822
rect 4892 7458 4926 7520
rect 5504 7458 5538 7520
rect 5134 7418 5150 7452
rect 5184 7418 5200 7452
rect 5326 7418 5342 7452
rect 5376 7418 5392 7452
rect 5006 7359 5040 7375
rect 5006 6967 5040 6983
rect 5102 7359 5136 7375
rect 5102 6967 5136 6983
rect 5198 7359 5232 7375
rect 5198 6967 5232 6983
rect 5294 7359 5328 7375
rect 5294 6967 5328 6983
rect 5390 7359 5424 7375
rect 5390 6967 5424 6983
rect 5038 6890 5054 6924
rect 5088 6890 5104 6924
rect 5230 6890 5246 6924
rect 5280 6890 5296 6924
rect 4892 6822 4926 6884
rect 6116 7458 6150 7520
rect 5746 7418 5762 7452
rect 5796 7418 5812 7452
rect 5938 7418 5954 7452
rect 5988 7418 6004 7452
rect 5618 7359 5652 7375
rect 5618 6967 5652 6983
rect 5714 7359 5748 7375
rect 5714 6967 5748 6983
rect 5810 7359 5844 7375
rect 5810 6967 5844 6983
rect 5906 7359 5940 7375
rect 5906 6967 5940 6983
rect 6002 7359 6036 7375
rect 6002 6967 6036 6983
rect 5650 6890 5666 6924
rect 5700 6890 5716 6924
rect 5842 6890 5858 6924
rect 5892 6890 5908 6924
rect 5504 6822 5538 6884
rect 6116 6822 6150 6884
rect 4892 6788 4988 6822
rect 5442 6788 5600 6822
rect 6054 6788 6150 6822
rect 6254 7502 6350 7536
rect 6804 7502 6962 7536
rect 7416 7502 7530 7536
rect 6254 7440 6288 7502
rect 6866 7440 6900 7502
rect 6496 7400 6512 7434
rect 6546 7400 6562 7434
rect 6688 7400 6704 7434
rect 6738 7400 6754 7434
rect 6368 7350 6402 7366
rect 6368 6958 6402 6974
rect 6464 7350 6498 7366
rect 6464 6958 6498 6974
rect 6560 7350 6594 7366
rect 6560 6958 6594 6974
rect 6656 7350 6690 7366
rect 6656 6958 6690 6974
rect 6752 7350 6786 7366
rect 6752 6958 6786 6974
rect 6400 6890 6416 6924
rect 6450 6890 6466 6924
rect 6592 6890 6608 6924
rect 6642 6890 6658 6924
rect 6254 6822 6288 6884
rect 7478 7440 7530 7502
rect 7108 7400 7124 7434
rect 7158 7400 7174 7434
rect 7300 7400 7316 7434
rect 7350 7400 7366 7434
rect 6980 7350 7014 7366
rect 6980 6958 7014 6974
rect 7076 7350 7110 7366
rect 7076 6958 7110 6974
rect 7172 7350 7206 7366
rect 7172 6958 7206 6974
rect 7268 7350 7302 7366
rect 7268 6958 7302 6974
rect 7364 7350 7398 7366
rect 7364 6958 7398 6974
rect 7012 6890 7028 6924
rect 7062 6890 7078 6924
rect 7204 6890 7220 6924
rect 7254 6890 7270 6924
rect 6866 6822 6900 6884
rect 7512 6884 7530 7440
rect 7478 6822 7530 6884
rect 6254 6788 6350 6822
rect 6804 6788 6962 6822
rect 7416 6788 7530 6822
rect 2400 6720 4480 6788
rect 6260 6750 7530 6788
rect 7570 6750 7620 9820
rect 6260 6720 7620 6750
rect -3490 6690 7620 6720
rect -3490 6630 -3400 6690
rect 7480 6630 7620 6690
rect -3490 6580 7620 6630
<< viali >>
rect -3390 9850 2640 9890
rect 2880 9840 7490 9890
rect -3460 7810 -3400 9790
rect -3204 9654 -3136 9688
rect -2932 9654 -2864 9688
rect -2660 9654 -2592 9688
rect -2388 9654 -2320 9688
rect -2116 9654 -2048 9688
rect -1844 9654 -1776 9688
rect -1572 9654 -1504 9688
rect -1300 9654 -1232 9688
rect -1028 9654 -960 9688
rect -756 9654 -688 9688
rect -484 9654 -416 9688
rect -212 9654 -144 9688
rect 60 9654 128 9688
rect -3266 8019 -3232 9595
rect -3108 8019 -3074 9595
rect -2994 8019 -2960 9595
rect -2836 8019 -2802 9595
rect -2722 8019 -2688 9595
rect -2564 8019 -2530 9595
rect -2450 8019 -2416 9595
rect -2292 8019 -2258 9595
rect -2178 8019 -2144 9595
rect -2020 8019 -1986 9595
rect -1906 8019 -1872 9595
rect -1748 8019 -1714 9595
rect -1634 8019 -1600 9595
rect -1476 8019 -1442 9595
rect -1362 8019 -1328 9595
rect -1204 8019 -1170 9595
rect -1090 8019 -1056 9595
rect -932 8019 -898 9595
rect -818 8019 -784 9595
rect -660 8019 -626 9595
rect -546 8019 -512 9595
rect -388 8019 -354 9595
rect -274 8019 -240 9595
rect -116 8019 -82 9595
rect -2 8019 32 9595
rect 156 8019 190 9595
rect -3204 7926 -3136 7960
rect -2932 7926 -2864 7960
rect -2660 7926 -2592 7960
rect -2388 7926 -2320 7960
rect -2116 7926 -2048 7960
rect -1844 7926 -1776 7960
rect -1572 7926 -1504 7960
rect -1300 7926 -1232 7960
rect -1028 7926 -960 7960
rect -756 7926 -688 7960
rect -484 7926 -416 7960
rect -212 7926 -144 7960
rect 60 7926 128 7960
rect 431 9654 465 9688
rect 627 9654 661 9688
rect 823 9654 857 9688
rect 1019 9654 1053 9688
rect 382 8419 416 9595
rect 480 8419 514 9595
rect 578 8419 612 9595
rect 676 8419 710 9595
rect 774 8419 808 9595
rect 872 8419 906 9595
rect 970 8419 1004 9595
rect 1068 8419 1102 9595
rect 1166 8419 1200 9595
rect 529 8326 563 8360
rect 725 8326 759 8360
rect 921 8326 955 8360
rect 1117 8326 1151 8360
rect 529 8218 563 8252
rect 725 8218 759 8252
rect 921 8218 955 8252
rect 1117 8218 1151 8252
rect -3351 7741 -3317 7775
rect -3259 7741 -3225 7775
rect -3167 7741 -3133 7775
rect -2600 7760 -2080 7820
rect -3230 7563 -3180 7570
rect -3230 7529 -3220 7563
rect -3220 7529 -3186 7563
rect -3186 7529 -3180 7563
rect -3230 7520 -3180 7529
rect -3314 7463 -3260 7477
rect -3314 7429 -3300 7463
rect -3300 7429 -3266 7463
rect -3266 7429 -3260 7463
rect -1942 7558 -1908 7734
rect -1684 7558 -1650 7734
rect -1426 7558 -1392 7734
rect -1880 7465 -1712 7499
rect -1622 7465 -1454 7499
rect -3351 7197 -3317 7231
rect -3259 7197 -3225 7231
rect -3167 7197 -3133 7231
rect -656 7592 -622 7626
rect -236 7592 -202 7626
rect -914 7166 -880 7542
rect -818 7166 -784 7542
rect -704 7166 -670 7542
rect -608 7166 -574 7542
rect -494 7166 -460 7542
rect -398 7166 -364 7542
rect -284 7166 -250 7542
rect -188 7166 -154 7542
rect -74 7166 -40 7542
rect 22 7166 56 7542
rect -866 7082 -832 7116
rect -446 7082 -412 7116
rect -26 7082 8 7116
rect 382 6983 416 8159
rect 480 6983 514 8159
rect 578 6983 612 8159
rect 676 6983 710 8159
rect 774 6983 808 8159
rect 872 6983 906 8159
rect 970 6983 1004 8159
rect 1068 6983 1102 8159
rect 1166 6983 1200 8159
rect 431 6890 465 6924
rect 627 6890 661 6924
rect 823 6890 857 6924
rect 1019 6890 1053 6924
rect 1443 9654 1477 9688
rect 1639 9654 1673 9688
rect 1835 9654 1869 9688
rect 2031 9654 2065 9688
rect 1394 8419 1428 9595
rect 1492 8419 1526 9595
rect 1590 8419 1624 9595
rect 1688 8419 1722 9595
rect 1786 8419 1820 9595
rect 1884 8419 1918 9595
rect 1982 8419 2016 9595
rect 2080 8419 2114 9595
rect 2178 8419 2212 9595
rect 1541 8326 1575 8360
rect 1737 8326 1771 8360
rect 1933 8326 1967 8360
rect 2129 8326 2163 8360
rect 1541 8218 1575 8252
rect 1737 8218 1771 8252
rect 1933 8218 1967 8252
rect 2129 8218 2163 8252
rect 1394 6983 1428 8159
rect 1492 6983 1526 8159
rect 1590 6983 1624 8159
rect 1688 6983 1722 8159
rect 1786 6983 1820 8159
rect 1884 6983 1918 8159
rect 1982 6983 2016 8159
rect 2080 6983 2114 8159
rect 2178 6983 2212 8159
rect 1443 6890 1477 6924
rect 1639 6890 1673 6924
rect 1835 6890 1869 6924
rect 2031 6890 2065 6924
rect 2512 9492 2546 9668
rect 2600 9492 2634 9668
rect 2556 9399 2590 9433
rect 2556 9052 2590 9086
rect 2512 8826 2546 9002
rect 2600 8826 2634 9002
rect 2556 8600 2590 8634
rect 2512 6974 2546 8550
rect 2600 6974 2634 8550
rect 2556 6890 2590 6924
rect 2968 9608 3365 9646
rect 6967 9608 7364 9646
rect 2968 9442 3365 9480
rect 6967 9442 7364 9480
rect 2968 9276 3365 9314
rect 6967 9276 7364 9314
rect 2968 9110 3365 9148
rect 6967 9110 7364 9148
rect 2968 8944 3365 8982
rect 6967 8944 7364 8982
rect 2968 8778 3365 8816
rect 6967 8778 7364 8816
rect 2968 8612 3365 8650
rect 6967 8612 7364 8650
rect 2968 8446 3365 8484
rect 6967 8446 7364 8484
rect 2968 8280 3365 8318
rect 6967 8280 7364 8318
rect 2968 8114 3365 8152
rect 6967 8114 7364 8152
rect 2968 7948 3365 7986
rect 6967 7948 7364 7986
rect 4940 7554 6080 7610
rect 4940 7550 4988 7554
rect 4988 7550 5442 7554
rect 5442 7550 5600 7554
rect 5600 7550 6054 7554
rect 6054 7550 6080 7554
rect 2954 7022 2988 7098
rect 3112 7022 3146 7098
rect 3270 7022 3304 7098
rect 3016 6938 3084 6972
rect 3174 6938 3242 6972
rect 4104 7380 4138 7414
rect 4296 7380 4330 7414
rect 3960 6974 3994 7330
rect 4056 6974 4090 7330
rect 4152 6974 4186 7330
rect 4248 6974 4282 7330
rect 4344 6974 4378 7330
rect 4008 6890 4042 6924
rect 4200 6890 4234 6924
rect 5150 7418 5184 7452
rect 5342 7418 5376 7452
rect 5006 6983 5040 7359
rect 5102 6983 5136 7359
rect 5198 6983 5232 7359
rect 5294 6983 5328 7359
rect 5390 6983 5424 7359
rect 5054 6890 5088 6924
rect 5246 6890 5280 6924
rect 5762 7418 5796 7452
rect 5954 7418 5988 7452
rect 5618 6983 5652 7359
rect 5714 6983 5748 7359
rect 5810 6983 5844 7359
rect 5906 6983 5940 7359
rect 6002 6983 6036 7359
rect 5666 6890 5700 6924
rect 5858 6890 5892 6924
rect 6512 7400 6546 7434
rect 6704 7400 6738 7434
rect 6368 6974 6402 7350
rect 6464 6974 6498 7350
rect 6560 6974 6594 7350
rect 6656 6974 6690 7350
rect 6752 6974 6786 7350
rect 6416 6890 6450 6924
rect 6608 6890 6642 6924
rect 7124 7400 7158 7434
rect 7316 7400 7350 7434
rect 6980 6974 7014 7350
rect 7076 6974 7110 7350
rect 7172 6974 7206 7350
rect 7268 6974 7302 7350
rect 7364 6974 7398 7350
rect 7028 6890 7062 6924
rect 7220 6890 7254 6924
rect 7530 6750 7570 9820
rect -3400 6630 7480 6690
<< metal1 >>
rect -3490 9890 2730 9930
rect -3490 9850 -3390 9890
rect 2640 9850 2730 9890
rect -3490 9790 2730 9850
rect -3600 8690 -3590 8750
rect -3530 8690 -3520 8750
rect -3580 7640 -3540 8690
rect -3490 7810 -3460 9790
rect -3400 9770 2730 9790
rect 2840 9890 7620 9930
rect 2840 9840 2880 9890
rect 7490 9840 7620 9890
rect 2840 9820 7620 9840
rect 2840 9770 7530 9820
rect -3400 9400 -3360 9770
rect -3230 9710 150 9720
rect -3230 9688 40 9710
rect 110 9688 150 9710
rect -3230 9654 -3204 9688
rect -3136 9654 -2932 9688
rect -2864 9654 -2660 9688
rect -2592 9654 -2388 9688
rect -2320 9654 -2116 9688
rect -2048 9654 -1844 9688
rect -1776 9654 -1572 9688
rect -1504 9654 -1300 9688
rect -1232 9654 -1028 9688
rect -960 9654 -756 9688
rect -688 9654 -484 9688
rect -416 9654 -212 9688
rect -144 9654 40 9688
rect 128 9654 150 9688
rect -3230 9640 40 9654
rect 110 9640 150 9654
rect -1480 9607 -1440 9640
rect -3272 9595 -3226 9607
rect -3272 9400 -3266 9595
rect -3400 9350 -3266 9400
rect -3400 7840 -3360 9350
rect -3272 8019 -3266 9350
rect -3232 9400 -3226 9595
rect -3114 9595 -3068 9607
rect -3114 9400 -3108 9595
rect -3232 9350 -3108 9400
rect -3232 8019 -3226 9350
rect -3272 8007 -3226 8019
rect -3114 8019 -3108 9350
rect -3074 8019 -3068 9595
rect -3000 9595 -2954 9607
rect -3000 9400 -2994 9595
rect -2960 9400 -2954 9595
rect -2842 9595 -2796 9607
rect -3020 9340 -3010 9400
rect -2950 9340 -2940 9400
rect -3000 8902 -2994 9340
rect -2960 8902 -2954 9340
rect -3024 8842 -3014 8902
rect -2954 8842 -2944 8902
rect -3000 8292 -2994 8842
rect -2960 8292 -2954 8842
rect -2842 8752 -2836 9595
rect -2802 8752 -2796 9595
rect -2728 9595 -2682 9607
rect -2728 9400 -2722 9595
rect -2688 9400 -2682 9595
rect -2570 9595 -2524 9607
rect -2750 9340 -2740 9400
rect -2680 9340 -2670 9400
rect -2728 8902 -2722 9340
rect -2688 8902 -2682 9340
rect -2754 8842 -2744 8902
rect -2684 8842 -2674 8902
rect -2864 8692 -2854 8752
rect -2794 8692 -2784 8752
rect -3024 8232 -3014 8292
rect -2954 8232 -2944 8292
rect -3114 8007 -3068 8019
rect -3000 8019 -2994 8232
rect -2960 8019 -2954 8232
rect -3000 8007 -2954 8019
rect -2842 8019 -2836 8692
rect -2802 8019 -2796 8692
rect -2728 8292 -2722 8842
rect -2688 8292 -2682 8842
rect -2570 8752 -2564 9595
rect -2530 8752 -2524 9595
rect -2456 9595 -2410 9607
rect -2456 9400 -2450 9595
rect -2416 9400 -2410 9595
rect -2298 9595 -2252 9607
rect -2470 9340 -2460 9400
rect -2400 9340 -2390 9400
rect -2456 8902 -2450 9340
rect -2416 8902 -2410 9340
rect -2474 8842 -2464 8902
rect -2404 8842 -2394 8902
rect -2594 8692 -2584 8752
rect -2524 8692 -2514 8752
rect -2754 8232 -2744 8292
rect -2684 8232 -2674 8292
rect -2842 8007 -2796 8019
rect -2728 8019 -2722 8232
rect -2688 8019 -2682 8232
rect -2728 8007 -2682 8019
rect -2570 8019 -2564 8692
rect -2530 8019 -2524 8692
rect -2456 8292 -2450 8842
rect -2416 8292 -2410 8842
rect -2298 8582 -2292 9595
rect -2258 8582 -2252 9595
rect -2184 9595 -2138 9607
rect -2184 9400 -2178 9595
rect -2144 9400 -2138 9595
rect -2026 9595 -1980 9607
rect -2200 9340 -2190 9400
rect -2130 9340 -2120 9400
rect -2184 8902 -2178 9340
rect -2144 8902 -2138 9340
rect -2204 8842 -2194 8902
rect -2134 8842 -2124 8902
rect -2314 8522 -2304 8582
rect -2244 8522 -2234 8582
rect -2474 8232 -2464 8292
rect -2404 8232 -2394 8292
rect -2570 8007 -2524 8019
rect -2456 8019 -2450 8232
rect -2416 8019 -2410 8232
rect -2298 8134 -2292 8522
rect -2258 8134 -2252 8522
rect -2184 8292 -2178 8842
rect -2144 8292 -2138 8842
rect -2026 8582 -2020 9595
rect -1986 8582 -1980 9595
rect -1912 9595 -1866 9607
rect -1912 9400 -1906 9595
rect -1872 9400 -1866 9595
rect -1754 9595 -1708 9607
rect -1930 9340 -1920 9400
rect -1860 9340 -1850 9400
rect -1912 8902 -1906 9340
rect -1872 8902 -1866 9340
rect -1934 8842 -1924 8902
rect -1864 8842 -1854 8902
rect -2044 8522 -2034 8582
rect -1974 8522 -1964 8582
rect -2204 8232 -2194 8292
rect -2134 8232 -2124 8292
rect -2318 8074 -2308 8134
rect -2248 8074 -2238 8134
rect -2456 8007 -2410 8019
rect -2298 8019 -2292 8074
rect -2258 8019 -2252 8074
rect -2298 8007 -2252 8019
rect -2184 8019 -2178 8232
rect -2144 8019 -2138 8232
rect -2026 8134 -2020 8522
rect -1986 8134 -1980 8522
rect -1912 8292 -1906 8842
rect -1872 8292 -1866 8842
rect -1754 8582 -1748 9595
rect -1714 8582 -1708 9595
rect -1640 9595 -1594 9607
rect -1640 9400 -1634 9595
rect -1600 9400 -1594 9595
rect -1482 9595 -1436 9607
rect -1660 9340 -1650 9400
rect -1590 9340 -1580 9400
rect -1640 8902 -1634 9340
rect -1600 8902 -1594 9340
rect -1664 8842 -1654 8902
rect -1594 8842 -1584 8902
rect -1774 8522 -1764 8582
rect -1704 8522 -1694 8582
rect -1934 8232 -1924 8292
rect -1864 8232 -1854 8292
rect -2048 8074 -2038 8134
rect -1978 8074 -1968 8134
rect -2184 8007 -2138 8019
rect -2026 8019 -2020 8074
rect -1986 8019 -1980 8074
rect -2026 8007 -1980 8019
rect -1912 8019 -1906 8232
rect -1872 8019 -1866 8232
rect -1754 8134 -1748 8522
rect -1714 8134 -1708 8522
rect -1640 8292 -1634 8842
rect -1600 8292 -1594 8842
rect -1664 8232 -1654 8292
rect -1594 8232 -1584 8292
rect -1778 8074 -1768 8134
rect -1708 8074 -1698 8134
rect -1912 8007 -1866 8019
rect -1754 8019 -1748 8074
rect -1714 8019 -1708 8074
rect -1754 8007 -1708 8019
rect -1640 8019 -1634 8232
rect -1600 8019 -1594 8232
rect -1640 8007 -1594 8019
rect -1482 8019 -1476 9595
rect -1442 8019 -1436 9595
rect -1368 9595 -1322 9607
rect -1368 9400 -1362 9595
rect -1328 9400 -1322 9595
rect -1210 9595 -1164 9607
rect -1390 9340 -1380 9400
rect -1320 9340 -1310 9400
rect -1368 8902 -1362 9340
rect -1328 8902 -1322 9340
rect -1394 8842 -1384 8902
rect -1324 8842 -1314 8902
rect -1368 8292 -1362 8842
rect -1328 8292 -1322 8842
rect -1210 8582 -1204 9595
rect -1170 8582 -1164 9595
rect -1096 9595 -1050 9607
rect -1096 9400 -1090 9595
rect -1056 9400 -1050 9595
rect -938 9595 -892 9607
rect -1110 9340 -1100 9400
rect -1040 9340 -1030 9400
rect -1096 8902 -1090 9340
rect -1056 8902 -1050 9340
rect -1114 8842 -1104 8902
rect -1044 8842 -1034 8902
rect -1234 8522 -1224 8582
rect -1164 8522 -1154 8582
rect -1394 8232 -1384 8292
rect -1324 8232 -1314 8292
rect -1482 8007 -1436 8019
rect -1368 8019 -1362 8232
rect -1328 8019 -1322 8232
rect -1210 8134 -1204 8522
rect -1170 8134 -1164 8522
rect -1096 8292 -1090 8842
rect -1056 8292 -1050 8842
rect -938 8582 -932 9595
rect -898 8582 -892 9595
rect -824 9595 -778 9607
rect -824 9400 -818 9595
rect -784 9400 -778 9595
rect -666 9595 -620 9607
rect -840 9340 -830 9400
rect -770 9340 -760 9400
rect -824 8902 -818 9340
rect -784 8902 -778 9340
rect -844 8842 -834 8902
rect -774 8842 -764 8902
rect -954 8522 -944 8582
rect -884 8522 -874 8582
rect -1114 8232 -1104 8292
rect -1044 8232 -1034 8292
rect -1238 8074 -1228 8134
rect -1168 8074 -1158 8134
rect -1368 8007 -1322 8019
rect -1210 8019 -1204 8074
rect -1170 8019 -1164 8074
rect -1210 8007 -1164 8019
rect -1096 8019 -1090 8232
rect -1056 8019 -1050 8232
rect -938 8134 -932 8522
rect -898 8134 -892 8522
rect -824 8292 -818 8842
rect -784 8292 -778 8842
rect -666 8582 -660 9595
rect -626 8582 -620 9595
rect -552 9595 -506 9607
rect -552 9400 -546 9595
rect -512 9400 -506 9595
rect -394 9595 -348 9607
rect -570 9340 -560 9400
rect -500 9340 -490 9400
rect -552 8902 -546 9340
rect -512 8902 -506 9340
rect -574 8842 -564 8902
rect -504 8842 -494 8902
rect -684 8522 -674 8582
rect -614 8522 -604 8582
rect -844 8232 -834 8292
rect -774 8232 -764 8292
rect -958 8074 -948 8134
rect -888 8074 -878 8134
rect -1096 8007 -1050 8019
rect -938 8019 -932 8074
rect -898 8019 -892 8074
rect -938 8007 -892 8019
rect -824 8019 -818 8232
rect -784 8019 -778 8232
rect -666 8134 -660 8522
rect -626 8134 -620 8522
rect -552 8292 -546 8842
rect -512 8292 -506 8842
rect -394 8462 -388 9595
rect -354 8462 -348 9595
rect -280 9595 -234 9607
rect -280 9400 -274 9595
rect -240 9400 -234 9595
rect -122 9595 -76 9607
rect -300 9340 -290 9400
rect -230 9340 -220 9400
rect -280 8902 -274 9340
rect -240 8902 -234 9340
rect -304 8842 -294 8902
rect -234 8842 -224 8902
rect -414 8402 -404 8462
rect -344 8402 -334 8462
rect -574 8232 -564 8292
rect -504 8232 -494 8292
rect -688 8074 -678 8134
rect -618 8074 -608 8134
rect -824 8007 -778 8019
rect -666 8019 -660 8074
rect -626 8019 -620 8074
rect -666 8007 -620 8019
rect -552 8019 -546 8232
rect -512 8019 -506 8232
rect -552 8007 -506 8019
rect -394 8019 -388 8402
rect -354 8019 -348 8402
rect -280 8292 -274 8842
rect -240 8292 -234 8842
rect -122 8750 -116 9595
rect -82 8750 -76 9595
rect -8 9595 38 9607
rect -140 8690 -130 8750
rect -70 8690 -60 8750
rect -304 8232 -294 8292
rect -234 8232 -224 8292
rect -394 8007 -348 8019
rect -280 8019 -274 8232
rect -240 8019 -234 8232
rect -280 8007 -234 8019
rect -122 8019 -116 8690
rect -82 8019 -76 8690
rect -122 8007 -76 8019
rect -8 8019 -2 9595
rect 32 9380 38 9595
rect 150 9595 196 9607
rect 150 9380 156 9595
rect 32 9330 156 9380
rect 32 8019 38 9330
rect -8 8007 38 8019
rect 150 8019 156 9330
rect 190 9380 196 9595
rect 230 9380 270 9770
rect 419 9690 477 9694
rect 615 9690 673 9694
rect 811 9690 869 9694
rect 1007 9690 1065 9694
rect 400 9688 1070 9690
rect 400 9685 431 9688
rect 190 9330 270 9380
rect 300 9655 431 9685
rect 190 8019 196 9330
rect 300 9250 330 9655
rect 400 9654 431 9655
rect 465 9654 627 9688
rect 661 9654 823 9688
rect 857 9654 1019 9688
rect 1053 9654 1070 9688
rect 1431 9688 1489 9694
rect 1431 9685 1443 9688
rect 400 9650 1070 9654
rect 1310 9655 1443 9685
rect 419 9648 477 9650
rect 615 9648 673 9650
rect 811 9648 869 9650
rect 1007 9648 1065 9650
rect 376 9595 422 9607
rect 260 9190 270 9250
rect 330 9190 340 9250
rect 300 8355 330 9190
rect 376 8590 382 9595
rect 416 8590 422 9595
rect 474 9595 520 9607
rect 474 8770 480 9595
rect 514 8770 520 9595
rect 572 9595 618 9607
rect 460 8710 470 8770
rect 530 8710 540 8770
rect 360 8530 370 8590
rect 430 8530 440 8590
rect 376 8419 382 8530
rect 416 8419 422 8530
rect 376 8407 422 8419
rect 474 8419 480 8710
rect 514 8419 520 8710
rect 572 8590 578 9595
rect 612 8590 618 9595
rect 670 9595 716 9607
rect 670 8770 676 9595
rect 710 8770 716 9595
rect 768 9595 814 9607
rect 650 8710 660 8770
rect 720 8710 730 8770
rect 550 8530 560 8590
rect 620 8530 630 8590
rect 474 8407 520 8419
rect 572 8419 578 8530
rect 612 8419 618 8530
rect 572 8407 618 8419
rect 670 8419 676 8710
rect 710 8419 716 8710
rect 768 8590 774 9595
rect 808 8590 814 9595
rect 866 9595 912 9607
rect 866 8770 872 9595
rect 906 8770 912 9595
rect 964 9595 1010 9607
rect 850 8710 860 8770
rect 920 8710 930 8770
rect 750 8530 760 8590
rect 820 8530 830 8590
rect 670 8407 716 8419
rect 768 8419 774 8530
rect 808 8419 814 8530
rect 768 8407 814 8419
rect 866 8419 872 8710
rect 906 8419 912 8710
rect 964 8590 970 9595
rect 1004 8590 1010 9595
rect 1062 9595 1108 9607
rect 1062 8770 1068 9595
rect 1102 8770 1108 9595
rect 1160 9595 1206 9607
rect 1050 8710 1060 8770
rect 1120 8710 1130 8770
rect 950 8530 960 8590
rect 1020 8530 1030 8590
rect 866 8407 912 8419
rect 964 8419 970 8530
rect 1004 8419 1010 8530
rect 964 8407 1010 8419
rect 1062 8419 1068 8710
rect 1102 8419 1108 8710
rect 1160 8590 1166 9595
rect 1200 8590 1206 9595
rect 1310 9130 1340 9655
rect 1431 9654 1443 9655
rect 1477 9685 1489 9688
rect 1627 9688 1685 9694
rect 1627 9685 1639 9688
rect 1477 9655 1639 9685
rect 1477 9654 1489 9655
rect 1431 9648 1489 9654
rect 1627 9654 1639 9655
rect 1673 9685 1685 9688
rect 1823 9688 1881 9694
rect 1823 9685 1835 9688
rect 1673 9655 1835 9685
rect 1673 9654 1685 9655
rect 1627 9648 1685 9654
rect 1823 9654 1835 9655
rect 1869 9685 1881 9688
rect 2019 9688 2077 9694
rect 2019 9685 2031 9688
rect 1869 9655 2031 9685
rect 1869 9654 1881 9655
rect 1823 9648 1881 9654
rect 2019 9654 2031 9655
rect 2065 9654 2077 9688
rect 2019 9648 2077 9654
rect 2390 9650 2400 9710
rect 2460 9650 2470 9710
rect 2506 9668 2552 9680
rect 1388 9595 1434 9607
rect 1280 9070 1290 9130
rect 1350 9070 1360 9130
rect 1140 8530 1150 8590
rect 1210 8530 1220 8590
rect 1062 8407 1108 8419
rect 1160 8419 1166 8530
rect 1200 8419 1206 8530
rect 1160 8407 1206 8419
rect 517 8360 575 8366
rect 517 8355 529 8360
rect 300 8326 529 8355
rect 563 8355 575 8360
rect 713 8360 771 8366
rect 713 8355 725 8360
rect 563 8326 725 8355
rect 759 8355 771 8360
rect 909 8360 967 8366
rect 909 8355 921 8360
rect 759 8326 921 8355
rect 955 8355 967 8360
rect 1090 8355 1100 8370
rect 955 8326 1100 8355
rect 300 8325 1100 8326
rect 517 8320 575 8325
rect 713 8320 771 8325
rect 909 8320 967 8325
rect 1090 8310 1100 8325
rect 1160 8310 1170 8370
rect 1310 8355 1340 9070
rect 1388 8590 1394 9595
rect 1428 8590 1434 9595
rect 1486 9595 1532 9607
rect 1486 8960 1492 9595
rect 1526 8960 1532 9595
rect 1584 9595 1630 9607
rect 1470 8900 1480 8960
rect 1540 8900 1550 8960
rect 1370 8530 1380 8590
rect 1440 8530 1450 8590
rect 1388 8419 1394 8530
rect 1428 8419 1434 8530
rect 1388 8407 1434 8419
rect 1486 8419 1492 8900
rect 1526 8419 1532 8900
rect 1584 8590 1590 9595
rect 1624 8590 1630 9595
rect 1682 9595 1728 9607
rect 1682 8960 1688 9595
rect 1722 8960 1728 9595
rect 1780 9595 1826 9607
rect 1660 8900 1670 8960
rect 1730 8900 1740 8960
rect 1570 8530 1580 8590
rect 1640 8530 1650 8590
rect 1486 8407 1532 8419
rect 1584 8419 1590 8530
rect 1624 8419 1630 8530
rect 1584 8407 1630 8419
rect 1682 8419 1688 8900
rect 1722 8419 1728 8900
rect 1780 8590 1786 9595
rect 1820 8590 1826 9595
rect 1878 9595 1924 9607
rect 1878 8960 1884 9595
rect 1918 8960 1924 9595
rect 1976 9595 2022 9607
rect 1860 8900 1870 8960
rect 1930 8900 1940 8960
rect 1770 8530 1780 8590
rect 1840 8530 1850 8590
rect 1682 8407 1728 8419
rect 1780 8419 1786 8530
rect 1820 8419 1826 8530
rect 1780 8407 1826 8419
rect 1878 8419 1884 8900
rect 1918 8419 1924 8900
rect 1976 8590 1982 9595
rect 2016 8590 2022 9595
rect 2074 9595 2120 9607
rect 2074 8960 2080 9595
rect 2114 8960 2120 9595
rect 2172 9595 2218 9607
rect 2060 8900 2070 8960
rect 2130 8900 2140 8960
rect 1960 8530 1970 8590
rect 2030 8530 2040 8590
rect 1878 8407 1924 8419
rect 1976 8419 1982 8530
rect 2016 8419 2022 8530
rect 1976 8407 2022 8419
rect 2074 8419 2080 8900
rect 2114 8419 2120 8900
rect 2172 8590 2178 9595
rect 2212 8590 2218 9595
rect 2410 9570 2440 9650
rect 2506 9570 2512 9668
rect 2410 9540 2512 9570
rect 2506 9492 2512 9540
rect 2546 9492 2552 9668
rect 2506 9480 2552 9492
rect 2594 9668 2640 9680
rect 2594 9492 2600 9668
rect 2634 9540 2640 9668
rect 2670 9540 2700 9770
rect 2970 9652 2980 9660
rect 2956 9646 2980 9652
rect 3050 9652 3060 9660
rect 3050 9646 3377 9652
rect 2956 9608 2968 9646
rect 3365 9608 3377 9646
rect 2956 9602 2980 9608
rect 2970 9590 2980 9602
rect 3050 9602 3377 9608
rect 6955 9646 7376 9652
rect 6955 9608 6967 9646
rect 7364 9608 7376 9646
rect 6955 9602 7376 9608
rect 3050 9590 3060 9602
rect 2634 9510 2700 9540
rect 2634 9492 2640 9510
rect 2594 9480 2640 9492
rect 6990 9486 7360 9602
rect 2956 9480 3377 9486
rect 6955 9480 7376 9486
rect 2956 9442 2968 9480
rect 3365 9442 3760 9480
rect 2956 9440 3760 9442
rect 2544 9433 2602 9439
rect 2956 9436 3377 9440
rect 2544 9399 2556 9433
rect 2590 9425 2602 9433
rect 2590 9399 2720 9425
rect 2544 9395 2720 9399
rect 2544 9393 2602 9395
rect 2544 9090 2602 9092
rect 2420 9086 2610 9090
rect 2420 9052 2556 9086
rect 2590 9052 2610 9086
rect 2420 9050 2610 9052
rect 2310 8900 2320 8960
rect 2380 8900 2390 8960
rect 2250 8710 2260 8770
rect 2320 8710 2330 8770
rect 2160 8530 2170 8590
rect 2230 8530 2240 8590
rect 2074 8407 2120 8419
rect 2172 8419 2178 8530
rect 2212 8419 2218 8530
rect 2172 8407 2218 8419
rect 1529 8360 1587 8366
rect 1529 8355 1541 8360
rect 1235 8326 1541 8355
rect 1575 8355 1587 8360
rect 1725 8360 1783 8366
rect 1725 8355 1737 8360
rect 1575 8326 1737 8355
rect 1771 8355 1783 8360
rect 1921 8360 1979 8366
rect 1921 8355 1933 8360
rect 1771 8326 1933 8355
rect 1967 8355 1979 8360
rect 2117 8360 2175 8366
rect 2117 8355 2129 8360
rect 1967 8326 2129 8355
rect 2163 8326 2175 8360
rect 1235 8325 2175 8326
rect 517 8255 575 8258
rect 713 8255 771 8258
rect 909 8255 967 8258
rect 1105 8255 1163 8258
rect 1235 8255 1265 8325
rect 1529 8320 1587 8325
rect 1725 8320 1783 8325
rect 1921 8320 1979 8325
rect 2117 8320 2175 8325
rect 1370 8255 1380 8280
rect 150 8007 196 8019
rect 300 8252 1265 8255
rect 300 8225 529 8252
rect -1480 7970 -1440 8007
rect -3230 7960 150 7970
rect -3230 7926 -3204 7960
rect -3136 7926 -2932 7960
rect -2864 7926 -2660 7960
rect -2592 7926 -2388 7960
rect -2320 7926 -2116 7960
rect -2048 7926 -1844 7960
rect -1776 7926 -1572 7960
rect -1504 7926 -1300 7960
rect -1232 7926 -1028 7960
rect -960 7926 -756 7960
rect -688 7926 -484 7960
rect -416 7926 -212 7960
rect -144 7926 60 7960
rect 128 7926 150 7960
rect -3230 7890 150 7926
rect -3400 7820 -2030 7840
rect -3400 7810 -2600 7820
rect -3490 7775 -2600 7810
rect -3490 7741 -3351 7775
rect -3317 7741 -3259 7775
rect -3225 7741 -3167 7775
rect -3133 7760 -2600 7775
rect -2080 7760 -2030 7820
rect -3133 7741 -2030 7760
rect -3490 7710 -2030 7741
rect -1948 7734 -1902 7746
rect -1948 7650 -1942 7734
rect -3600 7580 -3590 7640
rect -3530 7580 -3520 7640
rect -2010 7620 -1942 7650
rect -3242 7570 -3168 7576
rect -3242 7520 -3230 7570
rect -3180 7560 -3168 7570
rect -3180 7530 -2990 7560
rect -3180 7520 -3168 7530
rect -3242 7514 -3168 7520
rect -3326 7480 -3248 7483
rect -3330 7420 -3320 7480
rect -3260 7423 -3248 7480
rect -3260 7420 -3250 7423
rect -3380 7260 -3104 7262
rect -3490 7231 -3080 7260
rect -3490 7197 -3351 7231
rect -3317 7197 -3259 7231
rect -3225 7197 -3167 7231
rect -3133 7197 -3080 7231
rect -3020 7210 -2990 7530
rect -2740 7420 -2730 7480
rect -2670 7420 -2660 7480
rect -3490 6800 -3080 7197
rect -3050 7150 -3040 7210
rect -2980 7150 -2970 7210
rect -2720 6940 -2680 7420
rect -2010 7070 -1980 7620
rect -1948 7558 -1942 7620
rect -1908 7558 -1902 7734
rect -1690 7734 -1644 7746
rect -1690 7640 -1684 7734
rect -1650 7640 -1644 7734
rect -1432 7734 -1386 7746
rect -1432 7640 -1426 7734
rect -1392 7640 -1386 7734
rect -260 7700 -250 7760
rect -190 7700 -180 7760
rect -1710 7580 -1700 7640
rect -1640 7580 -1630 7640
rect -1450 7580 -1440 7640
rect -1380 7580 -1370 7640
rect -240 7632 -190 7700
rect -668 7630 -610 7632
rect -248 7630 -190 7632
rect -670 7626 -190 7630
rect -670 7592 -656 7626
rect -622 7592 -236 7626
rect -202 7592 -190 7626
rect -670 7590 -190 7592
rect -668 7586 -610 7590
rect -1948 7546 -1902 7558
rect -1690 7558 -1684 7580
rect -1650 7558 -1644 7580
rect -1690 7546 -1644 7558
rect -1432 7558 -1426 7580
rect -1392 7558 -1386 7580
rect -1432 7546 -1386 7558
rect -400 7554 -360 7590
rect -248 7586 -190 7590
rect -920 7542 -874 7554
rect -1892 7499 -1700 7505
rect -1892 7465 -1880 7499
rect -1712 7465 -1700 7499
rect -1892 7459 -1700 7465
rect -1634 7499 -1442 7505
rect -1634 7465 -1622 7499
rect -1454 7465 -1442 7499
rect -1634 7459 -1442 7465
rect -1820 7400 -1780 7459
rect -1840 7340 -1830 7400
rect -1770 7340 -1760 7400
rect -1560 7310 -1520 7459
rect -920 7320 -914 7542
rect -880 7400 -874 7542
rect -824 7542 -778 7554
rect -824 7400 -818 7542
rect -880 7370 -818 7400
rect -880 7320 -874 7370
rect -940 7310 -930 7320
rect -1580 7250 -1570 7310
rect -1510 7250 -1500 7310
rect -1030 7270 -930 7310
rect -2020 7010 -2010 7070
rect -1950 7010 -1940 7070
rect -2740 6880 -2730 6940
rect -2670 6880 -2660 6940
rect -1030 6800 -980 7270
rect -940 7260 -930 7270
rect -870 7310 -860 7320
rect -824 7310 -818 7370
rect -870 7270 -818 7310
rect -870 7260 -860 7270
rect -920 7166 -914 7260
rect -880 7166 -874 7260
rect -920 7154 -874 7166
rect -824 7166 -818 7270
rect -784 7166 -778 7542
rect -710 7542 -664 7554
rect -710 7320 -704 7542
rect -670 7320 -664 7542
rect -614 7542 -568 7554
rect -614 7410 -608 7542
rect -574 7410 -568 7542
rect -500 7542 -454 7554
rect -630 7350 -620 7410
rect -560 7350 -550 7410
rect -730 7260 -720 7320
rect -660 7260 -650 7320
rect -824 7154 -778 7166
rect -710 7166 -704 7260
rect -670 7166 -664 7260
rect -710 7154 -664 7166
rect -614 7166 -608 7350
rect -574 7166 -568 7350
rect -500 7320 -494 7542
rect -460 7320 -454 7542
rect -404 7542 -358 7554
rect -520 7260 -510 7320
rect -450 7260 -440 7320
rect -614 7154 -568 7166
rect -500 7166 -494 7260
rect -460 7166 -454 7260
rect -500 7154 -454 7166
rect -404 7166 -398 7542
rect -364 7166 -358 7542
rect -290 7542 -244 7554
rect -290 7320 -284 7542
rect -250 7320 -244 7542
rect -194 7542 -148 7554
rect -194 7410 -188 7542
rect -154 7410 -148 7542
rect -80 7542 -34 7554
rect -210 7350 -200 7410
rect -140 7350 -130 7410
rect -310 7260 -300 7320
rect -240 7260 -230 7320
rect -404 7154 -358 7166
rect -290 7166 -284 7260
rect -250 7166 -244 7260
rect -290 7154 -244 7166
rect -194 7166 -188 7350
rect -154 7166 -148 7350
rect -80 7320 -74 7542
rect -40 7390 -34 7542
rect 16 7542 62 7554
rect 16 7390 22 7542
rect -40 7360 22 7390
rect -40 7320 -34 7360
rect -100 7260 -90 7320
rect -30 7310 -20 7320
rect 16 7310 22 7360
rect -30 7270 22 7310
rect -30 7260 -20 7270
rect -194 7154 -148 7166
rect -80 7166 -74 7260
rect -40 7166 -34 7260
rect -80 7154 -34 7166
rect 16 7166 22 7270
rect 56 7166 62 7542
rect 16 7154 62 7166
rect -400 7122 -360 7154
rect -878 7120 -820 7122
rect -458 7120 -360 7122
rect -38 7120 20 7122
rect -890 7116 40 7120
rect -890 7082 -866 7116
rect -832 7082 -446 7116
rect -412 7082 -26 7116
rect 8 7082 40 7116
rect -890 7080 40 7082
rect -878 7076 -820 7080
rect -458 7076 -400 7080
rect -38 7076 20 7080
rect 300 6925 330 8225
rect 517 8218 529 8225
rect 563 8225 725 8252
rect 563 8218 575 8225
rect 517 8212 575 8218
rect 713 8218 725 8225
rect 759 8225 921 8252
rect 759 8218 771 8225
rect 713 8212 771 8218
rect 909 8218 921 8225
rect 955 8225 1117 8252
rect 955 8218 967 8225
rect 909 8212 967 8218
rect 1105 8218 1117 8225
rect 1151 8225 1265 8252
rect 1310 8225 1380 8255
rect 1151 8218 1163 8225
rect 1105 8212 1163 8218
rect 376 8159 422 8171
rect 376 8130 382 8159
rect 416 8130 422 8159
rect 474 8159 520 8171
rect 360 8070 370 8130
rect 430 8070 440 8130
rect 376 6983 382 8070
rect 416 6983 422 8070
rect 474 7600 480 8159
rect 514 7600 520 8159
rect 572 8159 618 8171
rect 572 8130 578 8159
rect 612 8130 618 8159
rect 670 8159 716 8171
rect 560 8070 570 8130
rect 630 8070 640 8130
rect 460 7540 470 7600
rect 530 7540 540 7600
rect 376 6971 422 6983
rect 474 6983 480 7540
rect 514 6983 520 7540
rect 474 6971 520 6983
rect 572 6983 578 8070
rect 612 6983 618 8070
rect 670 7600 676 8159
rect 710 7600 716 8159
rect 768 8159 814 8171
rect 768 8130 774 8159
rect 808 8130 814 8159
rect 866 8159 912 8171
rect 750 8070 760 8130
rect 820 8070 830 8130
rect 650 7540 660 7600
rect 720 7540 730 7600
rect 572 6971 618 6983
rect 670 6983 676 7540
rect 710 6983 716 7540
rect 670 6971 716 6983
rect 768 6983 774 8070
rect 808 6983 814 8070
rect 866 7600 872 8159
rect 906 7600 912 8159
rect 964 8159 1010 8171
rect 964 8130 970 8159
rect 1004 8130 1010 8159
rect 1062 8159 1108 8171
rect 950 8070 960 8130
rect 1020 8070 1030 8130
rect 850 7540 860 7600
rect 920 7540 930 7600
rect 768 6971 814 6983
rect 866 6983 872 7540
rect 906 6983 912 7540
rect 866 6971 912 6983
rect 964 6983 970 8070
rect 1004 6983 1010 8070
rect 1062 7600 1068 8159
rect 1102 7600 1108 8159
rect 1160 8159 1206 8171
rect 1160 8130 1166 8159
rect 1200 8130 1206 8159
rect 1140 8070 1150 8130
rect 1210 8070 1220 8130
rect 1050 7540 1060 7600
rect 1120 7540 1130 7600
rect 964 6971 1010 6983
rect 1062 6983 1068 7540
rect 1102 6983 1108 7540
rect 1062 6971 1108 6983
rect 1160 6983 1166 8070
rect 1200 6983 1206 8070
rect 1160 6971 1206 6983
rect 419 6925 477 6930
rect 615 6925 673 6930
rect 811 6925 869 6930
rect 1007 6925 1065 6930
rect 300 6924 1065 6925
rect 300 6895 431 6924
rect 419 6890 431 6895
rect 465 6895 627 6924
rect 465 6890 477 6895
rect 419 6884 477 6890
rect 615 6890 627 6895
rect 661 6895 823 6924
rect 661 6890 673 6895
rect 615 6884 673 6890
rect 811 6890 823 6895
rect 857 6895 1019 6924
rect 857 6890 869 6895
rect 811 6884 869 6890
rect 1007 6890 1019 6895
rect 1053 6890 1065 6924
rect 1310 6925 1340 8225
rect 1370 8220 1380 8225
rect 1440 8255 1450 8280
rect 1529 8255 1587 8258
rect 1725 8255 1783 8258
rect 1921 8255 1979 8258
rect 2117 8255 2175 8258
rect 1440 8252 2175 8255
rect 1440 8225 1541 8252
rect 1440 8220 1450 8225
rect 1529 8218 1541 8225
rect 1575 8225 1737 8252
rect 1575 8218 1587 8225
rect 1529 8212 1587 8218
rect 1725 8218 1737 8225
rect 1771 8225 1933 8252
rect 1771 8218 1783 8225
rect 1725 8212 1783 8218
rect 1921 8218 1933 8225
rect 1967 8225 2129 8252
rect 1967 8218 1979 8225
rect 1921 8212 1979 8218
rect 2117 8218 2129 8225
rect 2163 8218 2175 8252
rect 2117 8212 2175 8218
rect 1388 8159 1434 8171
rect 1388 8130 1394 8159
rect 1428 8130 1434 8159
rect 1486 8159 1532 8171
rect 1370 8070 1380 8130
rect 1440 8070 1450 8130
rect 1388 6983 1394 8070
rect 1428 6983 1434 8070
rect 1486 8000 1492 8159
rect 1526 8000 1532 8159
rect 1584 8159 1630 8171
rect 1584 8130 1590 8159
rect 1624 8130 1630 8159
rect 1682 8159 1728 8171
rect 1570 8070 1580 8130
rect 1640 8070 1650 8130
rect 1470 7940 1480 8000
rect 1540 7940 1550 8000
rect 1388 6971 1434 6983
rect 1486 6983 1492 7940
rect 1526 6983 1532 7940
rect 1486 6971 1532 6983
rect 1584 6983 1590 8070
rect 1624 6983 1630 8070
rect 1682 8000 1688 8159
rect 1722 8000 1728 8159
rect 1780 8159 1826 8171
rect 1780 8130 1786 8159
rect 1820 8130 1826 8159
rect 1878 8159 1924 8171
rect 1770 8070 1780 8130
rect 1840 8070 1850 8130
rect 1660 7940 1670 8000
rect 1730 7940 1740 8000
rect 1584 6971 1630 6983
rect 1682 6983 1688 7940
rect 1722 6983 1728 7940
rect 1682 6971 1728 6983
rect 1780 6983 1786 8070
rect 1820 6983 1826 8070
rect 1878 8000 1884 8159
rect 1918 8000 1924 8159
rect 1976 8159 2022 8171
rect 1976 8130 1982 8159
rect 2016 8130 2022 8159
rect 2074 8159 2120 8171
rect 1960 8070 1970 8130
rect 2030 8070 2040 8130
rect 1860 7940 1870 8000
rect 1930 7940 1940 8000
rect 1780 6971 1826 6983
rect 1878 6983 1884 7940
rect 1918 6983 1924 7940
rect 1878 6971 1924 6983
rect 1976 6983 1982 8070
rect 2016 6983 2022 8070
rect 2074 8000 2080 8159
rect 2114 8000 2120 8159
rect 2172 8159 2218 8171
rect 2172 8130 2178 8159
rect 2212 8130 2218 8159
rect 2160 8070 2170 8130
rect 2230 8070 2240 8130
rect 2060 7940 2070 8000
rect 2130 7940 2140 8000
rect 1976 6971 2022 6983
rect 2074 6983 2080 7940
rect 2114 6983 2120 7940
rect 2074 6971 2120 6983
rect 2172 6983 2178 8070
rect 2212 6983 2218 8070
rect 2270 8000 2310 8710
rect 2250 7940 2260 8000
rect 2320 7940 2330 8000
rect 2360 7600 2390 8900
rect 2310 7540 2320 7600
rect 2380 7540 2390 7600
rect 2420 7210 2450 9050
rect 2544 9046 2602 9050
rect 2506 9002 2552 9014
rect 2594 9010 2640 9014
rect 2506 8910 2512 9002
rect 2546 8910 2552 9002
rect 2580 8950 2590 9010
rect 2650 8950 2660 9010
rect 2480 8850 2490 8910
rect 2550 8850 2560 8910
rect 2506 8826 2512 8850
rect 2546 8826 2552 8850
rect 2506 8814 2552 8826
rect 2594 8826 2600 8950
rect 2634 8826 2640 8950
rect 2594 8814 2640 8826
rect 2544 8634 2602 8640
rect 2544 8630 2556 8634
rect 2540 8600 2556 8630
rect 2590 8630 2602 8634
rect 2690 8630 2720 9395
rect 3550 9320 3560 9380
rect 3620 9320 3630 9380
rect 2956 9314 3377 9320
rect 2956 9276 2968 9314
rect 3365 9276 3377 9314
rect 2956 9270 3377 9276
rect 3030 9154 3290 9270
rect 2956 9148 3377 9154
rect 2956 9110 2968 9148
rect 3365 9110 3377 9148
rect 2956 9104 3377 9110
rect 2830 8950 2840 9010
rect 2900 8950 2910 9010
rect 2956 8982 3377 8988
rect 2590 8600 2720 8630
rect 2544 8594 2602 8600
rect 2506 8550 2552 8562
rect 2390 7150 2400 7210
rect 2460 7150 2470 7210
rect 2506 7030 2512 8550
rect 2172 6971 2218 6983
rect 2400 6980 2512 7030
rect 1431 6925 1489 6930
rect 1627 6925 1685 6930
rect 1823 6925 1881 6930
rect 2019 6925 2077 6930
rect 1310 6924 2077 6925
rect 1310 6895 1443 6924
rect 1007 6884 1065 6890
rect 1431 6890 1443 6895
rect 1477 6895 1639 6924
rect 1477 6890 1489 6895
rect 1431 6884 1489 6890
rect 1627 6890 1639 6895
rect 1673 6895 1835 6924
rect 1673 6890 1685 6895
rect 1627 6884 1685 6890
rect 1823 6890 1835 6895
rect 1869 6895 2031 6924
rect 1869 6890 1881 6895
rect 1823 6884 1881 6890
rect 2019 6890 2031 6895
rect 2065 6890 2077 6924
rect 2019 6884 2077 6890
rect 2400 6800 2460 6980
rect 2506 6974 2512 6980
rect 2546 6974 2552 8550
rect 2594 8550 2640 8562
rect 2594 7880 2600 8550
rect 2634 7880 2640 8550
rect 2580 7820 2590 7880
rect 2650 7820 2660 7880
rect 2506 6962 2552 6974
rect 2594 6974 2600 7820
rect 2634 6974 2640 7820
rect 2594 6962 2640 6974
rect 2530 6870 2540 6930
rect 2600 6915 2610 6930
rect 2690 6915 2720 8600
rect 2600 6885 2720 6915
rect 2750 8850 2760 8910
rect 2820 8850 2830 8910
rect 2600 6870 2610 6885
rect 2750 6800 2780 8850
rect 2860 8460 2890 8950
rect 2956 8944 2968 8982
rect 3365 8944 3377 8982
rect 2956 8938 3377 8944
rect 3040 8822 3300 8938
rect 2956 8816 3377 8822
rect 2956 8778 2968 8816
rect 3365 8778 3377 8816
rect 2956 8772 3377 8778
rect 2956 8650 3377 8656
rect 2956 8612 2968 8650
rect 3365 8612 3377 8650
rect 2956 8606 3377 8612
rect 3060 8490 3320 8606
rect 2956 8484 3377 8490
rect 2840 8400 2850 8460
rect 2910 8400 2920 8460
rect 2956 8446 2968 8484
rect 3365 8446 3377 8484
rect 2956 8440 3377 8446
rect 2956 8318 3377 8324
rect 2956 8280 2968 8318
rect 3365 8280 3377 8318
rect 2956 8274 3377 8280
rect 2830 8160 2840 8220
rect 2900 8160 2910 8220
rect 2840 8000 2900 8160
rect 3040 8158 3300 8274
rect 2956 8152 3377 8158
rect 2956 8114 2968 8152
rect 3365 8114 3377 8152
rect 2956 8108 3377 8114
rect 2830 7940 2840 8000
rect 2900 7940 2910 8000
rect 2956 7986 3377 7992
rect 2956 7948 2968 7986
rect 3365 7948 3377 7986
rect 2956 7942 3377 7948
rect 2990 7940 3050 7942
rect 2990 7750 3020 7940
rect 3575 7885 3605 9320
rect 3120 7855 3605 7885
rect 3720 7880 3760 9440
rect 6955 9442 6967 9480
rect 7364 9442 7376 9480
rect 6955 9436 7376 9442
rect 5020 9400 5100 9410
rect 5020 9340 5030 9400
rect 5090 9340 5100 9400
rect 4770 8220 4850 8230
rect 4770 8160 4780 8220
rect 4840 8160 4850 8220
rect 2960 7690 2970 7750
rect 3030 7690 3040 7750
rect 2930 7110 2940 7170
rect 3000 7110 3010 7170
rect 3120 7110 3150 7855
rect 3700 7820 3710 7880
rect 3770 7820 3780 7880
rect 3350 7780 3410 7790
rect 3350 7710 3410 7720
rect 3470 7710 3530 7720
rect 3250 7110 3260 7170
rect 3320 7110 3330 7170
rect 2948 7098 2994 7110
rect 2948 7022 2954 7098
rect 2988 7022 2994 7098
rect 2948 7010 2994 7022
rect 3106 7098 3152 7110
rect 3106 7022 3112 7098
rect 3146 7022 3152 7098
rect 3106 7010 3152 7022
rect 3264 7098 3310 7110
rect 3264 7022 3270 7098
rect 3304 7022 3310 7098
rect 3264 7010 3310 7022
rect 3004 6972 3096 6978
rect 3004 6938 3016 6972
rect 3084 6938 3096 6972
rect 3004 6932 3096 6938
rect 3162 6975 3254 6978
rect 3370 6975 3400 7710
rect 3470 7640 3530 7650
rect 3162 6972 3400 6975
rect 3162 6938 3174 6972
rect 3242 6945 3400 6972
rect 3242 6938 3254 6945
rect 3162 6932 3254 6938
rect 3035 6895 3065 6932
rect 3490 6895 3520 7640
rect 4660 7540 4670 7600
rect 4730 7540 4740 7600
rect 4550 7430 4560 7490
rect 4620 7430 4630 7490
rect 3590 7360 3600 7420
rect 3660 7360 3670 7420
rect 4080 7370 4090 7430
rect 4150 7370 4160 7430
rect 4284 7414 4342 7420
rect 4284 7410 4296 7414
rect 4280 7380 4296 7410
rect 4330 7410 4342 7414
rect 4330 7380 4380 7410
rect 4280 7370 4380 7380
rect 3610 7170 3640 7360
rect 4350 7342 4380 7370
rect 3954 7330 4000 7342
rect 3954 7190 3960 7330
rect 3994 7190 4000 7330
rect 4050 7330 4096 7342
rect 3590 7110 3600 7170
rect 3660 7110 3670 7170
rect 3730 7130 3740 7190
rect 3800 7130 3810 7190
rect 3940 7130 3950 7190
rect 4010 7130 4020 7190
rect 3610 6930 3640 7110
rect 3730 6930 3810 7130
rect 3954 6974 3960 7130
rect 3994 6974 4000 7130
rect 4050 7070 4056 7330
rect 4090 7070 4096 7330
rect 4146 7330 4192 7342
rect 4146 7190 4152 7330
rect 4186 7190 4192 7330
rect 4242 7330 4288 7342
rect 4242 7300 4248 7330
rect 4282 7300 4288 7330
rect 4338 7330 4384 7342
rect 4230 7240 4240 7300
rect 4300 7240 4310 7300
rect 4130 7130 4140 7190
rect 4200 7130 4210 7190
rect 4030 7010 4040 7070
rect 4100 7010 4110 7070
rect 3954 6962 4000 6974
rect 4050 6974 4056 7010
rect 4090 6974 4096 7010
rect 4050 6962 4096 6974
rect 4146 6974 4152 7130
rect 4186 6974 4192 7130
rect 4146 6962 4192 6974
rect 4242 6974 4248 7240
rect 4282 6974 4288 7240
rect 4338 7190 4344 7330
rect 4378 7190 4384 7330
rect 4550 7300 4630 7430
rect 4550 7240 4560 7300
rect 4620 7240 4630 7300
rect 4320 7130 4330 7190
rect 4390 7130 4400 7190
rect 4242 6962 4288 6974
rect 4338 6974 4344 7130
rect 4378 6974 4384 7130
rect 4338 6962 4384 6974
rect 4550 7010 4560 7070
rect 4620 7010 4630 7070
rect 3035 6865 3520 6895
rect 3590 6870 3600 6930
rect 3660 6870 3670 6930
rect 3730 6924 4060 6930
rect 3730 6890 4008 6924
rect 4042 6890 4060 6924
rect 3730 6880 4060 6890
rect 3730 6800 3810 6880
rect 4180 6870 4190 6930
rect 4250 6870 4260 6930
rect 4550 6890 4630 7010
rect 4660 7020 4740 7540
rect 4770 7380 4850 8160
rect 5020 7640 5100 9340
rect 6955 9314 7376 9320
rect 6955 9310 6967 9314
rect 6230 9276 6967 9310
rect 7364 9276 7376 9314
rect 6230 9270 7376 9276
rect 6230 7690 6270 9270
rect 6955 9148 7376 9154
rect 6955 9110 6967 9148
rect 7364 9110 7376 9148
rect 6955 9104 7376 9110
rect 7060 8988 7320 9104
rect 6955 8982 7376 8988
rect 6955 8944 6967 8982
rect 7364 8944 7376 8982
rect 6955 8938 7376 8944
rect 6955 8816 7376 8822
rect 6955 8778 6967 8816
rect 7364 8778 7376 8816
rect 6955 8772 7376 8778
rect 7070 8656 7330 8772
rect 6955 8650 7376 8656
rect 6955 8612 6967 8650
rect 7364 8612 7376 8650
rect 6955 8606 7376 8612
rect 6955 8484 7376 8490
rect 6670 8400 6680 8460
rect 6740 8400 6750 8460
rect 6955 8446 6967 8484
rect 7364 8446 7376 8484
rect 6955 8440 7376 8446
rect 6700 7990 6730 8400
rect 7050 8324 7310 8440
rect 6955 8318 7376 8324
rect 6955 8280 6967 8318
rect 7364 8280 7376 8318
rect 6955 8274 7376 8280
rect 6955 8152 7376 8158
rect 6955 8114 6967 8152
rect 7364 8135 7376 8152
rect 7364 8114 7460 8135
rect 6955 8108 7460 8114
rect 7285 8105 7460 8108
rect 6955 7990 7376 7992
rect 6700 7986 7376 7990
rect 6700 7960 6967 7986
rect 4910 7610 6130 7640
rect 6210 7630 6220 7690
rect 6280 7630 6290 7690
rect 4910 7550 4940 7610
rect 6080 7550 6130 7610
rect 4910 7530 6130 7550
rect 5135 7452 6145 7465
rect 5135 7418 5150 7452
rect 5184 7418 5342 7452
rect 5376 7418 5762 7452
rect 5796 7418 5954 7452
rect 5988 7418 6145 7452
rect 5135 7415 6145 7418
rect 5138 7412 5196 7415
rect 5330 7412 5388 7415
rect 5750 7412 5808 7415
rect 5942 7412 6000 7415
rect 4770 7320 4780 7380
rect 4840 7320 4850 7380
rect 4770 7310 4850 7320
rect 5000 7359 5046 7371
rect 5000 7020 5006 7359
rect 5040 7020 5046 7359
rect 5096 7359 5142 7371
rect 5096 7130 5102 7359
rect 5136 7130 5142 7359
rect 5192 7359 5238 7371
rect 5080 7070 5090 7130
rect 5150 7070 5160 7130
rect 4660 6960 4670 7020
rect 4730 6960 4740 7020
rect 4980 6960 4990 7020
rect 5050 6960 5060 7020
rect 5096 6983 5102 7070
rect 5136 6983 5142 7070
rect 5192 7020 5198 7359
rect 5232 7020 5238 7359
rect 5288 7359 5334 7371
rect 5288 7130 5294 7359
rect 5328 7130 5334 7359
rect 5384 7359 5430 7371
rect 5270 7070 5280 7130
rect 5340 7070 5350 7130
rect 5096 6971 5142 6983
rect 5170 6960 5180 7020
rect 5240 6960 5250 7020
rect 5288 6983 5294 7070
rect 5328 6983 5334 7070
rect 5384 7020 5390 7359
rect 5424 7020 5430 7359
rect 5600 7320 5610 7380
rect 5670 7320 5680 7380
rect 5708 7359 5754 7371
rect 5288 6971 5334 6983
rect 5370 6960 5380 7020
rect 5440 6960 5450 7020
rect 5612 6983 5618 7320
rect 5652 6983 5658 7320
rect 5708 7250 5714 7359
rect 5748 7250 5754 7359
rect 5790 7320 5800 7380
rect 5860 7320 5870 7380
rect 5900 7359 5946 7371
rect 5690 7190 5700 7250
rect 5760 7190 5770 7250
rect 5612 6971 5658 6983
rect 5708 6983 5714 7190
rect 5748 6983 5754 7190
rect 5708 6971 5754 6983
rect 5804 6983 5810 7320
rect 5844 6983 5850 7320
rect 5900 7250 5906 7359
rect 5940 7250 5946 7359
rect 5980 7320 5990 7380
rect 6050 7320 6060 7380
rect 5880 7190 5890 7250
rect 5950 7190 5960 7250
rect 5804 6971 5850 6983
rect 5900 6983 5906 7190
rect 5940 6983 5946 7190
rect 5900 6971 5946 6983
rect 5996 6983 6002 7320
rect 6036 6983 6042 7320
rect 5996 6971 6042 6983
rect 6095 6930 6145 7415
rect 6230 7130 6270 7630
rect 6700 7440 6730 7960
rect 6955 7948 6967 7960
rect 7364 7948 7376 7986
rect 6955 7942 7376 7948
rect 7430 7790 7460 8105
rect 7380 7730 7390 7790
rect 7450 7730 7460 7790
rect 6490 7434 7362 7440
rect 6490 7400 6512 7434
rect 6546 7400 6704 7434
rect 6738 7400 7124 7434
rect 7158 7400 7316 7434
rect 7350 7400 7362 7434
rect 6490 7394 7362 7400
rect 6490 7390 7360 7394
rect 6362 7360 6408 7362
rect 6340 7300 6350 7360
rect 6410 7300 6420 7360
rect 6458 7350 6504 7362
rect 6554 7360 6600 7362
rect 6210 7070 6220 7130
rect 6280 7070 6290 7130
rect 6362 6974 6368 7300
rect 6402 6974 6408 7300
rect 6458 7130 6464 7350
rect 6498 7130 6504 7350
rect 6540 7300 6550 7360
rect 6610 7300 6620 7360
rect 6650 7350 6696 7362
rect 6746 7360 6792 7362
rect 6440 7070 6450 7130
rect 6510 7070 6520 7130
rect 6362 6962 6408 6974
rect 6458 6974 6464 7070
rect 6498 6974 6504 7070
rect 6458 6962 6504 6974
rect 6554 6974 6560 7300
rect 6594 6974 6600 7300
rect 6650 7130 6656 7350
rect 6690 7130 6696 7350
rect 6730 7300 6740 7360
rect 6800 7300 6810 7360
rect 6630 7070 6640 7130
rect 6700 7070 6710 7130
rect 6554 6962 6600 6974
rect 6650 6974 6656 7070
rect 6690 6974 6696 7070
rect 6650 6962 6696 6974
rect 6746 6974 6752 7300
rect 6786 6974 6792 7300
rect 6746 6962 6792 6974
rect 6840 6930 6880 7390
rect 6974 7350 7020 7362
rect 6974 7020 6980 7350
rect 7014 7020 7020 7350
rect 7070 7350 7116 7362
rect 7070 7250 7076 7350
rect 7110 7250 7116 7350
rect 7166 7350 7212 7362
rect 7050 7190 7060 7250
rect 7120 7190 7130 7250
rect 6960 6960 6970 7020
rect 7030 6960 7040 7020
rect 7070 6974 7076 7190
rect 7110 6974 7116 7190
rect 7166 7020 7172 7350
rect 7206 7020 7212 7350
rect 7262 7350 7308 7362
rect 7262 7250 7268 7350
rect 7302 7250 7308 7350
rect 7358 7350 7404 7362
rect 7250 7190 7260 7250
rect 7320 7190 7330 7250
rect 7070 6962 7116 6974
rect 7150 6960 7160 7020
rect 7220 6960 7230 7020
rect 7262 6974 7268 7190
rect 7302 6974 7308 7190
rect 7358 7020 7364 7350
rect 7398 7020 7404 7350
rect 7262 6962 7308 6974
rect 7340 6960 7350 7020
rect 7410 6960 7420 7020
rect 4550 6830 4560 6890
rect 4620 6830 4630 6890
rect 5035 6924 6145 6930
rect 5035 6890 5054 6924
rect 5088 6890 5246 6924
rect 5280 6890 5666 6924
rect 5700 6890 5858 6924
rect 5892 6890 6145 6924
rect 5035 6880 6145 6890
rect 6400 6924 7270 6930
rect 6400 6890 6416 6924
rect 6450 6890 6608 6924
rect 6642 6890 7028 6924
rect 7062 6890 7220 6924
rect 7254 6890 7270 6924
rect 6400 6880 7270 6890
rect -3490 6720 160 6800
rect 2400 6720 4480 6800
rect 5480 6720 5550 6880
rect 7490 6800 7530 9770
rect 6260 6750 7530 6800
rect 7570 6750 7620 9820
rect 6260 6720 7620 6750
rect -3490 6690 7620 6720
rect -3490 6630 -3400 6690
rect 7480 6630 7620 6690
rect -3490 6580 7620 6630
<< via1 >>
rect -3590 8690 -3530 8750
rect 40 9688 110 9710
rect 40 9654 60 9688
rect 60 9654 110 9688
rect 40 9640 110 9654
rect -3460 9340 -3400 9400
rect -3460 8840 -3400 8900
rect -3460 8230 -3400 8290
rect -3010 9340 -2994 9400
rect -2994 9340 -2960 9400
rect -2960 9340 -2950 9400
rect -3014 8842 -2994 8902
rect -2994 8842 -2960 8902
rect -2960 8842 -2954 8902
rect -2740 9340 -2722 9400
rect -2722 9340 -2688 9400
rect -2688 9340 -2680 9400
rect -2744 8842 -2722 8902
rect -2722 8842 -2688 8902
rect -2688 8842 -2684 8902
rect -2854 8692 -2836 8752
rect -2836 8692 -2802 8752
rect -2802 8692 -2794 8752
rect -3014 8232 -2994 8292
rect -2994 8232 -2960 8292
rect -2960 8232 -2954 8292
rect -2460 9340 -2450 9400
rect -2450 9340 -2416 9400
rect -2416 9340 -2400 9400
rect -2464 8842 -2450 8902
rect -2450 8842 -2416 8902
rect -2416 8842 -2404 8902
rect -2584 8692 -2564 8752
rect -2564 8692 -2530 8752
rect -2530 8692 -2524 8752
rect -2744 8232 -2722 8292
rect -2722 8232 -2688 8292
rect -2688 8232 -2684 8292
rect -2190 9340 -2178 9400
rect -2178 9340 -2144 9400
rect -2144 9340 -2130 9400
rect -2194 8842 -2178 8902
rect -2178 8842 -2144 8902
rect -2144 8842 -2134 8902
rect -2304 8522 -2292 8582
rect -2292 8522 -2258 8582
rect -2258 8522 -2244 8582
rect -2464 8232 -2450 8292
rect -2450 8232 -2416 8292
rect -2416 8232 -2404 8292
rect -1920 9340 -1906 9400
rect -1906 9340 -1872 9400
rect -1872 9340 -1860 9400
rect -1924 8842 -1906 8902
rect -1906 8842 -1872 8902
rect -1872 8842 -1864 8902
rect -2034 8522 -2020 8582
rect -2020 8522 -1986 8582
rect -1986 8522 -1974 8582
rect -2194 8232 -2178 8292
rect -2178 8232 -2144 8292
rect -2144 8232 -2134 8292
rect -2308 8074 -2292 8134
rect -2292 8074 -2258 8134
rect -2258 8074 -2248 8134
rect -1650 9340 -1634 9400
rect -1634 9340 -1600 9400
rect -1600 9340 -1590 9400
rect -1654 8842 -1634 8902
rect -1634 8842 -1600 8902
rect -1600 8842 -1594 8902
rect -1764 8522 -1748 8582
rect -1748 8522 -1714 8582
rect -1714 8522 -1704 8582
rect -1924 8232 -1906 8292
rect -1906 8232 -1872 8292
rect -1872 8232 -1864 8292
rect -2038 8074 -2020 8134
rect -2020 8074 -1986 8134
rect -1986 8074 -1978 8134
rect -1654 8232 -1634 8292
rect -1634 8232 -1600 8292
rect -1600 8232 -1594 8292
rect -1768 8074 -1748 8134
rect -1748 8074 -1714 8134
rect -1714 8074 -1708 8134
rect -1380 9340 -1362 9400
rect -1362 9340 -1328 9400
rect -1328 9340 -1320 9400
rect -1384 8842 -1362 8902
rect -1362 8842 -1328 8902
rect -1328 8842 -1324 8902
rect -1100 9340 -1090 9400
rect -1090 9340 -1056 9400
rect -1056 9340 -1040 9400
rect -1104 8842 -1090 8902
rect -1090 8842 -1056 8902
rect -1056 8842 -1044 8902
rect -1224 8522 -1204 8582
rect -1204 8522 -1170 8582
rect -1170 8522 -1164 8582
rect -1384 8232 -1362 8292
rect -1362 8232 -1328 8292
rect -1328 8232 -1324 8292
rect -830 9340 -818 9400
rect -818 9340 -784 9400
rect -784 9340 -770 9400
rect -834 8842 -818 8902
rect -818 8842 -784 8902
rect -784 8842 -774 8902
rect -944 8522 -932 8582
rect -932 8522 -898 8582
rect -898 8522 -884 8582
rect -1104 8232 -1090 8292
rect -1090 8232 -1056 8292
rect -1056 8232 -1044 8292
rect -1228 8074 -1204 8134
rect -1204 8074 -1170 8134
rect -1170 8074 -1168 8134
rect -560 9340 -546 9400
rect -546 9340 -512 9400
rect -512 9340 -500 9400
rect -564 8842 -546 8902
rect -546 8842 -512 8902
rect -512 8842 -504 8902
rect -674 8522 -660 8582
rect -660 8522 -626 8582
rect -626 8522 -614 8582
rect -834 8232 -818 8292
rect -818 8232 -784 8292
rect -784 8232 -774 8292
rect -948 8074 -932 8134
rect -932 8074 -898 8134
rect -898 8074 -888 8134
rect -290 9340 -274 9400
rect -274 9340 -240 9400
rect -240 9340 -230 9400
rect -294 8842 -274 8902
rect -274 8842 -240 8902
rect -240 8842 -234 8902
rect -404 8402 -388 8462
rect -388 8402 -354 8462
rect -354 8402 -344 8462
rect -564 8232 -546 8292
rect -546 8232 -512 8292
rect -512 8232 -504 8292
rect -678 8074 -660 8134
rect -660 8074 -626 8134
rect -626 8074 -618 8134
rect -130 8690 -116 8750
rect -116 8690 -82 8750
rect -82 8690 -70 8750
rect -294 8232 -274 8292
rect -274 8232 -240 8292
rect -240 8232 -234 8292
rect 270 9190 330 9250
rect 470 8710 480 8770
rect 480 8710 514 8770
rect 514 8710 530 8770
rect 370 8530 382 8590
rect 382 8530 416 8590
rect 416 8530 430 8590
rect 660 8710 676 8770
rect 676 8710 710 8770
rect 710 8710 720 8770
rect 560 8530 578 8590
rect 578 8530 612 8590
rect 612 8530 620 8590
rect 860 8710 872 8770
rect 872 8710 906 8770
rect 906 8710 920 8770
rect 760 8530 774 8590
rect 774 8530 808 8590
rect 808 8530 820 8590
rect 1060 8710 1068 8770
rect 1068 8710 1102 8770
rect 1102 8710 1120 8770
rect 960 8530 970 8590
rect 970 8530 1004 8590
rect 1004 8530 1020 8590
rect 2400 9650 2460 9710
rect 1290 9070 1350 9130
rect 1150 8530 1166 8590
rect 1166 8530 1200 8590
rect 1200 8530 1210 8590
rect 1100 8360 1160 8370
rect 1100 8326 1117 8360
rect 1117 8326 1151 8360
rect 1151 8326 1160 8360
rect 1100 8310 1160 8326
rect 1480 8900 1492 8960
rect 1492 8900 1526 8960
rect 1526 8900 1540 8960
rect 1380 8530 1394 8590
rect 1394 8530 1428 8590
rect 1428 8530 1440 8590
rect 1670 8900 1688 8960
rect 1688 8900 1722 8960
rect 1722 8900 1730 8960
rect 1580 8530 1590 8590
rect 1590 8530 1624 8590
rect 1624 8530 1640 8590
rect 1870 8900 1884 8960
rect 1884 8900 1918 8960
rect 1918 8900 1930 8960
rect 1780 8530 1786 8590
rect 1786 8530 1820 8590
rect 1820 8530 1840 8590
rect 2070 8900 2080 8960
rect 2080 8900 2114 8960
rect 2114 8900 2130 8960
rect 1970 8530 1982 8590
rect 1982 8530 2016 8590
rect 2016 8530 2030 8590
rect 2980 9646 3050 9660
rect 2980 9608 3050 9646
rect 2980 9590 3050 9608
rect 2320 8900 2380 8960
rect 2260 8710 2320 8770
rect 2170 8530 2178 8590
rect 2178 8530 2212 8590
rect 2212 8530 2230 8590
rect -3590 7580 -3530 7640
rect -3320 7477 -3260 7480
rect -3320 7429 -3314 7477
rect -3314 7429 -3260 7477
rect -3320 7420 -3260 7429
rect -2730 7420 -2670 7480
rect -3040 7150 -2980 7210
rect -250 7700 -190 7760
rect -1700 7580 -1684 7640
rect -1684 7580 -1650 7640
rect -1650 7580 -1640 7640
rect -1440 7580 -1426 7640
rect -1426 7580 -1392 7640
rect -1392 7580 -1380 7640
rect -1830 7340 -1770 7400
rect -1570 7250 -1510 7310
rect -2010 7010 -1950 7070
rect -2730 6880 -2670 6940
rect -930 7260 -914 7320
rect -914 7260 -880 7320
rect -880 7260 -870 7320
rect -620 7350 -608 7410
rect -608 7350 -574 7410
rect -574 7350 -560 7410
rect -720 7260 -704 7320
rect -704 7260 -670 7320
rect -670 7260 -660 7320
rect -510 7260 -494 7320
rect -494 7260 -460 7320
rect -460 7260 -450 7320
rect -200 7350 -188 7410
rect -188 7350 -154 7410
rect -154 7350 -140 7410
rect -300 7260 -284 7320
rect -284 7260 -250 7320
rect -250 7260 -240 7320
rect -90 7260 -74 7320
rect -74 7260 -40 7320
rect -40 7260 -30 7320
rect 370 8070 382 8130
rect 382 8070 416 8130
rect 416 8070 430 8130
rect 570 8070 578 8130
rect 578 8070 612 8130
rect 612 8070 630 8130
rect 470 7540 480 7600
rect 480 7540 514 7600
rect 514 7540 530 7600
rect 760 8070 774 8130
rect 774 8070 808 8130
rect 808 8070 820 8130
rect 660 7540 676 7600
rect 676 7540 710 7600
rect 710 7540 720 7600
rect 960 8070 970 8130
rect 970 8070 1004 8130
rect 1004 8070 1020 8130
rect 860 7540 872 7600
rect 872 7540 906 7600
rect 906 7540 920 7600
rect 1150 8070 1166 8130
rect 1166 8070 1200 8130
rect 1200 8070 1210 8130
rect 1060 7540 1068 7600
rect 1068 7540 1102 7600
rect 1102 7540 1120 7600
rect 1380 8220 1440 8280
rect 1380 8070 1394 8130
rect 1394 8070 1428 8130
rect 1428 8070 1440 8130
rect 1580 8070 1590 8130
rect 1590 8070 1624 8130
rect 1624 8070 1640 8130
rect 1480 7940 1492 8000
rect 1492 7940 1526 8000
rect 1526 7940 1540 8000
rect 1780 8070 1786 8130
rect 1786 8070 1820 8130
rect 1820 8070 1840 8130
rect 1670 7940 1688 8000
rect 1688 7940 1722 8000
rect 1722 7940 1730 8000
rect 1970 8070 1982 8130
rect 1982 8070 2016 8130
rect 2016 8070 2030 8130
rect 1870 7940 1884 8000
rect 1884 7940 1918 8000
rect 1918 7940 1930 8000
rect 2170 8070 2178 8130
rect 2178 8070 2212 8130
rect 2212 8070 2230 8130
rect 2070 7940 2080 8000
rect 2080 7940 2114 8000
rect 2114 7940 2130 8000
rect 2260 7940 2320 8000
rect 2320 7540 2380 7600
rect 2590 9002 2650 9010
rect 2590 8950 2600 9002
rect 2600 8950 2634 9002
rect 2634 8950 2650 9002
rect 2490 8850 2512 8910
rect 2512 8850 2546 8910
rect 2546 8850 2550 8910
rect 3560 9320 3620 9380
rect 2840 8950 2900 9010
rect 2400 7150 2460 7210
rect 2590 7820 2600 7880
rect 2600 7820 2634 7880
rect 2634 7820 2650 7880
rect 2540 6924 2600 6930
rect 2540 6890 2556 6924
rect 2556 6890 2590 6924
rect 2590 6890 2600 6924
rect 2540 6870 2600 6890
rect 2760 8850 2820 8910
rect 2850 8400 2910 8460
rect 2840 8160 2900 8220
rect 2840 7940 2900 8000
rect 5030 9340 5090 9400
rect 4780 8160 4840 8220
rect 2970 7690 3030 7750
rect 2940 7110 3000 7170
rect 3710 7820 3770 7880
rect 3350 7720 3410 7780
rect 3260 7110 3320 7170
rect 3470 7650 3530 7710
rect 4670 7540 4730 7600
rect 4560 7430 4620 7490
rect 3600 7360 3660 7420
rect 4090 7414 4150 7430
rect 4090 7380 4104 7414
rect 4104 7380 4138 7414
rect 4138 7380 4150 7414
rect 4090 7370 4150 7380
rect 3600 7110 3660 7170
rect 3740 7130 3800 7190
rect 3950 7130 3960 7190
rect 3960 7130 3994 7190
rect 3994 7130 4010 7190
rect 4240 7240 4248 7300
rect 4248 7240 4282 7300
rect 4282 7240 4300 7300
rect 4140 7130 4152 7190
rect 4152 7130 4186 7190
rect 4186 7130 4200 7190
rect 4040 7010 4056 7070
rect 4056 7010 4090 7070
rect 4090 7010 4100 7070
rect 4560 7240 4620 7300
rect 4330 7130 4344 7190
rect 4344 7130 4378 7190
rect 4378 7130 4390 7190
rect 4560 7010 4620 7070
rect 3600 6870 3660 6930
rect 4190 6924 4250 6930
rect 4190 6890 4200 6924
rect 4200 6890 4234 6924
rect 4234 6890 4250 6924
rect 4190 6870 4250 6890
rect 6680 8400 6740 8460
rect 6220 7630 6280 7690
rect 4780 7320 4840 7380
rect 5090 7070 5102 7130
rect 5102 7070 5136 7130
rect 5136 7070 5150 7130
rect 4670 6960 4730 7020
rect 4990 6983 5006 7020
rect 5006 6983 5040 7020
rect 5040 6983 5050 7020
rect 4990 6960 5050 6983
rect 5280 7070 5294 7130
rect 5294 7070 5328 7130
rect 5328 7070 5340 7130
rect 5180 6983 5198 7020
rect 5198 6983 5232 7020
rect 5232 6983 5240 7020
rect 5180 6960 5240 6983
rect 5610 7359 5670 7380
rect 5610 7320 5618 7359
rect 5618 7320 5652 7359
rect 5652 7320 5670 7359
rect 5380 6983 5390 7020
rect 5390 6983 5424 7020
rect 5424 6983 5440 7020
rect 5380 6960 5440 6983
rect 5800 7359 5860 7380
rect 5800 7320 5810 7359
rect 5810 7320 5844 7359
rect 5844 7320 5860 7359
rect 5700 7190 5714 7250
rect 5714 7190 5748 7250
rect 5748 7190 5760 7250
rect 5990 7359 6050 7380
rect 5990 7320 6002 7359
rect 6002 7320 6036 7359
rect 6036 7320 6050 7359
rect 5890 7190 5906 7250
rect 5906 7190 5940 7250
rect 5940 7190 5950 7250
rect 7390 7730 7450 7790
rect 6350 7350 6410 7360
rect 6350 7300 6368 7350
rect 6368 7300 6402 7350
rect 6402 7300 6410 7350
rect 6220 7070 6280 7130
rect 6550 7350 6610 7360
rect 6550 7300 6560 7350
rect 6560 7300 6594 7350
rect 6594 7300 6610 7350
rect 6450 7070 6464 7130
rect 6464 7070 6498 7130
rect 6498 7070 6510 7130
rect 6740 7350 6800 7360
rect 6740 7300 6752 7350
rect 6752 7300 6786 7350
rect 6786 7300 6800 7350
rect 6640 7070 6656 7130
rect 6656 7070 6690 7130
rect 6690 7070 6700 7130
rect 7060 7190 7076 7250
rect 7076 7190 7110 7250
rect 7110 7190 7120 7250
rect 6970 6974 6980 7020
rect 6980 6974 7014 7020
rect 7014 6974 7030 7020
rect 6970 6960 7030 6974
rect 7260 7190 7268 7250
rect 7268 7190 7302 7250
rect 7302 7190 7320 7250
rect 7160 6974 7172 7020
rect 7172 6974 7206 7020
rect 7206 6974 7220 7020
rect 7160 6960 7220 6974
rect 7350 6974 7364 7020
rect 7364 6974 7398 7020
rect 7398 6974 7410 7020
rect 7350 6960 7410 6974
rect 4560 6830 4620 6890
<< metal2 >>
rect 40 9710 110 9720
rect 2400 9710 2460 9720
rect 110 9650 2400 9710
rect 2460 9660 3050 9710
rect 2460 9650 2980 9660
rect 2400 9640 2460 9650
rect 40 9630 110 9640
rect 2980 9580 3050 9590
rect -3480 9400 5120 9420
rect -3480 9340 -3460 9400
rect -3400 9340 -3010 9400
rect -2950 9340 -2740 9400
rect -2680 9340 -2460 9400
rect -2400 9340 -2190 9400
rect -2130 9340 -1920 9400
rect -1860 9340 -1650 9400
rect -1590 9340 -1380 9400
rect -1320 9340 -1100 9400
rect -1040 9340 -830 9400
rect -770 9340 -560 9400
rect -500 9340 -290 9400
rect -230 9380 5030 9400
rect -230 9340 3560 9380
rect -3480 9320 3560 9340
rect 3620 9340 5030 9380
rect 5090 9340 5120 9400
rect 3620 9320 5120 9340
rect 3560 9310 3620 9320
rect 270 9250 330 9260
rect -3630 9200 270 9240
rect 270 9180 330 9190
rect 1290 9130 1350 9140
rect -3630 9080 1290 9120
rect 1290 9060 1350 9070
rect 2590 9010 2650 9020
rect 1470 8960 2390 8970
rect -3480 8902 -210 8920
rect -3480 8900 -3014 8902
rect -3480 8840 -3460 8900
rect -3400 8842 -3014 8900
rect -2954 8842 -2744 8902
rect -2684 8842 -2464 8902
rect -2404 8842 -2194 8902
rect -2134 8842 -1924 8902
rect -1864 8842 -1654 8902
rect -1594 8842 -1384 8902
rect -1324 8842 -1104 8902
rect -1044 8842 -834 8902
rect -774 8842 -564 8902
rect -504 8842 -294 8902
rect -234 8842 -210 8902
rect 1470 8900 1480 8960
rect 1540 8900 1670 8960
rect 1730 8900 1870 8960
rect 1930 8900 2070 8960
rect 2130 8900 2320 8960
rect 2380 8900 2390 8960
rect 2840 9010 2900 9020
rect 2650 8960 2840 8990
rect 2590 8940 2650 8950
rect 2840 8940 2900 8950
rect 1470 8890 2390 8900
rect 2490 8910 2550 8920
rect -3400 8840 -210 8842
rect 2760 8910 2820 8920
rect 2550 8860 2760 8890
rect 2490 8840 2550 8850
rect 2760 8840 2820 8850
rect -3480 8820 -210 8840
rect 460 8770 2320 8780
rect -3590 8750 -3530 8760
rect -2854 8752 -2794 8762
rect -3530 8692 -2854 8750
rect -2584 8752 -2524 8762
rect -2794 8692 -2584 8750
rect -130 8750 -70 8760
rect -2524 8692 -130 8750
rect -3530 8690 -130 8692
rect 460 8710 470 8770
rect 530 8710 660 8770
rect 720 8710 860 8770
rect 920 8710 1060 8770
rect 1120 8710 2260 8770
rect 460 8700 2320 8710
rect -3590 8680 -3530 8690
rect -2854 8682 -2794 8690
rect -2584 8682 -2524 8690
rect -130 8680 -70 8690
rect -2330 8590 2235 8610
rect -2330 8582 370 8590
rect -2330 8522 -2304 8582
rect -2244 8522 -2034 8582
rect -1974 8522 -1764 8582
rect -1704 8522 -1224 8582
rect -1164 8522 -944 8582
rect -884 8522 -674 8582
rect -614 8530 370 8582
rect 430 8530 560 8590
rect 620 8530 760 8590
rect 820 8530 960 8590
rect 1020 8530 1150 8590
rect 1210 8530 1380 8590
rect 1440 8530 1580 8590
rect 1640 8530 1780 8590
rect 1840 8530 1970 8590
rect 2030 8530 2170 8590
rect 2230 8530 2235 8590
rect -614 8522 2235 8530
rect -2330 8500 2235 8522
rect -404 8462 -344 8472
rect 2850 8460 2910 8470
rect -344 8410 2850 8450
rect -404 8392 -344 8402
rect 6680 8460 6740 8470
rect 2910 8410 6680 8450
rect 2850 8390 2910 8400
rect 6680 8390 6740 8400
rect 1100 8370 1160 8380
rect 1160 8320 1430 8360
rect -3480 8292 -210 8310
rect 1100 8300 1160 8310
rect -3480 8290 -3014 8292
rect -3480 8230 -3460 8290
rect -3400 8232 -3014 8290
rect -2954 8232 -2744 8292
rect -2684 8232 -2464 8292
rect -2404 8232 -2194 8292
rect -2134 8232 -1924 8292
rect -1864 8232 -1654 8292
rect -1594 8232 -1384 8292
rect -1324 8232 -1104 8292
rect -1044 8232 -834 8292
rect -774 8232 -564 8292
rect -504 8232 -294 8292
rect -234 8232 -210 8292
rect 1390 8290 1430 8320
rect -3400 8230 -210 8232
rect -3480 8210 -210 8230
rect 1380 8280 1440 8290
rect 1380 8210 1440 8220
rect 2840 8220 4840 8230
rect -2334 8134 2235 8162
rect 2900 8160 4780 8220
rect 2840 8150 4840 8160
rect -2334 8074 -2308 8134
rect -2248 8074 -2038 8134
rect -1978 8074 -1768 8134
rect -1708 8074 -1228 8134
rect -1168 8074 -948 8134
rect -888 8074 -678 8134
rect -618 8130 2235 8134
rect -618 8074 370 8130
rect -2334 8070 370 8074
rect 430 8070 570 8130
rect 630 8070 760 8130
rect 820 8070 960 8130
rect 1020 8070 1150 8130
rect 1210 8070 1380 8130
rect 1440 8070 1580 8130
rect 1640 8070 1780 8130
rect 1840 8070 1970 8130
rect 2030 8070 2170 8130
rect 2230 8070 2235 8130
rect -2334 8052 2235 8070
rect 1470 8000 2900 8010
rect 1470 7940 1480 8000
rect 1540 7940 1670 8000
rect 1730 7940 1870 8000
rect 1930 7940 2070 8000
rect 2130 7940 2260 8000
rect 2320 7940 2840 8000
rect 1470 7930 2900 7940
rect 2590 7880 2650 7890
rect 3710 7880 3770 7890
rect 2650 7830 3710 7870
rect 2590 7810 2650 7820
rect 3710 7810 3770 7820
rect 7390 7790 7450 7800
rect -250 7760 -190 7770
rect 2970 7750 3030 7760
rect -190 7710 2970 7740
rect -250 7690 -190 7700
rect 3340 7720 3350 7780
rect 3410 7740 7390 7780
rect 3410 7720 3420 7740
rect 2970 7680 3030 7690
rect 3460 7650 3470 7710
rect 3530 7700 3540 7710
rect 3530 7690 6280 7700
rect 3530 7660 6220 7690
rect 3530 7650 3540 7660
rect -3590 7640 -3530 7650
rect -1700 7640 -1640 7650
rect -3530 7590 -1700 7620
rect -3590 7570 -3530 7580
rect -1700 7570 -1640 7580
rect -1440 7640 -1380 7650
rect 6220 7620 6280 7630
rect -1440 7570 -1380 7580
rect 460 7600 4740 7610
rect -1425 7500 -1395 7570
rect 460 7540 470 7600
rect 530 7540 660 7600
rect 720 7540 860 7600
rect 920 7540 1060 7600
rect 1120 7540 2320 7600
rect 2380 7540 4670 7600
rect 4730 7540 4740 7600
rect 460 7530 4740 7540
rect -1425 7490 6210 7500
rect -3320 7480 -3260 7490
rect -3630 7430 -3320 7470
rect -2730 7480 -2670 7490
rect -3260 7430 -2730 7470
rect -3320 7410 -3260 7420
rect -1425 7470 4560 7490
rect 4090 7430 4150 7440
rect 3600 7420 3660 7430
rect -2730 7410 -2670 7420
rect -620 7410 -560 7420
rect -1830 7400 -1770 7410
rect -3630 7350 -1830 7380
rect -200 7410 -140 7420
rect -560 7360 -200 7400
rect -620 7340 -560 7350
rect -140 7360 3600 7400
rect 3660 7380 4090 7410
rect 4550 7430 4560 7470
rect 4620 7430 6210 7490
rect 4550 7420 6210 7430
rect 4090 7360 4150 7370
rect 4780 7380 6050 7390
rect 3600 7350 3660 7360
rect -200 7340 -140 7350
rect -1830 7330 -1770 7340
rect -930 7320 -870 7330
rect -1570 7310 -1510 7320
rect -3630 7260 -1570 7290
rect -720 7320 -660 7330
rect -870 7270 -720 7310
rect -930 7250 -870 7260
rect -510 7320 -450 7330
rect -660 7270 -510 7310
rect -720 7250 -660 7260
rect -300 7320 -240 7330
rect -450 7270 -300 7310
rect -510 7250 -450 7260
rect -90 7320 -30 7330
rect -240 7270 -90 7310
rect -300 7250 -240 7260
rect 4840 7320 5610 7380
rect 5670 7320 5800 7380
rect 5860 7320 5990 7380
rect 4780 7310 6050 7320
rect 6130 7370 6210 7420
rect 6130 7360 6800 7370
rect -90 7250 -30 7260
rect 4240 7300 4620 7310
rect -1570 7240 -1510 7250
rect 4300 7240 4560 7300
rect 6130 7300 6350 7360
rect 6410 7300 6550 7360
rect 6610 7300 6740 7360
rect 6130 7290 6800 7300
rect 6860 7260 6900 7740
rect 7390 7720 7450 7730
rect 4240 7230 4620 7240
rect 5700 7250 7330 7260
rect -3040 7210 -2980 7220
rect 2400 7210 2460 7220
rect -2980 7160 2400 7190
rect -3040 7140 -2980 7150
rect 3740 7190 4390 7200
rect 2400 7140 2460 7150
rect 2940 7170 3000 7180
rect 3260 7170 3320 7180
rect 3000 7120 3260 7150
rect 2940 7100 3000 7110
rect 3600 7170 3660 7180
rect 3320 7120 3600 7150
rect 3260 7100 3320 7110
rect 3800 7130 3950 7190
rect 4010 7130 4140 7190
rect 4200 7130 4330 7190
rect 5760 7190 5890 7250
rect 5950 7190 7060 7250
rect 7120 7190 7260 7250
rect 7320 7230 7330 7250
rect 7320 7200 7680 7230
rect 7320 7190 7330 7200
rect 5700 7180 7330 7190
rect 3740 7120 4390 7130
rect 5090 7130 6710 7140
rect 3600 7100 3660 7110
rect -2010 7070 -1950 7080
rect -2015 7020 -2010 7050
rect 4040 7070 4620 7080
rect -1950 7020 4040 7050
rect -2010 7000 -1950 7010
rect 4100 7010 4560 7070
rect 5150 7070 5280 7130
rect 5340 7070 6220 7130
rect 6280 7070 6450 7130
rect 6510 7070 6640 7130
rect 6700 7120 6710 7130
rect 6700 7090 7680 7120
rect 6700 7070 6710 7090
rect 5090 7060 6710 7070
rect 4040 7000 4620 7010
rect 4670 7020 5440 7030
rect 4730 6960 4990 7020
rect 5050 6960 5180 7020
rect 5240 6960 5380 7020
rect 4670 6950 5440 6960
rect 5520 7020 7420 7030
rect 5520 6960 6970 7020
rect 7030 6960 7160 7020
rect 7220 6960 7350 7020
rect 7410 6960 7420 7020
rect 5520 6950 7420 6960
rect -2730 6940 -2670 6950
rect 2540 6930 2600 6940
rect -2670 6890 2540 6930
rect -2730 6870 -2670 6880
rect 2540 6860 2600 6870
rect 3600 6930 3660 6940
rect 4190 6930 4250 6940
rect 3660 6880 4190 6910
rect 3600 6860 3660 6870
rect 5520 6900 5600 6950
rect 4190 6860 4250 6870
rect 4550 6890 5600 6900
rect 4550 6830 4560 6890
rect 4620 6830 5600 6890
rect 4550 6820 5600 6830
<< labels >>
rlabel metal2 -3630 9200 -3590 9240 1 IN_P
port 1 n
rlabel metal2 -3630 9080 -3590 9120 1 IN_N
port 2 n
rlabel metal2 7650 7200 7680 7230 1 OUT_N
port 3 n
rlabel metal2 7650 7090 7680 7120 1 OUT_P
port 4 n
rlabel metal2 -3630 7430 -3590 7470 1 EN
port 5 n
rlabel metal2 -3630 7350 -3600 7380 1 CAL_P
port 6 n
rlabel metal2 -3630 7260 -3600 7290 1 CAL_N
port 7 n
rlabel metal1 -3430 6730 -3190 6870 1 VSS
port 8 n
rlabel metal1 -3460 9780 -3220 9920 1 VDD
port 9 n
<< end >>
