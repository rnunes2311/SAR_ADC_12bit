magic
tech sky130A
magscale 1 2
timestamp 1711796880
<< error_p >>
rect -1951 881 -1889 887
rect -1823 881 -1761 887
rect -1695 881 -1633 887
rect -1567 881 -1505 887
rect -1439 881 -1377 887
rect -1311 881 -1249 887
rect -1183 881 -1121 887
rect -1055 881 -993 887
rect -927 881 -865 887
rect -799 881 -737 887
rect -671 881 -609 887
rect -543 881 -481 887
rect -415 881 -353 887
rect -287 881 -225 887
rect -159 881 -97 887
rect -31 881 31 887
rect 97 881 159 887
rect 225 881 287 887
rect 353 881 415 887
rect 481 881 543 887
rect 609 881 671 887
rect 737 881 799 887
rect 865 881 927 887
rect 993 881 1055 887
rect 1121 881 1183 887
rect 1249 881 1311 887
rect 1377 881 1439 887
rect 1505 881 1567 887
rect 1633 881 1695 887
rect 1761 881 1823 887
rect 1889 881 1951 887
rect -1951 847 -1939 881
rect -1823 847 -1811 881
rect -1695 847 -1683 881
rect -1567 847 -1555 881
rect -1439 847 -1427 881
rect -1311 847 -1299 881
rect -1183 847 -1171 881
rect -1055 847 -1043 881
rect -927 847 -915 881
rect -799 847 -787 881
rect -671 847 -659 881
rect -543 847 -531 881
rect -415 847 -403 881
rect -287 847 -275 881
rect -159 847 -147 881
rect -31 847 -19 881
rect 97 847 109 881
rect 225 847 237 881
rect 353 847 365 881
rect 481 847 493 881
rect 609 847 621 881
rect 737 847 749 881
rect 865 847 877 881
rect 993 847 1005 881
rect 1121 847 1133 881
rect 1249 847 1261 881
rect 1377 847 1389 881
rect 1505 847 1517 881
rect 1633 847 1645 881
rect 1761 847 1773 881
rect 1889 847 1901 881
rect -1951 841 -1889 847
rect -1823 841 -1761 847
rect -1695 841 -1633 847
rect -1567 841 -1505 847
rect -1439 841 -1377 847
rect -1311 841 -1249 847
rect -1183 841 -1121 847
rect -1055 841 -993 847
rect -927 841 -865 847
rect -799 841 -737 847
rect -671 841 -609 847
rect -543 841 -481 847
rect -415 841 -353 847
rect -287 841 -225 847
rect -159 841 -97 847
rect -31 841 31 847
rect 97 841 159 847
rect 225 841 287 847
rect 353 841 415 847
rect 481 841 543 847
rect 609 841 671 847
rect 737 841 799 847
rect 865 841 927 847
rect 993 841 1055 847
rect 1121 841 1183 847
rect 1249 841 1311 847
rect 1377 841 1439 847
rect 1505 841 1567 847
rect 1633 841 1695 847
rect 1761 841 1823 847
rect 1889 841 1951 847
rect -1951 -847 -1889 -841
rect -1823 -847 -1761 -841
rect -1695 -847 -1633 -841
rect -1567 -847 -1505 -841
rect -1439 -847 -1377 -841
rect -1311 -847 -1249 -841
rect -1183 -847 -1121 -841
rect -1055 -847 -993 -841
rect -927 -847 -865 -841
rect -799 -847 -737 -841
rect -671 -847 -609 -841
rect -543 -847 -481 -841
rect -415 -847 -353 -841
rect -287 -847 -225 -841
rect -159 -847 -97 -841
rect -31 -847 31 -841
rect 97 -847 159 -841
rect 225 -847 287 -841
rect 353 -847 415 -841
rect 481 -847 543 -841
rect 609 -847 671 -841
rect 737 -847 799 -841
rect 865 -847 927 -841
rect 993 -847 1055 -841
rect 1121 -847 1183 -841
rect 1249 -847 1311 -841
rect 1377 -847 1439 -841
rect 1505 -847 1567 -841
rect 1633 -847 1695 -841
rect 1761 -847 1823 -841
rect 1889 -847 1951 -841
rect -1951 -881 -1939 -847
rect -1823 -881 -1811 -847
rect -1695 -881 -1683 -847
rect -1567 -881 -1555 -847
rect -1439 -881 -1427 -847
rect -1311 -881 -1299 -847
rect -1183 -881 -1171 -847
rect -1055 -881 -1043 -847
rect -927 -881 -915 -847
rect -799 -881 -787 -847
rect -671 -881 -659 -847
rect -543 -881 -531 -847
rect -415 -881 -403 -847
rect -287 -881 -275 -847
rect -159 -881 -147 -847
rect -31 -881 -19 -847
rect 97 -881 109 -847
rect 225 -881 237 -847
rect 353 -881 365 -847
rect 481 -881 493 -847
rect 609 -881 621 -847
rect 737 -881 749 -847
rect 865 -881 877 -847
rect 993 -881 1005 -847
rect 1121 -881 1133 -847
rect 1249 -881 1261 -847
rect 1377 -881 1389 -847
rect 1505 -881 1517 -847
rect 1633 -881 1645 -847
rect 1761 -881 1773 -847
rect 1889 -881 1901 -847
rect -1951 -887 -1889 -881
rect -1823 -887 -1761 -881
rect -1695 -887 -1633 -881
rect -1567 -887 -1505 -881
rect -1439 -887 -1377 -881
rect -1311 -887 -1249 -881
rect -1183 -887 -1121 -881
rect -1055 -887 -993 -881
rect -927 -887 -865 -881
rect -799 -887 -737 -881
rect -671 -887 -609 -881
rect -543 -887 -481 -881
rect -415 -887 -353 -881
rect -287 -887 -225 -881
rect -159 -887 -97 -881
rect -31 -887 31 -881
rect 97 -887 159 -881
rect 225 -887 287 -881
rect 353 -887 415 -881
rect 481 -887 543 -881
rect 609 -887 671 -881
rect 737 -887 799 -881
rect 865 -887 927 -881
rect 993 -887 1055 -881
rect 1121 -887 1183 -881
rect 1249 -887 1311 -881
rect 1377 -887 1439 -881
rect 1505 -887 1567 -881
rect 1633 -887 1695 -881
rect 1761 -887 1823 -881
rect 1889 -887 1951 -881
<< nwell >>
rect -2151 -1019 3191 1019
<< pmoslvt >>
rect -1955 -800 -1885 800
rect -1827 -800 -1757 800
rect -1699 -800 -1629 800
rect -1571 -800 -1501 800
rect -1443 -800 -1373 800
rect -1315 -800 -1245 800
rect -1187 -800 -1117 800
rect -1059 -800 -989 800
rect -931 -800 -861 800
rect -803 -800 -733 800
rect -675 -800 -605 800
rect -547 -800 -477 800
rect -419 -800 -349 800
rect -291 -800 -221 800
rect -163 -800 -93 800
rect -35 -800 35 800
rect 93 -800 163 800
rect 221 -800 291 800
rect 349 -800 419 800
rect 477 -800 547 800
rect 605 -800 675 800
rect 733 -800 803 800
rect 861 -800 931 800
rect 989 -800 1059 800
rect 1117 -800 1187 800
rect 1245 -800 1315 800
rect 1373 -800 1443 800
rect 1501 -800 1571 800
rect 1629 -800 1699 800
rect 1757 -800 1827 800
rect 1885 -800 1955 800
<< pdiff >>
rect -2013 788 -1955 800
rect -2013 -788 -2001 788
rect -1967 -788 -1955 788
rect -2013 -800 -1955 -788
rect -1885 788 -1827 800
rect -1885 -788 -1873 788
rect -1839 -788 -1827 788
rect -1885 -800 -1827 -788
rect -1757 788 -1699 800
rect -1757 -788 -1745 788
rect -1711 -788 -1699 788
rect -1757 -800 -1699 -788
rect -1629 788 -1571 800
rect -1629 -788 -1617 788
rect -1583 -788 -1571 788
rect -1629 -800 -1571 -788
rect -1501 788 -1443 800
rect -1501 -788 -1489 788
rect -1455 -788 -1443 788
rect -1501 -800 -1443 -788
rect -1373 788 -1315 800
rect -1373 -788 -1361 788
rect -1327 -788 -1315 788
rect -1373 -800 -1315 -788
rect -1245 788 -1187 800
rect -1245 -788 -1233 788
rect -1199 -788 -1187 788
rect -1245 -800 -1187 -788
rect -1117 788 -1059 800
rect -1117 -788 -1105 788
rect -1071 -788 -1059 788
rect -1117 -800 -1059 -788
rect -989 788 -931 800
rect -989 -788 -977 788
rect -943 -788 -931 788
rect -989 -800 -931 -788
rect -861 788 -803 800
rect -861 -788 -849 788
rect -815 -788 -803 788
rect -861 -800 -803 -788
rect -733 788 -675 800
rect -733 -788 -721 788
rect -687 -788 -675 788
rect -733 -800 -675 -788
rect -605 788 -547 800
rect -605 -788 -593 788
rect -559 -788 -547 788
rect -605 -800 -547 -788
rect -477 788 -419 800
rect -477 -788 -465 788
rect -431 -788 -419 788
rect -477 -800 -419 -788
rect -349 788 -291 800
rect -349 -788 -337 788
rect -303 -788 -291 788
rect -349 -800 -291 -788
rect -221 788 -163 800
rect -221 -788 -209 788
rect -175 -788 -163 788
rect -221 -800 -163 -788
rect -93 788 -35 800
rect -93 -788 -81 788
rect -47 -788 -35 788
rect -93 -800 -35 -788
rect 35 788 93 800
rect 35 -788 47 788
rect 81 -788 93 788
rect 35 -800 93 -788
rect 163 788 221 800
rect 163 -788 175 788
rect 209 -788 221 788
rect 163 -800 221 -788
rect 291 788 349 800
rect 291 -788 303 788
rect 337 -788 349 788
rect 291 -800 349 -788
rect 419 788 477 800
rect 419 -788 431 788
rect 465 -788 477 788
rect 419 -800 477 -788
rect 547 788 605 800
rect 547 -788 559 788
rect 593 -788 605 788
rect 547 -800 605 -788
rect 675 788 733 800
rect 675 -788 687 788
rect 721 -788 733 788
rect 675 -800 733 -788
rect 803 788 861 800
rect 803 -788 815 788
rect 849 -788 861 788
rect 803 -800 861 -788
rect 931 788 989 800
rect 931 -788 943 788
rect 977 -788 989 788
rect 931 -800 989 -788
rect 1059 788 1117 800
rect 1059 -788 1071 788
rect 1105 -788 1117 788
rect 1059 -800 1117 -788
rect 1187 788 1245 800
rect 1187 -788 1199 788
rect 1233 -788 1245 788
rect 1187 -800 1245 -788
rect 1315 788 1373 800
rect 1315 -788 1327 788
rect 1361 -788 1373 788
rect 1315 -800 1373 -788
rect 1443 788 1501 800
rect 1443 -788 1455 788
rect 1489 -788 1501 788
rect 1443 -800 1501 -788
rect 1571 788 1629 800
rect 1571 -788 1583 788
rect 1617 -788 1629 788
rect 1571 -800 1629 -788
rect 1699 788 1757 800
rect 1699 -788 1711 788
rect 1745 -788 1757 788
rect 1699 -800 1757 -788
rect 1827 788 1885 800
rect 1827 -788 1839 788
rect 1873 -788 1885 788
rect 1827 -800 1885 -788
rect 1955 788 2013 800
rect 1955 -788 1967 788
rect 2001 -788 2013 788
rect 1955 -800 2013 -788
<< pdiffc >>
rect -2001 -788 -1967 788
rect -1873 -788 -1839 788
rect -1745 -788 -1711 788
rect -1617 -788 -1583 788
rect -1489 -788 -1455 788
rect -1361 -788 -1327 788
rect -1233 -788 -1199 788
rect -1105 -788 -1071 788
rect -977 -788 -943 788
rect -849 -788 -815 788
rect -721 -788 -687 788
rect -593 -788 -559 788
rect -465 -788 -431 788
rect -337 -788 -303 788
rect -209 -788 -175 788
rect -81 -788 -47 788
rect 47 -788 81 788
rect 175 -788 209 788
rect 303 -788 337 788
rect 431 -788 465 788
rect 559 -788 593 788
rect 687 -788 721 788
rect 815 -788 849 788
rect 943 -788 977 788
rect 1071 -788 1105 788
rect 1199 -788 1233 788
rect 1327 -788 1361 788
rect 1455 -788 1489 788
rect 1583 -788 1617 788
rect 1711 -788 1745 788
rect 1839 -788 1873 788
rect 1967 -788 2001 788
<< nsubdiff >>
rect -2115 949 -2019 983
rect 2019 949 3155 983
rect -2115 887 -2081 949
rect 3121 887 3155 949
rect -2115 -949 -2081 -887
rect 3121 -949 3155 -887
rect -2115 -983 -2019 -949
rect 2019 -983 3155 -949
<< nsubdiffcont >>
rect -2019 949 2019 983
rect -2115 -887 -2081 887
rect 3121 -887 3155 887
rect -2019 -983 2019 -949
<< poly >>
rect -1955 881 -1885 897
rect -1955 847 -1939 881
rect -1901 847 -1885 881
rect -1955 800 -1885 847
rect -1827 881 -1757 897
rect -1827 847 -1811 881
rect -1773 847 -1757 881
rect -1827 800 -1757 847
rect -1699 881 -1629 897
rect -1699 847 -1683 881
rect -1645 847 -1629 881
rect -1699 800 -1629 847
rect -1571 881 -1501 897
rect -1571 847 -1555 881
rect -1517 847 -1501 881
rect -1571 800 -1501 847
rect -1443 881 -1373 897
rect -1443 847 -1427 881
rect -1389 847 -1373 881
rect -1443 800 -1373 847
rect -1315 881 -1245 897
rect -1315 847 -1299 881
rect -1261 847 -1245 881
rect -1315 800 -1245 847
rect -1187 881 -1117 897
rect -1187 847 -1171 881
rect -1133 847 -1117 881
rect -1187 800 -1117 847
rect -1059 881 -989 897
rect -1059 847 -1043 881
rect -1005 847 -989 881
rect -1059 800 -989 847
rect -931 881 -861 897
rect -931 847 -915 881
rect -877 847 -861 881
rect -931 800 -861 847
rect -803 881 -733 897
rect -803 847 -787 881
rect -749 847 -733 881
rect -803 800 -733 847
rect -675 881 -605 897
rect -675 847 -659 881
rect -621 847 -605 881
rect -675 800 -605 847
rect -547 881 -477 897
rect -547 847 -531 881
rect -493 847 -477 881
rect -547 800 -477 847
rect -419 881 -349 897
rect -419 847 -403 881
rect -365 847 -349 881
rect -419 800 -349 847
rect -291 881 -221 897
rect -291 847 -275 881
rect -237 847 -221 881
rect -291 800 -221 847
rect -163 881 -93 897
rect -163 847 -147 881
rect -109 847 -93 881
rect -163 800 -93 847
rect -35 881 35 897
rect -35 847 -19 881
rect 19 847 35 881
rect -35 800 35 847
rect 93 881 163 897
rect 93 847 109 881
rect 147 847 163 881
rect 93 800 163 847
rect 221 881 291 897
rect 221 847 237 881
rect 275 847 291 881
rect 221 800 291 847
rect 349 881 419 897
rect 349 847 365 881
rect 403 847 419 881
rect 349 800 419 847
rect 477 881 547 897
rect 477 847 493 881
rect 531 847 547 881
rect 477 800 547 847
rect 605 881 675 897
rect 605 847 621 881
rect 659 847 675 881
rect 605 800 675 847
rect 733 881 803 897
rect 733 847 749 881
rect 787 847 803 881
rect 733 800 803 847
rect 861 881 931 897
rect 861 847 877 881
rect 915 847 931 881
rect 861 800 931 847
rect 989 881 1059 897
rect 989 847 1005 881
rect 1043 847 1059 881
rect 989 800 1059 847
rect 1117 881 1187 897
rect 1117 847 1133 881
rect 1171 847 1187 881
rect 1117 800 1187 847
rect 1245 881 1315 897
rect 1245 847 1261 881
rect 1299 847 1315 881
rect 1245 800 1315 847
rect 1373 881 1443 897
rect 1373 847 1389 881
rect 1427 847 1443 881
rect 1373 800 1443 847
rect 1501 881 1571 897
rect 1501 847 1517 881
rect 1555 847 1571 881
rect 1501 800 1571 847
rect 1629 881 1699 897
rect 1629 847 1645 881
rect 1683 847 1699 881
rect 1629 800 1699 847
rect 1757 881 1827 897
rect 1757 847 1773 881
rect 1811 847 1827 881
rect 1757 800 1827 847
rect 1885 881 1955 897
rect 1885 847 1901 881
rect 1939 847 1955 881
rect 1885 800 1955 847
rect -1955 -847 -1885 -800
rect -1955 -881 -1939 -847
rect -1901 -881 -1885 -847
rect -1955 -897 -1885 -881
rect -1827 -847 -1757 -800
rect -1827 -881 -1811 -847
rect -1773 -881 -1757 -847
rect -1827 -897 -1757 -881
rect -1699 -847 -1629 -800
rect -1699 -881 -1683 -847
rect -1645 -881 -1629 -847
rect -1699 -897 -1629 -881
rect -1571 -847 -1501 -800
rect -1571 -881 -1555 -847
rect -1517 -881 -1501 -847
rect -1571 -897 -1501 -881
rect -1443 -847 -1373 -800
rect -1443 -881 -1427 -847
rect -1389 -881 -1373 -847
rect -1443 -897 -1373 -881
rect -1315 -847 -1245 -800
rect -1315 -881 -1299 -847
rect -1261 -881 -1245 -847
rect -1315 -897 -1245 -881
rect -1187 -847 -1117 -800
rect -1187 -881 -1171 -847
rect -1133 -881 -1117 -847
rect -1187 -897 -1117 -881
rect -1059 -847 -989 -800
rect -1059 -881 -1043 -847
rect -1005 -881 -989 -847
rect -1059 -897 -989 -881
rect -931 -847 -861 -800
rect -931 -881 -915 -847
rect -877 -881 -861 -847
rect -931 -897 -861 -881
rect -803 -847 -733 -800
rect -803 -881 -787 -847
rect -749 -881 -733 -847
rect -803 -897 -733 -881
rect -675 -847 -605 -800
rect -675 -881 -659 -847
rect -621 -881 -605 -847
rect -675 -897 -605 -881
rect -547 -847 -477 -800
rect -547 -881 -531 -847
rect -493 -881 -477 -847
rect -547 -897 -477 -881
rect -419 -847 -349 -800
rect -419 -881 -403 -847
rect -365 -881 -349 -847
rect -419 -897 -349 -881
rect -291 -847 -221 -800
rect -291 -881 -275 -847
rect -237 -881 -221 -847
rect -291 -897 -221 -881
rect -163 -847 -93 -800
rect -163 -881 -147 -847
rect -109 -881 -93 -847
rect -163 -897 -93 -881
rect -35 -847 35 -800
rect -35 -881 -19 -847
rect 19 -881 35 -847
rect -35 -897 35 -881
rect 93 -847 163 -800
rect 93 -881 109 -847
rect 147 -881 163 -847
rect 93 -897 163 -881
rect 221 -847 291 -800
rect 221 -881 237 -847
rect 275 -881 291 -847
rect 221 -897 291 -881
rect 349 -847 419 -800
rect 349 -881 365 -847
rect 403 -881 419 -847
rect 349 -897 419 -881
rect 477 -847 547 -800
rect 477 -881 493 -847
rect 531 -881 547 -847
rect 477 -897 547 -881
rect 605 -847 675 -800
rect 605 -881 621 -847
rect 659 -881 675 -847
rect 605 -897 675 -881
rect 733 -847 803 -800
rect 733 -881 749 -847
rect 787 -881 803 -847
rect 733 -897 803 -881
rect 861 -847 931 -800
rect 861 -881 877 -847
rect 915 -881 931 -847
rect 861 -897 931 -881
rect 989 -847 1059 -800
rect 989 -881 1005 -847
rect 1043 -881 1059 -847
rect 989 -897 1059 -881
rect 1117 -847 1187 -800
rect 1117 -881 1133 -847
rect 1171 -881 1187 -847
rect 1117 -897 1187 -881
rect 1245 -847 1315 -800
rect 1245 -881 1261 -847
rect 1299 -881 1315 -847
rect 1245 -897 1315 -881
rect 1373 -847 1443 -800
rect 1373 -881 1389 -847
rect 1427 -881 1443 -847
rect 1373 -897 1443 -881
rect 1501 -847 1571 -800
rect 1501 -881 1517 -847
rect 1555 -881 1571 -847
rect 1501 -897 1571 -881
rect 1629 -847 1699 -800
rect 1629 -881 1645 -847
rect 1683 -881 1699 -847
rect 1629 -897 1699 -881
rect 1757 -847 1827 -800
rect 1757 -881 1773 -847
rect 1811 -881 1827 -847
rect 1757 -897 1827 -881
rect 1885 -847 1955 -800
rect 1885 -881 1901 -847
rect 1939 -881 1955 -847
rect 1885 -897 1955 -881
<< polycont >>
rect -1939 847 -1901 881
rect -1811 847 -1773 881
rect -1683 847 -1645 881
rect -1555 847 -1517 881
rect -1427 847 -1389 881
rect -1299 847 -1261 881
rect -1171 847 -1133 881
rect -1043 847 -1005 881
rect -915 847 -877 881
rect -787 847 -749 881
rect -659 847 -621 881
rect -531 847 -493 881
rect -403 847 -365 881
rect -275 847 -237 881
rect -147 847 -109 881
rect -19 847 19 881
rect 109 847 147 881
rect 237 847 275 881
rect 365 847 403 881
rect 493 847 531 881
rect 621 847 659 881
rect 749 847 787 881
rect 877 847 915 881
rect 1005 847 1043 881
rect 1133 847 1171 881
rect 1261 847 1299 881
rect 1389 847 1427 881
rect 1517 847 1555 881
rect 1645 847 1683 881
rect 1773 847 1811 881
rect 1901 847 1939 881
rect -1939 -881 -1901 -847
rect -1811 -881 -1773 -847
rect -1683 -881 -1645 -847
rect -1555 -881 -1517 -847
rect -1427 -881 -1389 -847
rect -1299 -881 -1261 -847
rect -1171 -881 -1133 -847
rect -1043 -881 -1005 -847
rect -915 -881 -877 -847
rect -787 -881 -749 -847
rect -659 -881 -621 -847
rect -531 -881 -493 -847
rect -403 -881 -365 -847
rect -275 -881 -237 -847
rect -147 -881 -109 -847
rect -19 -881 19 -847
rect 109 -881 147 -847
rect 237 -881 275 -847
rect 365 -881 403 -847
rect 493 -881 531 -847
rect 621 -881 659 -847
rect 749 -881 787 -847
rect 877 -881 915 -847
rect 1005 -881 1043 -847
rect 1133 -881 1171 -847
rect 1261 -881 1299 -847
rect 1389 -881 1427 -847
rect 1517 -881 1555 -847
rect 1645 -881 1683 -847
rect 1773 -881 1811 -847
rect 1901 -881 1939 -847
<< locali >>
rect -2115 949 -2019 983
rect 2019 949 3155 983
rect -2115 887 -2081 949
rect 3121 887 3155 949
rect -1955 847 -1939 881
rect -1901 847 -1885 881
rect -1827 847 -1811 881
rect -1773 847 -1757 881
rect -1699 847 -1683 881
rect -1645 847 -1629 881
rect -1571 847 -1555 881
rect -1517 847 -1501 881
rect -1443 847 -1427 881
rect -1389 847 -1373 881
rect -1315 847 -1299 881
rect -1261 847 -1245 881
rect -1187 847 -1171 881
rect -1133 847 -1117 881
rect -1059 847 -1043 881
rect -1005 847 -989 881
rect -931 847 -915 881
rect -877 847 -861 881
rect -803 847 -787 881
rect -749 847 -733 881
rect -675 847 -659 881
rect -621 847 -605 881
rect -547 847 -531 881
rect -493 847 -477 881
rect -419 847 -403 881
rect -365 847 -349 881
rect -291 847 -275 881
rect -237 847 -221 881
rect -163 847 -147 881
rect -109 847 -93 881
rect -35 847 -19 881
rect 19 847 35 881
rect 93 847 109 881
rect 147 847 163 881
rect 221 847 237 881
rect 275 847 291 881
rect 349 847 365 881
rect 403 847 419 881
rect 477 847 493 881
rect 531 847 547 881
rect 605 847 621 881
rect 659 847 675 881
rect 733 847 749 881
rect 787 847 803 881
rect 861 847 877 881
rect 915 847 931 881
rect 989 847 1005 881
rect 1043 847 1059 881
rect 1117 847 1133 881
rect 1171 847 1187 881
rect 1245 847 1261 881
rect 1299 847 1315 881
rect 1373 847 1389 881
rect 1427 847 1443 881
rect 1501 847 1517 881
rect 1555 847 1571 881
rect 1629 847 1645 881
rect 1683 847 1699 881
rect 1757 847 1773 881
rect 1811 847 1827 881
rect 1885 847 1901 881
rect 1939 847 1955 881
rect -2001 788 -1967 804
rect -2001 -804 -1967 -788
rect -1873 788 -1839 804
rect -1873 -804 -1839 -788
rect -1745 788 -1711 804
rect -1745 -804 -1711 -788
rect -1617 788 -1583 804
rect -1617 -804 -1583 -788
rect -1489 788 -1455 804
rect -1489 -804 -1455 -788
rect -1361 788 -1327 804
rect -1361 -804 -1327 -788
rect -1233 788 -1199 804
rect -1233 -804 -1199 -788
rect -1105 788 -1071 804
rect -1105 -804 -1071 -788
rect -977 788 -943 804
rect -977 -804 -943 -788
rect -849 788 -815 804
rect -849 -804 -815 -788
rect -721 788 -687 804
rect -721 -804 -687 -788
rect -593 788 -559 804
rect -593 -804 -559 -788
rect -465 788 -431 804
rect -465 -804 -431 -788
rect -337 788 -303 804
rect -337 -804 -303 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -81 788 -47 804
rect -81 -804 -47 -788
rect 47 788 81 804
rect 47 -804 81 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 303 788 337 804
rect 303 -804 337 -788
rect 431 788 465 804
rect 431 -804 465 -788
rect 559 788 593 804
rect 559 -804 593 -788
rect 687 788 721 804
rect 687 -804 721 -788
rect 815 788 849 804
rect 815 -804 849 -788
rect 943 788 977 804
rect 943 -804 977 -788
rect 1071 788 1105 804
rect 1071 -804 1105 -788
rect 1199 788 1233 804
rect 1199 -804 1233 -788
rect 1327 788 1361 804
rect 1327 -804 1361 -788
rect 1455 788 1489 804
rect 1455 -804 1489 -788
rect 1583 788 1617 804
rect 1583 -804 1617 -788
rect 1711 788 1745 804
rect 1711 -804 1745 -788
rect 1839 788 1873 804
rect 1839 -804 1873 -788
rect 1967 788 2001 804
rect 1967 -804 2001 -788
rect -1955 -881 -1939 -847
rect -1901 -881 -1885 -847
rect -1827 -881 -1811 -847
rect -1773 -881 -1757 -847
rect -1699 -881 -1683 -847
rect -1645 -881 -1629 -847
rect -1571 -881 -1555 -847
rect -1517 -881 -1501 -847
rect -1443 -881 -1427 -847
rect -1389 -881 -1373 -847
rect -1315 -881 -1299 -847
rect -1261 -881 -1245 -847
rect -1187 -881 -1171 -847
rect -1133 -881 -1117 -847
rect -1059 -881 -1043 -847
rect -1005 -881 -989 -847
rect -931 -881 -915 -847
rect -877 -881 -861 -847
rect -803 -881 -787 -847
rect -749 -881 -733 -847
rect -675 -881 -659 -847
rect -621 -881 -605 -847
rect -547 -881 -531 -847
rect -493 -881 -477 -847
rect -419 -881 -403 -847
rect -365 -881 -349 -847
rect -291 -881 -275 -847
rect -237 -881 -221 -847
rect -163 -881 -147 -847
rect -109 -881 -93 -847
rect -35 -881 -19 -847
rect 19 -881 35 -847
rect 93 -881 109 -847
rect 147 -881 163 -847
rect 221 -881 237 -847
rect 275 -881 291 -847
rect 349 -881 365 -847
rect 403 -881 419 -847
rect 477 -881 493 -847
rect 531 -881 547 -847
rect 605 -881 621 -847
rect 659 -881 675 -847
rect 733 -881 749 -847
rect 787 -881 803 -847
rect 861 -881 877 -847
rect 915 -881 931 -847
rect 989 -881 1005 -847
rect 1043 -881 1059 -847
rect 1117 -881 1133 -847
rect 1171 -881 1187 -847
rect 1245 -881 1261 -847
rect 1299 -881 1315 -847
rect 1373 -881 1389 -847
rect 1427 -881 1443 -847
rect 1501 -881 1517 -847
rect 1555 -881 1571 -847
rect 1629 -881 1645 -847
rect 1683 -881 1699 -847
rect 1757 -881 1773 -847
rect 1811 -881 1827 -847
rect 1885 -881 1901 -847
rect 1939 -881 1955 -847
rect -2115 -949 -2081 -887
rect 3121 -949 3155 -887
rect -2115 -983 -2019 -949
rect 2019 -983 3155 -949
<< viali >>
rect -1939 847 -1901 881
rect -1811 847 -1773 881
rect -1683 847 -1645 881
rect -1555 847 -1517 881
rect -1427 847 -1389 881
rect -1299 847 -1261 881
rect -1171 847 -1133 881
rect -1043 847 -1005 881
rect -915 847 -877 881
rect -787 847 -749 881
rect -659 847 -621 881
rect -531 847 -493 881
rect -403 847 -365 881
rect -275 847 -237 881
rect -147 847 -109 881
rect -19 847 19 881
rect 109 847 147 881
rect 237 847 275 881
rect 365 847 403 881
rect 493 847 531 881
rect 621 847 659 881
rect 749 847 787 881
rect 877 847 915 881
rect 1005 847 1043 881
rect 1133 847 1171 881
rect 1261 847 1299 881
rect 1389 847 1427 881
rect 1517 847 1555 881
rect 1645 847 1683 881
rect 1773 847 1811 881
rect 1901 847 1939 881
rect -2001 -788 -1967 788
rect -1873 -788 -1839 788
rect -1745 -788 -1711 788
rect -1617 -788 -1583 788
rect -1489 -788 -1455 788
rect -1361 -788 -1327 788
rect -1233 -788 -1199 788
rect -1105 -788 -1071 788
rect -977 -788 -943 788
rect -849 -788 -815 788
rect -721 -788 -687 788
rect -593 -788 -559 788
rect -465 -788 -431 788
rect -337 -788 -303 788
rect -209 -788 -175 788
rect -81 -788 -47 788
rect 47 -788 81 788
rect 175 -788 209 788
rect 303 -788 337 788
rect 431 -788 465 788
rect 559 -788 593 788
rect 687 -788 721 788
rect 815 -788 849 788
rect 943 -788 977 788
rect 1071 -788 1105 788
rect 1199 -788 1233 788
rect 1327 -788 1361 788
rect 1455 -788 1489 788
rect 1583 -788 1617 788
rect 1711 -788 1745 788
rect 1839 -788 1873 788
rect 1967 -788 2001 788
rect -1939 -881 -1901 -847
rect -1811 -881 -1773 -847
rect -1683 -881 -1645 -847
rect -1555 -881 -1517 -847
rect -1427 -881 -1389 -847
rect -1299 -881 -1261 -847
rect -1171 -881 -1133 -847
rect -1043 -881 -1005 -847
rect -915 -881 -877 -847
rect -787 -881 -749 -847
rect -659 -881 -621 -847
rect -531 -881 -493 -847
rect -403 -881 -365 -847
rect -275 -881 -237 -847
rect -147 -881 -109 -847
rect -19 -881 19 -847
rect 109 -881 147 -847
rect 237 -881 275 -847
rect 365 -881 403 -847
rect 493 -881 531 -847
rect 621 -881 659 -847
rect 749 -881 787 -847
rect 877 -881 915 -847
rect 1005 -881 1043 -847
rect 1133 -881 1171 -847
rect 1261 -881 1299 -847
rect 1389 -881 1427 -847
rect 1517 -881 1555 -847
rect 1645 -881 1683 -847
rect 1773 -881 1811 -847
rect 1901 -881 1939 -847
<< metal1 >>
rect -1951 881 -1889 887
rect -1951 847 -1939 881
rect -1901 847 -1889 881
rect -1951 841 -1889 847
rect -1823 881 -1761 887
rect -1823 847 -1811 881
rect -1773 847 -1761 881
rect -1823 841 -1761 847
rect -1695 881 -1633 887
rect -1695 847 -1683 881
rect -1645 847 -1633 881
rect -1695 841 -1633 847
rect -1567 881 -1505 887
rect -1567 847 -1555 881
rect -1517 847 -1505 881
rect -1567 841 -1505 847
rect -1439 881 -1377 887
rect -1439 847 -1427 881
rect -1389 847 -1377 881
rect -1439 841 -1377 847
rect -1311 881 -1249 887
rect -1311 847 -1299 881
rect -1261 847 -1249 881
rect -1311 841 -1249 847
rect -1183 881 -1121 887
rect -1183 847 -1171 881
rect -1133 847 -1121 881
rect -1183 841 -1121 847
rect -1055 881 -993 887
rect -1055 847 -1043 881
rect -1005 847 -993 881
rect -1055 841 -993 847
rect -927 881 -865 887
rect -927 847 -915 881
rect -877 847 -865 881
rect -927 841 -865 847
rect -799 881 -737 887
rect -799 847 -787 881
rect -749 847 -737 881
rect -799 841 -737 847
rect -671 881 -609 887
rect -671 847 -659 881
rect -621 847 -609 881
rect -671 841 -609 847
rect -543 881 -481 887
rect -543 847 -531 881
rect -493 847 -481 881
rect -543 841 -481 847
rect -415 881 -353 887
rect -415 847 -403 881
rect -365 847 -353 881
rect -415 841 -353 847
rect -287 881 -225 887
rect -287 847 -275 881
rect -237 847 -225 881
rect -287 841 -225 847
rect -159 881 -97 887
rect -159 847 -147 881
rect -109 847 -97 881
rect -159 841 -97 847
rect -31 881 31 887
rect -31 847 -19 881
rect 19 847 31 881
rect -31 841 31 847
rect 97 881 159 887
rect 97 847 109 881
rect 147 847 159 881
rect 97 841 159 847
rect 225 881 287 887
rect 225 847 237 881
rect 275 847 287 881
rect 225 841 287 847
rect 353 881 415 887
rect 353 847 365 881
rect 403 847 415 881
rect 353 841 415 847
rect 481 881 543 887
rect 481 847 493 881
rect 531 847 543 881
rect 481 841 543 847
rect 609 881 671 887
rect 609 847 621 881
rect 659 847 671 881
rect 609 841 671 847
rect 737 881 799 887
rect 737 847 749 881
rect 787 847 799 881
rect 737 841 799 847
rect 865 881 927 887
rect 865 847 877 881
rect 915 847 927 881
rect 865 841 927 847
rect 993 881 1055 887
rect 993 847 1005 881
rect 1043 847 1055 881
rect 993 841 1055 847
rect 1121 881 1183 887
rect 1121 847 1133 881
rect 1171 847 1183 881
rect 1121 841 1183 847
rect 1249 881 1311 887
rect 1249 847 1261 881
rect 1299 847 1311 881
rect 1249 841 1311 847
rect 1377 881 1439 887
rect 1377 847 1389 881
rect 1427 847 1439 881
rect 1377 841 1439 847
rect 1505 881 1567 887
rect 1505 847 1517 881
rect 1555 847 1567 881
rect 1505 841 1567 847
rect 1633 881 1695 887
rect 1633 847 1645 881
rect 1683 847 1695 881
rect 1633 841 1695 847
rect 1761 881 1823 887
rect 1761 847 1773 881
rect 1811 847 1823 881
rect 1761 841 1823 847
rect 1889 881 1951 887
rect 1889 847 1901 881
rect 1939 847 1951 881
rect 1889 841 1951 847
rect -2007 788 -1961 800
rect -2007 -788 -2001 788
rect -1967 -788 -1961 788
rect -2007 -800 -1961 -788
rect -1879 788 -1833 800
rect -1879 -788 -1873 788
rect -1839 -788 -1833 788
rect -1879 -800 -1833 -788
rect -1751 788 -1705 800
rect -1751 -788 -1745 788
rect -1711 -788 -1705 788
rect -1751 -800 -1705 -788
rect -1623 788 -1577 800
rect -1623 -788 -1617 788
rect -1583 -788 -1577 788
rect -1623 -800 -1577 -788
rect -1495 788 -1449 800
rect -1495 -788 -1489 788
rect -1455 -788 -1449 788
rect -1495 -800 -1449 -788
rect -1367 788 -1321 800
rect -1367 -788 -1361 788
rect -1327 -788 -1321 788
rect -1367 -800 -1321 -788
rect -1239 788 -1193 800
rect -1239 -788 -1233 788
rect -1199 -788 -1193 788
rect -1239 -800 -1193 -788
rect -1111 788 -1065 800
rect -1111 -788 -1105 788
rect -1071 -788 -1065 788
rect -1111 -800 -1065 -788
rect -983 788 -937 800
rect -983 -788 -977 788
rect -943 -788 -937 788
rect -983 -800 -937 -788
rect -855 788 -809 800
rect -855 -788 -849 788
rect -815 -788 -809 788
rect -855 -800 -809 -788
rect -727 788 -681 800
rect -727 -788 -721 788
rect -687 -788 -681 788
rect -727 -800 -681 -788
rect -599 788 -553 800
rect -599 -788 -593 788
rect -559 -788 -553 788
rect -599 -800 -553 -788
rect -471 788 -425 800
rect -471 -788 -465 788
rect -431 -788 -425 788
rect -471 -800 -425 -788
rect -343 788 -297 800
rect -343 -788 -337 788
rect -303 -788 -297 788
rect -343 -800 -297 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -87 788 -41 800
rect -87 -788 -81 788
rect -47 -788 -41 788
rect -87 -800 -41 -788
rect 41 788 87 800
rect 41 -788 47 788
rect 81 -788 87 788
rect 41 -800 87 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 297 788 343 800
rect 297 -788 303 788
rect 337 -788 343 788
rect 297 -800 343 -788
rect 425 788 471 800
rect 425 -788 431 788
rect 465 -788 471 788
rect 425 -800 471 -788
rect 553 788 599 800
rect 553 -788 559 788
rect 593 -788 599 788
rect 553 -800 599 -788
rect 681 788 727 800
rect 681 -788 687 788
rect 721 -788 727 788
rect 681 -800 727 -788
rect 809 788 855 800
rect 809 -788 815 788
rect 849 -788 855 788
rect 809 -800 855 -788
rect 937 788 983 800
rect 937 -788 943 788
rect 977 -788 983 788
rect 937 -800 983 -788
rect 1065 788 1111 800
rect 1065 -788 1071 788
rect 1105 -788 1111 788
rect 1065 -800 1111 -788
rect 1193 788 1239 800
rect 1193 -788 1199 788
rect 1233 -788 1239 788
rect 1193 -800 1239 -788
rect 1321 788 1367 800
rect 1321 -788 1327 788
rect 1361 -788 1367 788
rect 1321 -800 1367 -788
rect 1449 788 1495 800
rect 1449 -788 1455 788
rect 1489 -788 1495 788
rect 1449 -800 1495 -788
rect 1577 788 1623 800
rect 1577 -788 1583 788
rect 1617 -788 1623 788
rect 1577 -800 1623 -788
rect 1705 788 1751 800
rect 1705 -788 1711 788
rect 1745 -788 1751 788
rect 1705 -800 1751 -788
rect 1833 788 1879 800
rect 1833 -788 1839 788
rect 1873 -788 1879 788
rect 1833 -800 1879 -788
rect 1961 788 2007 800
rect 1961 -788 1967 788
rect 2001 -788 2007 788
rect 1961 -800 2007 -788
rect -1951 -847 -1889 -841
rect -1951 -881 -1939 -847
rect -1901 -881 -1889 -847
rect -1951 -887 -1889 -881
rect -1823 -847 -1761 -841
rect -1823 -881 -1811 -847
rect -1773 -881 -1761 -847
rect -1823 -887 -1761 -881
rect -1695 -847 -1633 -841
rect -1695 -881 -1683 -847
rect -1645 -881 -1633 -847
rect -1695 -887 -1633 -881
rect -1567 -847 -1505 -841
rect -1567 -881 -1555 -847
rect -1517 -881 -1505 -847
rect -1567 -887 -1505 -881
rect -1439 -847 -1377 -841
rect -1439 -881 -1427 -847
rect -1389 -881 -1377 -847
rect -1439 -887 -1377 -881
rect -1311 -847 -1249 -841
rect -1311 -881 -1299 -847
rect -1261 -881 -1249 -847
rect -1311 -887 -1249 -881
rect -1183 -847 -1121 -841
rect -1183 -881 -1171 -847
rect -1133 -881 -1121 -847
rect -1183 -887 -1121 -881
rect -1055 -847 -993 -841
rect -1055 -881 -1043 -847
rect -1005 -881 -993 -847
rect -1055 -887 -993 -881
rect -927 -847 -865 -841
rect -927 -881 -915 -847
rect -877 -881 -865 -847
rect -927 -887 -865 -881
rect -799 -847 -737 -841
rect -799 -881 -787 -847
rect -749 -881 -737 -847
rect -799 -887 -737 -881
rect -671 -847 -609 -841
rect -671 -881 -659 -847
rect -621 -881 -609 -847
rect -671 -887 -609 -881
rect -543 -847 -481 -841
rect -543 -881 -531 -847
rect -493 -881 -481 -847
rect -543 -887 -481 -881
rect -415 -847 -353 -841
rect -415 -881 -403 -847
rect -365 -881 -353 -847
rect -415 -887 -353 -881
rect -287 -847 -225 -841
rect -287 -881 -275 -847
rect -237 -881 -225 -847
rect -287 -887 -225 -881
rect -159 -847 -97 -841
rect -159 -881 -147 -847
rect -109 -881 -97 -847
rect -159 -887 -97 -881
rect -31 -847 31 -841
rect -31 -881 -19 -847
rect 19 -881 31 -847
rect -31 -887 31 -881
rect 97 -847 159 -841
rect 97 -881 109 -847
rect 147 -881 159 -847
rect 97 -887 159 -881
rect 225 -847 287 -841
rect 225 -881 237 -847
rect 275 -881 287 -847
rect 225 -887 287 -881
rect 353 -847 415 -841
rect 353 -881 365 -847
rect 403 -881 415 -847
rect 353 -887 415 -881
rect 481 -847 543 -841
rect 481 -881 493 -847
rect 531 -881 543 -847
rect 481 -887 543 -881
rect 609 -847 671 -841
rect 609 -881 621 -847
rect 659 -881 671 -847
rect 609 -887 671 -881
rect 737 -847 799 -841
rect 737 -881 749 -847
rect 787 -881 799 -847
rect 737 -887 799 -881
rect 865 -847 927 -841
rect 865 -881 877 -847
rect 915 -881 927 -847
rect 865 -887 927 -881
rect 993 -847 1055 -841
rect 993 -881 1005 -847
rect 1043 -881 1055 -847
rect 993 -887 1055 -881
rect 1121 -847 1183 -841
rect 1121 -881 1133 -847
rect 1171 -881 1183 -847
rect 1121 -887 1183 -881
rect 1249 -847 1311 -841
rect 1249 -881 1261 -847
rect 1299 -881 1311 -847
rect 1249 -887 1311 -881
rect 1377 -847 1439 -841
rect 1377 -881 1389 -847
rect 1427 -881 1439 -847
rect 1377 -887 1439 -881
rect 1505 -847 1567 -841
rect 1505 -881 1517 -847
rect 1555 -881 1567 -847
rect 1505 -887 1567 -881
rect 1633 -847 1695 -841
rect 1633 -881 1645 -847
rect 1683 -881 1695 -847
rect 1633 -887 1695 -881
rect 1761 -847 1823 -841
rect 1761 -881 1773 -847
rect 1811 -881 1823 -847
rect 1761 -887 1823 -881
rect 1889 -847 1951 -841
rect 1889 -881 1901 -847
rect 1939 -881 1951 -847
rect 1889 -887 1951 -881
<< properties >>
string FIXED_BBOX -2098 -966 2098 966
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.35 m 1 nf 31 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
