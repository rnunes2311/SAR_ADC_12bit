* NGSPICE file created from latched_comparator.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_7XK7PK a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_DTMSLK a_n182_n100# a_n348_n188# a_120_n100# a_28_n100#
+ a_n494_n274# a_n392_n100# a_330_n100# a_238_n100# a_n90_n100# a_n138_122# a_72_n188#
+ a_n300_n100# a_282_122#
X0 a_120_n100# a_72_n188# a_28_n100# a_n494_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1 a_330_n100# a_282_122# a_238_n100# a_n494_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2 a_n90_n100# a_n138_122# a_n182_n100# a_n494_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3 a_n300_n100# a_n348_n188# a_n392_n100# a_n494_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_UNYNRG a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGASDL a_n73_n400# a_15_n400# w_n211_n619# a_n33_n497#
X0 a_15_n400# a_n33_n497# a_n73_n400# w_n211_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_YRYNRG a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_KPCVAL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XG57AL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt latched_comparator VDD VIN_P VIN_N EN OUT_P OUT_N VSS
Xx1 EN VSS VSS VDD VDD x1/X sky130_fd_sc_hd__buf_4
Xx4 x4/A VSS VSS VDD VDD x7/A sky130_fd_sc_hd__inv_1
Xsky130_fd_pr__nfet_01v8_648S5X_0 m1_5800_n430# x4/A x5/A VSS sky130_fd_pr__nfet_01v8_648S5X
Xx5 x5/A VSS VSS VDD VDD x6/A sky130_fd_sc_hd__inv_1
Xx6 x6/A VSS VSS VDD VDD OUT_N sky130_fd_sc_hd__inv_4
XXM18 m1_6590_n1230# VSS VSS x1/X sky130_fd_pr__nfet_01v8_7XK7PK
Xx7 x7/A VSS VSS VDD VDD OUT_P sky130_fd_sc_hd__inv_4
XXM1 m1_5800_n430# m1_6590_n1230# m1_6380_n1050# m1_6590_n1230# VSS m1_6590_n1230#
+ m1_6590_n1230# m1_6590_n1230# m1_6590_n1230# VIN_P VIN_N m1_6590_n1230# m1_6590_n1230#
+ sky130_fd_pr__nfet_01v8_lvt_DTMSLK
XXM4 x4/A x5/A m1_6380_n1050# VSS sky130_fd_pr__nfet_01v8_648S5X
XXM5 VDD x5/A VDD x1/X sky130_fd_pr__pfet_01v8_UNYNRG
XXM6 VDD x5/A VDD x4/A sky130_fd_pr__pfet_01v8_XGASDL
XXM9 x4/A VDD VDD x5/A sky130_fd_pr__pfet_01v8_XGASDL
XXM10 VDD m1_5800_n430# VDD x1/X sky130_fd_pr__pfet_01v8_YRYNRG
Xsky130_fd_pr__pfet_01v8_KPCVAL_0 m1_6380_n1050# VDD VDD x1/X sky130_fd_pr__pfet_01v8_KPCVAL
XXM11 x4/A VDD VDD x1/X sky130_fd_pr__pfet_01v8_XG57AL
Xsky130_fd_pr__nfet_01v8_7XK7PK_0 m1_6590_n1230# VSS VSS x1/X sky130_fd_pr__nfet_01v8_7XK7PK
.ends

