magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -239 272 -181 278
rect 181 272 239 278
rect -239 238 -227 272
rect 181 238 193 272
rect -239 232 -181 238
rect 181 232 239 238
rect -449 -238 -391 -232
rect -29 -238 29 -232
rect 391 -238 449 -232
rect -449 -272 -437 -238
rect -29 -272 -17 -238
rect 391 -272 403 -238
rect -449 -278 -391 -272
rect -29 -278 29 -272
rect 391 -278 449 -272
<< pwell >>
rect -635 -410 635 410
<< nmos >>
rect -435 -200 -405 200
rect -225 -200 -195 200
rect -15 -200 15 200
rect 195 -200 225 200
rect 405 -200 435 200
<< ndiff >>
rect -497 188 -435 200
rect -497 -188 -485 188
rect -451 -188 -435 188
rect -497 -200 -435 -188
rect -405 188 -343 200
rect -405 -188 -389 188
rect -355 -188 -343 188
rect -405 -200 -343 -188
rect -287 188 -225 200
rect -287 -188 -275 188
rect -241 -188 -225 188
rect -287 -200 -225 -188
rect -195 188 -133 200
rect -195 -188 -179 188
rect -145 -188 -133 188
rect -195 -200 -133 -188
rect -77 188 -15 200
rect -77 -188 -65 188
rect -31 -188 -15 188
rect -77 -200 -15 -188
rect 15 188 77 200
rect 15 -188 31 188
rect 65 -188 77 188
rect 15 -200 77 -188
rect 133 188 195 200
rect 133 -188 145 188
rect 179 -188 195 188
rect 133 -200 195 -188
rect 225 188 287 200
rect 225 -188 241 188
rect 275 -188 287 188
rect 225 -200 287 -188
rect 343 188 405 200
rect 343 -188 355 188
rect 389 -188 405 188
rect 343 -200 405 -188
rect 435 188 497 200
rect 435 -188 451 188
rect 485 -188 497 188
rect 435 -200 497 -188
<< ndiffc >>
rect -485 -188 -451 188
rect -389 -188 -355 188
rect -275 -188 -241 188
rect -179 -188 -145 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 145 -188 179 188
rect 241 -188 275 188
rect 355 -188 389 188
rect 451 -188 485 188
<< psubdiff >>
rect -599 340 -503 374
rect 503 340 599 374
rect -599 278 -565 340
rect 565 278 599 340
rect -599 -340 -565 -278
rect 565 -340 599 -278
rect -599 -374 -503 -340
rect 503 -374 599 -340
<< psubdiffcont >>
rect -503 340 503 374
rect -599 -278 -565 278
rect 565 -278 599 278
rect -503 -374 503 -340
<< poly >>
rect -243 272 -177 288
rect -243 238 -227 272
rect -193 238 -177 272
rect -435 200 -405 226
rect -243 222 -177 238
rect 177 272 243 288
rect 177 238 193 272
rect 227 238 243 272
rect -225 200 -195 222
rect -15 200 15 226
rect 177 222 243 238
rect 195 200 225 222
rect 405 200 435 226
rect -435 -222 -405 -200
rect -453 -238 -387 -222
rect -225 -226 -195 -200
rect -15 -222 15 -200
rect -453 -272 -437 -238
rect -403 -272 -387 -238
rect -453 -288 -387 -272
rect -33 -238 33 -222
rect 195 -226 225 -200
rect 405 -222 435 -200
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
rect 387 -238 453 -222
rect 387 -272 403 -238
rect 437 -272 453 -238
rect 387 -288 453 -272
<< polycont >>
rect -227 238 -193 272
rect 193 238 227 272
rect -437 -272 -403 -238
rect -17 -272 17 -238
rect 403 -272 437 -238
<< locali >>
rect -599 340 -503 374
rect 503 340 599 374
rect -599 278 -565 340
rect 565 278 599 340
rect -243 238 -227 272
rect -193 238 -177 272
rect 177 238 193 272
rect 227 238 243 272
rect -485 188 -451 204
rect -485 -204 -451 -188
rect -389 188 -355 204
rect -389 -204 -355 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -179 188 -145 204
rect -179 -204 -145 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 145 188 179 204
rect 145 -204 179 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 355 188 389 204
rect 355 -204 389 -188
rect 451 188 485 204
rect 451 -204 485 -188
rect -453 -272 -437 -238
rect -403 -272 -387 -238
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 387 -272 403 -238
rect 437 -272 453 -238
rect -599 -340 -565 -278
rect 565 -340 599 -278
rect -599 -374 -503 -340
rect 503 -374 599 -340
<< viali >>
rect -227 238 -193 272
rect 193 238 227 272
rect -485 -188 -451 188
rect -389 -188 -355 188
rect -275 -188 -241 188
rect -179 -188 -145 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 145 -188 179 188
rect 241 -188 275 188
rect 355 -188 389 188
rect 451 -188 485 188
rect -437 -272 -403 -238
rect -17 -272 17 -238
rect 403 -272 437 -238
<< metal1 >>
rect -239 272 -181 278
rect -239 238 -227 272
rect -193 238 -181 272
rect -239 232 -181 238
rect 181 272 239 278
rect 181 238 193 272
rect 227 238 239 272
rect 181 232 239 238
rect -491 188 -445 200
rect -491 -188 -485 188
rect -451 -188 -445 188
rect -491 -200 -445 -188
rect -395 188 -349 200
rect -395 -188 -389 188
rect -355 -188 -349 188
rect -395 -200 -349 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -185 188 -139 200
rect -185 -188 -179 188
rect -145 -188 -139 188
rect -185 -200 -139 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 139 188 185 200
rect 139 -188 145 188
rect 179 -188 185 188
rect 139 -200 185 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 349 188 395 200
rect 349 -188 355 188
rect 389 -188 395 188
rect 349 -200 395 -188
rect 445 188 491 200
rect 445 -188 451 188
rect 485 -188 491 188
rect 445 -200 491 -188
rect -449 -238 -391 -232
rect -449 -272 -437 -238
rect -403 -272 -391 -238
rect -449 -278 -391 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 391 -238 449 -232
rect 391 -272 403 -238
rect 437 -272 449 -238
rect 391 -278 449 -272
<< properties >>
string FIXED_BBOX -582 -357 582 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
