magic
tech sky130A
magscale 1 2
timestamp 1711310191
<< metal3 >>
rect -1615 712 1615 740
rect -1615 -712 1531 712
rect 1595 -712 1615 712
rect -1615 -740 1615 -712
<< via3 >>
rect 1531 -712 1595 712
<< mimcap >>
rect -1575 660 1283 700
rect -1575 -660 -1535 660
rect 1243 -660 1283 660
rect -1575 -700 1283 -660
<< mimcapcontact >>
rect -1535 -660 1243 660
<< metal4 >>
rect 1515 712 1611 728
rect -1536 660 1244 661
rect -1536 -660 -1535 660
rect 1243 -660 1244 660
rect -1536 -661 1244 -660
rect 1515 -712 1531 712
rect 1595 -712 1611 712
rect 1515 -728 1611 -712
<< properties >>
string FIXED_BBOX -1615 -740 1323 740
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 14.29 l 7 val 208.15 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
