* NGSPICE file created from offset_calibration_flat.ext - technology: sky130A

.subckt offset_calibration VDD CAL_RESULT EN_COMP CAL_P CAL_N EN VSS CAL_CYCLE
X0 VSS LOAD_CAL_Z a_10288_1192# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 LOAD_CAL_Z a_10364_648# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X2 a_10640_648# CAL_CYCLE VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 a_10524_61# EN_COMP_Z a_10428_61# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 VDD CAL_RESULTi a_10524_n355# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 VDD CAL_CYCLE EN_COMP_Z VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=26.6508 ps=198.34 w=10 l=10
X7 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X8 VDD CAL_CYCLE CAL_RESULT_Z VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VSS EN_COMP_Z EN_COMPi VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_10364_648# EN_COMPi VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11 a_10428_61# LOAD_CAL_Z CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X12 a_10428_61# a_10288_1192# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X13 VDD EN LOAD_CAL_Z VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14 a_10524_n355# EN_COMP_Z a_10428_n355# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 VSS CAL_RESULT_Z CAL_RESULTi VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_10640_648# CAL_CYCLE VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_10428_n355# a_10288_1192# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X18 VSS CAL_CYCLE a_10599_1736# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VDD a_10640_648# LOAD_CAL_Z VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_10695_1512# a_10364_648# a_10599_1512# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 a_10364_648# EN_COMPi VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X22 EN_COMP_Z EN_COMP VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 a_10428_n355# LOAD_CAL_Z CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X25 VSS CAL_CYCLE a_10599_2600# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X27 CAL_RESULT_Z CAL_RESULT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 a_10536_n1060# EN_COMPi a_10428_61# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X29 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X30 a_10599_1512# EN LOAD_CAL_Z VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VDD LOAD_CAL_Z a_10288_1192# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X32 a_10536_n1458# EN_COMPi a_10428_n355# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X33 VSS CAL_RESULT_Z a_10536_n1060# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X34 VSS a_10640_648# a_10695_1512# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 CAL_P EN VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X36 a_10599_1736# EN_COMP EN_COMP_Z VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X37 CAL_N EN VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X38 VSS CAL_RESULTi a_10536_n1458# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X39 VDD EN_COMP_Z EN_COMPi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X40 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X41 a_10599_2600# CAL_RESULT CAL_RESULT_Z VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X42 VDD CAL_RESULT_Z CAL_RESULTi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X43 VDD CAL_RESULT_Z a_10524_61# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
C0 EN CAL_P 0.026947f
C1 EN_COMP EN 0.013548f
C2 a_10288_1192# CAL_P 0.024901f
C3 CAL_CYCLE EN 0.049117f
C4 a_10288_1192# EN 0.558498f
C5 CAL_RESULT EN 1.29e-20
C6 CAL_CYCLE EN_COMP 0.320018f
C7 CAL_N CAL_P 4.36627f
C8 a_10640_648# EN 0.093387f
C9 a_10288_1192# EN_COMP 0.001213f
C10 CAL_N EN 0.072224f
C11 CAL_RESULT EN_COMP 0.013171f
C12 VDD CAL_P 21.066301f
C13 a_10364_648# EN 0.253407f
C14 a_10640_648# EN_COMP 1.27e-19
C15 a_10288_1192# CAL_CYCLE 0.019601f
C16 LOAD_CAL_Z CAL_P 0.027034f
C17 VDD EN 0.83887f
C18 CAL_N EN_COMP 0.004981f
C19 CAL_RESULT CAL_CYCLE 0.55451f
C20 LOAD_CAL_Z EN 0.789507f
C21 a_10364_648# EN_COMP 5.47e-21
C22 a_10288_1192# CAL_RESULT 1.58e-20
C23 a_10640_648# CAL_CYCLE 0.136508f
C24 a_10536_n1458# CAL_P 9.62e-21
C25 VDD EN_COMP 0.125946f
C26 CAL_N CAL_CYCLE 0.00144f
C27 a_10640_648# a_10288_1192# 0.039734f
C28 a_10288_1192# CAL_N 0.024229f
C29 LOAD_CAL_Z EN_COMP 8.82e-19
C30 a_10640_648# CAL_RESULT 3.43e-20
C31 a_10364_648# CAL_CYCLE 0.038804f
C32 EN_COMPi CAL_P 0.005678f
C33 a_10536_n1060# CAL_P 1.35e-20
C34 VDD CAL_CYCLE 0.379163f
C35 CAL_N CAL_RESULT 0.005179f
C36 a_10364_648# a_10288_1192# 0.049703f
C37 EN_COMP_Z CAL_P 0.001469f
C38 a_10288_1192# VDD 0.356405f
C39 a_10640_648# CAL_N 2.99e-19
C40 EN_COMPi EN 0.666122f
C41 a_10599_1736# EN_COMP 4.3e-20
C42 a_10364_648# CAL_RESULT 2.05e-21
C43 LOAD_CAL_Z CAL_CYCLE 0.031209f
C44 a_10524_n355# CAL_P 1.58e-20
C45 VDD CAL_RESULT 0.093873f
C46 a_10364_648# a_10640_648# 0.235701f
C47 LOAD_CAL_Z a_10288_1192# 1.0295f
C48 a_10640_648# VDD 0.431879f
C49 a_10364_648# CAL_N 0.01247f
C50 EN_COMP_Z EN 0.213948f
C51 EN_COMPi EN_COMP 0.418198f
C52 LOAD_CAL_Z CAL_RESULT 6.33e-21
C53 a_10599_1736# CAL_CYCLE 1.96e-20
C54 a_10428_n355# CAL_P 0.205305f
C55 VDD CAL_N 20.9316f
C56 a_10524_n355# EN 1.35e-19
C57 a_10599_1736# a_10288_1192# 1.28e-20
C58 LOAD_CAL_Z a_10640_648# 0.112629f
C59 CAL_RESULTi CAL_P 0.001716f
C60 a_10364_648# VDD 0.536989f
C61 a_10288_1192# a_10536_n1458# 0.003149f
C62 LOAD_CAL_Z CAL_N 0.023597f
C63 EN_COMP_Z EN_COMP 0.260892f
C64 EN_COMPi CAL_CYCLE 0.242946f
C65 a_10428_n355# EN 3.5e-19
C66 EN_COMPi a_10288_1192# 0.353611f
C67 LOAD_CAL_Z a_10364_648# 0.27533f
C68 CAL_RESULT_Z CAL_P 6.35e-19
C69 LOAD_CAL_Z VDD 0.910209f
C70 a_10288_1192# a_10536_n1060# 0.002793f
C71 CAL_RESULTi EN 0.056594f
C72 EN_COMPi CAL_RESULT 6.22e-19
C73 EN_COMP_Z CAL_CYCLE 0.681137f
C74 a_10428_61# CAL_P 2.83e-19
C75 a_10524_n355# CAL_CYCLE 1.13e-20
C76 a_10524_61# EN 0.003319f
C77 EN_COMPi a_10640_648# 0.013073f
C78 EN_COMP_Z a_10288_1192# 0.037283f
C79 a_10599_1736# VDD 2.4e-19
C80 a_10288_1192# a_10524_n355# 3.12e-20
C81 EN_COMPi CAL_N 0.014789f
C82 CAL_RESULT_Z EN 0.072601f
C83 CAL_RESULTi EN_COMP 0.021292f
C84 EN_COMP_Z CAL_RESULT 1.09e-20
C85 a_10536_n1458# VDD 1.72e-20
C86 a_10536_n1060# CAL_N 7.87e-21
C87 a_10428_61# EN 0.20695f
C88 EN_COMPi a_10364_648# 0.121283f
C89 a_10599_1736# LOAD_CAL_Z 1.39e-19
C90 EN_COMP_Z a_10640_648# 0.131339f
C91 EN_COMPi VDD 0.666146f
C92 EN_COMP_Z CAL_N 6.29e-19
C93 CAL_RESULT_Z EN_COMP 0.021074f
C94 a_10599_2600# CAL_RESULT 3.7e-19
C95 CAL_RESULTi CAL_CYCLE 0.954497f
C96 a_10288_1192# a_10428_n355# 0.490939f
C97 a_10524_61# CAL_CYCLE 2.84e-20
C98 a_10536_n1060# VDD 3.6e-19
C99 CAL_RESULTi a_10288_1192# 0.604831f
C100 EN_COMPi LOAD_CAL_Z 0.126839f
C101 EN_COMP_Z a_10364_648# 0.004924f
C102 EN_COMP_Z VDD 1.04406f
C103 LOAD_CAL_Z a_10536_n1060# 2.12e-20
C104 CAL_RESULTi CAL_RESULT 0.069062f
C105 CAL_RESULT_Z CAL_CYCLE 0.131557f
C106 a_10428_61# CAL_CYCLE 1.37e-20
C107 a_10524_n355# VDD 0.085164f
C108 a_10428_n355# CAL_N 4.7e-20
C109 CAL_RESULTi a_10640_648# 0.002743f
C110 EN_COMP_Z LOAD_CAL_Z 0.457858f
C111 CAL_RESULT_Z a_10288_1192# 0.380006f
C112 a_10599_2600# VDD 1.38e-19
C113 LOAD_CAL_Z a_10524_n355# 0.004065f
C114 EN_COMPi a_10536_n1458# 0.011525f
C115 CAL_RESULTi CAL_N 0.007453f
C116 CAL_RESULT_Z CAL_RESULT 0.201616f
C117 a_10288_1192# a_10428_61# 0.198764f
C118 a_10536_n1060# a_10536_n1458# 0.003901f
C119 a_10428_n355# VDD 0.079488f
C120 a_10524_61# CAL_N 4.85e-21
C121 CAL_RESULTi a_10364_648# 9.26e-21
C122 EN_COMP_Z a_10599_1736# 0.010228f
C123 CAL_RESULT_Z a_10640_648# 0.002401f
C124 CAL_RESULTi VDD 0.563202f
C125 EN_COMPi a_10536_n1060# 0.012249f
C126 CAL_RESULT_Z CAL_N 0.006786f
C127 a_10640_648# a_10428_61# 8.2e-19
C128 a_10288_1192# a_10695_1512# 2.68e-19
C129 LOAD_CAL_Z a_10428_n355# 0.333805f
C130 a_10524_61# VDD 0.085998f
C131 a_10428_61# CAL_N 0.204621f
C132 CAL_RESULTi LOAD_CAL_Z 0.65678f
C133 EN_COMP_Z EN_COMPi 0.129251f
C134 CAL_RESULT_Z a_10364_648# 6.99e-20
C135 EN_COMPi a_10524_n355# 7.75e-19
C136 CAL_RESULT_Z VDD 0.802151f
C137 a_10364_648# a_10428_61# 2.17e-21
C138 a_10288_1192# a_10599_1512# 1.79e-19
C139 LOAD_CAL_Z a_10524_61# 0.004065f
C140 a_10524_n355# a_10536_n1060# 9.87e-19
C141 a_10428_61# VDD 0.317066f
C142 a_10428_n355# a_10536_n1458# 0.08947f
C143 CAL_RESULT_Z LOAD_CAL_Z 0.365591f
C144 CAL_RESULTi a_10536_n1458# 0.011861f
C145 EN_COMP_Z a_10524_n355# 0.016815f
C146 a_10364_648# a_10695_1512# 4.42e-19
C147 EN_COMPi a_10428_n355# 0.172129f
C148 LOAD_CAL_Z a_10428_61# 0.23688f
C149 a_10695_1512# VDD 3.12e-19
C150 CAL_RESULTi EN_COMPi 0.245891f
C151 CAL_RESULTi a_10536_n1060# 0.002464f
C152 CAL_RESULT_Z a_10536_n1458# 1.4e-19
C153 a_10364_648# a_10599_1512# 0.003614f
C154 EN_COMPi a_10524_61# 6.64e-21
C155 LOAD_CAL_Z a_10695_1512# 0.011942f
C156 EN_COMP_Z a_10428_n355# 0.234448f
C157 a_10428_n355# a_10524_n355# 0.087835f
C158 a_10599_1512# VDD 2.73e-20
C159 CAL_RESULTi EN_COMP_Z 0.076632f
C160 CAL_RESULT_Z EN_COMPi 1.41583f
C161 CAL_RESULTi a_10524_n355# 0.010408f
C162 CAL_RESULT_Z a_10536_n1060# 0.010048f
C163 EN_COMPi a_10428_61# 0.12318f
C164 LOAD_CAL_Z a_10599_1512# 0.01318f
C165 EN_COMP_Z a_10524_61# 0.010302f
C166 a_10524_61# a_10524_n355# 0.003483f
C167 a_10428_61# a_10536_n1060# 0.08753f
C168 CAL_RESULTi a_10599_2600# 4.21e-20
C169 CAL_RESULT_Z EN_COMP_Z 0.086402f
C170 CAL_RESULTi a_10428_n355# 0.130478f
C171 EN_COMP_Z a_10428_61# 0.1922f
C172 CAL_RESULT_Z a_10524_n355# 1.29e-19
C173 a_10428_61# a_10524_n355# 3.51e-20
C174 CAL_RESULT_Z a_10599_2600# 0.009658f
C175 CAL_RESULTi a_10524_61# 1.29e-19
C176 EN_COMP_Z a_10695_1512# 4.84e-19
C177 CAL_RESULT_Z a_10428_n355# 0.021352f
C178 a_10428_61# a_10428_n355# 0.32625f
C179 CAL_RESULT_Z CAL_RESULTi 1.99154f
C180 CAL_RESULTi a_10428_61# 0.066321f
C181 EN_COMP_Z a_10599_1512# 3.15e-19
C182 CAL_RESULT_Z a_10524_61# 0.008755f
C183 a_10428_61# a_10524_61# 0.090011f
C184 CAL_RESULT_Z a_10428_61# 0.032572f
C185 CAL_P VSS 7.04953f
C186 EN VSS 0.685064f
C187 EN_COMP VSS 0.371745f
C188 CAL_CYCLE VSS 1.15976f
C189 CAL_RESULT VSS 0.523258f
C190 CAL_N VSS 7.28241f
C191 VDD VSS 0.105798p
C192 a_10536_n1458# VSS 0.090949f 
C193 a_10536_n1060# VSS 0.088947f 
C194 a_10524_n355# VSS 0.004281f 
C195 a_10428_n355# VSS 0.394482f 
C196 a_10524_61# VSS 0.007525f 
C197 a_10428_61# VSS 0.448064f 
C198 a_10695_1512# VSS 9.64e-19 
C199 a_10599_1512# VSS 5.2e-19 
C200 a_10288_1192# VSS 2.52925f 
C201 a_10640_648# VSS 0.501057f 
C202 a_10364_648# VSS 0.287313f 
C203 LOAD_CAL_Z VSS 1.73056f 
C204 a_10599_1736# VSS 0.00198f 
C205 EN_COMPi VSS 2.11464f 
C206 EN_COMP_Z VSS 1.09989f 
C207 a_10599_2600# VSS 0.00202f 
C208 CAL_RESULTi VSS 1.54874f 
C209 CAL_RESULT_Z VSS 1.74553f 
.ends
