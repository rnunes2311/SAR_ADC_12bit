magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -734 -498 734 464
<< nwell >>
rect -734 -498 734 464
<< pmoslvt >>
rect -640 -436 -570 364
rect -398 -436 -328 364
rect -156 -436 -86 364
rect 86 -436 156 364
rect 328 -436 398 364
rect 570 -436 640 364
<< pdiff >>
rect -698 352 -640 364
rect -698 -424 -686 352
rect -652 -424 -640 352
rect -698 -436 -640 -424
rect -570 352 -512 364
rect -570 -424 -558 352
rect -524 -424 -512 352
rect -570 -436 -512 -424
rect -456 352 -398 364
rect -456 -424 -444 352
rect -410 -424 -398 352
rect -456 -436 -398 -424
rect -328 352 -270 364
rect -328 -424 -316 352
rect -282 -424 -270 352
rect -328 -436 -270 -424
rect -214 352 -156 364
rect -214 -424 -202 352
rect -168 -424 -156 352
rect -214 -436 -156 -424
rect -86 352 -28 364
rect -86 -424 -74 352
rect -40 -424 -28 352
rect -86 -436 -28 -424
rect 28 352 86 364
rect 28 -424 40 352
rect 74 -424 86 352
rect 28 -436 86 -424
rect 156 352 214 364
rect 156 -424 168 352
rect 202 -424 214 352
rect 156 -436 214 -424
rect 270 352 328 364
rect 270 -424 282 352
rect 316 -424 328 352
rect 270 -436 328 -424
rect 398 352 456 364
rect 398 -424 410 352
rect 444 -424 456 352
rect 398 -436 456 -424
rect 512 352 570 364
rect 512 -424 524 352
rect 558 -424 570 352
rect 512 -436 570 -424
rect 640 352 698 364
rect 640 -424 652 352
rect 686 -424 698 352
rect 640 -436 698 -424
<< pdiffc >>
rect -686 -424 -652 352
rect -558 -424 -524 352
rect -444 -424 -410 352
rect -316 -424 -282 352
rect -202 -424 -168 352
rect -74 -424 -40 352
rect 40 -424 74 352
rect 168 -424 202 352
rect 282 -424 316 352
rect 410 -424 444 352
rect 524 -424 558 352
rect 652 -424 686 352
<< poly >>
rect -640 445 -570 461
rect -640 411 -624 445
rect -586 411 -570 445
rect -640 364 -570 411
rect -398 445 -328 461
rect -398 411 -382 445
rect -344 411 -328 445
rect -398 364 -328 411
rect -156 445 -86 461
rect -156 411 -140 445
rect -102 411 -86 445
rect -156 364 -86 411
rect 86 445 156 461
rect 86 411 102 445
rect 140 411 156 445
rect 86 364 156 411
rect 328 445 398 461
rect 328 411 344 445
rect 382 411 398 445
rect 328 364 398 411
rect 570 445 640 461
rect 570 411 586 445
rect 624 411 640 445
rect 570 364 640 411
rect -640 -462 -570 -436
rect -398 -462 -328 -436
rect -156 -462 -86 -436
rect 86 -462 156 -436
rect 328 -462 398 -436
rect 570 -462 640 -436
<< polycont >>
rect -624 411 -586 445
rect -382 411 -344 445
rect -140 411 -102 445
rect 102 411 140 445
rect 344 411 382 445
rect 586 411 624 445
<< locali >>
rect -640 411 -624 445
rect -586 411 -570 445
rect -398 411 -382 445
rect -344 411 -328 445
rect -156 411 -140 445
rect -102 411 -86 445
rect 86 411 102 445
rect 140 411 156 445
rect 328 411 344 445
rect 382 411 398 445
rect 570 411 586 445
rect 624 411 640 445
rect -686 352 -652 368
rect -686 -440 -652 -424
rect -558 352 -524 368
rect -558 -440 -524 -424
rect -444 352 -410 368
rect -444 -440 -410 -424
rect -316 352 -282 368
rect -316 -440 -282 -424
rect -202 352 -168 368
rect -202 -440 -168 -424
rect -74 352 -40 368
rect -74 -440 -40 -424
rect 40 352 74 368
rect 40 -440 74 -424
rect 168 352 202 368
rect 168 -440 202 -424
rect 282 352 316 368
rect 282 -440 316 -424
rect 410 352 444 368
rect 410 -440 444 -424
rect 524 352 558 368
rect 524 -440 558 -424
rect 652 352 686 368
rect 652 -440 686 -424
<< viali >>
rect -624 411 -586 445
rect -382 411 -344 445
rect -140 411 -102 445
rect 102 411 140 445
rect 344 411 382 445
rect 586 411 624 445
rect -686 -424 -652 352
rect -558 -424 -524 352
rect -444 -424 -410 352
rect -316 -424 -282 352
rect -202 -424 -168 352
rect -74 -424 -40 352
rect 40 -424 74 352
rect 168 -424 202 352
rect 282 -424 316 352
rect 410 -424 444 352
rect 524 -424 558 352
rect 652 -424 686 352
<< metal1 >>
rect -636 445 -574 451
rect -636 411 -624 445
rect -586 411 -574 445
rect -636 405 -574 411
rect -394 445 -332 451
rect -394 411 -382 445
rect -344 411 -332 445
rect -394 405 -332 411
rect -152 445 -90 451
rect -152 411 -140 445
rect -102 411 -90 445
rect -152 405 -90 411
rect 90 445 152 451
rect 90 411 102 445
rect 140 411 152 445
rect 90 405 152 411
rect 332 445 394 451
rect 332 411 344 445
rect 382 411 394 445
rect 332 405 394 411
rect 574 445 636 451
rect 574 411 586 445
rect 624 411 636 445
rect 574 405 636 411
rect -692 352 -646 364
rect -692 -424 -686 352
rect -652 -424 -646 352
rect -692 -436 -646 -424
rect -564 352 -518 364
rect -564 -424 -558 352
rect -524 -424 -518 352
rect -564 -436 -518 -424
rect -450 352 -404 364
rect -450 -424 -444 352
rect -410 -424 -404 352
rect -450 -436 -404 -424
rect -322 352 -276 364
rect -322 -424 -316 352
rect -282 -424 -276 352
rect -322 -436 -276 -424
rect -208 352 -162 364
rect -208 -424 -202 352
rect -168 -424 -162 352
rect -208 -436 -162 -424
rect -80 352 -34 364
rect -80 -424 -74 352
rect -40 -424 -34 352
rect -80 -436 -34 -424
rect 34 352 80 364
rect 34 -424 40 352
rect 74 -424 80 352
rect 34 -436 80 -424
rect 162 352 208 364
rect 162 -424 168 352
rect 202 -424 208 352
rect 162 -436 208 -424
rect 276 352 322 364
rect 276 -424 282 352
rect 316 -424 322 352
rect 276 -436 322 -424
rect 404 352 450 364
rect 404 -424 410 352
rect 444 -424 450 352
rect 404 -436 450 -424
rect 518 352 564 364
rect 518 -424 524 352
rect 558 -424 564 352
rect 518 -436 564 -424
rect 646 352 692 364
rect 646 -424 652 352
rect 686 -424 692 352
rect 646 -436 692 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 0.35 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
