magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< nwell >>
rect -3545 -1017 3545 1017
<< pmos >>
rect -3349 118 -29 798
rect 29 118 3349 798
rect -3349 -798 -29 -118
rect 29 -798 3349 -118
<< pdiff >>
rect -3407 786 -3349 798
rect -3407 130 -3395 786
rect -3361 130 -3349 786
rect -3407 118 -3349 130
rect -29 786 29 798
rect -29 130 -17 786
rect 17 130 29 786
rect -29 118 29 130
rect 3349 786 3407 798
rect 3349 130 3361 786
rect 3395 130 3407 786
rect 3349 118 3407 130
rect -3407 -130 -3349 -118
rect -3407 -786 -3395 -130
rect -3361 -786 -3349 -130
rect -3407 -798 -3349 -786
rect -29 -130 29 -118
rect -29 -786 -17 -130
rect 17 -786 29 -130
rect -29 -798 29 -786
rect 3349 -130 3407 -118
rect 3349 -786 3361 -130
rect 3395 -786 3407 -130
rect 3349 -798 3407 -786
<< pdiffc >>
rect -3395 130 -3361 786
rect -17 130 17 786
rect 3361 130 3395 786
rect -3395 -786 -3361 -130
rect -17 -786 17 -130
rect 3361 -786 3395 -130
<< nsubdiff >>
rect -3509 947 -3413 981
rect 3413 947 3509 981
rect -3509 885 -3475 947
rect 3475 885 3509 947
rect -3509 -947 -3475 -885
rect 3475 -947 3509 -885
rect -3509 -981 -3413 -947
rect 3413 -981 3509 -947
<< nsubdiffcont >>
rect -3413 947 3413 981
rect -3509 -885 -3475 885
rect 3475 -885 3509 885
rect -3413 -981 3413 -947
<< poly >>
rect -3349 879 -29 895
rect -3349 845 -3333 879
rect -45 845 -29 879
rect -3349 798 -29 845
rect 29 879 3349 895
rect 29 845 45 879
rect 3333 845 3349 879
rect 29 798 3349 845
rect -3349 71 -29 118
rect -3349 37 -3333 71
rect -45 37 -29 71
rect -3349 21 -29 37
rect 29 71 3349 118
rect 29 37 45 71
rect 3333 37 3349 71
rect 29 21 3349 37
rect -3349 -37 -29 -21
rect -3349 -71 -3333 -37
rect -45 -71 -29 -37
rect -3349 -118 -29 -71
rect 29 -37 3349 -21
rect 29 -71 45 -37
rect 3333 -71 3349 -37
rect 29 -118 3349 -71
rect -3349 -845 -29 -798
rect -3349 -879 -3333 -845
rect -45 -879 -29 -845
rect -3349 -895 -29 -879
rect 29 -845 3349 -798
rect 29 -879 45 -845
rect 3333 -879 3349 -845
rect 29 -895 3349 -879
<< polycont >>
rect -3333 845 -45 879
rect 45 845 3333 879
rect -3333 37 -45 71
rect 45 37 3333 71
rect -3333 -71 -45 -37
rect 45 -71 3333 -37
rect -3333 -879 -45 -845
rect 45 -879 3333 -845
<< locali >>
rect -3509 947 -3413 981
rect 3413 947 3509 981
rect -3509 885 -3475 947
rect 3475 885 3509 947
rect -3349 845 -3333 879
rect -45 845 -29 879
rect 29 845 45 879
rect 3333 845 3349 879
rect -3395 786 -3361 802
rect -3395 114 -3361 130
rect -17 786 17 802
rect -17 114 17 130
rect 3361 786 3395 802
rect 3361 114 3395 130
rect -3349 37 -3333 71
rect -45 37 -29 71
rect 29 37 45 71
rect 3333 37 3349 71
rect -3349 -71 -3333 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 3333 -71 3349 -37
rect -3395 -130 -3361 -114
rect -3395 -802 -3361 -786
rect -17 -130 17 -114
rect -17 -802 17 -786
rect 3361 -130 3395 -114
rect 3361 -802 3395 -786
rect -3349 -879 -3333 -845
rect -45 -879 -29 -845
rect 29 -879 45 -845
rect 3333 -879 3349 -845
rect -3509 -947 -3475 -885
rect 3475 -947 3509 -885
rect -3509 -981 -3413 -947
rect 3413 -981 3509 -947
<< viali >>
rect -3333 845 -45 879
rect 45 845 3333 879
rect -3395 130 -3361 786
rect -17 130 17 786
rect 3361 130 3395 786
rect -3333 37 -45 71
rect 45 37 3333 71
rect -3333 -71 -45 -37
rect 45 -71 3333 -37
rect -3395 -786 -3361 -130
rect -17 -786 17 -130
rect 3361 -786 3395 -130
rect -3333 -879 -45 -845
rect 45 -879 3333 -845
<< metal1 >>
rect -3345 879 -33 885
rect -3345 845 -3333 879
rect -45 845 -33 879
rect -3345 839 -33 845
rect 33 879 3345 885
rect 33 845 45 879
rect 3333 845 3345 879
rect 33 839 3345 845
rect -3401 786 -3355 798
rect -3401 130 -3395 786
rect -3361 130 -3355 786
rect -3401 118 -3355 130
rect -23 786 23 798
rect -23 130 -17 786
rect 17 130 23 786
rect -23 118 23 130
rect 3355 786 3401 798
rect 3355 130 3361 786
rect 3395 130 3401 786
rect 3355 118 3401 130
rect -3345 71 -33 77
rect -3345 37 -3333 71
rect -45 37 -33 71
rect -3345 31 -33 37
rect 33 71 3345 77
rect 33 37 45 71
rect 3333 37 3345 71
rect 33 31 3345 37
rect -3345 -37 -33 -31
rect -3345 -71 -3333 -37
rect -45 -71 -33 -37
rect -3345 -77 -33 -71
rect 33 -37 3345 -31
rect 33 -71 45 -37
rect 3333 -71 3345 -37
rect 33 -77 3345 -71
rect -3401 -130 -3355 -118
rect -3401 -786 -3395 -130
rect -3361 -786 -3355 -130
rect -3401 -798 -3355 -786
rect -23 -130 23 -118
rect -23 -786 -17 -130
rect 17 -786 23 -130
rect -23 -798 23 -786
rect 3355 -130 3401 -118
rect 3355 -786 3361 -130
rect 3395 -786 3401 -130
rect 3355 -798 3401 -786
rect -3345 -845 -33 -839
rect -3345 -879 -3333 -845
rect -45 -879 -33 -845
rect -3345 -885 -33 -879
rect 33 -845 3345 -839
rect 33 -879 45 -845
rect 3333 -879 3345 -845
rect 33 -885 3345 -879
<< properties >>
string FIXED_BBOX -3492 -964 3492 964
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4 l 16.6 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
