magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< nwell >>
rect -246 -5609 246 5609
<< pmos >>
rect -50 3790 50 5390
rect -50 1954 50 3554
rect -50 118 50 1718
rect -50 -1718 50 -118
rect -50 -3554 50 -1954
rect -50 -5390 50 -3790
<< pdiff >>
rect -108 5378 -50 5390
rect -108 3802 -96 5378
rect -62 3802 -50 5378
rect -108 3790 -50 3802
rect 50 5378 108 5390
rect 50 3802 62 5378
rect 96 3802 108 5378
rect 50 3790 108 3802
rect -108 3542 -50 3554
rect -108 1966 -96 3542
rect -62 1966 -50 3542
rect -108 1954 -50 1966
rect 50 3542 108 3554
rect 50 1966 62 3542
rect 96 1966 108 3542
rect 50 1954 108 1966
rect -108 1706 -50 1718
rect -108 130 -96 1706
rect -62 130 -50 1706
rect -108 118 -50 130
rect 50 1706 108 1718
rect 50 130 62 1706
rect 96 130 108 1706
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -1706 -96 -130
rect -62 -1706 -50 -130
rect -108 -1718 -50 -1706
rect 50 -130 108 -118
rect 50 -1706 62 -130
rect 96 -1706 108 -130
rect 50 -1718 108 -1706
rect -108 -1966 -50 -1954
rect -108 -3542 -96 -1966
rect -62 -3542 -50 -1966
rect -108 -3554 -50 -3542
rect 50 -1966 108 -1954
rect 50 -3542 62 -1966
rect 96 -3542 108 -1966
rect 50 -3554 108 -3542
rect -108 -3802 -50 -3790
rect -108 -5378 -96 -3802
rect -62 -5378 -50 -3802
rect -108 -5390 -50 -5378
rect 50 -3802 108 -3790
rect 50 -5378 62 -3802
rect 96 -5378 108 -3802
rect 50 -5390 108 -5378
<< pdiffc >>
rect -96 3802 -62 5378
rect 62 3802 96 5378
rect -96 1966 -62 3542
rect 62 1966 96 3542
rect -96 130 -62 1706
rect 62 130 96 1706
rect -96 -1706 -62 -130
rect 62 -1706 96 -130
rect -96 -3542 -62 -1966
rect 62 -3542 96 -1966
rect -96 -5378 -62 -3802
rect 62 -5378 96 -3802
<< nsubdiff >>
rect -210 5539 -114 5573
rect 114 5539 210 5573
rect -210 5477 -176 5539
rect 176 5477 210 5539
rect -210 -5539 -176 -5477
rect 176 -5539 210 -5477
rect -210 -5573 -114 -5539
rect 114 -5573 210 -5539
<< nsubdiffcont >>
rect -114 5539 114 5573
rect -210 -5477 -176 5477
rect 176 -5477 210 5477
rect -114 -5573 114 -5539
<< poly >>
rect -50 5471 50 5487
rect -50 5437 -34 5471
rect 34 5437 50 5471
rect -50 5390 50 5437
rect -50 3743 50 3790
rect -50 3709 -34 3743
rect 34 3709 50 3743
rect -50 3693 50 3709
rect -50 3635 50 3651
rect -50 3601 -34 3635
rect 34 3601 50 3635
rect -50 3554 50 3601
rect -50 1907 50 1954
rect -50 1873 -34 1907
rect 34 1873 50 1907
rect -50 1857 50 1873
rect -50 1799 50 1815
rect -50 1765 -34 1799
rect 34 1765 50 1799
rect -50 1718 50 1765
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -1765 50 -1718
rect -50 -1799 -34 -1765
rect 34 -1799 50 -1765
rect -50 -1815 50 -1799
rect -50 -1873 50 -1857
rect -50 -1907 -34 -1873
rect 34 -1907 50 -1873
rect -50 -1954 50 -1907
rect -50 -3601 50 -3554
rect -50 -3635 -34 -3601
rect 34 -3635 50 -3601
rect -50 -3651 50 -3635
rect -50 -3709 50 -3693
rect -50 -3743 -34 -3709
rect 34 -3743 50 -3709
rect -50 -3790 50 -3743
rect -50 -5437 50 -5390
rect -50 -5471 -34 -5437
rect 34 -5471 50 -5437
rect -50 -5487 50 -5471
<< polycont >>
rect -34 5437 34 5471
rect -34 3709 34 3743
rect -34 3601 34 3635
rect -34 1873 34 1907
rect -34 1765 34 1799
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1799 34 -1765
rect -34 -1907 34 -1873
rect -34 -3635 34 -3601
rect -34 -3743 34 -3709
rect -34 -5471 34 -5437
<< locali >>
rect -210 5539 -114 5573
rect 114 5539 210 5573
rect -210 5477 -176 5539
rect 176 5477 210 5539
rect -50 5437 -34 5471
rect 34 5437 50 5471
rect -96 5378 -62 5394
rect -96 3786 -62 3802
rect 62 5378 96 5394
rect 62 3786 96 3802
rect -50 3709 -34 3743
rect 34 3709 50 3743
rect -50 3601 -34 3635
rect 34 3601 50 3635
rect -96 3542 -62 3558
rect -96 1950 -62 1966
rect 62 3542 96 3558
rect 62 1950 96 1966
rect -50 1873 -34 1907
rect 34 1873 50 1907
rect -50 1765 -34 1799
rect 34 1765 50 1799
rect -96 1706 -62 1722
rect -96 114 -62 130
rect 62 1706 96 1722
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -1722 -62 -1706
rect 62 -130 96 -114
rect 62 -1722 96 -1706
rect -50 -1799 -34 -1765
rect 34 -1799 50 -1765
rect -50 -1907 -34 -1873
rect 34 -1907 50 -1873
rect -96 -1966 -62 -1950
rect -96 -3558 -62 -3542
rect 62 -1966 96 -1950
rect 62 -3558 96 -3542
rect -50 -3635 -34 -3601
rect 34 -3635 50 -3601
rect -50 -3743 -34 -3709
rect 34 -3743 50 -3709
rect -96 -3802 -62 -3786
rect -96 -5394 -62 -5378
rect 62 -3802 96 -3786
rect 62 -5394 96 -5378
rect -50 -5471 -34 -5437
rect 34 -5471 50 -5437
rect -210 -5539 -176 -5477
rect 176 -5539 210 -5477
rect -210 -5573 -114 -5539
rect 114 -5573 210 -5539
<< viali >>
rect -34 5437 34 5471
rect -96 3802 -62 5378
rect 62 3802 96 5378
rect -34 3709 34 3743
rect -34 3601 34 3635
rect -96 1966 -62 3542
rect 62 1966 96 3542
rect -34 1873 34 1907
rect -34 1765 34 1799
rect -96 130 -62 1706
rect 62 130 96 1706
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1706 -62 -130
rect 62 -1706 96 -130
rect -34 -1799 34 -1765
rect -34 -1907 34 -1873
rect -96 -3542 -62 -1966
rect 62 -3542 96 -1966
rect -34 -3635 34 -3601
rect -34 -3743 34 -3709
rect -96 -5378 -62 -3802
rect 62 -5378 96 -3802
rect -34 -5471 34 -5437
<< metal1 >>
rect -46 5471 46 5477
rect -46 5437 -34 5471
rect 34 5437 46 5471
rect -46 5431 46 5437
rect -102 5378 -56 5390
rect -102 3802 -96 5378
rect -62 3802 -56 5378
rect -102 3790 -56 3802
rect 56 5378 102 5390
rect 56 3802 62 5378
rect 96 3802 102 5378
rect 56 3790 102 3802
rect -46 3743 46 3749
rect -46 3709 -34 3743
rect 34 3709 46 3743
rect -46 3703 46 3709
rect -46 3635 46 3641
rect -46 3601 -34 3635
rect 34 3601 46 3635
rect -46 3595 46 3601
rect -102 3542 -56 3554
rect -102 1966 -96 3542
rect -62 1966 -56 3542
rect -102 1954 -56 1966
rect 56 3542 102 3554
rect 56 1966 62 3542
rect 96 1966 102 3542
rect 56 1954 102 1966
rect -46 1907 46 1913
rect -46 1873 -34 1907
rect 34 1873 46 1907
rect -46 1867 46 1873
rect -46 1799 46 1805
rect -46 1765 -34 1799
rect 34 1765 46 1799
rect -46 1759 46 1765
rect -102 1706 -56 1718
rect -102 130 -96 1706
rect -62 130 -56 1706
rect -102 118 -56 130
rect 56 1706 102 1718
rect 56 130 62 1706
rect 96 130 102 1706
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -1706 -96 -130
rect -62 -1706 -56 -130
rect -102 -1718 -56 -1706
rect 56 -130 102 -118
rect 56 -1706 62 -130
rect 96 -1706 102 -130
rect 56 -1718 102 -1706
rect -46 -1765 46 -1759
rect -46 -1799 -34 -1765
rect 34 -1799 46 -1765
rect -46 -1805 46 -1799
rect -46 -1873 46 -1867
rect -46 -1907 -34 -1873
rect 34 -1907 46 -1873
rect -46 -1913 46 -1907
rect -102 -1966 -56 -1954
rect -102 -3542 -96 -1966
rect -62 -3542 -56 -1966
rect -102 -3554 -56 -3542
rect 56 -1966 102 -1954
rect 56 -3542 62 -1966
rect 96 -3542 102 -1966
rect 56 -3554 102 -3542
rect -46 -3601 46 -3595
rect -46 -3635 -34 -3601
rect 34 -3635 46 -3601
rect -46 -3641 46 -3635
rect -46 -3709 46 -3703
rect -46 -3743 -34 -3709
rect 34 -3743 46 -3709
rect -46 -3749 46 -3743
rect -102 -3802 -56 -3790
rect -102 -5378 -96 -3802
rect -62 -5378 -56 -3802
rect -102 -5390 -56 -5378
rect 56 -3802 102 -3790
rect 56 -5378 62 -3802
rect 96 -5378 102 -3802
rect 56 -5390 102 -5378
rect -46 -5437 46 -5431
rect -46 -5471 -34 -5437
rect 34 -5471 46 -5437
rect -46 -5477 46 -5471
<< properties >>
string FIXED_BBOX -193 -5556 193 5556
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
