magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< error_p >>
rect -372 2835 -314 2841
rect -176 2835 -118 2841
rect 20 2835 78 2841
rect 216 2835 274 2841
rect -372 2801 -360 2835
rect -176 2801 -164 2835
rect 20 2801 32 2835
rect 216 2801 228 2835
rect -372 2795 -314 2801
rect -176 2795 -118 2801
rect 20 2795 78 2801
rect 216 2795 274 2801
rect -274 1507 -216 1513
rect -78 1507 -20 1513
rect 118 1507 176 1513
rect 314 1507 372 1513
rect -274 1473 -262 1507
rect -78 1473 -66 1507
rect 118 1473 130 1507
rect 314 1473 326 1507
rect -274 1467 -216 1473
rect -78 1467 -20 1473
rect 118 1467 176 1473
rect 314 1467 372 1473
rect -274 1399 -216 1405
rect -78 1399 -20 1405
rect 118 1399 176 1405
rect 314 1399 372 1405
rect -274 1365 -262 1399
rect -78 1365 -66 1399
rect 118 1365 130 1399
rect 314 1365 326 1399
rect -274 1359 -216 1365
rect -78 1359 -20 1365
rect 118 1359 176 1365
rect 314 1359 372 1365
rect -372 71 -314 77
rect -176 71 -118 77
rect 20 71 78 77
rect 216 71 274 77
rect -372 37 -360 71
rect -176 37 -164 71
rect 20 37 32 71
rect 216 37 228 71
rect -372 31 -314 37
rect -176 31 -118 37
rect 20 31 78 37
rect 216 31 274 37
rect -372 -37 -314 -31
rect -176 -37 -118 -31
rect 20 -37 78 -31
rect 216 -37 274 -31
rect -372 -71 -360 -37
rect -176 -71 -164 -37
rect 20 -71 32 -37
rect 216 -71 228 -37
rect -372 -77 -314 -71
rect -176 -77 -118 -71
rect 20 -77 78 -71
rect 216 -77 274 -71
rect -274 -1365 -216 -1359
rect -78 -1365 -20 -1359
rect 118 -1365 176 -1359
rect 314 -1365 372 -1359
rect -274 -1399 -262 -1365
rect -78 -1399 -66 -1365
rect 118 -1399 130 -1365
rect 314 -1399 326 -1365
rect -274 -1405 -216 -1399
rect -78 -1405 -20 -1399
rect 118 -1405 176 -1399
rect 314 -1405 372 -1399
rect -274 -1473 -216 -1467
rect -78 -1473 -20 -1467
rect 118 -1473 176 -1467
rect 314 -1473 372 -1467
rect -274 -1507 -262 -1473
rect -78 -1507 -66 -1473
rect 118 -1507 130 -1473
rect 314 -1507 326 -1473
rect -274 -1513 -216 -1507
rect -78 -1513 -20 -1507
rect 118 -1513 176 -1507
rect 314 -1513 372 -1507
rect -372 -2801 -314 -2795
rect -176 -2801 -118 -2795
rect 20 -2801 78 -2795
rect 216 -2801 274 -2795
rect -372 -2835 -360 -2801
rect -176 -2835 -164 -2801
rect 20 -2835 32 -2801
rect 216 -2835 228 -2801
rect -372 -2841 -314 -2835
rect -176 -2841 -118 -2835
rect 20 -2841 78 -2835
rect 216 -2841 274 -2835
<< nwell >>
rect -559 -2973 559 2973
<< pmos >>
rect -363 1554 -323 2754
rect -265 1554 -225 2754
rect -167 1554 -127 2754
rect -69 1554 -29 2754
rect 29 1554 69 2754
rect 127 1554 167 2754
rect 225 1554 265 2754
rect 323 1554 363 2754
rect -363 118 -323 1318
rect -265 118 -225 1318
rect -167 118 -127 1318
rect -69 118 -29 1318
rect 29 118 69 1318
rect 127 118 167 1318
rect 225 118 265 1318
rect 323 118 363 1318
rect -363 -1318 -323 -118
rect -265 -1318 -225 -118
rect -167 -1318 -127 -118
rect -69 -1318 -29 -118
rect 29 -1318 69 -118
rect 127 -1318 167 -118
rect 225 -1318 265 -118
rect 323 -1318 363 -118
rect -363 -2754 -323 -1554
rect -265 -2754 -225 -1554
rect -167 -2754 -127 -1554
rect -69 -2754 -29 -1554
rect 29 -2754 69 -1554
rect 127 -2754 167 -1554
rect 225 -2754 265 -1554
rect 323 -2754 363 -1554
<< pdiff >>
rect -421 2742 -363 2754
rect -421 1566 -409 2742
rect -375 1566 -363 2742
rect -421 1554 -363 1566
rect -323 2742 -265 2754
rect -323 1566 -311 2742
rect -277 1566 -265 2742
rect -323 1554 -265 1566
rect -225 2742 -167 2754
rect -225 1566 -213 2742
rect -179 1566 -167 2742
rect -225 1554 -167 1566
rect -127 2742 -69 2754
rect -127 1566 -115 2742
rect -81 1566 -69 2742
rect -127 1554 -69 1566
rect -29 2742 29 2754
rect -29 1566 -17 2742
rect 17 1566 29 2742
rect -29 1554 29 1566
rect 69 2742 127 2754
rect 69 1566 81 2742
rect 115 1566 127 2742
rect 69 1554 127 1566
rect 167 2742 225 2754
rect 167 1566 179 2742
rect 213 1566 225 2742
rect 167 1554 225 1566
rect 265 2742 323 2754
rect 265 1566 277 2742
rect 311 1566 323 2742
rect 265 1554 323 1566
rect 363 2742 421 2754
rect 363 1566 375 2742
rect 409 1566 421 2742
rect 363 1554 421 1566
rect -421 1306 -363 1318
rect -421 130 -409 1306
rect -375 130 -363 1306
rect -421 118 -363 130
rect -323 1306 -265 1318
rect -323 130 -311 1306
rect -277 130 -265 1306
rect -323 118 -265 130
rect -225 1306 -167 1318
rect -225 130 -213 1306
rect -179 130 -167 1306
rect -225 118 -167 130
rect -127 1306 -69 1318
rect -127 130 -115 1306
rect -81 130 -69 1306
rect -127 118 -69 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 69 1306 127 1318
rect 69 130 81 1306
rect 115 130 127 1306
rect 69 118 127 130
rect 167 1306 225 1318
rect 167 130 179 1306
rect 213 130 225 1306
rect 167 118 225 130
rect 265 1306 323 1318
rect 265 130 277 1306
rect 311 130 323 1306
rect 265 118 323 130
rect 363 1306 421 1318
rect 363 130 375 1306
rect 409 130 421 1306
rect 363 118 421 130
rect -421 -130 -363 -118
rect -421 -1306 -409 -130
rect -375 -1306 -363 -130
rect -421 -1318 -363 -1306
rect -323 -130 -265 -118
rect -323 -1306 -311 -130
rect -277 -1306 -265 -130
rect -323 -1318 -265 -1306
rect -225 -130 -167 -118
rect -225 -1306 -213 -130
rect -179 -1306 -167 -130
rect -225 -1318 -167 -1306
rect -127 -130 -69 -118
rect -127 -1306 -115 -130
rect -81 -1306 -69 -130
rect -127 -1318 -69 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 69 -130 127 -118
rect 69 -1306 81 -130
rect 115 -1306 127 -130
rect 69 -1318 127 -1306
rect 167 -130 225 -118
rect 167 -1306 179 -130
rect 213 -1306 225 -130
rect 167 -1318 225 -1306
rect 265 -130 323 -118
rect 265 -1306 277 -130
rect 311 -1306 323 -130
rect 265 -1318 323 -1306
rect 363 -130 421 -118
rect 363 -1306 375 -130
rect 409 -1306 421 -130
rect 363 -1318 421 -1306
rect -421 -1566 -363 -1554
rect -421 -2742 -409 -1566
rect -375 -2742 -363 -1566
rect -421 -2754 -363 -2742
rect -323 -1566 -265 -1554
rect -323 -2742 -311 -1566
rect -277 -2742 -265 -1566
rect -323 -2754 -265 -2742
rect -225 -1566 -167 -1554
rect -225 -2742 -213 -1566
rect -179 -2742 -167 -1566
rect -225 -2754 -167 -2742
rect -127 -1566 -69 -1554
rect -127 -2742 -115 -1566
rect -81 -2742 -69 -1566
rect -127 -2754 -69 -2742
rect -29 -1566 29 -1554
rect -29 -2742 -17 -1566
rect 17 -2742 29 -1566
rect -29 -2754 29 -2742
rect 69 -1566 127 -1554
rect 69 -2742 81 -1566
rect 115 -2742 127 -1566
rect 69 -2754 127 -2742
rect 167 -1566 225 -1554
rect 167 -2742 179 -1566
rect 213 -2742 225 -1566
rect 167 -2754 225 -2742
rect 265 -1566 323 -1554
rect 265 -2742 277 -1566
rect 311 -2742 323 -1566
rect 265 -2754 323 -2742
rect 363 -1566 421 -1554
rect 363 -2742 375 -1566
rect 409 -2742 421 -1566
rect 363 -2754 421 -2742
<< pdiffc >>
rect -409 1566 -375 2742
rect -311 1566 -277 2742
rect -213 1566 -179 2742
rect -115 1566 -81 2742
rect -17 1566 17 2742
rect 81 1566 115 2742
rect 179 1566 213 2742
rect 277 1566 311 2742
rect 375 1566 409 2742
rect -409 130 -375 1306
rect -311 130 -277 1306
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect 277 130 311 1306
rect 375 130 409 1306
rect -409 -1306 -375 -130
rect -311 -1306 -277 -130
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect 277 -1306 311 -130
rect 375 -1306 409 -130
rect -409 -2742 -375 -1566
rect -311 -2742 -277 -1566
rect -213 -2742 -179 -1566
rect -115 -2742 -81 -1566
rect -17 -2742 17 -1566
rect 81 -2742 115 -1566
rect 179 -2742 213 -1566
rect 277 -2742 311 -1566
rect 375 -2742 409 -1566
<< nsubdiff >>
rect -523 2903 -427 2937
rect 427 2903 523 2937
rect -523 2841 -489 2903
rect 489 2841 523 2903
rect -523 -2903 -489 -2841
rect 489 -2903 523 -2841
rect -523 -2937 -427 -2903
rect 427 -2937 523 -2903
<< nsubdiffcont >>
rect -427 2903 427 2937
rect -523 -2841 -489 2841
rect 489 -2841 523 2841
rect -427 -2937 427 -2903
<< poly >>
rect -376 2835 -310 2851
rect -376 2801 -360 2835
rect -326 2801 -310 2835
rect -376 2785 -310 2801
rect -180 2835 -114 2851
rect -180 2801 -164 2835
rect -130 2801 -114 2835
rect -180 2785 -114 2801
rect 16 2835 82 2851
rect 16 2801 32 2835
rect 66 2801 82 2835
rect 16 2785 82 2801
rect 212 2835 278 2851
rect 212 2801 228 2835
rect 262 2801 278 2835
rect 212 2785 278 2801
rect -363 2754 -323 2785
rect -265 2754 -225 2780
rect -167 2754 -127 2785
rect -69 2754 -29 2780
rect 29 2754 69 2785
rect 127 2754 167 2780
rect 225 2754 265 2785
rect 323 2754 363 2780
rect -363 1528 -323 1554
rect -265 1523 -225 1554
rect -167 1528 -127 1554
rect -69 1523 -29 1554
rect 29 1528 69 1554
rect 127 1523 167 1554
rect 225 1528 265 1554
rect 323 1523 363 1554
rect -278 1507 -212 1523
rect -278 1473 -262 1507
rect -228 1473 -212 1507
rect -278 1457 -212 1473
rect -82 1507 -16 1523
rect -82 1473 -66 1507
rect -32 1473 -16 1507
rect -82 1457 -16 1473
rect 114 1507 180 1523
rect 114 1473 130 1507
rect 164 1473 180 1507
rect 114 1457 180 1473
rect 310 1507 376 1523
rect 310 1473 326 1507
rect 360 1473 376 1507
rect 310 1457 376 1473
rect -278 1399 -212 1415
rect -278 1365 -262 1399
rect -228 1365 -212 1399
rect -278 1349 -212 1365
rect -82 1399 -16 1415
rect -82 1365 -66 1399
rect -32 1365 -16 1399
rect -82 1349 -16 1365
rect 114 1399 180 1415
rect 114 1365 130 1399
rect 164 1365 180 1399
rect 114 1349 180 1365
rect 310 1399 376 1415
rect 310 1365 326 1399
rect 360 1365 376 1399
rect 310 1349 376 1365
rect -363 1318 -323 1344
rect -265 1318 -225 1349
rect -167 1318 -127 1344
rect -69 1318 -29 1349
rect 29 1318 69 1344
rect 127 1318 167 1349
rect 225 1318 265 1344
rect 323 1318 363 1349
rect -363 87 -323 118
rect -265 92 -225 118
rect -167 87 -127 118
rect -69 92 -29 118
rect 29 87 69 118
rect 127 92 167 118
rect 225 87 265 118
rect 323 92 363 118
rect -376 71 -310 87
rect -376 37 -360 71
rect -326 37 -310 71
rect -376 21 -310 37
rect -180 71 -114 87
rect -180 37 -164 71
rect -130 37 -114 71
rect -180 21 -114 37
rect 16 71 82 87
rect 16 37 32 71
rect 66 37 82 71
rect 16 21 82 37
rect 212 71 278 87
rect 212 37 228 71
rect 262 37 278 71
rect 212 21 278 37
rect -376 -37 -310 -21
rect -376 -71 -360 -37
rect -326 -71 -310 -37
rect -376 -87 -310 -71
rect -180 -37 -114 -21
rect -180 -71 -164 -37
rect -130 -71 -114 -37
rect -180 -87 -114 -71
rect 16 -37 82 -21
rect 16 -71 32 -37
rect 66 -71 82 -37
rect 16 -87 82 -71
rect 212 -37 278 -21
rect 212 -71 228 -37
rect 262 -71 278 -37
rect 212 -87 278 -71
rect -363 -118 -323 -87
rect -265 -118 -225 -92
rect -167 -118 -127 -87
rect -69 -118 -29 -92
rect 29 -118 69 -87
rect 127 -118 167 -92
rect 225 -118 265 -87
rect 323 -118 363 -92
rect -363 -1344 -323 -1318
rect -265 -1349 -225 -1318
rect -167 -1344 -127 -1318
rect -69 -1349 -29 -1318
rect 29 -1344 69 -1318
rect 127 -1349 167 -1318
rect 225 -1344 265 -1318
rect 323 -1349 363 -1318
rect -278 -1365 -212 -1349
rect -278 -1399 -262 -1365
rect -228 -1399 -212 -1365
rect -278 -1415 -212 -1399
rect -82 -1365 -16 -1349
rect -82 -1399 -66 -1365
rect -32 -1399 -16 -1365
rect -82 -1415 -16 -1399
rect 114 -1365 180 -1349
rect 114 -1399 130 -1365
rect 164 -1399 180 -1365
rect 114 -1415 180 -1399
rect 310 -1365 376 -1349
rect 310 -1399 326 -1365
rect 360 -1399 376 -1365
rect 310 -1415 376 -1399
rect -278 -1473 -212 -1457
rect -278 -1507 -262 -1473
rect -228 -1507 -212 -1473
rect -278 -1523 -212 -1507
rect -82 -1473 -16 -1457
rect -82 -1507 -66 -1473
rect -32 -1507 -16 -1473
rect -82 -1523 -16 -1507
rect 114 -1473 180 -1457
rect 114 -1507 130 -1473
rect 164 -1507 180 -1473
rect 114 -1523 180 -1507
rect 310 -1473 376 -1457
rect 310 -1507 326 -1473
rect 360 -1507 376 -1473
rect 310 -1523 376 -1507
rect -363 -1554 -323 -1528
rect -265 -1554 -225 -1523
rect -167 -1554 -127 -1528
rect -69 -1554 -29 -1523
rect 29 -1554 69 -1528
rect 127 -1554 167 -1523
rect 225 -1554 265 -1528
rect 323 -1554 363 -1523
rect -363 -2785 -323 -2754
rect -265 -2780 -225 -2754
rect -167 -2785 -127 -2754
rect -69 -2780 -29 -2754
rect 29 -2785 69 -2754
rect 127 -2780 167 -2754
rect 225 -2785 265 -2754
rect 323 -2780 363 -2754
rect -376 -2801 -310 -2785
rect -376 -2835 -360 -2801
rect -326 -2835 -310 -2801
rect -376 -2851 -310 -2835
rect -180 -2801 -114 -2785
rect -180 -2835 -164 -2801
rect -130 -2835 -114 -2801
rect -180 -2851 -114 -2835
rect 16 -2801 82 -2785
rect 16 -2835 32 -2801
rect 66 -2835 82 -2801
rect 16 -2851 82 -2835
rect 212 -2801 278 -2785
rect 212 -2835 228 -2801
rect 262 -2835 278 -2801
rect 212 -2851 278 -2835
<< polycont >>
rect -360 2801 -326 2835
rect -164 2801 -130 2835
rect 32 2801 66 2835
rect 228 2801 262 2835
rect -262 1473 -228 1507
rect -66 1473 -32 1507
rect 130 1473 164 1507
rect 326 1473 360 1507
rect -262 1365 -228 1399
rect -66 1365 -32 1399
rect 130 1365 164 1399
rect 326 1365 360 1399
rect -360 37 -326 71
rect -164 37 -130 71
rect 32 37 66 71
rect 228 37 262 71
rect -360 -71 -326 -37
rect -164 -71 -130 -37
rect 32 -71 66 -37
rect 228 -71 262 -37
rect -262 -1399 -228 -1365
rect -66 -1399 -32 -1365
rect 130 -1399 164 -1365
rect 326 -1399 360 -1365
rect -262 -1507 -228 -1473
rect -66 -1507 -32 -1473
rect 130 -1507 164 -1473
rect 326 -1507 360 -1473
rect -360 -2835 -326 -2801
rect -164 -2835 -130 -2801
rect 32 -2835 66 -2801
rect 228 -2835 262 -2801
<< locali >>
rect -523 2903 -427 2937
rect 427 2903 523 2937
rect -523 2841 -489 2903
rect 489 2841 523 2903
rect -376 2801 -360 2835
rect -326 2801 -310 2835
rect -180 2801 -164 2835
rect -130 2801 -114 2835
rect 16 2801 32 2835
rect 66 2801 82 2835
rect 212 2801 228 2835
rect 262 2801 278 2835
rect -409 2742 -375 2758
rect -409 1550 -375 1566
rect -311 2742 -277 2758
rect -311 1550 -277 1566
rect -213 2742 -179 2758
rect -213 1550 -179 1566
rect -115 2742 -81 2758
rect -115 1550 -81 1566
rect -17 2742 17 2758
rect -17 1550 17 1566
rect 81 2742 115 2758
rect 81 1550 115 1566
rect 179 2742 213 2758
rect 179 1550 213 1566
rect 277 2742 311 2758
rect 277 1550 311 1566
rect 375 2742 409 2758
rect 375 1550 409 1566
rect -278 1473 -262 1507
rect -228 1473 -212 1507
rect -82 1473 -66 1507
rect -32 1473 -16 1507
rect 114 1473 130 1507
rect 164 1473 180 1507
rect 310 1473 326 1507
rect 360 1473 376 1507
rect -278 1365 -262 1399
rect -228 1365 -212 1399
rect -82 1365 -66 1399
rect -32 1365 -16 1399
rect 114 1365 130 1399
rect 164 1365 180 1399
rect 310 1365 326 1399
rect 360 1365 376 1399
rect -409 1306 -375 1322
rect -409 114 -375 130
rect -311 1306 -277 1322
rect -311 114 -277 130
rect -213 1306 -179 1322
rect -213 114 -179 130
rect -115 1306 -81 1322
rect -115 114 -81 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 81 1306 115 1322
rect 81 114 115 130
rect 179 1306 213 1322
rect 179 114 213 130
rect 277 1306 311 1322
rect 277 114 311 130
rect 375 1306 409 1322
rect 375 114 409 130
rect -376 37 -360 71
rect -326 37 -310 71
rect -180 37 -164 71
rect -130 37 -114 71
rect 16 37 32 71
rect 66 37 82 71
rect 212 37 228 71
rect 262 37 278 71
rect -376 -71 -360 -37
rect -326 -71 -310 -37
rect -180 -71 -164 -37
rect -130 -71 -114 -37
rect 16 -71 32 -37
rect 66 -71 82 -37
rect 212 -71 228 -37
rect 262 -71 278 -37
rect -409 -130 -375 -114
rect -409 -1322 -375 -1306
rect -311 -130 -277 -114
rect -311 -1322 -277 -1306
rect -213 -130 -179 -114
rect -213 -1322 -179 -1306
rect -115 -130 -81 -114
rect -115 -1322 -81 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 81 -130 115 -114
rect 81 -1322 115 -1306
rect 179 -130 213 -114
rect 179 -1322 213 -1306
rect 277 -130 311 -114
rect 277 -1322 311 -1306
rect 375 -130 409 -114
rect 375 -1322 409 -1306
rect -278 -1399 -262 -1365
rect -228 -1399 -212 -1365
rect -82 -1399 -66 -1365
rect -32 -1399 -16 -1365
rect 114 -1399 130 -1365
rect 164 -1399 180 -1365
rect 310 -1399 326 -1365
rect 360 -1399 376 -1365
rect -278 -1507 -262 -1473
rect -228 -1507 -212 -1473
rect -82 -1507 -66 -1473
rect -32 -1507 -16 -1473
rect 114 -1507 130 -1473
rect 164 -1507 180 -1473
rect 310 -1507 326 -1473
rect 360 -1507 376 -1473
rect -409 -1566 -375 -1550
rect -409 -2758 -375 -2742
rect -311 -1566 -277 -1550
rect -311 -2758 -277 -2742
rect -213 -1566 -179 -1550
rect -213 -2758 -179 -2742
rect -115 -1566 -81 -1550
rect -115 -2758 -81 -2742
rect -17 -1566 17 -1550
rect -17 -2758 17 -2742
rect 81 -1566 115 -1550
rect 81 -2758 115 -2742
rect 179 -1566 213 -1550
rect 179 -2758 213 -2742
rect 277 -1566 311 -1550
rect 277 -2758 311 -2742
rect 375 -1566 409 -1550
rect 375 -2758 409 -2742
rect -376 -2835 -360 -2801
rect -326 -2835 -310 -2801
rect -180 -2835 -164 -2801
rect -130 -2835 -114 -2801
rect 16 -2835 32 -2801
rect 66 -2835 82 -2801
rect 212 -2835 228 -2801
rect 262 -2835 278 -2801
rect -523 -2903 -489 -2841
rect 489 -2903 523 -2841
rect -523 -2937 -427 -2903
rect 427 -2937 523 -2903
<< viali >>
rect -360 2801 -326 2835
rect -164 2801 -130 2835
rect 32 2801 66 2835
rect 228 2801 262 2835
rect -409 1566 -375 2742
rect -311 1566 -277 2742
rect -213 1566 -179 2742
rect -115 1566 -81 2742
rect -17 1566 17 2742
rect 81 1566 115 2742
rect 179 1566 213 2742
rect 277 1566 311 2742
rect 375 1566 409 2742
rect -262 1473 -228 1507
rect -66 1473 -32 1507
rect 130 1473 164 1507
rect 326 1473 360 1507
rect -262 1365 -228 1399
rect -66 1365 -32 1399
rect 130 1365 164 1399
rect 326 1365 360 1399
rect -409 130 -375 1306
rect -311 130 -277 1306
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect 277 130 311 1306
rect 375 130 409 1306
rect -360 37 -326 71
rect -164 37 -130 71
rect 32 37 66 71
rect 228 37 262 71
rect -360 -71 -326 -37
rect -164 -71 -130 -37
rect 32 -71 66 -37
rect 228 -71 262 -37
rect -409 -1306 -375 -130
rect -311 -1306 -277 -130
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect 277 -1306 311 -130
rect 375 -1306 409 -130
rect -262 -1399 -228 -1365
rect -66 -1399 -32 -1365
rect 130 -1399 164 -1365
rect 326 -1399 360 -1365
rect -262 -1507 -228 -1473
rect -66 -1507 -32 -1473
rect 130 -1507 164 -1473
rect 326 -1507 360 -1473
rect -409 -2742 -375 -1566
rect -311 -2742 -277 -1566
rect -213 -2742 -179 -1566
rect -115 -2742 -81 -1566
rect -17 -2742 17 -1566
rect 81 -2742 115 -1566
rect 179 -2742 213 -1566
rect 277 -2742 311 -1566
rect 375 -2742 409 -1566
rect -360 -2835 -326 -2801
rect -164 -2835 -130 -2801
rect 32 -2835 66 -2801
rect 228 -2835 262 -2801
<< metal1 >>
rect -372 2835 -314 2841
rect -372 2801 -360 2835
rect -326 2801 -314 2835
rect -372 2795 -314 2801
rect -176 2835 -118 2841
rect -176 2801 -164 2835
rect -130 2801 -118 2835
rect -176 2795 -118 2801
rect 20 2835 78 2841
rect 20 2801 32 2835
rect 66 2801 78 2835
rect 20 2795 78 2801
rect 216 2835 274 2841
rect 216 2801 228 2835
rect 262 2801 274 2835
rect 216 2795 274 2801
rect -415 2742 -369 2754
rect -415 1566 -409 2742
rect -375 1566 -369 2742
rect -415 1554 -369 1566
rect -317 2742 -271 2754
rect -317 1566 -311 2742
rect -277 1566 -271 2742
rect -317 1554 -271 1566
rect -219 2742 -173 2754
rect -219 1566 -213 2742
rect -179 1566 -173 2742
rect -219 1554 -173 1566
rect -121 2742 -75 2754
rect -121 1566 -115 2742
rect -81 1566 -75 2742
rect -121 1554 -75 1566
rect -23 2742 23 2754
rect -23 1566 -17 2742
rect 17 1566 23 2742
rect -23 1554 23 1566
rect 75 2742 121 2754
rect 75 1566 81 2742
rect 115 1566 121 2742
rect 75 1554 121 1566
rect 173 2742 219 2754
rect 173 1566 179 2742
rect 213 1566 219 2742
rect 173 1554 219 1566
rect 271 2742 317 2754
rect 271 1566 277 2742
rect 311 1566 317 2742
rect 271 1554 317 1566
rect 369 2742 415 2754
rect 369 1566 375 2742
rect 409 1566 415 2742
rect 369 1554 415 1566
rect -274 1507 -216 1513
rect -274 1473 -262 1507
rect -228 1473 -216 1507
rect -274 1467 -216 1473
rect -78 1507 -20 1513
rect -78 1473 -66 1507
rect -32 1473 -20 1507
rect -78 1467 -20 1473
rect 118 1507 176 1513
rect 118 1473 130 1507
rect 164 1473 176 1507
rect 118 1467 176 1473
rect 314 1507 372 1513
rect 314 1473 326 1507
rect 360 1473 372 1507
rect 314 1467 372 1473
rect -274 1399 -216 1405
rect -274 1365 -262 1399
rect -228 1365 -216 1399
rect -274 1359 -216 1365
rect -78 1399 -20 1405
rect -78 1365 -66 1399
rect -32 1365 -20 1399
rect -78 1359 -20 1365
rect 118 1399 176 1405
rect 118 1365 130 1399
rect 164 1365 176 1399
rect 118 1359 176 1365
rect 314 1399 372 1405
rect 314 1365 326 1399
rect 360 1365 372 1399
rect 314 1359 372 1365
rect -415 1306 -369 1318
rect -415 130 -409 1306
rect -375 130 -369 1306
rect -415 118 -369 130
rect -317 1306 -271 1318
rect -317 130 -311 1306
rect -277 130 -271 1306
rect -317 118 -271 130
rect -219 1306 -173 1318
rect -219 130 -213 1306
rect -179 130 -173 1306
rect -219 118 -173 130
rect -121 1306 -75 1318
rect -121 130 -115 1306
rect -81 130 -75 1306
rect -121 118 -75 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 75 1306 121 1318
rect 75 130 81 1306
rect 115 130 121 1306
rect 75 118 121 130
rect 173 1306 219 1318
rect 173 130 179 1306
rect 213 130 219 1306
rect 173 118 219 130
rect 271 1306 317 1318
rect 271 130 277 1306
rect 311 130 317 1306
rect 271 118 317 130
rect 369 1306 415 1318
rect 369 130 375 1306
rect 409 130 415 1306
rect 369 118 415 130
rect -372 71 -314 77
rect -372 37 -360 71
rect -326 37 -314 71
rect -372 31 -314 37
rect -176 71 -118 77
rect -176 37 -164 71
rect -130 37 -118 71
rect -176 31 -118 37
rect 20 71 78 77
rect 20 37 32 71
rect 66 37 78 71
rect 20 31 78 37
rect 216 71 274 77
rect 216 37 228 71
rect 262 37 274 71
rect 216 31 274 37
rect -372 -37 -314 -31
rect -372 -71 -360 -37
rect -326 -71 -314 -37
rect -372 -77 -314 -71
rect -176 -37 -118 -31
rect -176 -71 -164 -37
rect -130 -71 -118 -37
rect -176 -77 -118 -71
rect 20 -37 78 -31
rect 20 -71 32 -37
rect 66 -71 78 -37
rect 20 -77 78 -71
rect 216 -37 274 -31
rect 216 -71 228 -37
rect 262 -71 274 -37
rect 216 -77 274 -71
rect -415 -130 -369 -118
rect -415 -1306 -409 -130
rect -375 -1306 -369 -130
rect -415 -1318 -369 -1306
rect -317 -130 -271 -118
rect -317 -1306 -311 -130
rect -277 -1306 -271 -130
rect -317 -1318 -271 -1306
rect -219 -130 -173 -118
rect -219 -1306 -213 -130
rect -179 -1306 -173 -130
rect -219 -1318 -173 -1306
rect -121 -130 -75 -118
rect -121 -1306 -115 -130
rect -81 -1306 -75 -130
rect -121 -1318 -75 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 75 -130 121 -118
rect 75 -1306 81 -130
rect 115 -1306 121 -130
rect 75 -1318 121 -1306
rect 173 -130 219 -118
rect 173 -1306 179 -130
rect 213 -1306 219 -130
rect 173 -1318 219 -1306
rect 271 -130 317 -118
rect 271 -1306 277 -130
rect 311 -1306 317 -130
rect 271 -1318 317 -1306
rect 369 -130 415 -118
rect 369 -1306 375 -130
rect 409 -1306 415 -130
rect 369 -1318 415 -1306
rect -274 -1365 -216 -1359
rect -274 -1399 -262 -1365
rect -228 -1399 -216 -1365
rect -274 -1405 -216 -1399
rect -78 -1365 -20 -1359
rect -78 -1399 -66 -1365
rect -32 -1399 -20 -1365
rect -78 -1405 -20 -1399
rect 118 -1365 176 -1359
rect 118 -1399 130 -1365
rect 164 -1399 176 -1365
rect 118 -1405 176 -1399
rect 314 -1365 372 -1359
rect 314 -1399 326 -1365
rect 360 -1399 372 -1365
rect 314 -1405 372 -1399
rect -274 -1473 -216 -1467
rect -274 -1507 -262 -1473
rect -228 -1507 -216 -1473
rect -274 -1513 -216 -1507
rect -78 -1473 -20 -1467
rect -78 -1507 -66 -1473
rect -32 -1507 -20 -1473
rect -78 -1513 -20 -1507
rect 118 -1473 176 -1467
rect 118 -1507 130 -1473
rect 164 -1507 176 -1473
rect 118 -1513 176 -1507
rect 314 -1473 372 -1467
rect 314 -1507 326 -1473
rect 360 -1507 372 -1473
rect 314 -1513 372 -1507
rect -415 -1566 -369 -1554
rect -415 -2742 -409 -1566
rect -375 -2742 -369 -1566
rect -415 -2754 -369 -2742
rect -317 -1566 -271 -1554
rect -317 -2742 -311 -1566
rect -277 -2742 -271 -1566
rect -317 -2754 -271 -2742
rect -219 -1566 -173 -1554
rect -219 -2742 -213 -1566
rect -179 -2742 -173 -1566
rect -219 -2754 -173 -2742
rect -121 -1566 -75 -1554
rect -121 -2742 -115 -1566
rect -81 -2742 -75 -1566
rect -121 -2754 -75 -2742
rect -23 -1566 23 -1554
rect -23 -2742 -17 -1566
rect 17 -2742 23 -1566
rect -23 -2754 23 -2742
rect 75 -1566 121 -1554
rect 75 -2742 81 -1566
rect 115 -2742 121 -1566
rect 75 -2754 121 -2742
rect 173 -1566 219 -1554
rect 173 -2742 179 -1566
rect 213 -2742 219 -1566
rect 173 -2754 219 -2742
rect 271 -1566 317 -1554
rect 271 -2742 277 -1566
rect 311 -2742 317 -1566
rect 271 -2754 317 -2742
rect 369 -1566 415 -1554
rect 369 -2742 375 -1566
rect 409 -2742 415 -1566
rect 369 -2754 415 -2742
rect -372 -2801 -314 -2795
rect -372 -2835 -360 -2801
rect -326 -2835 -314 -2801
rect -372 -2841 -314 -2835
rect -176 -2801 -118 -2795
rect -176 -2835 -164 -2801
rect -130 -2835 -118 -2801
rect -176 -2841 -118 -2835
rect 20 -2801 78 -2795
rect 20 -2835 32 -2801
rect 66 -2835 78 -2801
rect 20 -2841 78 -2835
rect 216 -2801 274 -2795
rect 216 -2835 228 -2801
rect 262 -2835 274 -2801
rect 216 -2841 274 -2835
<< properties >>
string FIXED_BBOX -506 -2920 506 2920
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.2 m 4 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
