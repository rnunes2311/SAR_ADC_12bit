magic
tech sky130A
magscale 1 2
timestamp 1711984062
<< nwell >>
rect 5524 978 6894 986
rect 5524 657 7668 978
rect 5524 135 6894 657
rect 5524 -252 7668 135
rect 7040 -431 7668 -252
<< pwell >>
rect 6936 417 7122 599
rect 7181 417 7619 599
rect 6936 413 6957 417
rect 6923 379 6957 413
rect 6936 375 6957 379
rect 7199 375 7233 417
rect 6936 193 7122 375
rect 7181 193 7619 375
rect 5523 -872 6893 -252
rect 7107 -671 7629 -489
rect 7566 -709 7600 -671
rect 5523 -966 5945 -872
rect 6471 -966 6893 -872
rect 5523 -1072 6893 -966
rect 5686 -1586 6746 -1072
<< nmos >>
rect 5719 -862 5749 -462
rect 6035 -662 6065 -462
rect 6351 -662 6381 -462
rect 6667 -862 6697 -462
<< scnmos >>
rect 7014 443 7044 573
rect 7259 443 7289 573
rect 7343 443 7373 573
rect 7427 443 7457 573
rect 7511 443 7541 573
rect 7014 219 7044 349
rect 7259 219 7289 349
rect 7343 219 7373 349
rect 7427 219 7457 349
rect 7511 219 7541 349
rect 7185 -645 7215 -515
rect 7269 -645 7299 -515
rect 7353 -645 7383 -515
rect 7437 -645 7467 -515
rect 7521 -645 7551 -515
<< pmos >>
rect 5720 567 5750 767
rect 5720 -33 5750 167
rect 6036 -33 6066 767
rect 6352 -33 6382 767
rect 6668 567 6698 767
rect 6668 -33 6698 167
<< scpmoshvt >>
rect 7014 693 7044 893
rect 7259 693 7289 893
rect 7343 693 7373 893
rect 7427 693 7457 893
rect 7511 693 7541 893
rect 7014 -101 7044 99
rect 7259 -101 7289 99
rect 7343 -101 7373 99
rect 7427 -101 7457 99
rect 7511 -101 7541 99
rect 7185 -395 7215 -195
rect 7269 -395 7299 -195
rect 7353 -395 7383 -195
rect 7437 -395 7467 -195
rect 7521 -395 7551 -195
<< nmoslvt >>
rect 5886 -1376 5916 -1176
rect 6096 -1376 6126 -1176
rect 6306 -1376 6336 -1176
rect 6516 -1376 6546 -1176
<< ndiff >>
rect 6962 561 7014 573
rect 6962 527 6970 561
rect 7004 527 7014 561
rect 6962 493 7014 527
rect 6962 459 6970 493
rect 7004 459 7014 493
rect 6962 443 7014 459
rect 7044 561 7096 573
rect 7044 527 7054 561
rect 7088 527 7096 561
rect 7044 493 7096 527
rect 7044 459 7054 493
rect 7088 459 7096 493
rect 7044 443 7096 459
rect 7207 489 7259 573
rect 7207 455 7215 489
rect 7249 455 7259 489
rect 7207 443 7259 455
rect 7289 497 7343 573
rect 7289 463 7299 497
rect 7333 463 7343 497
rect 7289 443 7343 463
rect 7373 489 7427 573
rect 7373 455 7383 489
rect 7417 455 7427 489
rect 7373 443 7427 455
rect 7457 497 7511 573
rect 7457 463 7467 497
rect 7501 463 7511 497
rect 7457 443 7511 463
rect 7541 490 7593 573
rect 7541 456 7551 490
rect 7585 456 7593 490
rect 7541 443 7593 456
rect 6962 333 7014 349
rect 6962 299 6970 333
rect 7004 299 7014 333
rect 6962 265 7014 299
rect 6962 231 6970 265
rect 7004 231 7014 265
rect 6962 219 7014 231
rect 7044 333 7096 349
rect 7044 299 7054 333
rect 7088 299 7096 333
rect 7044 265 7096 299
rect 7044 231 7054 265
rect 7088 231 7096 265
rect 7044 219 7096 231
rect 7207 337 7259 349
rect 7207 303 7215 337
rect 7249 303 7259 337
rect 7207 219 7259 303
rect 7289 329 7343 349
rect 7289 295 7299 329
rect 7333 295 7343 329
rect 7289 219 7343 295
rect 7373 337 7427 349
rect 7373 303 7383 337
rect 7417 303 7427 337
rect 7373 219 7427 303
rect 7457 329 7511 349
rect 7457 295 7467 329
rect 7501 295 7511 329
rect 7457 219 7511 295
rect 7541 336 7593 349
rect 7541 302 7551 336
rect 7585 302 7593 336
rect 7541 219 7593 302
rect 5661 -474 5719 -462
rect 5661 -850 5673 -474
rect 5707 -850 5719 -474
rect 5661 -862 5719 -850
rect 5749 -474 5807 -462
rect 5749 -850 5761 -474
rect 5795 -850 5807 -474
rect 5749 -862 5807 -850
rect 5977 -474 6035 -462
rect 5977 -650 5989 -474
rect 6023 -650 6035 -474
rect 5977 -662 6035 -650
rect 6065 -474 6123 -462
rect 6065 -650 6077 -474
rect 6111 -650 6123 -474
rect 6065 -662 6123 -650
rect 6293 -474 6351 -462
rect 6293 -650 6305 -474
rect 6339 -650 6351 -474
rect 6293 -662 6351 -650
rect 6381 -474 6439 -462
rect 6381 -650 6393 -474
rect 6427 -650 6439 -474
rect 6381 -662 6439 -650
rect 6609 -474 6667 -462
rect 6609 -850 6621 -474
rect 6655 -850 6667 -474
rect 6609 -862 6667 -850
rect 6697 -474 6755 -462
rect 6697 -850 6709 -474
rect 6743 -850 6755 -474
rect 6697 -862 6755 -850
rect 7133 -531 7185 -515
rect 7133 -565 7141 -531
rect 7175 -565 7185 -531
rect 7133 -599 7185 -565
rect 7133 -633 7141 -599
rect 7175 -633 7185 -599
rect 7133 -645 7185 -633
rect 7215 -563 7269 -515
rect 7215 -597 7225 -563
rect 7259 -597 7269 -563
rect 7215 -645 7269 -597
rect 7299 -595 7353 -515
rect 7299 -629 7309 -595
rect 7343 -629 7353 -595
rect 7299 -645 7353 -629
rect 7383 -563 7437 -515
rect 7383 -597 7393 -563
rect 7427 -597 7437 -563
rect 7383 -645 7437 -597
rect 7467 -595 7521 -515
rect 7467 -629 7477 -595
rect 7511 -629 7521 -595
rect 7467 -645 7521 -629
rect 7551 -563 7603 -515
rect 7551 -597 7561 -563
rect 7595 -597 7603 -563
rect 7551 -645 7603 -597
rect 5824 -1188 5886 -1176
rect 5824 -1364 5836 -1188
rect 5870 -1364 5886 -1188
rect 5824 -1376 5886 -1364
rect 5916 -1188 5978 -1176
rect 5916 -1364 5932 -1188
rect 5966 -1364 5978 -1188
rect 5916 -1376 5978 -1364
rect 6034 -1188 6096 -1176
rect 6034 -1364 6046 -1188
rect 6080 -1364 6096 -1188
rect 6034 -1376 6096 -1364
rect 6126 -1188 6188 -1176
rect 6126 -1364 6142 -1188
rect 6176 -1364 6188 -1188
rect 6126 -1376 6188 -1364
rect 6244 -1188 6306 -1176
rect 6244 -1364 6256 -1188
rect 6290 -1364 6306 -1188
rect 6244 -1376 6306 -1364
rect 6336 -1188 6398 -1176
rect 6336 -1364 6352 -1188
rect 6386 -1364 6398 -1188
rect 6336 -1376 6398 -1364
rect 6454 -1188 6516 -1176
rect 6454 -1364 6466 -1188
rect 6500 -1364 6516 -1188
rect 6454 -1376 6516 -1364
rect 6546 -1188 6608 -1176
rect 6546 -1364 6562 -1188
rect 6596 -1364 6608 -1188
rect 6546 -1376 6608 -1364
<< pdiff >>
rect 5662 755 5720 767
rect 5662 579 5674 755
rect 5708 579 5720 755
rect 5662 567 5720 579
rect 5750 755 5808 767
rect 5750 579 5762 755
rect 5796 579 5808 755
rect 5750 567 5808 579
rect 5662 155 5720 167
rect 5662 -21 5674 155
rect 5708 -21 5720 155
rect 5662 -33 5720 -21
rect 5750 155 5808 167
rect 5750 -21 5762 155
rect 5796 -21 5808 155
rect 5750 -33 5808 -21
rect 5978 755 6036 767
rect 5978 -21 5990 755
rect 6024 -21 6036 755
rect 5978 -33 6036 -21
rect 6066 755 6124 767
rect 6066 -21 6078 755
rect 6112 -21 6124 755
rect 6066 -33 6124 -21
rect 6294 755 6352 767
rect 6294 -21 6306 755
rect 6340 -21 6352 755
rect 6294 -33 6352 -21
rect 6382 755 6440 767
rect 6382 -21 6394 755
rect 6428 -21 6440 755
rect 6382 -33 6440 -21
rect 6610 755 6668 767
rect 6610 579 6622 755
rect 6656 579 6668 755
rect 6610 567 6668 579
rect 6698 755 6756 767
rect 6698 579 6710 755
rect 6744 579 6756 755
rect 6698 567 6756 579
rect 6962 881 7014 893
rect 6962 847 6970 881
rect 7004 847 7014 881
rect 6962 813 7014 847
rect 6962 779 6970 813
rect 7004 779 7014 813
rect 6962 745 7014 779
rect 6962 711 6970 745
rect 7004 711 7014 745
rect 6962 693 7014 711
rect 7044 881 7096 893
rect 7044 847 7054 881
rect 7088 847 7096 881
rect 7044 813 7096 847
rect 7044 779 7054 813
rect 7088 779 7096 813
rect 7044 745 7096 779
rect 7044 711 7054 745
rect 7088 711 7096 745
rect 7044 693 7096 711
rect 7207 881 7259 893
rect 7207 847 7215 881
rect 7249 847 7259 881
rect 7207 813 7259 847
rect 7207 779 7215 813
rect 7249 779 7259 813
rect 7207 745 7259 779
rect 7207 711 7215 745
rect 7249 711 7259 745
rect 7207 693 7259 711
rect 7289 881 7343 893
rect 7289 847 7299 881
rect 7333 847 7343 881
rect 7289 813 7343 847
rect 7289 779 7299 813
rect 7333 779 7343 813
rect 7289 745 7343 779
rect 7289 711 7299 745
rect 7333 711 7343 745
rect 7289 693 7343 711
rect 7373 881 7427 893
rect 7373 847 7383 881
rect 7417 847 7427 881
rect 7373 813 7427 847
rect 7373 779 7383 813
rect 7417 779 7427 813
rect 7373 693 7427 779
rect 7457 881 7511 893
rect 7457 847 7467 881
rect 7501 847 7511 881
rect 7457 813 7511 847
rect 7457 779 7467 813
rect 7501 779 7511 813
rect 7457 745 7511 779
rect 7457 711 7467 745
rect 7501 711 7511 745
rect 7457 693 7511 711
rect 7541 881 7593 893
rect 7541 847 7551 881
rect 7585 847 7593 881
rect 7541 693 7593 847
rect 6610 155 6668 167
rect 6610 -21 6622 155
rect 6656 -21 6668 155
rect 6610 -33 6668 -21
rect 6698 155 6756 167
rect 6698 -21 6710 155
rect 6744 -21 6756 155
rect 6698 -33 6756 -21
rect 6962 81 7014 99
rect 6962 47 6970 81
rect 7004 47 7014 81
rect 6962 13 7014 47
rect 6962 -21 6970 13
rect 7004 -21 7014 13
rect 6962 -55 7014 -21
rect 6962 -89 6970 -55
rect 7004 -89 7014 -55
rect 6962 -101 7014 -89
rect 7044 81 7096 99
rect 7044 47 7054 81
rect 7088 47 7096 81
rect 7044 13 7096 47
rect 7044 -21 7054 13
rect 7088 -21 7096 13
rect 7044 -55 7096 -21
rect 7044 -89 7054 -55
rect 7088 -89 7096 -55
rect 7044 -101 7096 -89
rect 7207 81 7259 99
rect 7207 47 7215 81
rect 7249 47 7259 81
rect 7207 13 7259 47
rect 7207 -21 7215 13
rect 7249 -21 7259 13
rect 7207 -55 7259 -21
rect 7207 -89 7215 -55
rect 7249 -89 7259 -55
rect 7207 -101 7259 -89
rect 7289 81 7343 99
rect 7289 47 7299 81
rect 7333 47 7343 81
rect 7289 13 7343 47
rect 7289 -21 7299 13
rect 7333 -21 7343 13
rect 7289 -55 7343 -21
rect 7289 -89 7299 -55
rect 7333 -89 7343 -55
rect 7289 -101 7343 -89
rect 7373 13 7427 99
rect 7373 -21 7383 13
rect 7417 -21 7427 13
rect 7373 -55 7427 -21
rect 7373 -89 7383 -55
rect 7417 -89 7427 -55
rect 7373 -101 7427 -89
rect 7457 81 7511 99
rect 7457 47 7467 81
rect 7501 47 7511 81
rect 7457 13 7511 47
rect 7457 -21 7467 13
rect 7501 -21 7511 13
rect 7457 -55 7511 -21
rect 7457 -89 7467 -55
rect 7501 -89 7511 -55
rect 7457 -101 7511 -89
rect 7541 -55 7593 99
rect 7541 -89 7551 -55
rect 7585 -89 7593 -55
rect 7541 -101 7593 -89
rect 7133 -207 7185 -195
rect 7133 -241 7141 -207
rect 7175 -241 7185 -207
rect 7133 -275 7185 -241
rect 7133 -309 7141 -275
rect 7175 -309 7185 -275
rect 7133 -343 7185 -309
rect 7133 -377 7141 -343
rect 7175 -377 7185 -343
rect 7133 -395 7185 -377
rect 7215 -229 7269 -195
rect 7215 -263 7225 -229
rect 7259 -263 7269 -229
rect 7215 -324 7269 -263
rect 7215 -358 7225 -324
rect 7259 -358 7269 -324
rect 7215 -395 7269 -358
rect 7299 -207 7353 -195
rect 7299 -241 7309 -207
rect 7343 -241 7353 -207
rect 7299 -275 7353 -241
rect 7299 -309 7309 -275
rect 7343 -309 7353 -275
rect 7299 -395 7353 -309
rect 7383 -229 7437 -195
rect 7383 -263 7393 -229
rect 7427 -263 7437 -229
rect 7383 -324 7437 -263
rect 7383 -358 7393 -324
rect 7427 -358 7437 -324
rect 7383 -395 7437 -358
rect 7467 -207 7521 -195
rect 7467 -241 7477 -207
rect 7511 -241 7521 -207
rect 7467 -275 7521 -241
rect 7467 -309 7477 -275
rect 7511 -309 7521 -275
rect 7467 -395 7521 -309
rect 7551 -213 7603 -195
rect 7551 -247 7561 -213
rect 7595 -247 7603 -213
rect 7551 -281 7603 -247
rect 7551 -315 7561 -281
rect 7595 -315 7603 -281
rect 7551 -349 7603 -315
rect 7551 -383 7561 -349
rect 7595 -383 7603 -349
rect 7551 -395 7603 -383
<< ndiffc >>
rect 6970 527 7004 561
rect 6970 459 7004 493
rect 7054 527 7088 561
rect 7054 459 7088 493
rect 7215 455 7249 489
rect 7299 463 7333 497
rect 7383 455 7417 489
rect 7467 463 7501 497
rect 7551 456 7585 490
rect 6970 299 7004 333
rect 6970 231 7004 265
rect 7054 299 7088 333
rect 7054 231 7088 265
rect 7215 303 7249 337
rect 7299 295 7333 329
rect 7383 303 7417 337
rect 7467 295 7501 329
rect 7551 302 7585 336
rect 5673 -850 5707 -474
rect 5761 -850 5795 -474
rect 5989 -650 6023 -474
rect 6077 -650 6111 -474
rect 6305 -650 6339 -474
rect 6393 -650 6427 -474
rect 6621 -850 6655 -474
rect 6709 -850 6743 -474
rect 7141 -565 7175 -531
rect 7141 -633 7175 -599
rect 7225 -597 7259 -563
rect 7309 -629 7343 -595
rect 7393 -597 7427 -563
rect 7477 -629 7511 -595
rect 7561 -597 7595 -563
rect 5836 -1364 5870 -1188
rect 5932 -1364 5966 -1188
rect 6046 -1364 6080 -1188
rect 6142 -1364 6176 -1188
rect 6256 -1364 6290 -1188
rect 6352 -1364 6386 -1188
rect 6466 -1364 6500 -1188
rect 6562 -1364 6596 -1188
<< pdiffc >>
rect 5674 579 5708 755
rect 5762 579 5796 755
rect 5674 -21 5708 155
rect 5762 -21 5796 155
rect 5990 -21 6024 755
rect 6078 -21 6112 755
rect 6306 -21 6340 755
rect 6394 -21 6428 755
rect 6622 579 6656 755
rect 6710 579 6744 755
rect 6970 847 7004 881
rect 6970 779 7004 813
rect 6970 711 7004 745
rect 7054 847 7088 881
rect 7054 779 7088 813
rect 7054 711 7088 745
rect 7215 847 7249 881
rect 7215 779 7249 813
rect 7215 711 7249 745
rect 7299 847 7333 881
rect 7299 779 7333 813
rect 7299 711 7333 745
rect 7383 847 7417 881
rect 7383 779 7417 813
rect 7467 847 7501 881
rect 7467 779 7501 813
rect 7467 711 7501 745
rect 7551 847 7585 881
rect 6622 -21 6656 155
rect 6710 -21 6744 155
rect 6970 47 7004 81
rect 6970 -21 7004 13
rect 6970 -89 7004 -55
rect 7054 47 7088 81
rect 7054 -21 7088 13
rect 7054 -89 7088 -55
rect 7215 47 7249 81
rect 7215 -21 7249 13
rect 7215 -89 7249 -55
rect 7299 47 7333 81
rect 7299 -21 7333 13
rect 7299 -89 7333 -55
rect 7383 -21 7417 13
rect 7383 -89 7417 -55
rect 7467 47 7501 81
rect 7467 -21 7501 13
rect 7467 -89 7501 -55
rect 7551 -89 7585 -55
rect 7141 -241 7175 -207
rect 7141 -309 7175 -275
rect 7141 -377 7175 -343
rect 7225 -263 7259 -229
rect 7225 -358 7259 -324
rect 7309 -241 7343 -207
rect 7309 -309 7343 -275
rect 7393 -263 7427 -229
rect 7393 -358 7427 -324
rect 7477 -241 7511 -207
rect 7477 -309 7511 -275
rect 7561 -247 7595 -213
rect 7561 -315 7595 -281
rect 7561 -383 7595 -349
<< psubdiff >>
rect 5559 -322 5655 -288
rect 5813 -322 5971 -288
rect 6129 -322 6287 -288
rect 6445 -322 6603 -288
rect 6761 -322 6857 -288
rect 5559 -384 5593 -322
rect 5875 -384 5909 -322
rect 6191 -384 6225 -322
rect 5875 -802 5909 -740
rect 6507 -384 6541 -322
rect 6191 -802 6225 -740
rect 6823 -384 6857 -322
rect 6507 -802 6541 -740
rect 5875 -836 5971 -802
rect 6129 -836 6287 -802
rect 6445 -836 6541 -802
rect 5559 -1002 5593 -940
rect 5875 -1002 5909 -836
rect 6507 -1002 6541 -836
rect 6823 -1002 6857 -940
rect 5559 -1036 5818 -1002
rect 6614 -1036 6857 -1002
rect 5722 -1098 5756 -1036
rect 6676 -1098 6710 -1036
rect 5722 -1516 5756 -1454
rect 6676 -1516 6710 -1454
rect 5722 -1550 5818 -1516
rect 6614 -1550 6710 -1516
<< nsubdiff >>
rect 5560 916 5656 950
rect 5814 916 5972 950
rect 6130 916 6288 950
rect 6446 916 6604 950
rect 6762 916 6858 950
rect 5560 854 5594 916
rect 5876 854 5910 916
rect 5560 418 5594 480
rect 5560 384 5656 418
rect 5814 384 5876 418
rect 5560 316 5876 384
rect 5560 254 5594 316
rect 5560 -182 5594 -120
rect 6192 854 6226 916
rect 5876 -182 5910 -120
rect 6508 854 6542 916
rect 6192 -182 6226 -120
rect 6824 854 6858 916
rect 6824 420 6858 480
rect 6542 418 6858 420
rect 6542 384 6604 418
rect 6762 384 6858 418
rect 6542 316 6858 384
rect 6824 254 6858 316
rect 6508 -182 6542 -120
rect 6824 -182 6858 -120
rect 5560 -216 5656 -182
rect 5814 -216 5972 -182
rect 6130 -216 6288 -182
rect 6446 -216 6604 -182
rect 6762 -216 6858 -182
<< psubdiffcont >>
rect 5655 -322 5813 -288
rect 5971 -322 6129 -288
rect 6287 -322 6445 -288
rect 6603 -322 6761 -288
rect 5559 -940 5593 -384
rect 5875 -740 5909 -384
rect 6191 -740 6225 -384
rect 6507 -740 6541 -384
rect 5971 -836 6129 -802
rect 6287 -836 6445 -802
rect 6823 -940 6857 -384
rect 5818 -1036 6614 -1002
rect 5722 -1454 5756 -1098
rect 6676 -1454 6710 -1098
rect 5818 -1550 6614 -1516
<< nsubdiffcont >>
rect 5656 916 5814 950
rect 5972 916 6130 950
rect 6288 916 6446 950
rect 6604 916 6762 950
rect 5560 480 5594 854
rect 5656 384 5814 418
rect 5560 -120 5594 254
rect 5876 -120 5910 854
rect 6192 -120 6226 854
rect 6508 -120 6542 854
rect 6824 480 6858 854
rect 6604 384 6762 418
rect 6824 -120 6858 254
rect 5656 -216 5814 -182
rect 5972 -216 6130 -182
rect 6288 -216 6446 -182
rect 6604 -216 6762 -182
<< poly >>
rect 5702 848 5768 864
rect 5702 814 5718 848
rect 5752 814 5768 848
rect 5702 798 5768 814
rect 5720 767 5750 798
rect 5720 536 5750 567
rect 5702 520 5768 536
rect 5702 486 5718 520
rect 5752 486 5768 520
rect 5702 470 5768 486
rect 5702 248 5768 264
rect 5702 214 5718 248
rect 5752 214 5768 248
rect 5702 198 5768 214
rect 5720 167 5750 198
rect 5720 -64 5750 -33
rect 5702 -80 5768 -64
rect 5702 -114 5718 -80
rect 5752 -114 5768 -80
rect 5702 -130 5768 -114
rect 6018 848 6084 864
rect 6018 814 6034 848
rect 6068 814 6084 848
rect 6018 798 6084 814
rect 6036 767 6066 798
rect 6036 -64 6066 -33
rect 6018 -80 6084 -64
rect 6018 -114 6034 -80
rect 6068 -114 6084 -80
rect 6018 -130 6084 -114
rect 6334 848 6400 864
rect 6334 814 6350 848
rect 6384 814 6400 848
rect 6334 798 6400 814
rect 6352 767 6382 798
rect 6352 -64 6382 -33
rect 6334 -80 6400 -64
rect 6334 -114 6350 -80
rect 6384 -114 6400 -80
rect 6334 -130 6400 -114
rect 6650 848 6716 864
rect 6650 814 6666 848
rect 6700 814 6716 848
rect 6650 798 6716 814
rect 7014 893 7044 919
rect 7259 893 7289 919
rect 7343 893 7373 919
rect 7427 893 7457 919
rect 7511 893 7541 919
rect 6668 767 6698 798
rect 6668 536 6698 567
rect 6650 520 6716 536
rect 6650 486 6666 520
rect 6700 486 6716 520
rect 6650 470 6716 486
rect 7014 661 7044 693
rect 7259 661 7289 693
rect 7343 661 7373 693
rect 7427 661 7457 693
rect 7511 661 7541 693
rect 6958 645 7044 661
rect 6958 611 6974 645
rect 7008 611 7044 645
rect 6958 595 7044 611
rect 7191 645 7541 661
rect 7191 611 7207 645
rect 7241 611 7299 645
rect 7333 611 7383 645
rect 7417 611 7467 645
rect 7501 611 7541 645
rect 7191 595 7541 611
rect 7014 573 7044 595
rect 7259 573 7289 595
rect 7343 573 7373 595
rect 7427 573 7457 595
rect 7511 573 7541 595
rect 7014 417 7044 443
rect 7259 417 7289 443
rect 7343 417 7373 443
rect 7427 417 7457 443
rect 7511 417 7541 443
rect 7014 349 7044 375
rect 7259 349 7289 375
rect 7343 349 7373 375
rect 7427 349 7457 375
rect 7511 349 7541 375
rect 6650 248 6716 264
rect 6650 214 6666 248
rect 6700 214 6716 248
rect 6650 198 6716 214
rect 6668 167 6698 198
rect 6668 -64 6698 -33
rect 6650 -80 6716 -64
rect 6650 -114 6666 -80
rect 6700 -114 6716 -80
rect 6650 -130 6716 -114
rect 7014 197 7044 219
rect 7259 197 7289 219
rect 7343 197 7373 219
rect 7427 197 7457 219
rect 7511 197 7541 219
rect 6958 181 7044 197
rect 6958 147 6974 181
rect 7008 147 7044 181
rect 6958 131 7044 147
rect 7191 181 7541 197
rect 7191 147 7207 181
rect 7241 147 7299 181
rect 7333 147 7383 181
rect 7417 147 7467 181
rect 7501 147 7541 181
rect 7191 131 7541 147
rect 7014 99 7044 131
rect 7259 99 7289 131
rect 7343 99 7373 131
rect 7427 99 7457 131
rect 7511 99 7541 131
rect 7014 -127 7044 -101
rect 7259 -127 7289 -101
rect 7343 -127 7373 -101
rect 7427 -127 7457 -101
rect 7511 -127 7541 -101
rect 7185 -195 7215 -169
rect 7269 -195 7299 -169
rect 7353 -195 7383 -169
rect 7437 -195 7467 -169
rect 7521 -195 7551 -169
rect 5701 -390 5767 -374
rect 5701 -424 5717 -390
rect 5751 -424 5767 -390
rect 5701 -440 5767 -424
rect 5719 -462 5749 -440
rect 6017 -390 6083 -374
rect 6017 -424 6033 -390
rect 6067 -424 6083 -390
rect 6017 -440 6083 -424
rect 6035 -462 6065 -440
rect 6035 -684 6065 -662
rect 6017 -700 6083 -684
rect 6017 -734 6033 -700
rect 6067 -734 6083 -700
rect 6017 -750 6083 -734
rect 6333 -390 6399 -374
rect 6333 -424 6349 -390
rect 6383 -424 6399 -390
rect 6333 -440 6399 -424
rect 6351 -462 6381 -440
rect 6351 -684 6381 -662
rect 6333 -700 6399 -684
rect 6333 -734 6349 -700
rect 6383 -734 6399 -700
rect 6333 -750 6399 -734
rect 6649 -390 6715 -374
rect 6649 -424 6665 -390
rect 6699 -424 6715 -390
rect 6649 -440 6715 -424
rect 6667 -462 6697 -440
rect 5719 -884 5749 -862
rect 5701 -900 5767 -884
rect 5701 -934 5717 -900
rect 5751 -934 5767 -900
rect 5701 -950 5767 -934
rect 6667 -884 6697 -862
rect 6649 -900 6715 -884
rect 6649 -934 6665 -900
rect 6699 -934 6715 -900
rect 6649 -950 6715 -934
rect 7185 -433 7215 -395
rect 7269 -433 7299 -395
rect 7353 -433 7383 -395
rect 7437 -433 7467 -395
rect 7521 -431 7551 -395
rect 7185 -443 7468 -433
rect 7185 -477 7418 -443
rect 7452 -477 7468 -443
rect 7185 -487 7468 -477
rect 7521 -443 7602 -431
rect 7521 -477 7552 -443
rect 7586 -477 7602 -443
rect 7185 -515 7215 -487
rect 7269 -515 7299 -487
rect 7353 -515 7383 -487
rect 7437 -515 7467 -487
rect 7521 -489 7602 -477
rect 7521 -515 7551 -489
rect 7185 -671 7215 -645
rect 7269 -671 7299 -645
rect 7353 -671 7383 -645
rect 7437 -671 7467 -645
rect 7521 -671 7551 -645
rect 6078 -1104 6144 -1088
rect 6078 -1138 6094 -1104
rect 6128 -1138 6144 -1104
rect 5886 -1176 5916 -1150
rect 6078 -1154 6144 -1138
rect 6498 -1104 6564 -1088
rect 6498 -1138 6514 -1104
rect 6548 -1138 6564 -1104
rect 6096 -1176 6126 -1154
rect 6306 -1176 6336 -1150
rect 6498 -1154 6564 -1138
rect 6516 -1176 6546 -1154
rect 5886 -1398 5916 -1376
rect 5868 -1414 5934 -1398
rect 6096 -1402 6126 -1376
rect 6306 -1398 6336 -1376
rect 5868 -1448 5884 -1414
rect 5918 -1448 5934 -1414
rect 5868 -1464 5934 -1448
rect 6288 -1414 6354 -1398
rect 6516 -1402 6546 -1376
rect 6288 -1448 6304 -1414
rect 6338 -1448 6354 -1414
rect 6288 -1464 6354 -1448
<< polycont >>
rect 5718 814 5752 848
rect 5718 486 5752 520
rect 5718 214 5752 248
rect 5718 -114 5752 -80
rect 6034 814 6068 848
rect 6034 -114 6068 -80
rect 6350 814 6384 848
rect 6350 -114 6384 -80
rect 6666 814 6700 848
rect 6666 486 6700 520
rect 6974 611 7008 645
rect 7207 611 7241 645
rect 7299 611 7333 645
rect 7383 611 7417 645
rect 7467 611 7501 645
rect 6666 214 6700 248
rect 6666 -114 6700 -80
rect 6974 147 7008 181
rect 7207 147 7241 181
rect 7299 147 7333 181
rect 7383 147 7417 181
rect 7467 147 7501 181
rect 5717 -424 5751 -390
rect 6033 -424 6067 -390
rect 6033 -734 6067 -700
rect 6349 -424 6383 -390
rect 6349 -734 6383 -700
rect 6665 -424 6699 -390
rect 5717 -934 5751 -900
rect 6665 -934 6699 -900
rect 7418 -477 7452 -443
rect 7552 -477 7586 -443
rect 6094 -1138 6128 -1104
rect 6514 -1138 6548 -1104
rect 5884 -1448 5918 -1414
rect 6304 -1448 6338 -1414
<< locali >>
rect 5540 1070 7820 1100
rect 5540 1010 5600 1070
rect 7730 1010 7820 1070
rect 5540 957 7820 1010
rect 5540 950 6923 957
rect 5540 940 5656 950
rect 5560 916 5656 940
rect 5814 916 5972 950
rect 6130 916 6288 950
rect 6446 916 6604 950
rect 6762 940 6923 950
rect 6762 916 6858 940
rect 6894 923 6923 940
rect 6957 923 7015 957
rect 7049 923 7107 957
rect 7141 923 7199 957
rect 7233 923 7291 957
rect 7325 923 7383 957
rect 7417 923 7475 957
rect 7509 923 7567 957
rect 7601 940 7820 957
rect 7601 923 7630 940
rect 5560 854 5594 916
rect 5876 854 5910 916
rect 5702 814 5718 848
rect 5752 814 5768 848
rect 5674 755 5708 771
rect 5674 563 5708 579
rect 5762 755 5796 771
rect 5762 563 5796 579
rect 5702 486 5718 520
rect 5752 486 5768 520
rect 5560 418 5594 480
rect 5560 384 5656 418
rect 5814 384 5876 418
rect 5560 316 5876 384
rect 5560 254 5594 316
rect 5702 214 5718 248
rect 5752 214 5768 248
rect 5674 155 5708 171
rect 5674 -37 5708 -21
rect 5762 155 5796 171
rect 5762 -37 5796 -21
rect 5702 -114 5718 -80
rect 5752 -114 5768 -80
rect 5560 -182 5594 -120
rect 6192 854 6226 916
rect 6018 814 6034 848
rect 6068 814 6084 848
rect 5990 755 6024 771
rect 5990 -37 6024 -21
rect 6078 755 6112 771
rect 6078 -37 6112 -21
rect 6018 -114 6034 -80
rect 6068 -114 6084 -80
rect 5876 -182 5910 -120
rect 6508 854 6542 916
rect 6334 814 6350 848
rect 6384 814 6400 848
rect 6306 755 6340 771
rect 6306 -37 6340 -21
rect 6394 755 6428 771
rect 6394 -37 6428 -21
rect 6334 -114 6350 -80
rect 6384 -114 6400 -80
rect 6192 -182 6226 -120
rect 6824 854 6858 916
rect 6650 814 6666 848
rect 6700 814 6716 848
rect 6622 755 6656 771
rect 6622 563 6656 579
rect 6710 755 6744 771
rect 6710 563 6744 579
rect 6650 486 6666 520
rect 6700 486 6716 520
rect 6962 881 7004 923
rect 6962 847 6970 881
rect 6962 813 7004 847
rect 6962 779 6970 813
rect 6962 745 7004 779
rect 6962 711 6970 745
rect 6962 695 7004 711
rect 7038 881 7104 889
rect 7038 847 7054 881
rect 7088 847 7104 881
rect 7038 813 7104 847
rect 7038 779 7054 813
rect 7088 779 7104 813
rect 7038 745 7104 779
rect 7038 711 7054 745
rect 7088 711 7104 745
rect 7038 693 7104 711
rect 7196 881 7249 923
rect 7196 847 7215 881
rect 7196 813 7249 847
rect 7196 779 7215 813
rect 7196 745 7249 779
rect 7196 711 7215 745
rect 7196 695 7249 711
rect 7283 881 7349 889
rect 7283 847 7299 881
rect 7333 847 7349 881
rect 7283 813 7349 847
rect 7283 779 7299 813
rect 7333 779 7349 813
rect 7283 745 7349 779
rect 7383 881 7417 923
rect 7383 813 7417 847
rect 7383 763 7417 779
rect 7451 881 7517 889
rect 7451 847 7467 881
rect 7501 847 7517 881
rect 7451 813 7517 847
rect 7551 881 7593 923
rect 7585 847 7593 881
rect 7551 831 7593 847
rect 7451 779 7467 813
rect 7501 779 7517 813
rect 7283 711 7299 745
rect 7333 729 7349 745
rect 7451 745 7517 779
rect 7451 729 7467 745
rect 7333 711 7467 729
rect 7501 733 7517 745
rect 7501 711 7604 733
rect 7283 695 7604 711
rect 7058 660 7104 693
rect 7191 660 7517 661
rect 6958 658 7024 659
rect 6958 611 6959 658
rect 7022 611 7024 658
rect 7058 645 7517 660
rect 7058 611 7207 645
rect 7241 611 7299 645
rect 7333 611 7383 645
rect 7417 611 7467 645
rect 7501 611 7517 645
rect 7551 660 7604 695
rect 7058 610 7200 611
rect 6824 420 6858 480
rect 6542 418 6858 420
rect 6542 384 6604 418
rect 6762 384 6858 418
rect 6958 561 7004 577
rect 7058 573 7104 610
rect 7551 600 7560 660
rect 7551 577 7604 600
rect 6958 527 6970 561
rect 6958 493 7004 527
rect 6958 459 6970 493
rect 6958 413 7004 459
rect 7038 561 7104 573
rect 7038 527 7054 561
rect 7088 527 7104 561
rect 7038 493 7104 527
rect 7283 541 7604 577
rect 7038 459 7054 493
rect 7088 459 7104 493
rect 7038 447 7104 459
rect 7196 489 7249 505
rect 7196 455 7215 489
rect 7196 413 7249 455
rect 7283 497 7349 541
rect 7283 463 7299 497
rect 7333 463 7349 497
rect 7283 447 7349 463
rect 7383 489 7417 505
rect 7383 413 7417 455
rect 7451 497 7517 541
rect 7451 463 7467 497
rect 7501 463 7517 497
rect 7451 447 7517 463
rect 7551 490 7601 506
rect 7585 456 7601 490
rect 7551 413 7601 456
rect 6542 316 6858 384
rect 6894 379 6923 413
rect 6957 379 7015 413
rect 7049 379 7107 413
rect 7141 379 7199 413
rect 7233 379 7291 413
rect 7325 379 7383 413
rect 7417 379 7475 413
rect 7509 379 7567 413
rect 7601 379 7630 413
rect 6824 254 6858 316
rect 6650 214 6666 248
rect 6700 214 6716 248
rect 6622 155 6656 171
rect 6622 -37 6656 -21
rect 6710 155 6744 171
rect 6710 -37 6744 -21
rect 6650 -114 6666 -80
rect 6700 -114 6716 -80
rect 6508 -182 6542 -120
rect 6958 333 7004 379
rect 6958 299 6970 333
rect 6958 265 7004 299
rect 6958 231 6970 265
rect 6958 215 7004 231
rect 7038 333 7104 345
rect 7038 299 7054 333
rect 7088 299 7104 333
rect 7038 265 7104 299
rect 7196 337 7249 379
rect 7196 303 7215 337
rect 7196 287 7249 303
rect 7283 329 7349 345
rect 7283 295 7299 329
rect 7333 295 7349 329
rect 7038 231 7054 265
rect 7088 231 7104 265
rect 7038 219 7104 231
rect 7058 181 7104 219
rect 7283 251 7349 295
rect 7383 337 7417 379
rect 7383 287 7417 303
rect 7451 329 7517 345
rect 7451 295 7467 329
rect 7501 295 7517 329
rect 7451 251 7517 295
rect 7551 336 7601 379
rect 7585 302 7601 336
rect 7551 286 7601 302
rect 7283 215 7604 251
rect 7551 190 7604 215
rect 7058 147 7207 181
rect 7241 147 7299 181
rect 7333 147 7383 181
rect 7417 147 7467 181
rect 7501 147 7517 181
rect 7058 131 7517 147
rect 7058 99 7104 131
rect 6824 -182 6858 -120
rect 6962 81 7004 97
rect 6962 47 6970 81
rect 6962 13 7004 47
rect 6962 -21 6970 13
rect 6962 -55 7004 -21
rect 6962 -89 6970 -55
rect 6962 -131 7004 -89
rect 7038 81 7104 99
rect 7551 130 7560 190
rect 7551 97 7604 130
rect 7038 47 7054 81
rect 7088 47 7104 81
rect 7038 13 7104 47
rect 7038 -21 7054 13
rect 7088 -21 7104 13
rect 7038 -55 7104 -21
rect 7038 -89 7054 -55
rect 7088 -89 7104 -55
rect 7038 -97 7104 -89
rect 7196 81 7249 97
rect 7196 47 7215 81
rect 7196 13 7249 47
rect 7196 -21 7215 13
rect 7196 -55 7249 -21
rect 7196 -89 7215 -55
rect 7196 -131 7249 -89
rect 7283 81 7604 97
rect 7283 47 7299 81
rect 7333 63 7467 81
rect 7333 47 7349 63
rect 7283 13 7349 47
rect 7451 47 7467 63
rect 7501 59 7604 81
rect 7501 47 7517 59
rect 7283 -21 7299 13
rect 7333 -21 7349 13
rect 7283 -55 7349 -21
rect 7283 -89 7299 -55
rect 7333 -89 7349 -55
rect 7283 -97 7349 -89
rect 7383 13 7417 29
rect 7383 -55 7417 -21
rect 7383 -131 7417 -89
rect 7451 13 7517 47
rect 7451 -21 7467 13
rect 7501 -21 7517 13
rect 7451 -55 7517 -21
rect 7451 -89 7467 -55
rect 7501 -89 7517 -55
rect 7451 -97 7517 -89
rect 7551 -55 7593 -39
rect 7585 -89 7593 -55
rect 7551 -131 7593 -89
rect 6894 -165 6923 -131
rect 6957 -165 7015 -131
rect 7049 -165 7107 -131
rect 7141 -165 7199 -131
rect 7233 -165 7291 -131
rect 7325 -165 7383 -131
rect 7417 -165 7475 -131
rect 7509 -165 7567 -131
rect 7601 -165 7630 -131
rect 5560 -216 5656 -182
rect 5814 -216 5972 -182
rect 6130 -216 6288 -182
rect 6446 -216 6604 -182
rect 6762 -216 6858 -182
rect 7125 -207 7191 -165
rect 7125 -241 7141 -207
rect 7175 -241 7191 -207
rect 7125 -275 7191 -241
rect 5559 -290 5655 -288
rect 5540 -322 5655 -290
rect 5813 -322 5971 -288
rect 6129 -322 6287 -288
rect 6445 -322 6603 -288
rect 6761 -290 6857 -288
rect 6761 -322 6880 -290
rect 5540 -384 5593 -322
rect 5540 -940 5559 -384
rect 5875 -384 5909 -322
rect 5701 -424 5717 -390
rect 5751 -424 5767 -390
rect 5673 -474 5707 -458
rect 5673 -866 5707 -850
rect 5761 -474 5795 -458
rect 5761 -866 5795 -850
rect 6191 -384 6225 -322
rect 6017 -424 6033 -390
rect 6067 -424 6083 -390
rect 5989 -474 6023 -458
rect 5989 -666 6023 -650
rect 6077 -474 6111 -458
rect 6077 -666 6111 -650
rect 6017 -734 6033 -700
rect 6067 -734 6083 -700
rect 5875 -802 5909 -740
rect 6507 -384 6541 -322
rect 6333 -424 6349 -390
rect 6383 -424 6399 -390
rect 6305 -474 6339 -458
rect 6305 -666 6339 -650
rect 6393 -474 6427 -458
rect 6393 -666 6427 -650
rect 6333 -734 6349 -700
rect 6383 -734 6399 -700
rect 6191 -802 6225 -740
rect 6823 -384 6880 -322
rect 6649 -424 6665 -390
rect 6699 -424 6715 -390
rect 6507 -802 6541 -740
rect 5875 -836 5971 -802
rect 6129 -836 6287 -802
rect 6445 -836 6541 -802
rect 5701 -934 5717 -900
rect 5751 -934 5767 -900
rect 5540 -1002 5593 -940
rect 5875 -1002 6541 -836
rect 6621 -474 6655 -458
rect 6621 -866 6655 -850
rect 6709 -474 6743 -458
rect 6709 -866 6743 -850
rect 6649 -934 6665 -900
rect 6699 -934 6715 -900
rect 6857 -940 6880 -384
rect 7125 -309 7141 -275
rect 7175 -309 7191 -275
rect 7125 -343 7191 -309
rect 7125 -377 7141 -343
rect 7175 -377 7191 -343
rect 7125 -395 7191 -377
rect 7225 -229 7259 -199
rect 7225 -324 7259 -263
rect 7293 -207 7359 -165
rect 7293 -241 7309 -207
rect 7343 -241 7359 -207
rect 7293 -275 7359 -241
rect 7293 -309 7309 -275
rect 7343 -309 7359 -275
rect 7293 -325 7359 -309
rect 7393 -229 7427 -199
rect 7393 -324 7427 -263
rect 7225 -369 7259 -358
rect 7463 -207 7511 -165
rect 7463 -241 7477 -207
rect 7463 -275 7511 -241
rect 7463 -309 7477 -275
rect 7463 -325 7511 -309
rect 7545 -213 7611 -199
rect 7545 -247 7561 -213
rect 7595 -247 7611 -213
rect 7545 -281 7611 -247
rect 7545 -315 7561 -281
rect 7595 -315 7611 -281
rect 7393 -369 7427 -358
rect 7545 -349 7611 -315
rect 7545 -361 7561 -349
rect 7225 -403 7427 -369
rect 7468 -383 7561 -361
rect 7595 -383 7611 -349
rect 7468 -395 7611 -383
rect 7225 -430 7324 -403
rect 7225 -490 7240 -430
rect 7300 -490 7324 -430
rect 7468 -443 7502 -395
rect 7402 -477 7418 -443
rect 7452 -477 7502 -443
rect 7536 -477 7540 -429
rect 7607 -477 7612 -429
rect 7225 -511 7324 -490
rect 7468 -511 7502 -477
rect 7125 -531 7191 -515
rect 7125 -565 7141 -531
rect 7175 -565 7191 -531
rect 7125 -599 7191 -565
rect 7125 -633 7141 -599
rect 7175 -633 7191 -599
rect 7125 -675 7191 -633
rect 7225 -545 7427 -511
rect 7468 -545 7595 -511
rect 7225 -563 7259 -545
rect 7393 -563 7427 -545
rect 7225 -641 7259 -597
rect 7293 -595 7359 -579
rect 7293 -629 7309 -595
rect 7343 -629 7359 -595
rect 7293 -675 7359 -629
rect 7561 -563 7595 -545
rect 7393 -641 7427 -597
rect 7477 -595 7525 -579
rect 7511 -629 7525 -595
rect 7477 -675 7525 -629
rect 7561 -641 7595 -597
rect 7078 -709 7107 -675
rect 7141 -709 7199 -675
rect 7233 -709 7291 -675
rect 7325 -709 7383 -675
rect 7417 -709 7475 -675
rect 7509 -709 7567 -675
rect 7601 -709 7630 -675
rect 6823 -1002 6880 -940
rect 5540 -1036 5818 -1002
rect 6614 -1036 6880 -1002
rect 5540 -1098 5756 -1036
rect 5540 -1454 5722 -1098
rect 6676 -1098 6880 -1036
rect 6078 -1138 6094 -1104
rect 6128 -1138 6144 -1104
rect 6498 -1138 6514 -1104
rect 6548 -1138 6564 -1104
rect 5836 -1188 5870 -1172
rect 5836 -1380 5870 -1364
rect 5932 -1188 5966 -1172
rect 5932 -1380 5966 -1364
rect 6046 -1188 6080 -1172
rect 6046 -1380 6080 -1364
rect 6142 -1188 6176 -1172
rect 6142 -1380 6176 -1364
rect 6256 -1188 6290 -1172
rect 6256 -1380 6290 -1364
rect 6352 -1188 6386 -1172
rect 6352 -1380 6386 -1364
rect 6466 -1188 6500 -1172
rect 6466 -1380 6500 -1364
rect 6562 -1188 6596 -1172
rect 6562 -1380 6596 -1364
rect 5868 -1448 5884 -1414
rect 5918 -1448 5934 -1414
rect 6288 -1448 6304 -1414
rect 6338 -1448 6354 -1414
rect 5540 -1516 5756 -1454
rect 6710 -1454 6880 -1098
rect 6676 -1516 6880 -1454
rect 5540 -1550 5818 -1516
rect 6614 -1520 6880 -1516
rect 6614 -1550 7820 -1520
rect 5540 -1630 7820 -1550
rect 5540 -1690 5600 -1630
rect 7730 -1690 7820 -1630
rect 5540 -1740 7820 -1690
<< viali >>
rect 5600 1010 7730 1070
rect 6923 923 6957 957
rect 7015 923 7049 957
rect 7107 923 7141 957
rect 7199 923 7233 957
rect 7291 923 7325 957
rect 7383 923 7417 957
rect 7475 923 7509 957
rect 7567 923 7601 957
rect 5718 814 5752 848
rect 5674 579 5708 755
rect 5762 579 5796 755
rect 5718 486 5752 520
rect 5718 214 5752 248
rect 5674 -21 5708 155
rect 5762 -21 5796 155
rect 5718 -114 5752 -80
rect 6034 814 6068 848
rect 5990 -21 6024 755
rect 6078 -21 6112 755
rect 6034 -114 6068 -80
rect 6350 814 6384 848
rect 6306 -21 6340 755
rect 6394 -21 6428 755
rect 6350 -114 6384 -80
rect 6666 814 6700 848
rect 6622 579 6656 755
rect 6710 579 6744 755
rect 6666 486 6700 520
rect 6959 645 7022 658
rect 6959 611 6974 645
rect 6974 611 7008 645
rect 7008 611 7022 645
rect 7560 600 7620 660
rect 6923 379 6957 413
rect 7015 379 7049 413
rect 7107 379 7141 413
rect 7199 379 7233 413
rect 7291 379 7325 413
rect 7383 379 7417 413
rect 7475 379 7509 413
rect 7567 379 7601 413
rect 6666 214 6700 248
rect 6622 -21 6656 155
rect 6710 -21 6744 155
rect 6666 -114 6700 -80
rect 6958 147 6974 181
rect 6974 147 7008 181
rect 7008 147 7024 181
rect 6958 133 7024 147
rect 7560 130 7620 190
rect 6923 -165 6957 -131
rect 7015 -165 7049 -131
rect 7107 -165 7141 -131
rect 7199 -165 7233 -131
rect 7291 -165 7325 -131
rect 7383 -165 7417 -131
rect 7475 -165 7509 -131
rect 7567 -165 7601 -131
rect 5717 -424 5751 -390
rect 5673 -850 5707 -474
rect 5761 -850 5795 -474
rect 6033 -424 6067 -390
rect 5989 -650 6023 -474
rect 6077 -650 6111 -474
rect 6033 -734 6067 -700
rect 6349 -424 6383 -390
rect 6305 -650 6339 -474
rect 6393 -650 6427 -474
rect 6349 -734 6383 -700
rect 6665 -424 6699 -390
rect 5717 -934 5751 -900
rect 6621 -850 6655 -474
rect 6709 -850 6743 -474
rect 6665 -934 6699 -900
rect 7240 -490 7300 -430
rect 7540 -443 7607 -429
rect 7540 -477 7552 -443
rect 7552 -477 7586 -443
rect 7586 -477 7607 -443
rect 7107 -709 7141 -675
rect 7199 -709 7233 -675
rect 7291 -709 7325 -675
rect 7383 -709 7417 -675
rect 7475 -709 7509 -675
rect 7567 -709 7601 -675
rect 6094 -1138 6128 -1104
rect 6514 -1138 6548 -1104
rect 5836 -1364 5870 -1188
rect 5932 -1364 5966 -1188
rect 6046 -1364 6080 -1188
rect 6142 -1364 6176 -1188
rect 6256 -1364 6290 -1188
rect 6352 -1364 6386 -1188
rect 6466 -1364 6500 -1188
rect 6562 -1364 6596 -1188
rect 5884 -1448 5918 -1414
rect 6304 -1448 6338 -1414
rect 5600 -1690 7730 -1630
<< metal1 >>
rect 5540 1070 7820 1100
rect 5540 1010 5600 1070
rect 7730 1010 7820 1070
rect 5540 990 5650 1010
rect 5710 990 5900 1010
rect 5970 990 6040 1010
rect 6110 990 6320 1010
rect 6390 990 6450 1010
rect 6520 990 6710 1010
rect 6770 990 7320 1010
rect 7380 990 7420 1010
rect 7480 990 7820 1010
rect 5540 957 7820 990
rect 5540 940 6923 957
rect 6894 923 6923 940
rect 6957 923 7015 957
rect 7049 923 7107 957
rect 7141 923 7199 957
rect 7233 923 7291 957
rect 7325 923 7383 957
rect 7417 923 7475 957
rect 7509 923 7567 957
rect 7601 940 7820 957
rect 7601 923 7630 940
rect 6894 892 7630 923
rect 5706 850 5764 854
rect 5560 848 5770 850
rect 5560 814 5718 848
rect 5752 814 5770 848
rect 6022 848 6080 854
rect 6022 845 6034 848
rect 5560 810 5770 814
rect 5880 815 6034 845
rect 5560 520 5600 810
rect 5706 808 5764 810
rect 5668 755 5714 767
rect 5668 740 5674 755
rect 5708 740 5714 755
rect 5756 755 5802 767
rect 5640 680 5650 740
rect 5710 680 5720 740
rect 5668 579 5674 680
rect 5708 579 5714 680
rect 5668 567 5714 579
rect 5756 579 5762 755
rect 5796 595 5802 755
rect 5796 579 5850 595
rect 5756 567 5850 579
rect 5775 565 5850 567
rect 5706 520 5764 526
rect 5560 486 5718 520
rect 5752 486 5770 520
rect 5560 480 5770 486
rect 5560 250 5600 480
rect 5820 410 5850 565
rect 5770 350 5780 410
rect 5840 350 5850 410
rect 5706 250 5764 254
rect 5560 248 5770 250
rect 5560 214 5718 248
rect 5752 214 5770 248
rect 5560 210 5770 214
rect 5560 -80 5600 210
rect 5706 208 5764 210
rect 5668 155 5714 167
rect 5668 130 5674 155
rect 5708 130 5714 155
rect 5756 155 5802 167
rect 5640 70 5650 130
rect 5710 70 5720 130
rect 5668 -21 5674 70
rect 5708 -21 5714 70
rect 5668 -33 5714 -21
rect 5756 -21 5762 155
rect 5796 20 5802 155
rect 5796 -21 5830 20
rect 5756 -33 5830 -21
rect 5706 -80 5764 -74
rect 5560 -114 5718 -80
rect 5752 -114 5770 -80
rect 5560 -120 5770 -114
rect 5560 -390 5600 -120
rect 5800 -350 5830 -33
rect 5880 -85 5910 815
rect 6022 814 6034 815
rect 6068 814 6080 848
rect 6022 808 6080 814
rect 6338 848 6396 854
rect 6338 814 6350 848
rect 6384 845 6396 848
rect 6654 850 6712 854
rect 6654 848 6860 850
rect 6384 815 6540 845
rect 6384 814 6396 815
rect 6338 808 6396 814
rect 5984 755 6030 767
rect 5984 740 5990 755
rect 6024 740 6030 755
rect 6072 755 6118 767
rect 5960 680 5970 740
rect 6030 680 6040 740
rect 5984 640 5990 680
rect 6024 640 6030 680
rect 5960 580 5970 640
rect 6030 580 6040 640
rect 5984 550 5990 580
rect 6024 550 6030 580
rect 5960 490 5970 550
rect 6030 490 6040 550
rect 5984 -21 5990 490
rect 6024 -21 6030 490
rect 6072 410 6078 755
rect 6112 410 6118 755
rect 6300 755 6346 767
rect 6300 410 6306 755
rect 6340 410 6346 755
rect 6388 755 6434 767
rect 6388 740 6394 755
rect 6428 740 6434 755
rect 6380 680 6390 740
rect 6450 680 6460 740
rect 6388 640 6394 680
rect 6428 640 6434 680
rect 6380 580 6390 640
rect 6450 580 6460 640
rect 6388 550 6394 580
rect 6428 550 6434 580
rect 6380 490 6390 550
rect 6450 490 6460 550
rect 6060 350 6070 410
rect 6130 350 6140 410
rect 6280 350 6290 410
rect 6350 350 6360 410
rect 5984 -33 6030 -21
rect 6072 -21 6078 350
rect 6112 115 6118 350
rect 6300 115 6306 350
rect 6112 85 6180 115
rect 6112 -21 6118 85
rect 6072 -33 6118 -21
rect 6150 -70 6180 85
rect 6240 85 6306 115
rect 6022 -80 6080 -74
rect 6022 -85 6034 -80
rect 5880 -114 6034 -85
rect 6068 -114 6080 -80
rect 5880 -115 6080 -114
rect 5880 -180 5910 -115
rect 6022 -120 6080 -115
rect 6120 -130 6130 -70
rect 6190 -130 6200 -70
rect 5860 -240 5870 -180
rect 5930 -240 5940 -180
rect 5800 -360 5860 -350
rect 5705 -390 5763 -384
rect 5560 -424 5717 -390
rect 5751 -424 5763 -390
rect 5560 -430 5763 -424
rect 5800 -430 5860 -420
rect 5900 -395 5930 -240
rect 6021 -390 6079 -384
rect 6021 -395 6033 -390
rect 5900 -424 6033 -395
rect 6067 -424 6079 -390
rect 5900 -425 6079 -424
rect 5560 -900 5590 -430
rect 5667 -474 5713 -462
rect 5667 -480 5673 -474
rect 5630 -540 5640 -480
rect 5667 -640 5673 -540
rect 5630 -700 5640 -640
rect 5667 -850 5673 -700
rect 5707 -850 5713 -474
rect 5667 -862 5713 -850
rect 5755 -474 5801 -462
rect 5755 -850 5761 -474
rect 5795 -750 5801 -474
rect 5900 -705 5930 -425
rect 6021 -430 6079 -425
rect 5983 -474 6029 -462
rect 5983 -580 5989 -474
rect 5960 -590 5989 -580
rect 6023 -590 6029 -474
rect 6071 -474 6117 -462
rect 6023 -650 6030 -590
rect 6071 -650 6077 -474
rect 6111 -530 6117 -474
rect 6150 -530 6180 -130
rect 6240 -180 6270 85
rect 6300 -21 6306 85
rect 6340 -21 6346 350
rect 6300 -33 6346 -21
rect 6388 -21 6394 490
rect 6428 -21 6434 490
rect 6388 -33 6434 -21
rect 6510 -70 6540 815
rect 6654 814 6666 848
rect 6700 814 6860 848
rect 6654 810 6860 814
rect 6654 808 6712 810
rect 6616 755 6662 767
rect 6616 595 6622 755
rect 6570 579 6622 595
rect 6656 579 6662 755
rect 6704 755 6750 767
rect 6704 740 6710 755
rect 6744 740 6750 755
rect 6700 680 6710 740
rect 6770 680 6780 740
rect 6570 567 6662 579
rect 6704 579 6710 680
rect 6744 579 6750 680
rect 6704 567 6750 579
rect 6570 565 6645 567
rect 6570 410 6600 565
rect 6820 530 6860 810
rect 6950 664 6960 670
rect 6947 658 6960 664
rect 7020 664 7030 670
rect 7020 658 7034 664
rect 6947 611 6959 658
rect 7022 611 7034 658
rect 6947 610 6960 611
rect 7020 610 7034 611
rect 6947 605 7034 610
rect 7548 660 7632 666
rect 7548 600 7560 660
rect 7620 600 7632 660
rect 7548 594 7632 600
rect 6660 526 6870 530
rect 6654 520 6870 526
rect 6654 486 6666 520
rect 6700 490 6870 520
rect 6700 486 6712 490
rect 6654 480 6712 486
rect 6570 350 6580 410
rect 6640 350 6650 410
rect 6654 250 6712 254
rect 6820 250 6860 490
rect 7540 444 7820 460
rect 6894 413 7820 444
rect 6894 379 6923 413
rect 6957 379 7015 413
rect 7049 379 7107 413
rect 7141 379 7199 413
rect 7233 379 7291 413
rect 7325 379 7383 413
rect 7417 379 7475 413
rect 7509 379 7567 413
rect 7601 379 7820 413
rect 6894 348 7820 379
rect 7540 340 7820 348
rect 6654 248 6870 250
rect 6654 214 6666 248
rect 6700 214 6870 248
rect 6654 210 6870 214
rect 6654 208 6712 210
rect 6616 155 6662 167
rect 6616 20 6622 155
rect 6590 -21 6622 20
rect 6656 -21 6662 155
rect 6704 155 6750 167
rect 6704 130 6710 155
rect 6744 130 6750 155
rect 6700 70 6710 130
rect 6770 70 6780 130
rect 6590 -33 6662 -21
rect 6704 -21 6710 70
rect 6744 -21 6750 70
rect 6704 -33 6750 -21
rect 6338 -80 6396 -74
rect 6338 -114 6350 -80
rect 6384 -85 6396 -80
rect 6480 -85 6490 -70
rect 6384 -114 6490 -85
rect 6338 -115 6490 -114
rect 6338 -120 6396 -115
rect 6480 -130 6490 -115
rect 6550 -130 6560 -70
rect 6220 -240 6230 -180
rect 6290 -240 6300 -180
rect 6111 -560 6180 -530
rect 6240 -530 6270 -240
rect 6337 -390 6395 -384
rect 6490 -390 6520 -130
rect 6590 -350 6620 -33
rect 6654 -80 6712 -74
rect 6820 -80 6860 210
rect 7548 190 7632 196
rect 6950 187 6960 190
rect 6946 181 6960 187
rect 7020 187 7030 190
rect 7020 181 7036 187
rect 6946 133 6958 181
rect 7024 133 7036 181
rect 6946 130 6960 133
rect 7020 130 7036 133
rect 6946 127 7036 130
rect 7548 130 7560 190
rect 7620 130 7632 190
rect 7548 124 7632 130
rect 6650 -114 6666 -80
rect 6700 -114 6860 -80
rect 6650 -120 6860 -114
rect 6337 -424 6349 -390
rect 6383 -424 6520 -390
rect 6337 -430 6520 -424
rect 6560 -360 6620 -350
rect 6820 -380 6860 -120
rect 6894 -120 7630 -100
rect 6894 -131 7320 -120
rect 7380 -131 7420 -120
rect 7480 -131 7630 -120
rect 6894 -165 6923 -131
rect 6957 -165 7015 -131
rect 7049 -165 7107 -131
rect 7141 -165 7199 -131
rect 7233 -165 7291 -131
rect 7380 -165 7383 -131
rect 7417 -165 7420 -131
rect 7509 -165 7567 -131
rect 7601 -165 7630 -131
rect 6894 -180 7320 -165
rect 7380 -180 7420 -165
rect 7480 -180 7630 -165
rect 6894 -196 7630 -180
rect 6650 -390 6860 -380
rect 6650 -420 6665 -390
rect 6560 -430 6620 -420
rect 6653 -424 6665 -420
rect 6699 -420 6860 -390
rect 6699 -424 6711 -420
rect 6653 -430 6711 -424
rect 6299 -474 6345 -462
rect 6299 -530 6305 -474
rect 6240 -560 6305 -530
rect 6111 -650 6117 -560
rect 5960 -660 6029 -650
rect 5983 -662 6029 -660
rect 6071 -662 6117 -650
rect 6299 -650 6305 -560
rect 6339 -650 6345 -474
rect 6387 -474 6433 -462
rect 6387 -590 6393 -474
rect 6427 -590 6433 -474
rect 6380 -650 6390 -590
rect 6450 -650 6460 -590
rect 6299 -662 6345 -650
rect 6387 -662 6433 -650
rect 6021 -700 6079 -694
rect 6021 -705 6033 -700
rect 5900 -734 6033 -705
rect 6067 -734 6079 -700
rect 5900 -735 6079 -734
rect 5900 -740 5930 -735
rect 6021 -740 6079 -735
rect 6337 -700 6395 -694
rect 6490 -700 6520 -430
rect 6337 -734 6349 -700
rect 6383 -734 6520 -700
rect 6337 -740 6520 -734
rect 6615 -474 6661 -462
rect 6615 -750 6621 -474
rect 5840 -810 5850 -750
rect 6580 -810 6590 -750
rect 5795 -850 5801 -810
rect 5755 -862 5801 -850
rect 6615 -850 6621 -810
rect 6655 -850 6661 -474
rect 6703 -474 6749 -462
rect 6703 -480 6709 -474
rect 6743 -480 6749 -474
rect 6690 -540 6700 -480
rect 6760 -540 6770 -480
rect 6703 -640 6709 -540
rect 6743 -640 6749 -540
rect 6690 -700 6700 -640
rect 6760 -700 6770 -640
rect 6615 -862 6661 -850
rect 6703 -850 6709 -700
rect 6743 -850 6749 -700
rect 6703 -862 6749 -850
rect 5705 -900 5763 -894
rect 6653 -900 6711 -894
rect 6820 -900 6854 -420
rect 7220 -424 7310 -420
rect 7220 -430 7312 -424
rect 7220 -490 7240 -430
rect 7300 -490 7312 -430
rect 7528 -429 7619 -423
rect 7528 -477 7540 -429
rect 7607 -430 7619 -429
rect 7528 -483 7550 -477
rect 7540 -490 7550 -483
rect 7610 -490 7620 -430
rect 7220 -496 7312 -490
rect 7220 -500 7310 -496
rect 7700 -640 7820 340
rect 7540 -644 7820 -640
rect 7078 -675 7820 -644
rect 7078 -709 7107 -675
rect 7141 -709 7199 -675
rect 7233 -709 7291 -675
rect 7325 -709 7383 -675
rect 7417 -709 7475 -675
rect 7509 -709 7567 -675
rect 7601 -709 7820 -675
rect 7078 -740 7820 -709
rect 7540 -760 7820 -740
rect 7220 -900 7230 -880
rect 5560 -934 5717 -900
rect 5751 -934 6665 -900
rect 6699 -934 7230 -900
rect 5560 -940 7230 -934
rect 7290 -940 7300 -880
rect 5630 -1040 5640 -980
rect 5700 -1040 5710 -980
rect 5630 -1520 5710 -1040
rect 5770 -1050 5780 -990
rect 5840 -1050 5850 -990
rect 5950 -1050 5960 -990
rect 6020 -1025 6030 -990
rect 6020 -1050 6040 -1025
rect 6380 -1050 6390 -990
rect 6450 -1050 6460 -990
rect 6580 -1050 6590 -990
rect 6650 -1050 6660 -990
rect 6690 -1040 6700 -980
rect 6760 -1040 6770 -980
rect 6010 -1176 6040 -1050
rect 6070 -1140 6080 -1080
rect 6140 -1140 6150 -1080
rect 6082 -1144 6140 -1140
rect 6390 -1176 6420 -1050
rect 6502 -1100 6560 -1098
rect 6500 -1104 6560 -1100
rect 6500 -1138 6514 -1104
rect 6548 -1138 6560 -1104
rect 6500 -1176 6560 -1138
rect 6590 -1176 6620 -1050
rect 5830 -1188 5876 -1176
rect 5830 -1364 5836 -1188
rect 5870 -1310 5876 -1188
rect 5926 -1188 5972 -1176
rect 5926 -1310 5932 -1188
rect 5830 -1370 5870 -1364
rect 5930 -1364 5932 -1310
rect 5966 -1364 5972 -1188
rect 6010 -1188 6086 -1176
rect 6010 -1220 6046 -1188
rect 5930 -1370 5972 -1364
rect 5830 -1376 5972 -1370
rect 6040 -1364 6046 -1220
rect 6080 -1364 6086 -1188
rect 6040 -1376 6086 -1364
rect 6136 -1188 6182 -1176
rect 6136 -1364 6142 -1188
rect 6176 -1310 6182 -1188
rect 6250 -1188 6296 -1176
rect 6176 -1364 6190 -1310
rect 6136 -1370 6190 -1364
rect 6250 -1364 6256 -1188
rect 6290 -1364 6296 -1188
rect 6136 -1376 6182 -1370
rect 6250 -1376 6296 -1364
rect 6346 -1188 6420 -1176
rect 6346 -1364 6352 -1188
rect 6386 -1220 6420 -1188
rect 6460 -1188 6620 -1176
rect 6386 -1364 6392 -1220
rect 6346 -1376 6392 -1364
rect 6460 -1364 6466 -1188
rect 6500 -1240 6562 -1188
rect 6500 -1310 6506 -1240
rect 6556 -1310 6562 -1240
rect 6460 -1370 6500 -1364
rect 6560 -1364 6562 -1310
rect 6596 -1240 6620 -1188
rect 6596 -1364 6602 -1240
rect 6560 -1370 6602 -1364
rect 6460 -1376 6506 -1370
rect 6556 -1376 6602 -1370
rect 5870 -1414 5930 -1376
rect 6292 -1410 6350 -1408
rect 5870 -1448 5884 -1414
rect 5918 -1448 5930 -1414
rect 5870 -1460 5930 -1448
rect 6280 -1470 6290 -1410
rect 6350 -1470 6360 -1410
rect 6690 -1520 6770 -1040
rect 7700 -1520 7820 -760
rect 5540 -1630 7820 -1520
rect 5540 -1690 5600 -1630
rect 7730 -1690 7820 -1630
rect 5540 -1740 7820 -1690
<< via1 >>
rect 5650 1010 5710 1050
rect 5900 1010 5970 1050
rect 6040 1010 6110 1050
rect 6320 1010 6390 1050
rect 6450 1010 6520 1050
rect 6710 1010 6770 1050
rect 7320 1010 7380 1050
rect 7420 1010 7480 1050
rect 5650 990 5710 1010
rect 5900 990 5970 1010
rect 6040 990 6110 1010
rect 6320 990 6390 1010
rect 6450 990 6520 1010
rect 6710 990 6770 1010
rect 7320 990 7380 1010
rect 7420 990 7480 1010
rect 5650 680 5674 740
rect 5674 680 5708 740
rect 5708 680 5710 740
rect 5780 350 5840 410
rect 5650 70 5674 130
rect 5674 70 5708 130
rect 5708 70 5710 130
rect 5970 680 5990 740
rect 5990 680 6024 740
rect 6024 680 6030 740
rect 5970 580 5990 640
rect 5990 580 6024 640
rect 6024 580 6030 640
rect 5970 490 5990 550
rect 5990 490 6024 550
rect 6024 490 6030 550
rect 6390 680 6394 740
rect 6394 680 6428 740
rect 6428 680 6450 740
rect 6390 580 6394 640
rect 6394 580 6428 640
rect 6428 580 6450 640
rect 6390 490 6394 550
rect 6394 490 6428 550
rect 6428 490 6450 550
rect 6070 350 6078 410
rect 6078 350 6112 410
rect 6112 350 6130 410
rect 6290 350 6306 410
rect 6306 350 6340 410
rect 6340 350 6350 410
rect 6130 -130 6190 -70
rect 5870 -240 5930 -180
rect 5800 -420 5860 -360
rect 5640 -540 5673 -480
rect 5673 -540 5700 -480
rect 5640 -700 5673 -640
rect 5673 -700 5700 -640
rect 5960 -650 5989 -590
rect 5989 -650 6020 -590
rect 6710 680 6744 740
rect 6744 680 6770 740
rect 6960 658 7020 670
rect 6960 611 7020 658
rect 6960 610 7020 611
rect 7560 600 7620 660
rect 6580 350 6640 410
rect 6710 70 6744 130
rect 6744 70 6770 130
rect 6490 -130 6550 -70
rect 6230 -240 6290 -180
rect 6960 181 7020 190
rect 6960 133 7020 181
rect 6960 130 7020 133
rect 7560 130 7620 190
rect 6560 -420 6620 -360
rect 7320 -131 7380 -120
rect 7420 -131 7480 -120
rect 7320 -165 7325 -131
rect 7325 -165 7380 -131
rect 7420 -165 7475 -131
rect 7475 -165 7480 -131
rect 7320 -180 7380 -165
rect 7420 -180 7480 -165
rect 6390 -650 6393 -590
rect 6393 -650 6427 -590
rect 6427 -650 6450 -590
rect 5780 -810 5795 -750
rect 5795 -810 5840 -750
rect 6590 -810 6621 -750
rect 6621 -810 6650 -750
rect 6700 -540 6709 -480
rect 6709 -540 6743 -480
rect 6743 -540 6760 -480
rect 6700 -700 6709 -640
rect 6709 -700 6743 -640
rect 6743 -700 6760 -640
rect 7240 -490 7300 -430
rect 7550 -477 7607 -430
rect 7607 -477 7610 -430
rect 7550 -490 7610 -477
rect 7230 -940 7290 -880
rect 5640 -1040 5700 -980
rect 5780 -1050 5840 -990
rect 5960 -1050 6020 -990
rect 6390 -1050 6450 -990
rect 6590 -1050 6650 -990
rect 6700 -1040 6760 -980
rect 6080 -1104 6140 -1080
rect 6080 -1138 6094 -1104
rect 6094 -1138 6128 -1104
rect 6128 -1138 6140 -1104
rect 6080 -1140 6140 -1138
rect 5870 -1370 5930 -1310
rect 6190 -1370 6250 -1310
rect 6500 -1370 6560 -1310
rect 6290 -1414 6350 -1410
rect 6290 -1448 6304 -1414
rect 6304 -1448 6338 -1414
rect 6338 -1448 6350 -1414
rect 6290 -1470 6350 -1448
<< metal2 >>
rect 5650 1050 5710 1060
rect 5650 740 5710 990
rect 5900 1050 6520 1060
rect 5970 990 6040 1050
rect 6110 990 6320 1050
rect 6390 990 6450 1050
rect 5900 980 6520 990
rect 6710 1050 6770 1060
rect 5650 130 5710 680
rect 5970 740 6040 980
rect 6030 680 6040 740
rect 5970 640 6040 680
rect 6030 580 6040 640
rect 5970 550 6040 580
rect 6030 490 6040 550
rect 5970 480 6040 490
rect 6390 740 6450 980
rect 6390 640 6450 680
rect 6390 550 6450 580
rect 6390 480 6450 490
rect 6710 740 6770 990
rect 7320 1050 7480 1060
rect 7380 990 7420 1050
rect 5780 410 5840 420
rect 6070 410 6130 420
rect 5840 360 6070 400
rect 5780 340 5840 350
rect 6070 340 6130 350
rect 6290 410 6350 420
rect 6580 410 6640 420
rect 6350 360 6580 400
rect 6290 340 6350 350
rect 6580 340 6640 350
rect 5650 60 5710 70
rect 6710 130 6770 680
rect 6960 670 7020 680
rect 7020 615 7115 645
rect 6960 600 7020 610
rect 6960 190 7020 200
rect 6960 120 7020 130
rect 6710 60 6770 70
rect 6130 -70 6190 -60
rect 6490 -70 6550 -60
rect 6190 -120 6490 -90
rect 6130 -140 6190 -130
rect 6975 -90 7005 120
rect 6550 -120 7005 -90
rect 6490 -140 6550 -130
rect 5870 -180 5930 -170
rect 6230 -180 6290 -170
rect 5930 -230 6230 -200
rect 5870 -250 5930 -240
rect 7085 -200 7115 615
rect 7320 -120 7480 990
rect 7560 660 7620 670
rect 7620 610 7860 650
rect 7560 590 7620 600
rect 7560 190 7620 200
rect 7620 140 7860 180
rect 7560 120 7620 130
rect 7380 -180 7420 -120
rect 7320 -190 7480 -180
rect 6290 -230 7115 -200
rect 6230 -250 6290 -240
rect 5800 -360 5860 -350
rect 6560 -360 6620 -350
rect 5860 -415 6000 -385
rect 5800 -430 5860 -420
rect 5640 -480 5700 -470
rect 5640 -640 5700 -540
rect 5970 -580 6000 -415
rect 6415 -420 6560 -390
rect 6415 -580 6445 -420
rect 6560 -430 6620 -420
rect 7240 -430 7300 -420
rect 6700 -480 6760 -470
rect 5960 -590 6020 -580
rect 5960 -660 6020 -650
rect 6390 -590 6450 -580
rect 6390 -660 6450 -650
rect 6700 -640 6760 -540
rect 5640 -980 5700 -700
rect 5780 -750 5840 -740
rect 5780 -820 5840 -810
rect 5790 -980 5820 -820
rect 5970 -980 6010 -660
rect 6400 -980 6440 -660
rect 6590 -750 6650 -740
rect 6590 -820 6650 -810
rect 6610 -980 6640 -820
rect 6700 -980 6760 -700
rect 7240 -500 7300 -490
rect 7550 -430 7610 -420
rect 7610 -480 7860 -440
rect 7550 -500 7610 -490
rect 7240 -870 7280 -500
rect 7230 -880 7290 -870
rect 7230 -950 7290 -940
rect 5640 -1050 5700 -1040
rect 5780 -990 5840 -980
rect 5780 -1060 5840 -1050
rect 5960 -990 6020 -980
rect 5960 -1060 6020 -1050
rect 6390 -990 6450 -980
rect 6390 -1060 6450 -1050
rect 6590 -990 6650 -980
rect 6700 -1050 6760 -1040
rect 6590 -1060 6650 -1050
rect 6080 -1080 6140 -1070
rect 5450 -1130 6080 -1090
rect 6080 -1150 6140 -1140
rect 5870 -1310 5930 -1300
rect 6190 -1310 6250 -1300
rect 5930 -1360 6190 -1320
rect 5870 -1380 5930 -1370
rect 6500 -1310 6560 -1300
rect 6250 -1360 6500 -1320
rect 6190 -1380 6250 -1370
rect 6500 -1380 6560 -1370
rect 6290 -1410 6350 -1400
rect 5450 -1460 6290 -1420
rect 6290 -1480 6350 -1470
<< labels >>
rlabel metal2 7820 -480 7860 -440 1 EN
port 3 n
rlabel metal2 5450 -1130 5490 -1090 1 VIN_P
port 1 n
rlabel metal2 5450 -1460 5490 -1420 1 VIN_N
port 2 n
rlabel metal2 7820 140 7860 180 1 OUT_N
port 5 n
rlabel metal2 7820 610 7860 650 1 OUT_P
port 4 n
rlabel locali 5570 970 5830 1080 1 VDD
port 0 n
rlabel metal1 5580 -1710 5840 -1600 1 VSS
port 6 n
<< end >>
