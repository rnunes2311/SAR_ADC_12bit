** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12b/delay_cell/delay_cell.sch

.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt delay_cell VDD t_10ns t_8p5ns t_7ns t_5p3ns t_3p7ns t_2p1ns OUT IN VSS
*.PININFO OUT:O t_10ns:B t_8p5ns:B t_7ns:B t_5p3ns:B t_3p7ns:B t_2p1ns:B VSS:I IN:I VDD:I
XM1 RAMP IN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 t_10ns IN_Z VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=12 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 t_8p5ns t_10ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
XR2 t_7ns t_8p5ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
XR3 t_5p3ns t_7ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
XR4 t_3p7ns t_5p3ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
XR5 t_2p1ns t_3p7ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
x1 IN VSS VSS VDD VDD IN_Z sky130_fd_sc_hd__inv_2
XM4 ST_OUT RAMP VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 RAMP VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 ST_OUT n1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 ST_OUT IN_Z VSS VSS VDD VDD n1 sky130_fd_sc_hd__nor2_2
x3 n1 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_2
x4 net1 VSS VSS VDD VDD OUT sky130_fd_sc_hd__inv_4
XR6 RAMP t_2p1ns VSS sky130_fd_pr__res_high_po_0p35 L=12.5 mult=1 m=1
XM7 ST_OUT n1 net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC2 RAMP VSS sky130_fd_pr__cap_mim_m3_1 W=12.5 L=8 MF=1 m=1
.ends
.end
