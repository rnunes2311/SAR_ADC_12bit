magic
tech sky130A
magscale 1 2
timestamp 1717107273
<< locali >>
rect -3490 9890 2730 9930
rect -3490 9850 -3390 9890
rect 2640 9850 2730 9890
rect -3490 9790 2730 9850
rect -3490 7810 -3460 9790
rect -3400 9770 2730 9790
rect 2840 9890 7620 9930
rect 2840 9840 2880 9890
rect 7490 9840 7620 9890
rect 2840 9820 7620 9840
rect 2840 9770 7530 9820
rect -3400 7840 -3360 9770
rect -3400 7820 -2040 7840
rect -3400 7810 -2600 7820
rect -3490 7770 -2600 7810
rect -3490 7710 -3360 7770
rect -3150 7760 -2600 7770
rect -2080 7760 -2040 7820
rect -3150 7740 -2040 7760
rect 4910 7610 6130 7640
rect 4910 7550 4940 7610
rect 6080 7550 6130 7610
rect 4910 7530 6130 7550
rect -3490 6800 -3110 7220
rect -1020 6800 160 7000
rect -3490 6720 160 6800
rect 2400 6970 2530 7030
rect 2400 6800 2460 6970
rect 7490 6800 7530 9770
rect 2400 6720 4480 6800
rect 6260 6750 7530 6800
rect 7570 6750 7620 9820
rect 6260 6720 7620 6750
rect -3490 6690 7620 6720
rect -3490 6630 -3400 6690
rect 7480 6630 7620 6690
rect -3490 6580 7620 6630
<< viali >>
rect -3390 9850 2640 9890
rect -3460 7810 -3400 9790
rect 2880 9840 7490 9890
rect -2600 7760 -2080 7820
rect -3230 7520 -3180 7570
rect 4940 7550 6080 7610
rect -3314 7429 -3260 7477
rect 7530 6750 7570 9820
rect -3400 6630 7480 6690
<< metal1 >>
rect -3490 9890 2730 9930
rect -3490 9850 -3390 9890
rect 2640 9850 2730 9890
rect -3490 9790 2730 9850
rect -3600 8690 -3590 8750
rect -3530 8690 -3520 8750
rect -3580 7640 -3540 8690
rect -3490 7810 -3460 9790
rect -3400 9770 2730 9790
rect 2840 9890 7620 9930
rect 2840 9840 2880 9890
rect 7490 9840 7620 9890
rect 2840 9820 7620 9840
rect 2840 9770 7530 9820
rect -3400 9400 -3360 9770
rect -3230 9710 150 9720
rect -3230 9640 40 9710
rect 110 9640 150 9710
rect -1480 9580 -1440 9640
rect -3400 9350 -3090 9400
rect -3400 7840 -3360 9350
rect -3020 9340 -3010 9400
rect -2950 9340 -2940 9400
rect -2750 9340 -2740 9400
rect -2680 9340 -2670 9400
rect -2470 9340 -2460 9400
rect -2400 9340 -2390 9400
rect -2200 9340 -2190 9400
rect -2130 9340 -2120 9400
rect -1930 9340 -1920 9400
rect -1860 9340 -1850 9400
rect -1660 9340 -1650 9400
rect -1590 9340 -1580 9400
rect -1390 9340 -1380 9400
rect -1320 9340 -1310 9400
rect -1110 9340 -1100 9400
rect -1040 9340 -1030 9400
rect -840 9340 -830 9400
rect -770 9340 -760 9400
rect -570 9340 -560 9400
rect -500 9340 -490 9400
rect -300 9340 -290 9400
rect -230 9340 -220 9400
rect 230 9380 270 9770
rect 400 9685 1070 9690
rect 10 9330 270 9380
rect 300 9655 1070 9685
rect 300 9250 330 9655
rect 400 9650 1070 9655
rect 1310 9655 2075 9685
rect 260 9190 270 9250
rect 330 9190 340 9250
rect -3024 8842 -3014 8902
rect -2954 8842 -2944 8902
rect -2754 8842 -2744 8902
rect -2684 8842 -2674 8902
rect -2474 8842 -2464 8902
rect -2404 8842 -2394 8902
rect -2204 8842 -2194 8902
rect -2134 8842 -2124 8902
rect -1934 8842 -1924 8902
rect -1864 8842 -1854 8902
rect -1664 8842 -1654 8902
rect -1594 8842 -1584 8902
rect -1394 8842 -1384 8902
rect -1324 8842 -1314 8902
rect -1114 8842 -1104 8902
rect -1044 8842 -1034 8902
rect -844 8842 -834 8902
rect -774 8842 -764 8902
rect -574 8842 -564 8902
rect -504 8842 -494 8902
rect -304 8842 -294 8902
rect -234 8842 -224 8902
rect -2864 8692 -2854 8752
rect -2794 8692 -2784 8752
rect -2594 8692 -2584 8752
rect -2524 8692 -2514 8752
rect -140 8690 -130 8750
rect -70 8690 -60 8750
rect -2314 8522 -2304 8582
rect -2244 8522 -2234 8582
rect -2044 8522 -2034 8582
rect -1974 8522 -1964 8582
rect -1774 8522 -1764 8582
rect -1704 8522 -1694 8582
rect -1234 8522 -1224 8582
rect -1164 8522 -1154 8582
rect -954 8522 -944 8582
rect -884 8522 -874 8582
rect -684 8522 -674 8582
rect -614 8522 -604 8582
rect -414 8402 -404 8462
rect -344 8402 -334 8462
rect 300 8355 330 9190
rect 1310 9130 1340 9655
rect 2390 9650 2400 9710
rect 2460 9650 2470 9710
rect 2410 9570 2440 9650
rect 2410 9540 2520 9570
rect 2670 9540 2700 9770
rect 2970 9590 2980 9660
rect 3050 9590 3060 9660
rect 2620 9510 2700 9540
rect 3350 9440 3760 9480
rect 6990 9470 7360 9630
rect 2565 9395 2720 9425
rect 1280 9070 1290 9130
rect 1350 9070 1360 9130
rect 460 8710 470 8770
rect 530 8710 540 8770
rect 650 8710 660 8770
rect 720 8710 730 8770
rect 850 8710 860 8770
rect 920 8710 930 8770
rect 1050 8710 1060 8770
rect 1120 8710 1130 8770
rect 360 8530 370 8590
rect 430 8530 440 8590
rect 550 8530 560 8590
rect 620 8530 630 8590
rect 750 8530 760 8590
rect 820 8530 830 8590
rect 950 8530 960 8590
rect 1020 8530 1030 8590
rect 1140 8530 1150 8590
rect 1210 8530 1220 8590
rect 1090 8355 1100 8370
rect 300 8325 1100 8355
rect 1090 8310 1100 8325
rect 1160 8310 1170 8370
rect 1310 8355 1340 9070
rect 2420 9050 2610 9090
rect 1470 8900 1480 8960
rect 1540 8900 1550 8960
rect 1660 8900 1670 8960
rect 1730 8900 1740 8960
rect 1860 8900 1870 8960
rect 1930 8900 1940 8960
rect 2060 8900 2070 8960
rect 2130 8900 2140 8960
rect 2310 8900 2320 8960
rect 2380 8900 2390 8960
rect 2250 8710 2260 8770
rect 2320 8710 2330 8770
rect 1370 8530 1380 8590
rect 1440 8530 1450 8590
rect 1570 8530 1580 8590
rect 1640 8530 1650 8590
rect 1770 8530 1780 8590
rect 1840 8530 1850 8590
rect 1960 8530 1970 8590
rect 2030 8530 2040 8590
rect 2160 8530 2170 8590
rect 2230 8530 2240 8590
rect 1235 8325 2175 8355
rect -3024 8232 -3014 8292
rect -2954 8232 -2944 8292
rect -2754 8232 -2744 8292
rect -2684 8232 -2674 8292
rect -2474 8232 -2464 8292
rect -2404 8232 -2394 8292
rect -2204 8232 -2194 8292
rect -2134 8232 -2124 8292
rect -1934 8232 -1924 8292
rect -1864 8232 -1854 8292
rect -1664 8232 -1654 8292
rect -1594 8232 -1584 8292
rect -1394 8232 -1384 8292
rect -1324 8232 -1314 8292
rect -1114 8232 -1104 8292
rect -1044 8232 -1034 8292
rect -844 8232 -834 8292
rect -774 8232 -764 8292
rect -574 8232 -564 8292
rect -504 8232 -494 8292
rect -304 8232 -294 8292
rect -234 8232 -224 8292
rect 1235 8255 1265 8325
rect 1370 8255 1380 8280
rect 300 8225 1265 8255
rect 1310 8225 1380 8255
rect -2318 8074 -2308 8134
rect -2248 8074 -2238 8134
rect -2048 8074 -2038 8134
rect -1978 8074 -1968 8134
rect -1778 8074 -1768 8134
rect -1708 8074 -1698 8134
rect -1238 8074 -1228 8134
rect -1168 8074 -1158 8134
rect -958 8074 -948 8134
rect -888 8074 -878 8134
rect -688 8074 -678 8134
rect -618 8074 -608 8134
rect -1480 7970 -1440 8040
rect -3230 7890 150 7970
rect -3400 7820 -2030 7840
rect -3400 7810 -2600 7820
rect -3490 7760 -2600 7810
rect -2080 7760 -2030 7820
rect -3490 7710 -2030 7760
rect -260 7700 -250 7760
rect -190 7700 -180 7760
rect -3600 7580 -3590 7640
rect -3530 7580 -3520 7640
rect -2010 7620 -1930 7650
rect -3242 7570 -3168 7576
rect -3242 7520 -3230 7570
rect -3180 7560 -3168 7570
rect -3180 7530 -2990 7560
rect -3180 7520 -3168 7530
rect -3242 7514 -3168 7520
rect -3326 7480 -3248 7483
rect -3330 7420 -3320 7480
rect -3260 7423 -3248 7480
rect -3260 7420 -3250 7423
rect -3490 6800 -3080 7260
rect -3020 7210 -2990 7530
rect -2740 7420 -2730 7480
rect -2670 7420 -2660 7480
rect -3050 7150 -3040 7210
rect -2980 7150 -2970 7210
rect -2720 6940 -2680 7420
rect -2010 7070 -1980 7620
rect -1710 7580 -1700 7640
rect -1640 7580 -1630 7640
rect -1450 7580 -1440 7640
rect -1380 7580 -1370 7640
rect -240 7630 -190 7700
rect -670 7590 -190 7630
rect -400 7540 -360 7590
rect -1820 7400 -1780 7480
rect -1840 7340 -1830 7400
rect -1770 7340 -1760 7400
rect -1560 7310 -1520 7480
rect -890 7370 -884 7400
rect -630 7350 -620 7410
rect -560 7350 -550 7410
rect -210 7350 -200 7410
rect -140 7350 -130 7410
rect -940 7310 -930 7320
rect -1580 7250 -1570 7310
rect -1510 7250 -1500 7310
rect -1030 7270 -930 7310
rect -2020 7010 -2010 7070
rect -1950 7010 -1940 7070
rect -2740 6880 -2730 6940
rect -2670 6880 -2660 6940
rect -1030 6800 -980 7270
rect -940 7260 -930 7270
rect -870 7310 -860 7320
rect -870 7270 -800 7310
rect -870 7260 -860 7270
rect -730 7260 -720 7320
rect -660 7260 -650 7320
rect -520 7260 -510 7320
rect -450 7260 -440 7320
rect -310 7260 -300 7320
rect -240 7260 -230 7320
rect -100 7260 -90 7320
rect -30 7310 -20 7320
rect -30 7270 40 7310
rect -30 7260 -20 7270
rect -400 7180 -370 7200
rect -400 7120 -360 7180
rect -890 7080 40 7120
rect 300 6925 330 8225
rect 360 8070 370 8130
rect 430 8070 440 8130
rect 560 8070 570 8130
rect 630 8070 640 8130
rect 750 8070 760 8130
rect 820 8070 830 8130
rect 950 8070 960 8130
rect 1020 8070 1030 8130
rect 1140 8070 1150 8130
rect 1210 8070 1220 8130
rect 460 7540 470 7600
rect 530 7540 540 7600
rect 650 7540 660 7600
rect 720 7540 730 7600
rect 850 7540 860 7600
rect 920 7540 930 7600
rect 1050 7540 1060 7600
rect 1120 7540 1130 7600
rect 1310 6925 1340 8225
rect 1370 8220 1380 8225
rect 1440 8255 1450 8280
rect 1440 8225 2175 8255
rect 1440 8220 1450 8225
rect 1370 8070 1380 8130
rect 1440 8070 1450 8130
rect 1570 8070 1580 8130
rect 1640 8070 1650 8130
rect 1770 8070 1780 8130
rect 1840 8070 1850 8130
rect 1960 8070 1970 8130
rect 2030 8070 2040 8130
rect 2160 8070 2170 8130
rect 2230 8070 2240 8130
rect 2270 8000 2310 8710
rect 1470 7940 1480 8000
rect 1540 7940 1550 8000
rect 1660 7940 1670 8000
rect 1730 7940 1740 8000
rect 1860 7940 1870 8000
rect 1930 7940 1940 8000
rect 2060 7940 2070 8000
rect 2130 7940 2140 8000
rect 2250 7940 2260 8000
rect 2320 7940 2330 8000
rect 2360 7600 2390 8900
rect 2310 7540 2320 7600
rect 2380 7540 2390 7600
rect 2420 7210 2450 9050
rect 2580 8950 2590 9010
rect 2650 8950 2660 9010
rect 2480 8850 2490 8910
rect 2550 8850 2560 8910
rect 2690 8630 2720 9395
rect 3550 9320 3560 9380
rect 3620 9320 3630 9380
rect 3030 9130 3290 9310
rect 2830 8950 2840 9010
rect 2900 8950 2910 9010
rect 2540 8600 2720 8630
rect 2580 7820 2590 7880
rect 2650 7820 2660 7880
rect 2390 7150 2400 7210
rect 2460 7150 2470 7210
rect 2400 6980 2540 7030
rect 300 6895 1065 6925
rect 1310 6895 2075 6925
rect 2400 6800 2460 6980
rect 2530 6870 2540 6930
rect 2600 6915 2610 6930
rect 2690 6915 2720 8600
rect 2600 6885 2720 6915
rect 2750 8850 2760 8910
rect 2820 8850 2830 8910
rect 2600 6870 2610 6885
rect 2750 6800 2780 8850
rect 2860 8460 2890 8950
rect 3040 8790 3300 8970
rect 3060 8460 3320 8640
rect 2840 8400 2850 8460
rect 2910 8400 2920 8460
rect 2830 8160 2840 8220
rect 2900 8160 2910 8220
rect 2840 8000 2900 8160
rect 3040 8130 3300 8310
rect 2830 7940 2840 8000
rect 2900 7940 2910 8000
rect 2990 7940 3050 7990
rect 2990 7750 3020 7940
rect 3575 7885 3605 9320
rect 3120 7855 3605 7885
rect 3720 7880 3760 9440
rect 5020 9400 5100 9410
rect 5020 9340 5030 9400
rect 5090 9340 5100 9400
rect 4770 8220 4850 8230
rect 4770 8160 4780 8220
rect 4840 8160 4850 8220
rect 2960 7690 2970 7750
rect 3030 7690 3040 7750
rect 2930 7110 2940 7170
rect 3000 7110 3010 7170
rect 3120 7090 3150 7855
rect 3700 7820 3710 7880
rect 3770 7820 3780 7880
rect 3350 7780 3410 7790
rect 3350 7710 3410 7720
rect 3470 7710 3530 7720
rect 3250 7110 3260 7170
rect 3320 7110 3330 7170
rect 3370 6975 3400 7710
rect 3470 7640 3530 7650
rect 3035 6895 3065 6955
rect 3205 6945 3400 6975
rect 3490 6895 3520 7640
rect 4660 7540 4670 7600
rect 4730 7540 4740 7600
rect 4550 7430 4560 7490
rect 4620 7430 4630 7490
rect 3590 7360 3600 7420
rect 3660 7360 3670 7420
rect 4080 7370 4090 7430
rect 4150 7370 4160 7430
rect 4280 7370 4380 7410
rect 3610 7170 3640 7360
rect 4350 7340 4380 7370
rect 4550 7300 4630 7430
rect 4230 7240 4240 7300
rect 4300 7240 4310 7300
rect 4550 7240 4560 7300
rect 4620 7240 4630 7300
rect 3590 7110 3600 7170
rect 3660 7110 3670 7170
rect 3730 7130 3740 7190
rect 3800 7130 3810 7190
rect 3940 7130 3950 7190
rect 4010 7130 4020 7190
rect 4130 7130 4140 7190
rect 4200 7130 4210 7190
rect 4320 7130 4330 7190
rect 4390 7130 4400 7190
rect 3610 6930 3640 7110
rect 3730 6930 3810 7130
rect 4030 7010 4040 7070
rect 4100 7010 4110 7070
rect 4550 7010 4560 7070
rect 4620 7010 4630 7070
rect 3035 6865 3520 6895
rect 3590 6870 3600 6930
rect 3660 6870 3670 6930
rect 3730 6880 4060 6930
rect 3730 6800 3810 6880
rect 4180 6870 4190 6930
rect 4250 6870 4260 6930
rect 4550 6890 4630 7010
rect 4660 7020 4740 7540
rect 4770 7380 4850 8160
rect 5020 7640 5100 9340
rect 6230 9270 7140 9310
rect 6230 7690 6270 9270
rect 7060 8960 7320 9140
rect 7070 8630 7330 8810
rect 6670 8400 6680 8460
rect 6740 8400 6750 8460
rect 6700 7990 6730 8400
rect 7050 8300 7310 8480
rect 7285 8105 7460 8135
rect 6700 7960 7070 7990
rect 4910 7610 6130 7640
rect 6210 7630 6220 7690
rect 6280 7630 6290 7690
rect 4910 7550 4940 7610
rect 6080 7550 6130 7610
rect 4910 7530 6130 7550
rect 5135 7415 6145 7465
rect 4770 7320 4780 7380
rect 4840 7320 4850 7380
rect 5600 7320 5610 7380
rect 5670 7320 5680 7380
rect 5790 7320 5800 7380
rect 5860 7320 5870 7380
rect 5980 7320 5990 7380
rect 6050 7320 6060 7380
rect 4770 7310 4850 7320
rect 5690 7190 5700 7250
rect 5760 7190 5770 7250
rect 5880 7190 5890 7250
rect 5950 7190 5960 7250
rect 5080 7070 5090 7130
rect 5150 7070 5160 7130
rect 5270 7070 5280 7130
rect 5340 7070 5350 7130
rect 4660 6960 4670 7020
rect 4730 6960 4740 7020
rect 4980 6960 4990 7020
rect 5050 6960 5060 7020
rect 5170 6960 5180 7020
rect 5240 6960 5250 7020
rect 5370 6960 5380 7020
rect 5440 6960 5450 7020
rect 6095 6930 6145 7415
rect 6230 7130 6270 7630
rect 6700 7440 6730 7960
rect 7430 7790 7460 8105
rect 7380 7730 7390 7790
rect 7450 7730 7460 7790
rect 6490 7390 7360 7440
rect 6340 7300 6350 7360
rect 6410 7300 6420 7360
rect 6540 7300 6550 7360
rect 6610 7300 6620 7360
rect 6730 7300 6740 7360
rect 6800 7300 6810 7360
rect 6210 7070 6220 7130
rect 6280 7070 6290 7130
rect 6440 7070 6450 7130
rect 6510 7070 6520 7130
rect 6630 7070 6640 7130
rect 6700 7070 6710 7130
rect 6840 6930 6880 7390
rect 7050 7190 7060 7250
rect 7120 7190 7130 7250
rect 7250 7190 7260 7250
rect 7320 7190 7330 7250
rect 6960 6960 6970 7020
rect 7030 6960 7040 7020
rect 7150 6960 7160 7020
rect 7220 6960 7230 7020
rect 7340 6960 7350 7020
rect 7410 6960 7420 7020
rect 4550 6830 4560 6890
rect 4620 6830 4630 6890
rect 5035 6880 6145 6930
rect 6400 6880 7270 6930
rect -3490 6720 160 6800
rect 2400 6720 4480 6800
rect 5480 6720 5550 6880
rect 7490 6800 7530 9770
rect 6260 6750 7530 6800
rect 7570 6750 7620 9820
rect 6260 6720 7620 6750
rect -3490 6690 7620 6720
rect -3490 6630 -3400 6690
rect 7480 6630 7620 6690
rect -3490 6580 7620 6630
<< via1 >>
rect -3590 8690 -3530 8750
rect 40 9640 110 9710
rect -3460 9340 -3400 9400
rect -3460 8840 -3400 8900
rect -3460 8230 -3400 8290
rect -3010 9340 -2950 9400
rect -2740 9340 -2680 9400
rect -2460 9340 -2400 9400
rect -2190 9340 -2130 9400
rect -1920 9340 -1860 9400
rect -1650 9340 -1590 9400
rect -1380 9340 -1320 9400
rect -1100 9340 -1040 9400
rect -830 9340 -770 9400
rect -560 9340 -500 9400
rect -290 9340 -230 9400
rect 270 9190 330 9250
rect -3014 8842 -2954 8902
rect -2744 8842 -2684 8902
rect -2464 8842 -2404 8902
rect -2194 8842 -2134 8902
rect -1924 8842 -1864 8902
rect -1654 8842 -1594 8902
rect -1384 8842 -1324 8902
rect -1104 8842 -1044 8902
rect -834 8842 -774 8902
rect -564 8842 -504 8902
rect -294 8842 -234 8902
rect -2854 8692 -2794 8752
rect -2584 8692 -2524 8752
rect -130 8690 -70 8750
rect -2304 8522 -2244 8582
rect -2034 8522 -1974 8582
rect -1764 8522 -1704 8582
rect -1224 8522 -1164 8582
rect -944 8522 -884 8582
rect -674 8522 -614 8582
rect -404 8402 -344 8462
rect 2400 9650 2460 9710
rect 2980 9590 3050 9660
rect 1290 9070 1350 9130
rect 470 8710 530 8770
rect 660 8710 720 8770
rect 860 8710 920 8770
rect 1060 8710 1120 8770
rect 370 8530 430 8590
rect 560 8530 620 8590
rect 760 8530 820 8590
rect 960 8530 1020 8590
rect 1150 8530 1210 8590
rect 1100 8310 1160 8370
rect 1480 8900 1540 8960
rect 1670 8900 1730 8960
rect 1870 8900 1930 8960
rect 2070 8900 2130 8960
rect 2320 8900 2380 8960
rect 2260 8710 2320 8770
rect 1380 8530 1440 8590
rect 1580 8530 1640 8590
rect 1780 8530 1840 8590
rect 1970 8530 2030 8590
rect 2170 8530 2230 8590
rect -3014 8232 -2954 8292
rect -2744 8232 -2684 8292
rect -2464 8232 -2404 8292
rect -2194 8232 -2134 8292
rect -1924 8232 -1864 8292
rect -1654 8232 -1594 8292
rect -1384 8232 -1324 8292
rect -1104 8232 -1044 8292
rect -834 8232 -774 8292
rect -564 8232 -504 8292
rect -294 8232 -234 8292
rect -2308 8074 -2248 8134
rect -2038 8074 -1978 8134
rect -1768 8074 -1708 8134
rect -1228 8074 -1168 8134
rect -948 8074 -888 8134
rect -678 8074 -618 8134
rect -250 7700 -190 7760
rect -3590 7580 -3530 7640
rect -3320 7477 -3260 7480
rect -3320 7429 -3314 7477
rect -3314 7429 -3260 7477
rect -3320 7420 -3260 7429
rect -2730 7420 -2670 7480
rect -3040 7150 -2980 7210
rect -1700 7580 -1640 7640
rect -1440 7580 -1380 7640
rect -1830 7340 -1770 7400
rect -620 7350 -560 7410
rect -200 7350 -140 7410
rect -1570 7250 -1510 7310
rect -2010 7010 -1950 7070
rect -2730 6880 -2670 6940
rect -930 7260 -870 7320
rect -720 7260 -660 7320
rect -510 7260 -450 7320
rect -300 7260 -240 7320
rect -90 7260 -30 7320
rect 370 8070 430 8130
rect 570 8070 630 8130
rect 760 8070 820 8130
rect 960 8070 1020 8130
rect 1150 8070 1210 8130
rect 470 7540 530 7600
rect 660 7540 720 7600
rect 860 7540 920 7600
rect 1060 7540 1120 7600
rect 1380 8220 1440 8280
rect 1380 8070 1440 8130
rect 1580 8070 1640 8130
rect 1780 8070 1840 8130
rect 1970 8070 2030 8130
rect 2170 8070 2230 8130
rect 1480 7940 1540 8000
rect 1670 7940 1730 8000
rect 1870 7940 1930 8000
rect 2070 7940 2130 8000
rect 2260 7940 2320 8000
rect 2320 7540 2380 7600
rect 2590 8950 2650 9010
rect 2490 8850 2550 8910
rect 3560 9320 3620 9380
rect 2840 8950 2900 9010
rect 2590 7820 2650 7880
rect 2400 7150 2460 7210
rect 2540 6870 2600 6930
rect 2760 8850 2820 8910
rect 2850 8400 2910 8460
rect 2840 8160 2900 8220
rect 2840 7940 2900 8000
rect 5030 9340 5090 9400
rect 4780 8160 4840 8220
rect 2970 7690 3030 7750
rect 2940 7110 3000 7170
rect 3710 7820 3770 7880
rect 3350 7720 3410 7780
rect 3260 7110 3320 7170
rect 3470 7650 3530 7710
rect 4670 7540 4730 7600
rect 4560 7430 4620 7490
rect 3600 7360 3660 7420
rect 4090 7370 4150 7430
rect 4240 7240 4300 7300
rect 4560 7240 4620 7300
rect 3600 7110 3660 7170
rect 3740 7130 3800 7190
rect 3950 7130 4010 7190
rect 4140 7130 4200 7190
rect 4330 7130 4390 7190
rect 4040 7010 4100 7070
rect 4560 7010 4620 7070
rect 3600 6870 3660 6930
rect 4190 6870 4250 6930
rect 6680 8400 6740 8460
rect 6220 7630 6280 7690
rect 4780 7320 4840 7380
rect 5610 7320 5670 7380
rect 5800 7320 5860 7380
rect 5990 7320 6050 7380
rect 5700 7190 5760 7250
rect 5890 7190 5950 7250
rect 5090 7070 5150 7130
rect 5280 7070 5340 7130
rect 4670 6960 4730 7020
rect 4990 6960 5050 7020
rect 5180 6960 5240 7020
rect 5380 6960 5440 7020
rect 7390 7730 7450 7790
rect 6350 7300 6410 7360
rect 6550 7300 6610 7360
rect 6740 7300 6800 7360
rect 6220 7070 6280 7130
rect 6450 7070 6510 7130
rect 6640 7070 6700 7130
rect 7060 7190 7120 7250
rect 7260 7190 7320 7250
rect 6970 6960 7030 7020
rect 7160 6960 7220 7020
rect 7350 6960 7410 7020
rect 4560 6830 4620 6890
<< metal2 >>
rect 40 9710 110 9720
rect 2400 9710 2460 9720
rect 110 9650 2400 9710
rect 2460 9660 3050 9710
rect 2460 9650 2980 9660
rect 2400 9640 2460 9650
rect 40 9630 110 9640
rect 2980 9580 3050 9590
rect -3480 9400 5120 9420
rect -3480 9340 -3460 9400
rect -3400 9340 -3010 9400
rect -2950 9340 -2740 9400
rect -2680 9340 -2460 9400
rect -2400 9340 -2190 9400
rect -2130 9340 -1920 9400
rect -1860 9340 -1650 9400
rect -1590 9340 -1380 9400
rect -1320 9340 -1100 9400
rect -1040 9340 -830 9400
rect -770 9340 -560 9400
rect -500 9340 -290 9400
rect -230 9380 5030 9400
rect -230 9340 3560 9380
rect -3480 9320 3560 9340
rect 3620 9340 5030 9380
rect 5090 9340 5120 9400
rect 3620 9320 5120 9340
rect 3560 9310 3620 9320
rect 270 9250 330 9260
rect -3630 9200 270 9240
rect 270 9180 330 9190
rect 1290 9130 1350 9140
rect -3630 9080 1290 9120
rect 1290 9060 1350 9070
rect 2590 9010 2650 9020
rect 1470 8960 2390 8970
rect -3480 8902 -210 8920
rect -3480 8900 -3014 8902
rect -3480 8840 -3460 8900
rect -3400 8842 -3014 8900
rect -2954 8842 -2744 8902
rect -2684 8842 -2464 8902
rect -2404 8842 -2194 8902
rect -2134 8842 -1924 8902
rect -1864 8842 -1654 8902
rect -1594 8842 -1384 8902
rect -1324 8842 -1104 8902
rect -1044 8842 -834 8902
rect -774 8842 -564 8902
rect -504 8842 -294 8902
rect -234 8842 -210 8902
rect 1470 8900 1480 8960
rect 1540 8900 1670 8960
rect 1730 8900 1870 8960
rect 1930 8900 2070 8960
rect 2130 8900 2320 8960
rect 2380 8900 2390 8960
rect 2840 9010 2900 9020
rect 2650 8960 2840 8990
rect 2590 8940 2650 8950
rect 2840 8940 2900 8950
rect 1470 8890 2390 8900
rect 2490 8910 2550 8920
rect -3400 8840 -210 8842
rect 2760 8910 2820 8920
rect 2550 8860 2760 8890
rect 2490 8840 2550 8850
rect 2760 8840 2820 8850
rect -3480 8820 -210 8840
rect 460 8770 2320 8780
rect -3590 8750 -3530 8760
rect -2854 8752 -2794 8762
rect -3530 8692 -2854 8750
rect -2584 8752 -2524 8762
rect -2794 8692 -2584 8750
rect -130 8750 -70 8760
rect -2524 8692 -130 8750
rect -3530 8690 -130 8692
rect 460 8710 470 8770
rect 530 8710 660 8770
rect 720 8710 860 8770
rect 920 8710 1060 8770
rect 1120 8710 2260 8770
rect 460 8700 2320 8710
rect -3590 8680 -3530 8690
rect -2854 8682 -2794 8690
rect -2584 8682 -2524 8690
rect -130 8680 -70 8690
rect -2330 8590 2235 8610
rect -2330 8582 370 8590
rect -2330 8522 -2304 8582
rect -2244 8522 -2034 8582
rect -1974 8522 -1764 8582
rect -1704 8522 -1224 8582
rect -1164 8522 -944 8582
rect -884 8522 -674 8582
rect -614 8530 370 8582
rect 430 8530 560 8590
rect 620 8530 760 8590
rect 820 8530 960 8590
rect 1020 8530 1150 8590
rect 1210 8530 1380 8590
rect 1440 8530 1580 8590
rect 1640 8530 1780 8590
rect 1840 8530 1970 8590
rect 2030 8530 2170 8590
rect 2230 8530 2235 8590
rect -614 8522 2235 8530
rect -2330 8500 2235 8522
rect -404 8462 -344 8472
rect 2850 8460 2910 8470
rect -344 8410 2850 8450
rect -404 8392 -344 8402
rect 6680 8460 6740 8470
rect 2910 8410 6680 8450
rect 2850 8390 2910 8400
rect 6680 8390 6740 8400
rect 1100 8370 1160 8380
rect 1160 8320 1430 8360
rect -3480 8292 -210 8310
rect 1100 8300 1160 8310
rect -3480 8290 -3014 8292
rect -3480 8230 -3460 8290
rect -3400 8232 -3014 8290
rect -2954 8232 -2744 8292
rect -2684 8232 -2464 8292
rect -2404 8232 -2194 8292
rect -2134 8232 -1924 8292
rect -1864 8232 -1654 8292
rect -1594 8232 -1384 8292
rect -1324 8232 -1104 8292
rect -1044 8232 -834 8292
rect -774 8232 -564 8292
rect -504 8232 -294 8292
rect -234 8232 -210 8292
rect 1390 8290 1430 8320
rect -3400 8230 -210 8232
rect -3480 8210 -210 8230
rect 1380 8280 1440 8290
rect 1380 8210 1440 8220
rect 2840 8220 4840 8230
rect -2334 8134 2235 8162
rect 2900 8160 4780 8220
rect 2840 8150 4840 8160
rect -2334 8074 -2308 8134
rect -2248 8074 -2038 8134
rect -1978 8074 -1768 8134
rect -1708 8074 -1228 8134
rect -1168 8074 -948 8134
rect -888 8074 -678 8134
rect -618 8130 2235 8134
rect -618 8074 370 8130
rect -2334 8070 370 8074
rect 430 8070 570 8130
rect 630 8070 760 8130
rect 820 8070 960 8130
rect 1020 8070 1150 8130
rect 1210 8070 1380 8130
rect 1440 8070 1580 8130
rect 1640 8070 1780 8130
rect 1840 8070 1970 8130
rect 2030 8070 2170 8130
rect 2230 8070 2235 8130
rect -2334 8052 2235 8070
rect 1470 8000 2900 8010
rect 1470 7940 1480 8000
rect 1540 7940 1670 8000
rect 1730 7940 1870 8000
rect 1930 7940 2070 8000
rect 2130 7940 2260 8000
rect 2320 7940 2840 8000
rect 1470 7930 2900 7940
rect 2590 7880 2650 7890
rect 3710 7880 3770 7890
rect 2650 7830 3710 7870
rect 2590 7810 2650 7820
rect 3710 7810 3770 7820
rect 7390 7790 7450 7800
rect -250 7760 -190 7770
rect 2970 7750 3030 7760
rect -190 7710 2970 7740
rect -250 7690 -190 7700
rect 3340 7720 3350 7780
rect 3410 7740 7390 7780
rect 3410 7720 3420 7740
rect 2970 7680 3030 7690
rect 3460 7650 3470 7710
rect 3530 7700 3540 7710
rect 3530 7690 6280 7700
rect 3530 7660 6220 7690
rect 3530 7650 3540 7660
rect -3590 7640 -3530 7650
rect -1700 7640 -1640 7650
rect -3530 7590 -1700 7620
rect -3590 7570 -3530 7580
rect -1700 7570 -1640 7580
rect -1440 7640 -1380 7650
rect 6220 7620 6280 7630
rect -1440 7570 -1380 7580
rect 460 7600 4740 7610
rect -1425 7500 -1395 7570
rect 460 7540 470 7600
rect 530 7540 660 7600
rect 720 7540 860 7600
rect 920 7540 1060 7600
rect 1120 7540 2320 7600
rect 2380 7540 4670 7600
rect 4730 7540 4740 7600
rect 460 7530 4740 7540
rect -1425 7490 6210 7500
rect -3320 7480 -3260 7490
rect -3630 7430 -3320 7470
rect -2730 7480 -2670 7490
rect -3260 7430 -2730 7470
rect -3320 7410 -3260 7420
rect -1425 7470 4560 7490
rect 4090 7430 4150 7440
rect 3600 7420 3660 7430
rect -2730 7410 -2670 7420
rect -620 7410 -560 7420
rect -1830 7400 -1770 7410
rect -3630 7350 -1830 7380
rect -200 7410 -140 7420
rect -560 7360 -200 7400
rect -620 7340 -560 7350
rect -140 7360 3600 7400
rect 3660 7380 4090 7410
rect 4550 7430 4560 7470
rect 4620 7430 6210 7490
rect 4550 7420 6210 7430
rect 4090 7360 4150 7370
rect 4780 7380 6050 7390
rect 3600 7350 3660 7360
rect -200 7340 -140 7350
rect -1830 7330 -1770 7340
rect -930 7320 -870 7330
rect -1570 7310 -1510 7320
rect -3630 7260 -1570 7290
rect -720 7320 -660 7330
rect -870 7270 -720 7310
rect -930 7250 -870 7260
rect -510 7320 -450 7330
rect -660 7270 -510 7310
rect -720 7250 -660 7260
rect -300 7320 -240 7330
rect -450 7270 -300 7310
rect -510 7250 -450 7260
rect -90 7320 -30 7330
rect -240 7270 -90 7310
rect -300 7250 -240 7260
rect 4840 7320 5610 7380
rect 5670 7320 5800 7380
rect 5860 7320 5990 7380
rect 4780 7310 6050 7320
rect 6130 7370 6210 7420
rect 6130 7360 6800 7370
rect -90 7250 -30 7260
rect 4240 7300 4620 7310
rect -1570 7240 -1510 7250
rect 4300 7240 4560 7300
rect 6130 7300 6350 7360
rect 6410 7300 6550 7360
rect 6610 7300 6740 7360
rect 6130 7290 6800 7300
rect 6860 7260 6900 7740
rect 7390 7720 7450 7730
rect 4240 7230 4620 7240
rect 5700 7250 7330 7260
rect -3040 7210 -2980 7220
rect 2400 7210 2460 7220
rect -2980 7160 2400 7190
rect -3040 7140 -2980 7150
rect 3740 7190 4390 7200
rect 2400 7140 2460 7150
rect 2940 7170 3000 7180
rect 3260 7170 3320 7180
rect 3000 7120 3260 7150
rect 2940 7100 3000 7110
rect 3600 7170 3660 7180
rect 3320 7120 3600 7150
rect 3260 7100 3320 7110
rect 3800 7130 3950 7190
rect 4010 7130 4140 7190
rect 4200 7130 4330 7190
rect 5760 7190 5890 7250
rect 5950 7190 7060 7250
rect 7120 7190 7260 7250
rect 7320 7230 7330 7250
rect 7320 7200 7680 7230
rect 7320 7190 7330 7200
rect 5700 7180 7330 7190
rect 3740 7120 4390 7130
rect 5090 7130 6710 7140
rect 3600 7100 3660 7110
rect -2010 7070 -1950 7080
rect -2015 7020 -2010 7050
rect 4040 7070 4620 7080
rect -1950 7020 4040 7050
rect -2010 7000 -1950 7010
rect 4100 7010 4560 7070
rect 5150 7070 5280 7130
rect 5340 7070 6220 7130
rect 6280 7070 6450 7130
rect 6510 7070 6640 7130
rect 6700 7120 6710 7130
rect 6700 7090 7680 7120
rect 6700 7070 6710 7090
rect 5090 7060 6710 7070
rect 4040 7000 4620 7010
rect 4670 7020 5440 7030
rect 4730 6960 4990 7020
rect 5050 6960 5180 7020
rect 5240 6960 5380 7020
rect 4670 6950 5440 6960
rect 5520 7020 7420 7030
rect 5520 6960 6970 7020
rect 7030 6960 7160 7020
rect 7220 6960 7350 7020
rect 7410 6960 7420 7020
rect 5520 6950 7420 6960
rect -2730 6940 -2670 6950
rect 2540 6930 2600 6940
rect -2670 6890 2540 6930
rect -2730 6870 -2670 6880
rect 2540 6860 2600 6870
rect 3600 6930 3660 6940
rect 4190 6930 4250 6940
rect 3660 6880 4190 6910
rect 3600 6860 3660 6870
rect 5520 6900 5600 6950
rect 4190 6860 4250 6870
rect 4550 6890 5600 6900
rect 4550 6830 4560 6890
rect 4620 6830 5600 6890
rect 4550 6820 5600 6830
use sky130_fd_pr__nfet_01v8_7CP4KT  sky130_fd_pr__nfet_01v8_7CP4KT_0
timestamp 1717106919
transform 1 0 -429 0 1 7354
box -635 -410 635 410
use sky130_fd_pr__nfet_01v8_F5PS5H  sky130_fd_pr__nfet_01v8_F5PS5H_0
timestamp 1717106919
transform 1 0 7189 0 1 7162
box -359 -410 359 410
use sky130_fd_pr__pfet_01v8_3QWEX8  sky130_fd_pr__pfet_01v8_3QWEX8_0
timestamp 1717106919
transform 1 0 791 0 1 8289
box -559 -1537 559 1537
use sky130_fd_pr__pfet_01v8_GCK2T6  sky130_fd_pr__pfet_01v8_GCK2T6_0
timestamp 1717106919
transform 1 0 -1538 0 1 8807
box -1878 -1019 1878 1019
use sky130_fd_pr__pfet_01v8_hvt_U47ZGH  sky130_fd_pr__pfet_01v8_hvt_U47ZGH_0
timestamp 1717106919
transform 1 0 5827 0 1 7171
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_hvt_U47ZGH  sky130_fd_pr__pfet_01v8_hvt_U47ZGH_1
timestamp 1717106919
transform 1 0 5215 0 1 7171
box -359 -419 359 419
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1717106919
transform 1 0 2573 0 1 9544
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_XPKDX6  sky130_fd_pr__pfet_01v8_XPKDX6_0
timestamp 1717106919
transform 1 0 1803 0 1 8289
box -559 -1537 559 1537
use sky130_fd_pr__res_high_po_0p35_699HP9  sky130_fd_pr__res_high_po_0p35_699HP9_0
timestamp 1717106919
transform 0 -1 5166 1 0 8797
box -1031 -2382 1031 2382
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -3380 0 1 7214
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_lvt_56HSEP  XM8
timestamp 1717106919
transform 1 0 4169 0 1 7152
box -359 -400 359 400
use sky130_fd_pr__nfet_01v8_F5PS5H  XM12
timestamp 1717106919
transform 1 0 6577 0 1 7162
box -359 -410 359 410
use sky130_fd_pr__pfet_01v8_lvt_6VC8VM  XM15
timestamp 1717106919
transform 1 0 -1667 0 1 7610
box -425 -284 425 284
use sky130_fd_pr__nfet_01v8_VGBCTM  XM16
timestamp 1717106919
transform 1 0 2573 0 1 7762
box -211 -1010 211 1010
use sky130_fd_pr__nfet_01v8_64Z3AY  XM18
timestamp 1717106919
transform 1 0 2573 0 1 8945
box -211 -279 211 279
use sky130_fd_pr__nfet_03v3_nvt_Y5TA2C  XM19
timestamp 1717106919
transform 1 0 3129 0 1 7029
box -357 -277 357 277
<< labels >>
rlabel metal2 -3630 9200 -3590 9240 1 IN_P
port 1 n
rlabel metal2 -3630 9080 -3590 9120 1 IN_N
port 2 n
rlabel metal2 7650 7200 7680 7230 1 OUT_N
port 3 n
rlabel metal2 7650 7090 7680 7120 1 OUT_P
port 4 n
rlabel metal2 -3630 7430 -3590 7470 1 EN
port 5 n
rlabel metal2 -3630 7350 -3600 7380 1 CAL_P
port 6 n
rlabel metal2 -3630 7260 -3600 7290 1 CAL_N
port 7 n
rlabel metal1 -3430 6730 -3190 6870 1 VSS
port 8 n
rlabel metal1 -3460 9780 -3220 9920 1 VDD
port 9 n
<< end >>
