magic
tech sky130A
magscale 1 2
timestamp 1711813427
<< error_p >>
rect 19 272 77 278
rect 19 238 31 272
rect 19 232 77 238
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -77 -278 -19 -272
<< nmos >>
rect -63 -200 -33 200
rect 33 -200 63 200
<< ndiff >>
rect -125 188 -63 200
rect -125 -188 -113 188
rect -79 -188 -63 188
rect -125 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 125 200
rect 63 -188 79 188
rect 113 -188 125 188
rect 63 -200 125 -188
<< ndiffc >>
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
<< poly >>
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -63 200 -33 226
rect 15 222 81 238
rect 33 200 63 222
rect -63 -222 -33 -200
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
<< polycont >>
rect 31 238 65 272
rect -65 -272 -31 -238
<< locali >>
rect 15 238 31 272
rect 65 238 81 272
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect -81 -272 -65 -238
rect -31 -272 -15 -238
<< viali >>
rect 31 238 65 272
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect -65 -272 -31 -238
<< metal1 >>
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
