* SPICE3 file created from SAR_ADC_12bit_flat.ext - technology: sky130A

.subckt SAR_ADC_12bit_flat CLK_DATA DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5]
+ RST_Z START EN_OFFSET_CAL VDD CLK SINGLE_ENDED VIN_P VIN_N VCM VREF VREF_GND VSS
X0 a_13076_44458# a_13259_45724# a_13296_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2 VSS a_12427_45724# a_10490_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=361.2627 ps=3.22652k w=0.87 l=2.89
X5 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X7 VDD a_2903_42308# a_3080_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8 VDD a_12861_44030# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VSS a_1209_43370# a_n1557_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_16237_45028# a_16147_45260# a_16019_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VDD a_n755_45592# a_1176_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X13 a_6756_44260# a_5937_45572# a_6453_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X14 a_15868_43402# a_15681_43442# a_15781_43660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X15 a_n1533_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X16 a_8103_44636# a_8375_44464# a_8333_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 VSS a_16327_47482# a_16377_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 a_2437_43646# a_n443_46116# a_2437_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X20 a_n2810_45028# a_n2840_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X21 a_2113_38308# VDAC_Ni a_2112_39137# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X22 VDD a_3626_43646# a_19647_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 VSS a_10334_44484# a_10440_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_1576_42282# a_1755_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X25 a_10933_46660# a_10554_47026# a_10861_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 a_14021_43940# a_13483_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X27 a_16867_43762# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X29 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_n2840_43370# a_n2661_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X32 a_3457_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X33 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_14180_46482# a_14035_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X35 VSS a_18989_43940# a_19006_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X36 VSS a_9672_43914# a_2107_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X37 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VSS a_10695_43548# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X39 a_n2104_42282# a_n1925_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X40 a_20749_43396# a_12549_44172# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X41 VDD a_3877_44458# a_2382_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_n1699_44726# a_n1917_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X43 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X44 a_9241_45822# a_5066_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X45 VDD a_12883_44458# a_n2293_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X46 a_11909_44484# a_3232_43370# a_11827_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X47 a_835_46155# a_584_46384# a_376_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X48 a_5210_46155# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X49 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X50 VDD a_167_45260# a_1609_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 VSS a_526_44458# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 a_19268_43646# a_19319_43548# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X53 VSS a_22959_44484# a_19237_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X54 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X55 a_n2216_39072# a_n2312_39304# a_n2302_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X56 a_19987_42826# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X57 a_6151_47436# a_14311_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X58 a_8145_46902# a_7927_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X59 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X60 a_14275_46494# a_13925_46122# a_14180_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X61 a_20512_43084# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X62 a_14539_43914# a_17701_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X64 a_644_44056# a_626_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X65 a_10949_43914# a_12429_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X66 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X67 VSS a_21811_47423# a_20916_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X68 VDD a_3699_46634# a_3686_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X70 a_8035_47026# a_7411_46660# a_7927_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X71 a_5691_45260# a_5111_44636# a_5837_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X72 VDD a_1307_43914# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X73 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X74 a_18249_42858# a_18083_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 VDD a_104_43370# a_n971_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X76 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X77 a_3363_44484# a_1823_45246# a_3232_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X78 a_n1331_43914# a_n1549_44318# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X79 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X80 VSS a_n3565_39590# a_n3607_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X81 VSS a_12281_43396# a_12563_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X82 VSS a_22400_42852# a_22780_40081# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X83 VSS a_18780_47178# a_13661_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X84 a_n4318_39768# a_n2840_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X85 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X86 a_7230_45938# a_6472_45840# a_6667_45809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X87 VDD a_8049_45260# a_22959_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X88 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X89 a_8746_45002# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X90 a_15004_44636# a_11691_44458# a_15146_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X91 a_16223_45938# a_15599_45572# a_16115_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X92 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X93 a_n809_44244# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X94 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X95 a_17124_42282# a_17303_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X96 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X97 VSS a_3065_45002# a_2680_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X98 a_5193_42852# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X99 VDD a_6969_46634# a_6999_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X100 VDD a_10623_46897# a_10554_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X101 a_16137_43396# a_15781_43660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X102 VDD a_n2472_46634# a_n2442_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X103 VDD a_4185_45028# a_22959_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X104 a_15225_45822# a_15037_45618# a_15143_45578# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X105 VSS a_3537_45260# a_4640_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 a_n2012_43396# a_n2129_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X107 VDD a_n13_43084# a_n1853_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X108 a_5068_46348# a_n1151_42308# a_5210_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X109 a_873_42968# a_685_42968# a_791_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X110 a_17730_32519# a_22591_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X111 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X112 VDD a_22485_44484# a_20974_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X113 a_n1021_46688# a_n1151_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X114 VSS a_11599_46634# a_11735_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X115 a_13163_45724# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X116 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X117 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X118 a_n2012_44484# a_n2129_44697# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X119 a_13940_44484# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X120 VSS a_1414_42308# a_1525_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X121 a_8487_44056# a_4223_44672# a_8415_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X122 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X123 a_16434_46660# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X124 a_3315_47570# a_n1151_42308# a_2952_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X125 a_2680_45002# a_1823_45246# a_2903_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X126 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X127 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 a_22731_47423# SMPL_ON_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X129 VDD a_1307_43914# a_3681_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X130 a_n863_45724# a_1667_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 a_22521_40599# COMP_P VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X132 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X133 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X134 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X135 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=218.18214 ps=2.11206k w=0.55 l=0.59
X136 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X137 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X138 a_10467_46802# a_11599_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X139 VDD a_13747_46662# a_19862_44208# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X140 a_n2946_39866# a_n2956_39768# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X141 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X142 VSS a_15279_43071# a_14579_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X143 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X144 VSS a_8049_45260# a_22959_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X145 a_7584_44260# a_7542_44172# a_7281_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X146 a_n97_42460# a_19700_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X147 VDD a_19647_42308# a_13258_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X148 a_3754_39466# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X149 VSS a_2952_47436# a_2747_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X150 VDD a_16751_45260# a_6171_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X151 a_18326_43940# a_18079_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X152 a_9248_44260# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X153 a_3503_45724# a_3775_45552# a_3733_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X154 a_n2017_45002# a_19987_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X155 a_288_46660# a_171_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X156 a_10037_46155# a_9804_47204# a_9823_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X157 a_20075_46420# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X158 VDD a_196_42282# a_n3674_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X159 VSS a_14513_46634# a_14447_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X160 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X161 a_1149_42558# a_961_42354# a_1067_42314# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X162 a_13569_47204# a_13381_47204# a_13487_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X163 VDD a_14840_46494# a_15015_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X164 C6_P_btm a_n3565_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X165 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X166 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X167 a_14537_43396# a_14358_43442# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X168 VDD a_14955_47212# a_10227_46804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X169 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X170 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X171 a_n901_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X172 a_17668_45572# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X173 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X174 a_15493_43396# a_14955_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X175 a_7309_43172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X176 VDD a_1138_42852# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X177 a_1427_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X178 a_18184_42460# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X179 VDD a_13351_46090# a_10903_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X180 a_8379_46155# a_8128_46384# a_7920_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X181 VSS a_3483_46348# a_17325_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X182 VDD a_9290_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X183 VSS a_11823_42460# a_14358_43442# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X184 a_18310_42308# a_10193_42453# a_18220_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X185 VDD a_n2288_47178# a_n2312_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X186 a_17719_45144# a_16375_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VDD a_5891_43370# a_5147_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X188 a_7287_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X189 a_22609_38406# a_22469_39537# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X190 a_11173_44260# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X191 a_11897_42308# a_11823_42460# a_11551_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X192 VDD a_12861_44030# a_13759_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X193 a_19466_46812# a_19778_44110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X194 a_9049_44484# a_8701_44490# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X195 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X196 VDD a_16588_47582# a_16763_47508# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 a_9396_43370# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X198 C0_P_btm a_n784_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X199 a_n1736_42282# a_n1557_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X200 VDD a_14113_42308# a_16522_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X201 a_10651_43940# a_3090_45724# a_10555_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X202 VDD a_8667_46634# a_n237_47217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X203 a_6123_31319# a_7227_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X204 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X205 VSS a_n755_45592# a_1145_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X206 C7_P_btm a_5534_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X207 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X208 VSS a_n4064_37984# a_n2302_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X209 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X210 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X211 a_3581_42558# a_3539_42460# a_3497_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 a_n3674_38680# a_n2840_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X213 VSS a_5907_45546# a_5937_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X214 a_18783_43370# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X215 VSS a_1799_45572# a_1983_46706# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X216 VDD a_22959_46660# a_21076_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X217 VDD a_1736_39043# a_1239_39043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X218 a_13467_32519# a_21487_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X219 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X220 a_2864_46660# a_2747_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X221 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X222 a_8199_44636# a_10355_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X223 a_14403_45348# a_13259_45724# a_14309_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X224 a_556_44484# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X225 VSS a_15433_44458# a_15367_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X226 a_n1630_35242# a_564_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X227 a_n2840_43370# a_n2661_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X228 VSS a_13747_46662# a_13693_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X229 a_18245_44484# a_17767_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X230 a_19741_43940# a_19862_44208# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X231 a_16855_43396# a_16409_43396# a_16759_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X232 a_13113_42826# a_12895_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X233 VSS a_22365_46825# a_20202_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X234 a_n1079_45724# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X235 a_19386_47436# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X236 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X237 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X238 a_n89_47570# a_n237_47217# a_n452_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X239 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X240 a_1176_45822# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X241 a_10341_43396# a_9803_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X242 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=10.615 ps=76.96 w=3.75 l=15
X243 VDD a_n4209_38502# a_n4334_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X244 a_5111_42852# a_4905_42826# a_5193_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X245 a_13887_32519# a_22223_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X246 a_5437_45600# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X247 a_18953_45572# a_18909_45814# a_18787_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X248 VDD a_4791_45118# a_6165_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X249 VDD a_3429_45260# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X250 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X251 a_n3607_39616# a_n3674_39768# a_n3690_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X252 a_4842_47570# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X253 a_1337_46116# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X254 a_11136_45572# a_11322_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X255 a_n2661_42834# a_10809_44734# a_12189_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X256 VSS a_10249_46116# a_11186_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X257 a_16655_46660# a_n743_46660# a_16292_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X258 a_n1991_46122# a_n2157_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X259 VREF_GND a_n3420_39072# C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X260 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X261 VDD a_1576_42282# a_1606_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X262 a_5159_47243# a_n443_46116# a_4700_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X263 VSS a_5891_43370# a_8375_44464# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X264 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VDD a_13076_44458# a_12883_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X266 VSS a_14539_43914# a_14485_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X267 VDD en_comp a_1177_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X268 C0_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X269 a_15297_45822# a_11823_42460# a_15225_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X270 a_18479_47436# a_20075_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X271 a_1423_45028# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X272 a_2382_45260# a_3877_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X273 a_8103_44636# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X274 a_n1899_43946# a_n2065_43946# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 a_6765_43638# a_6547_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X276 a_n2293_43922# a_12741_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X277 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X278 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X279 a_945_42968# a_n1059_45260# a_873_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X280 VDD a_3785_47178# a_3815_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X281 VDD a_14084_46812# a_14035_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X282 a_765_45546# a_12549_44172# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X283 VDD a_20974_43370# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X284 a_14275_46494# a_13759_46122# a_14180_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X285 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 a_1609_45822# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X287 a_17517_44484# a_16979_44734# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X288 VDD a_4915_47217# a_12891_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 a_20679_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X290 VSS a_1423_45028# a_9838_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X291 a_13921_42308# a_13259_45724# a_13575_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X292 VCM a_n784_42308# C0_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X293 VSS a_11599_46634# a_13759_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X294 a_14127_45572# a_11823_42460# a_14033_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X295 a_13569_43230# a_12379_42858# a_13460_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X296 a_5072_46660# a_4955_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X297 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X298 a_8037_42858# a_7871_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X299 VSS a_22591_46660# a_20820_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X301 a_3686_47026# a_2609_46660# a_3524_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X302 a_9672_43914# a_10057_43914# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X303 VDD a_18429_43548# a_16823_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X304 a_17339_46660# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 VSS a_1606_42308# a_2351_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X306 a_16409_43396# a_16243_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 VSS a_9625_46129# a_10044_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X308 VDD a_n4209_37414# a_n4334_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X309 a_13468_44734# a_768_44030# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X310 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_2124_47436# a_584_46384# a_2266_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X312 VDD a_n971_45724# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X313 a_10809_44734# a_2063_45854# a_10809_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X314 a_7577_46660# a_7411_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4921_42308# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_16023_47582# a_15507_47210# a_15928_47570# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X317 a_12791_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X318 a_10193_42453# a_20712_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X319 VSS a_n881_46662# a_n659_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 a_6481_42558# a_n913_45002# a_1755_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X321 a_n2956_38680# a_n2472_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X322 a_14955_43940# a_14537_43396# a_15037_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X323 VREF_GND a_14097_32519# C4_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X324 VDD a_21188_45572# a_21363_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X326 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 a_18907_42674# a_18727_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X328 a_12545_42858# a_12379_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X330 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X331 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X332 a_13720_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X333 a_15125_43396# a_15095_43370# a_15037_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X334 VREF a_20692_30879# C6_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X335 a_2998_44172# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X336 a_20974_43370# a_22485_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X337 a_18548_42308# a_18494_42460# a_18057_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X338 a_n875_44318# a_n2065_43946# a_n984_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X339 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X340 a_n2293_42834# a_8049_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X341 VSS a_4743_44484# a_4791_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X342 a_3626_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X343 VSS a_n2438_43548# a_n2433_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X344 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X345 VDD a_17973_43940# a_18079_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X346 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X347 VREF_GND a_17538_32519# C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X348 VDD a_22223_46124# a_20205_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X349 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X350 a_4704_46090# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X351 a_5815_47464# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X352 a_17478_45572# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X353 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X354 a_22609_38406# a_22521_39511# CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X355 VSS a_19864_35138# a_21589_35634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X356 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X357 a_17034_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X358 VSS a_n3420_39616# a_n2946_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X359 a_133_42852# a_n97_42460# a_n13_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X360 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X361 a_n1925_46634# a_8162_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X362 a_21350_47026# a_20273_46660# a_21188_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X363 VDD a_2713_42308# a_2903_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X364 a_n3674_39304# a_n2840_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X365 a_13565_43940# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X366 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VDD a_1823_45246# a_2202_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X368 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X369 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X370 a_2211_45572# a_2063_45854# a_1848_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X371 VSS a_16112_44458# a_14673_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X372 VSS a_3316_45546# a_3260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X373 VDD a_n443_46116# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X374 a_n310_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X375 a_21177_47436# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X376 VSS a_9290_44172# a_13943_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X377 a_n3674_37592# a_196_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X378 a_18780_47178# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X379 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X380 VSS a_8791_42308# a_5934_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X381 a_421_43172# a_n97_42460# a_n13_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X382 VDD a_17339_46660# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X383 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X384 VSS a_n2840_46090# a_n2956_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X385 a_n2661_43370# a_10907_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X386 a_9396_43370# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X387 VDD a_19333_46634# a_19123_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X388 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X389 a_5755_42852# a_n97_42460# a_5837_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X390 a_n4251_39392# a_n4318_39304# a_n4334_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X391 a_805_46414# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X392 VDD a_n1076_43230# a_n901_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X393 a_21845_43940# a_12549_44172# a_19692_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X394 VDD a_4520_42826# a_4093_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X395 a_12469_46902# a_12251_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X396 a_15415_45028# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X397 a_19479_31679# a_22223_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X398 a_7542_44172# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X399 a_3080_42308# a_2903_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X400 VSS a_22165_42308# a_22223_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X401 VDD a_10249_46116# a_11186_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X402 a_3905_42558# a_2382_45260# a_3823_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X403 a_12347_46660# a_11901_46660# a_12251_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X404 VSS a_16137_43396# a_16414_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X405 a_5066_45546# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X406 a_14581_44484# a_13249_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X407 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X408 a_2113_38308# a_1343_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X409 a_n473_42460# a_n755_45592# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X410 VDD a_n1699_43638# a_n1809_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X411 a_13759_47204# a_13717_47436# a_13675_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X412 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X413 C4_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X414 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X415 a_2779_44458# a_1423_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X416 VDD a_19319_43548# a_19268_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X417 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X418 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X419 a_1123_46634# a_948_46660# a_1302_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X420 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 a_2952_47436# a_3160_47472# a_3094_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X422 a_5807_45002# a_16763_47508# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X423 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X424 a_6293_42852# a_5755_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X425 a_8120_45572# a_8034_45724# a_n1925_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X426 a_11541_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X427 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X428 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X429 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 a_5257_43370# a_5907_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X432 a_4880_45572# a_5066_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X433 VIN_P EN_VIN_BSTR_P C0_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X434 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X435 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X436 a_3497_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X437 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X438 a_16223_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X439 a_4883_46098# a_21363_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X440 a_2711_45572# a_768_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X441 VSS a_2553_47502# a_2487_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X442 VDD a_12469_46902# a_12359_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X443 a_6453_43914# a_6109_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X444 a_7765_42852# a_7227_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X445 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X446 a_17786_45822# a_15861_45028# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X447 a_18450_45144# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X448 a_6765_43638# a_6547_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X449 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X450 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X451 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X452 a_12089_42308# a_11551_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X453 a_16547_43609# a_16414_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X454 a_3221_46660# a_3177_46902# a_3055_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X455 a_6667_45809# a_6472_45840# a_6977_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X456 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X457 a_6643_43396# a_6197_43396# a_6547_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X458 a_5837_45348# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X459 a_5565_43396# a_4905_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X460 a_7418_45067# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X461 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X462 a_1793_42852# a_742_44458# a_1709_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 VDD a_10227_46804# a_10083_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X464 a_11301_43218# a_10922_42852# a_11229_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X465 VSS a_13291_42460# a_13249_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X466 a_18341_45572# a_18175_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X467 a_19113_45348# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X468 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X469 a_8696_44636# a_16855_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X470 a_12189_44484# a_8975_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X471 a_n1736_46482# a_n1853_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X472 a_1239_47204# a_1209_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X473 VDD VDAC_Ni a_6886_37412# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X474 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X475 a_1606_42308# a_1576_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X476 VDD a_n443_42852# a_6481_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X477 VDD a_12005_46116# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X478 a_18315_45260# a_18587_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X479 VSS a_768_44030# a_3600_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X480 VDD a_4958_30871# a_17531_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X481 a_16795_42852# a_n97_42460# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X482 a_18900_46660# a_18834_46812# a_18285_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X483 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X484 a_17973_43940# a_17737_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X485 VSS a_22821_38993# a_22876_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X486 a_6419_46155# a_5257_43370# a_6347_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X487 a_18597_46090# a_19431_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X488 a_3737_43940# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X489 VDD a_1823_45246# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X490 EN_VIN_BSTR_P VDD a_n1386_35608# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X491 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X492 VSS a_21496_47436# a_13507_46334# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X493 VSS a_10723_42308# a_5742_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X494 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X495 VSS a_n4209_38216# a_n4251_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X496 a_12891_46348# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X497 VSS a_20679_44626# a_20640_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X498 a_21115_43940# a_20935_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X499 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X500 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X501 VDD a_10951_45334# a_10775_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X502 a_20850_46155# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X503 VDD a_13661_43548# a_18587_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X504 a_11649_44734# a_3232_43370# a_n2661_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X505 a_20820_30879# a_22591_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X506 VSS a_21359_45002# a_21101_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X507 a_17364_32525# a_22959_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X508 a_18989_43940# a_18451_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X509 a_6197_43396# a_6031_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X510 EN_VIN_BSTR_P VDD a_n83_35174# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X511 VDD a_12891_46348# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X512 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X513 VREF_GND a_13467_32519# C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X514 VDD a_584_46384# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X515 a_8873_43396# a_5891_43370# a_8791_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X516 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X517 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X518 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X519 a_10809_44484# a_10057_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X520 C6_N_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X521 a_6545_47178# a_6419_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X522 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X523 a_6109_44484# a_5518_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X524 a_n4318_38216# a_n2472_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X525 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X526 a_13258_32519# a_19647_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X527 VDD a_11599_46634# a_18819_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X528 a_n1435_47204# a_n1605_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X529 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X530 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X531 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X532 a_14113_42308# a_13575_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X533 VSS a_4646_46812# a_4651_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X534 a_13381_47204# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X535 VSS a_n2472_46090# a_n2956_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X536 a_4958_30871# a_17124_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X537 VSS a_22223_42860# a_22400_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X538 C0_P_btm a_n3565_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X539 VDD a_1208_46090# a_472_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X540 VSS a_18479_47436# a_19452_47524# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X541 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X542 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X543 a_22545_38993# a_22459_39145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X544 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X545 a_20623_45572# a_20107_45572# a_20528_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X546 a_12281_43396# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X547 C1_P_btm a_n4209_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X548 VSS a_n3565_39304# a_n3607_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X549 a_15486_42560# a_15764_42576# a_15720_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X550 VSS a_n1613_43370# a_8649_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X551 a_15765_45572# a_15599_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X552 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X553 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X554 VSS a_14495_45572# a_n881_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X555 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X556 a_10617_44484# a_10440_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X557 VDD a_5111_44636# a_8487_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X558 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X559 VCM a_5932_42308# C3_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X560 a_20708_46348# a_15227_44166# a_20850_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X561 a_n2267_44484# a_n2433_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X562 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X563 a_1115_44172# a_453_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X564 VSS COMP_P a_n1329_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X565 VSS a_1847_42826# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X566 VSS a_15861_45028# a_17023_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X567 a_16292_46812# a_5807_45002# a_16434_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X568 a_17325_44484# a_15227_44166# a_16979_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X569 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X570 a_15803_42450# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X571 a_5534_30871# a_12563_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X572 VSS a_3381_47502# a_3315_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X573 VDD a_9863_46634# a_2063_45854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X574 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X575 VDD a_n2840_43370# a_n4318_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X576 VSS a_584_46384# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X577 VIN_N EN_VIN_BSTR_N C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X578 a_3863_42891# a_3681_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X579 VDD a_9049_44484# a_9313_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X580 VDD a_376_46348# a_171_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X581 a_11541_44484# a_11453_44696# a_n2661_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X582 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X583 a_19553_46090# a_19335_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X584 a_21589_35634# a_19864_35138# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X585 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X586 a_18727_42674# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X587 a_n1925_42282# a_4185_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X588 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X589 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X590 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X591 VDD a_19164_43230# a_19339_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X592 a_2479_44172# a_2905_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X593 VSS a_4361_42308# a_21855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X594 a_n1741_47186# a_12891_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X595 VDD a_8103_44636# a_7640_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X596 a_8192_45572# a_8162_45546# a_8120_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X597 a_5009_45028# a_3090_45724# a_4927_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X598 a_12549_44172# a_20567_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X599 VSS a_n2840_42282# a_n3674_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 a_5129_47502# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X601 a_14840_46494# a_13759_46122# a_14493_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X602 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X603 VSS a_n913_45002# a_2713_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X604 VDD a_n863_45724# a_1221_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X605 a_8601_46660# a_7411_46660# a_8492_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X606 a_2307_45899# a_n237_47217# a_1848_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X607 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X608 VDD a_n4209_39304# a_n4334_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X609 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X610 a_n2946_39072# a_n2956_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X611 a_15861_45028# a_15595_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X612 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X613 VSS a_n1613_43370# a_3221_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X614 a_1756_43548# a_768_44030# a_1987_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X615 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X616 a_3754_39134# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X617 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X618 a_n4318_40392# a_n2840_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X619 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X620 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X621 a_19332_42282# a_19511_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X622 VSS a_17583_46090# a_13259_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X623 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X624 a_20623_43914# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X625 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X626 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X627 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X628 a_4185_45348# a_3065_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X629 a_n2661_46634# a_13017_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X630 VDD a_19321_45002# a_20567_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X631 VDD a_6545_47178# a_6575_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 VDD a_18285_46348# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X633 a_2864_46660# a_2747_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X634 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X635 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X636 VDD a_1307_43914# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X637 a_13351_46090# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X638 a_18374_44850# a_18248_44752# a_17970_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X639 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X640 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X641 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X642 a_13657_42308# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X643 a_375_42282# a_413_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X644 a_3090_45724# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X645 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X646 a_10334_44484# a_10157_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X647 VSS a_10903_43370# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X648 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X649 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X650 VSS a_n2438_43548# a_n133_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X651 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X652 VSS a_22959_46124# a_20692_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X653 a_n3674_39768# a_n2472_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X654 VREF a_n4209_39304# C7_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X655 VSS a_20107_42308# a_7174_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X656 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X657 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X658 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X659 a_20301_43646# a_19692_46634# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X660 VDD a_n901_46420# a_n914_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X661 a_n971_45724# a_104_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X662 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X663 a_20447_31679# a_22959_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X664 VSS a_13348_45260# a_13159_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X665 a_n4334_38304# a_n4318_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X666 VSS a_n881_46662# a_6517_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X667 a_8685_42308# a_8515_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X668 VSS a_6491_46660# a_6851_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X669 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X670 VDD a_14493_46090# a_14383_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X671 a_n327_42308# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X672 a_22485_44484# a_22315_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X673 a_15673_47210# a_15507_47210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X674 a_8605_42826# a_8387_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X675 a_1709_42852# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X676 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X677 VDD a_n1736_42282# a_n4318_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X678 VREF a_19721_31679# C2_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X679 VSS a_895_43940# a_2537_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X680 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X681 a_17609_46634# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 VDD a_11599_46634# a_18175_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X683 a_8945_43396# a_3537_45260# a_8873_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X684 a_13249_42308# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X685 a_601_46902# a_383_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X686 a_4640_45348# a_4574_45260# a_4558_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X687 a_n467_45028# a_n745_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X688 a_1208_46090# a_765_45546# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X689 a_3820_44260# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X690 VSS a_n863_45724# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 VSS a_16721_46634# a_16655_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X692 C5_P_btm a_n4064_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X693 a_21588_30879# a_22223_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X694 a_16877_42852# a_16823_43084# a_16795_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X695 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X696 VSS a_17715_44484# a_17737_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X697 a_16241_47178# a_16023_47582# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X698 a_12359_47026# a_11735_46660# a_12251_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X699 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X700 a_5883_43914# a_8333_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X701 a_16759_43396# a_16409_43396# a_16664_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X702 a_22876_39857# a_22545_38993# a_22780_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X703 VDD a_n3565_39590# a_n3690_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X704 a_17665_42852# a_17595_43084# a_14539_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X705 VSS a_n2438_43548# a_n2157_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X706 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X707 a_1990_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X708 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X709 a_5072_46660# a_4955_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X710 VDD a_3357_43084# a_22591_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X711 VSS a_3815_47204# a_4007_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X712 a_1736_39587# a_1736_39043# a_2112_39137# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X713 a_15803_42450# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X714 a_20528_46660# a_20411_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X715 a_n1838_35608# a_n1386_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X716 a_n3607_39392# a_n3674_39304# a_n3690_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X717 VDD a_n4064_39616# a_n2216_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X718 a_21421_42336# a_16327_47482# a_21335_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X719 a_6655_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X720 a_14371_46494# a_13925_46122# a_14275_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X721 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X722 VDD a_3503_45724# a_3218_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X723 VDD a_n2840_43914# a_n4318_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X724 a_15037_43940# a_13556_45296# a_14955_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X725 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X726 VDD a_10467_46802# a_10428_46928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X727 a_15060_45348# a_13661_43548# a_14976_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X728 a_9895_44260# a_9290_44172# a_9801_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X729 VDD a_6171_42473# a_5379_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X730 a_5009_45028# a_5147_45002# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X731 a_13904_45546# a_10903_43370# a_14127_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X732 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X733 a_19900_46494# a_18985_46122# a_19553_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X734 VDD a_8696_44636# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X735 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X736 a_3935_42891# a_3905_42865# a_3863_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X737 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X738 VSS a_n881_46662# a_11117_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X739 C3_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X740 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X741 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X742 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X743 a_1057_46660# a_n133_46660# a_948_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X744 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X745 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X746 VSS a_2982_43646# a_21487_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X747 a_21363_45546# a_21188_45572# a_21542_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X748 VSS a_11823_42460# a_11322_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 a_18204_44850# a_17767_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X750 a_n447_43370# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X751 a_17324_43396# a_16409_43396# a_16977_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X752 VSS a_n4064_38528# a_n2302_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X753 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X754 a_15095_43370# a_15567_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X755 a_10150_46912# a_10428_46928# a_10384_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X756 VSS a_n2472_42282# a_n4318_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X757 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X758 a_8492_46660# a_7577_46660# a_8145_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X759 a_5649_42852# a_5111_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X760 VDD a_18287_44626# a_18248_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X761 a_20894_47436# a_20990_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X762 a_19636_46660# a_19594_46812# a_19333_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X763 a_10249_46116# a_9823_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X764 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X765 a_10227_46804# a_14955_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X766 a_739_46482# a_n743_46660# a_376_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X767 VSS a_10775_45002# a_10180_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X768 a_2896_43646# a_2479_44172# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X769 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X770 a_12791_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X771 VSS a_5807_45002# a_11691_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X772 VSS a_3357_43084# a_22591_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X773 VSS a_2382_45260# a_2304_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X774 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X775 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X776 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X777 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X778 VDD a_2277_45546# a_2307_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X779 a_10053_45546# a_8746_45002# a_10306_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X780 a_n2956_39768# a_n2840_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X781 VDD a_4361_42308# a_21855_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X782 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X783 VSS a_6945_45028# a_22223_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X784 VDD a_5257_43370# a_5263_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X787 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X788 a_18494_42460# a_18907_42674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X789 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X790 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X791 a_n1151_42308# a_n1329_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X792 a_16763_47508# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X793 a_21259_43561# a_4190_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X794 a_8349_46414# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X795 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X796 a_17970_44736# a_18287_44626# a_18245_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X797 a_1123_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X798 a_n237_47217# a_8667_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X799 a_5837_42852# a_3537_45260# a_5755_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X800 VSS a_19692_46634# a_19636_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X801 a_8697_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X802 a_1145_45348# a_n863_45724# a_626_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X803 VSS a_5934_30871# a_8515_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X804 VSS a_1239_47204# a_1431_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X805 a_22705_38406# a_22521_40055# a_22609_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X806 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X807 a_11173_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X808 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X809 a_22165_42308# a_21887_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X810 a_5244_44056# a_5147_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X811 VSS a_n4064_37440# a_n2302_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X812 VDD a_8952_43230# a_9127_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X813 a_n2956_37592# a_n2472_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X814 VSS a_2127_44172# a_n2661_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X815 VSS a_15493_43940# a_22959_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X816 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X817 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X818 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X819 a_19339_43156# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X820 VDD a_n1920_47178# a_n2312_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X821 VDD a_n1177_44458# a_n1190_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X822 VDD a_16292_46812# a_15811_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X823 a_5164_46348# a_4927_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X824 a_9482_43914# a_9838_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X825 a_20835_44721# a_20679_44626# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X826 VSS a_5937_45572# a_8781_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X827 a_5837_42852# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X828 a_10037_47542# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X829 a_7221_43396# a_6031_43396# a_7112_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X830 VSS a_5937_45572# a_8560_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X831 C7_N_btm a_20820_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X832 VSS a_15559_46634# a_13059_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X833 a_5385_46902# a_5167_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X834 VDD a_10334_44484# a_10440_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X835 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X836 a_19597_46482# a_19553_46090# a_19431_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X837 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X838 a_18051_46116# a_18189_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X839 a_15493_43940# a_14955_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X840 a_16414_43172# a_n1059_45260# a_16328_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X841 a_21297_46660# a_20107_46660# a_21188_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X842 a_11813_46116# a_11387_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X843 VSS SMPL_ON_P a_n1605_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X844 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X845 a_5894_47026# a_4817_46660# a_5732_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X846 VDD a_4699_43561# a_3539_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X847 VSS a_n3420_39072# a_n2946_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X848 VDD a_n97_42460# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X849 VDD a_13163_45724# a_11962_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X850 a_15433_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X851 VDD a_16327_47482# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X852 a_18114_32519# a_22223_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X853 a_n452_44636# a_n1151_42308# a_n310_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X854 VDD a_22959_43396# a_17364_32525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X855 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X856 VDD a_1307_43914# a_4149_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X857 VSS a_n357_42282# a_7573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X858 VDD a_9863_47436# a_9804_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X859 a_22821_38993# a_22400_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X860 a_3754_39134# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X861 a_4649_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X862 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X863 VSS a_1848_45724# a_1799_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X864 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X865 a_20885_45572# a_20841_45814# a_20719_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X866 a_10554_47026# a_10428_46928# a_10150_46912# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X867 a_n746_45260# a_n1177_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X868 a_7_44811# a_n1151_42308# a_n452_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X869 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X870 VDD a_10355_46116# a_8199_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X871 a_4181_43396# a_4093_43548# a_n2661_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X872 VDD a_2437_43646# a_22223_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X873 a_21005_45260# a_21101_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X874 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X875 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X876 a_3754_38802# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X877 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X878 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X879 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X880 VSS a_12861_44030# a_17339_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X881 VDD a_n2840_45002# a_n2810_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X882 a_10057_43914# a_10807_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X883 a_5343_44458# a_7963_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X884 a_n1423_42826# a_n1641_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X885 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X886 VDD a_11827_44484# a_22223_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X887 VDD a_n2472_43914# a_n3674_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X888 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X889 a_6945_45028# a_5937_45572# a_6945_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X890 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X891 a_20301_43646# a_13661_43548# a_743_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X892 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X893 a_n2216_39866# a_n2442_46660# a_n2302_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X894 VDD a_22000_46634# a_15227_44166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X895 VSS a_2889_44172# a_413_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X896 VSS a_n97_42460# a_n144_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X897 a_n3674_38216# a_n2104_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X898 a_16321_45348# a_1307_43914# a_16019_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X899 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X900 VDD a_9290_44172# a_13070_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X901 a_133_42852# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X902 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X903 VDD a_22465_38105# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X904 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X905 a_n2860_38778# a_n2956_38680# a_n2946_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X906 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X907 a_6517_45366# a_5937_45572# a_6431_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X908 a_10555_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X909 VDD a_5111_44636# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X910 a_14401_32519# a_22223_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X911 VSS a_9290_44172# a_13070_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X912 VSS a_5068_46348# a_4955_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X913 VDD a_9290_44172# a_10586_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X914 a_16751_45260# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X915 a_1736_39587# a_1736_39043# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X916 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X917 VSS a_11599_46634# a_15507_47210# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X918 VSS a_768_44030# a_644_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X919 a_12465_44636# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X920 VDD a_n357_42282# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X921 a_5193_43172# a_3905_42865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X922 VSS a_18783_43370# a_18525_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X923 a_3540_43646# a_1414_42308# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X924 a_21363_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X925 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X926 a_5421_42558# a_5379_42460# a_5337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X927 VDD a_12861_44030# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X928 a_n2956_38216# a_n2472_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X929 a_13885_46660# a_13607_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X930 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X931 a_2232_45348# a_1609_45822# a_n2293_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X932 a_5691_45260# a_6171_45002# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X933 a_9801_44260# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X934 VCM a_3080_42308# C2_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X935 a_327_44734# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X936 VSS a_7499_43078# a_8746_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X937 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X938 a_15743_43084# a_19339_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X939 VSS a_22591_43396# a_14209_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X940 VSS a_2437_43646# a_22223_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X941 a_6547_43396# a_6197_43396# a_6452_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X942 a_20556_43646# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X943 a_1987_43646# a_742_44458# a_1891_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X944 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X945 a_648_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X946 VDD a_n23_47502# a_7_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X947 a_17609_46634# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X948 a_3602_45348# a_3537_45260# a_3495_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X949 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X950 VDD a_2982_43646# a_21487_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X951 a_13661_43548# a_18780_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X952 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X953 a_9313_44734# a_3232_43370# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X954 C6_P_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X955 a_11323_42473# a_5742_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X956 a_14383_46116# a_13759_46122# a_14275_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X957 a_2813_43396# a_2479_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X958 a_16721_46634# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X959 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X960 VDD a_526_44458# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X961 VREF a_20820_30879# C7_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X962 VDD a_15681_43442# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X963 a_6125_45348# a_3232_43370# a_5691_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X964 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X965 a_10907_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X966 a_14955_43396# a_9145_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X967 a_8128_46384# a_7903_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X968 a_3429_45260# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X969 VDD a_15227_44166# a_17969_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X970 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X971 a_n2860_37690# a_n2956_37592# a_n2946_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X972 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X973 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X974 C4_P_btm a_n3420_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X975 a_18599_43230# a_18083_42858# a_18504_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X976 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X977 a_18057_42282# a_18494_42460# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X978 a_11117_47542# a_4915_47217# a_11031_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X979 VDD a_22400_42852# a_22521_40599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X980 a_7112_43396# a_6197_43396# a_6765_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X981 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X982 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X983 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X984 a_19240_46482# a_19123_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X985 VCM a_5742_30871# C6_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X986 VSS a_10193_42453# a_10149_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X987 VDD a_10193_42453# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X988 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X989 VSS a_n967_45348# a_n961_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X990 a_564_42282# a_743_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X991 a_21195_42852# a_20922_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X992 VDD a_6575_47204# a_9067_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X993 a_22612_30879# a_22959_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X994 a_21188_46660# a_20273_46660# a_20841_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X995 a_13749_43396# a_13661_43548# a_13667_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X996 VSS a_n2840_45546# a_n2810_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X997 a_13490_45394# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X998 a_n2840_43914# a_n2661_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X999 a_n822_43940# a_n1899_43946# a_n984_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1000 a_21613_42308# a_21335_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1001 a_7112_43396# a_6031_43396# a_6765_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1002 a_14537_43396# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1003 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1004 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1005 a_n23_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1006 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1007 a_14543_43071# a_5534_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1008 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1009 VDD a_19900_46494# a_20075_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1010 VDD a_7227_45028# a_7230_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1011 VSS a_16327_47482# a_19597_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1012 a_9823_46155# a_n743_46660# a_9751_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1013 VDD a_22959_43948# a_17538_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1014 a_18214_42558# a_16137_43396# a_18057_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1015 a_n3690_38304# a_n3674_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1016 a_15009_46634# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1017 a_17591_47464# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1018 VSS a_10227_46804# a_15521_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1019 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1020 a_22485_44484# a_22315_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1021 a_n1644_44306# a_n1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1022 VDD RST_Z a_8530_39574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1023 VDD a_n1329_42308# a_n1151_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1024 VSS a_13507_46334# a_18184_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1025 a_n630_44306# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1026 a_18783_43370# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1027 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1028 VSS a_22521_40599# a_22469_40625# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1029 a_8325_42308# a_n913_45002# a_8337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1030 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X1031 a_21973_42336# a_20202_43084# a_21887_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1032 VSS a_n1613_43370# a_645_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1033 a_10341_42308# a_9803_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1034 a_n1920_47178# a_n1741_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1035 VSS a_16327_47482# a_20885_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1036 VSS a_10807_43548# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1037 VSS a_5257_43370# a_3905_42865# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1038 a_9127_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1039 VDD a_n2472_45002# a_n2956_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1040 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1041 a_13259_45724# a_17583_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1042 VSS a_10586_45546# a_10544_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X1043 a_16751_45260# a_17023_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1044 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1045 VSS a_n4209_38502# a_n4251_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1046 VSS a_7227_42308# a_6123_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1047 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1048 a_n2840_42826# a_n2661_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1049 a_1302_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1050 a_5907_45546# a_6194_45824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1051 a_13059_46348# a_15559_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1052 a_n2302_37984# a_n2810_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1053 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1054 VREF_GND a_14209_32519# C5_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1055 a_3065_45002# a_3318_42354# a_3581_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1056 a_16023_47582# a_15673_47210# a_15928_47570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1057 VSS a_n881_46662# a_n935_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1058 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1059 C6_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1060 VDD a_21487_43396# a_13467_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1061 a_2553_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1062 VDD a_n443_42852# a_997_45618# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 a_8568_45546# a_8199_44636# a_8791_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1064 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1065 a_13635_43156# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1066 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1067 VDD a_564_42282# a_n1630_35242# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1068 a_n473_42460# a_n971_45724# a_n327_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1069 a_16335_44484# a_13661_43548# a_16241_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1070 VDD a_15861_45028# a_17023_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1071 a_5205_44734# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1072 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1073 VSS a_1123_46634# a_1057_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1074 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1075 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1076 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1077 VSS a_13259_45724# a_18315_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1078 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1079 VSS a_22223_43396# a_13887_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1080 a_11682_45822# a_11322_45546# a_11525_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1081 VDD a_22591_45572# a_19963_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1082 a_5934_30871# a_8791_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1083 a_18429_43548# a_18525_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1084 a_509_45822# a_n1099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1085 a_20980_44850# a_20766_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1086 a_4190_30871# a_19332_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1087 a_3381_47502# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1088 VDD a_3537_45260# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1089 a_6682_46660# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1090 a_20273_45572# a_20107_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1091 VDD a_11963_45334# a_11787_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1092 VDD a_1423_45028# a_9838_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1093 a_19256_45572# a_18175_45572# a_18909_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1094 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1095 VSS a_3699_46634# a_3633_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1096 VSS a_5937_45572# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1097 a_14226_46987# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1098 VSS a_n2438_43548# a_n2157_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1099 VSS a_8953_45546# a_9241_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1100 a_n2840_45002# a_n2661_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1101 a_n722_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1102 a_12005_46436# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1103 a_9885_43396# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1104 VSS a_n4209_37414# a_n4251_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1105 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1106 a_18817_42826# a_18599_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1107 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1108 VDD a_167_45260# a_1423_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1109 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1110 VSS a_4704_46090# a_1823_45246# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1111 a_16886_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X1112 a_11688_45572# a_11652_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X1113 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1114 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1115 a_4520_42826# a_1823_45246# a_4743_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1116 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1117 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1118 VDD a_n2104_42282# a_n3674_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1119 VDD RST_Z a_14311_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1120 a_19721_31679# a_22959_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1121 a_458_43396# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X1122 a_19339_43156# a_19164_43230# a_19518_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1123 a_11453_44696# a_17719_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1124 a_22717_36887# a_22459_39145# a_22609_37990# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1125 VDD a_n3420_37984# a_n2860_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1126 a_13711_45394# a_12891_46348# a_13348_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1127 a_16664_43396# a_16547_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1128 a_1138_42852# a_791_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1129 a_21259_43561# a_4190_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1130 a_10586_45546# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1131 VSS a_11599_46634# a_15599_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1132 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1133 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1134 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1135 a_196_42282# a_375_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1136 VSS a_n881_46662# a_7989_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1137 a_7832_46660# a_7715_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1138 VDD a_n2109_45247# en_comp VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1139 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1140 a_15928_47570# a_15811_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1141 a_3633_46660# a_2443_46660# a_3524_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1142 VSS a_n2472_45546# a_n2956_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1143 a_2127_44172# a_2675_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1144 a_9885_43646# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1145 a_n2472_43914# a_n2293_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1146 VDD a_12991_46634# a_12978_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1147 VDD a_1667_45002# a_n863_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1148 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1149 a_14084_46812# a_n1151_42308# a_14226_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1150 a_5837_45028# a_3232_43370# a_5691_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X1151 VDD a_21195_42852# a_21671_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1152 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1153 a_12427_45724# a_12791_45546# a_12749_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1154 VSS a_n913_45002# a_4921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 a_14209_32519# a_22591_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1156 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1157 a_12553_44484# a_12465_44636# a_n2661_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1159 a_5829_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1160 a_16237_45028# a_n743_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1161 VDD a_22959_45036# a_19721_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1162 a_14761_44260# a_14673_44172# a_n2293_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1163 VSS a_n1613_43370# a_5429_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1164 VSS a_21363_46634# a_21297_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1165 VDD a_n452_45724# a_n1853_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1166 VDD a_584_46384# a_2998_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1167 VSS a_4699_43561# a_3539_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1168 VDD a_15959_42545# a_15890_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1169 VSS a_10227_46804# a_13157_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1170 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1171 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1172 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1173 a_17538_32519# a_22959_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1174 a_n144_43396# a_n971_45724# a_n447_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1175 a_16680_45572# a_15599_45572# a_16333_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1176 VSS a_5937_45572# a_6101_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1177 a_9672_43914# a_8199_44636# a_9895_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1178 a_15231_43396# a_9145_43396# a_15125_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1179 a_8387_43230# a_7871_42858# a_8292_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1180 VDD a_22731_47423# a_13717_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1181 VDD a_9290_44172# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1182 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1183 VDD a_10903_43370# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X1184 VDD a_17767_44458# a_17715_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1185 VDD a_7845_44172# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X1186 a_n2840_44458# a_n2661_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1187 a_22400_42852# a_22223_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1188 VDD a_n863_45724# a_945_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1189 VSS a_9482_43914# a_10157_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1190 VDD a_12549_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X1191 a_4933_42558# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_19333_46634# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1193 a_13565_44260# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1194 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1195 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1196 a_n2293_46098# a_5663_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1197 VSS a_11453_44696# a_22959_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1198 VSS a_12563_42308# a_5534_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1199 a_n2472_42826# a_n2293_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1200 a_7920_46348# a_8128_46384# a_8062_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1201 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1202 a_n13_43084# a_n443_42852# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1203 a_2698_46116# a_2521_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1204 a_15785_43172# a_15743_43084# a_15095_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1205 a_8654_47026# a_7577_46660# a_8492_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1206 VDD a_21363_46634# a_21350_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1207 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1208 VDD a_n809_44244# a_n822_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1209 a_766_43646# a_626_44172# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X1210 a_n784_42308# a_n961_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1211 a_12895_43230# a_12379_42858# a_12800_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1212 VSS a_805_46414# a_739_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1213 VSS a_8191_45002# a_8137_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1214 a_15959_42545# a_15803_42450# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1215 a_5210_46482# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1216 a_11341_43940# a_3232_43370# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1217 VDD a_7705_45326# a_7735_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1218 a_13720_44458# a_13661_43548# a_13940_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1219 a_2162_46660# a_2107_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1220 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1221 a_n1423_42826# a_n1641_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1222 a_n2956_39304# a_n2840_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1223 VDD a_11415_45002# a_n2661_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1224 a_15037_43940# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1225 VDD a_1606_42308# a_2351_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1226 a_2277_45546# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1227 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1228 a_6903_46660# a_6755_46942# a_6540_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1229 VDD a_14180_45002# a_13017_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1230 a_3232_43370# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1231 a_22521_40055# en_comp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1232 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1233 VDD a_8199_44636# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1234 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1235 a_1576_42282# a_1755_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1236 a_7573_43172# a_7499_43078# a_7227_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1237 VSS a_21855_43396# a_13678_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1238 VDD a_18989_43940# a_19006_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1239 VSS a_6540_46812# a_6491_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1240 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1241 VDD a_22223_45572# a_19479_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1242 VIN_N EN_VIN_BSTR_N C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1243 VSS a_2903_42308# a_3080_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 VSS a_n863_45724# a_n906_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1245 a_n2840_44458# a_n2661_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1246 a_3823_42558# a_3065_45002# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1247 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1248 VSS a_5263_45724# a_5204_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1249 VDD a_2124_47436# a_1209_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1250 a_12925_46660# a_11735_46660# a_12816_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1251 VSS a_2957_45546# a_2905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1252 a_376_46348# a_n743_46660# a_518_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1253 a_11415_45002# a_4915_47217# a_14581_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1254 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X1255 a_n2104_42282# a_n1925_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1256 a_n2472_45002# a_n2293_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1257 a_21398_44850# a_20679_44626# a_20835_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1258 VDD a_22521_40599# a_22705_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1259 VDD a_16333_45814# a_16223_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1260 a_16241_44484# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1261 a_3905_42865# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1262 VSS a_8685_43396# a_15231_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1263 VSS a_10623_46897# a_10554_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1264 a_13485_45572# a_12549_44172# a_13385_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1265 C3_P_btm a_n4209_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1266 VSS a_22959_45572# a_20447_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 a_19120_35138# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1268 VDD a_19987_42826# a_n2017_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X1269 a_9028_43914# a_9482_43914# a_9420_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1270 VSS a_17973_43940# a_18079_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1271 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1272 a_n2860_39072# a_n2956_39304# a_n2946_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1273 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1274 a_3059_42968# a_742_44458# a_2987_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1275 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1276 a_n452_44636# a_n467_45028# a_n310_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1277 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1278 VDD a_768_44030# a_2711_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1279 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1280 VDD a_12281_43396# a_12563_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1281 VDD a_12741_44636# a_22959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1282 a_8333_44734# a_3537_45260# a_8238_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1283 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1284 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1285 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1286 a_17124_42282# a_17303_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1287 a_12156_46660# a_11813_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1288 VDD a_10809_44734# a_22959_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1289 VSS a_1115_44172# a_n2293_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1290 a_5013_44260# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1291 VDD a_n447_43370# a_n2129_43609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1292 a_3357_43084# a_5257_43370# a_5565_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1293 a_1568_43370# a_1847_42826# a_1793_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1294 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1295 a_11682_45822# a_10586_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1296 a_18315_45260# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1297 a_n2012_44484# a_n2129_44697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1298 a_14543_43071# a_5534_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1299 a_16147_45260# a_17478_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1300 a_19963_31679# a_22591_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1301 a_n967_45348# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1302 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1303 VDD a_11599_46634# a_20107_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1304 VSS a_7276_45260# a_7227_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1305 a_1241_44260# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1306 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1307 VSS a_n815_47178# a_n785_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1308 a_n4334_40480# a_n4318_40392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1309 a_3175_45822# a_3090_45724# a_2957_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1310 a_14621_43646# a_14579_43548# a_14537_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1311 VDD a_n1386_35608# a_n1838_35608# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1312 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1313 VREF a_20205_31679# C4_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1314 VSS a_15227_44166# a_18900_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1315 a_n310_44811# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1316 VDD a_16977_43638# a_16867_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1317 VDD a_15227_44166# a_17749_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1318 a_3147_46376# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1319 a_12638_46436# a_12594_46348# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1320 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1321 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1322 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1323 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1324 a_21071_46482# a_15227_44166# a_20708_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1325 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1326 VDD a_1343_38525# a_2684_37794# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1327 a_961_42354# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1328 a_9127_43156# a_8952_43230# a_9306_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1329 VSS a_12741_44636# a_22959_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1330 VSS a_8349_46414# a_8283_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1331 VSS a_11787_45002# a_11652_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1332 a_4223_44672# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1333 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1334 a_509_45822# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1335 a_16119_47582# a_15673_47210# a_16023_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1336 a_6452_43396# a_6293_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1337 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1338 a_6194_45824# a_6472_45840# a_6428_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1339 a_3754_38802# a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1340 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1341 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1342 VDD a_n881_46662# a_11031_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1343 VSS a_1209_47178# a_1239_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1344 a_15559_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1345 a_12429_44172# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1346 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1347 a_11229_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1348 a_16020_45572# a_15903_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1349 C3_P_btm a_5932_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1350 a_10149_42308# a_9290_44172# a_9803_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1351 VSS a_20708_46348# a_20411_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1352 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1353 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1354 a_10793_43218# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1355 a_n863_45724# a_1667_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1356 a_13635_43156# a_13460_43230# a_13814_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1357 a_12379_46436# a_12594_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1358 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1359 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1360 a_1209_43370# a_1049_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1361 a_2982_43646# a_3232_43370# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1362 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1363 a_21542_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1364 VSS a_19647_42308# a_13258_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1365 a_18985_46122# a_18819_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1366 a_12839_46116# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1367 VDD a_n2438_43548# a_2443_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1368 VDD a_9028_43914# a_8975_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1369 VDD a_17124_42282# a_4958_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1370 VSS a_10053_45546# a_9625_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X1371 a_17639_46660# a_17609_46634# a_765_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1372 VSS a_380_45546# a_n356_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1373 VSS a_20193_45348# a_21973_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1374 VSS a_196_42282# a_n3674_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1375 VDD a_5257_43370# a_5826_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X1376 a_9803_42558# a_n97_42460# a_9885_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1377 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1378 VSS a_10227_46804# a_10553_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1379 VSS a_18597_46090# a_16375_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1380 VSS a_n913_45002# a_12281_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1381 a_12816_46660# a_11901_46660# a_12469_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1382 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1383 a_20205_45028# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1384 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1385 VDD a_13259_45724# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1386 a_n1736_42282# a_n1557_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1387 a_13747_46662# a_19386_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1388 VSS a_4791_45118# a_6165_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X1389 a_261_44278# a_n863_45724# a_175_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1390 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1391 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1392 a_8325_42308# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1393 a_10623_46897# a_10467_46802# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1394 a_17957_46116# a_765_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1395 a_2675_43914# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1396 a_18695_43230# a_18249_42858# a_18599_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1397 a_17613_45144# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1398 a_n4318_39304# a_n2840_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1399 a_18799_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1400 VSS a_19862_44208# a_20922_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1401 a_6151_47436# a_14311_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1402 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1403 VSS a_5129_47502# a_5063_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1404 VSS a_167_45260# a_2521_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1405 a_3733_45822# a_n755_45592# a_3638_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1406 a_16333_45814# a_16115_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1407 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1408 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1409 a_1337_46116# a_1176_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1410 a_13163_45724# a_13527_45546# a_13485_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1411 a_8605_42826# a_8387_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1412 VDD a_4419_46090# a_n1925_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1413 a_n83_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1414 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1415 a_20712_42282# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1416 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1417 a_1241_43940# a_1467_44172# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1418 a_9145_43396# a_8791_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1419 VDD a_n961_42308# a_n784_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1420 a_7227_42852# a_n97_42460# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1421 a_14976_45348# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1422 a_9863_47436# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1423 a_743_42282# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1424 a_4915_47217# a_12991_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1425 VSS a_12891_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1426 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1427 a_n3674_38680# a_n2840_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1428 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1429 VSS a_3539_42460# a_3065_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1430 a_17801_45144# a_17613_45144# a_17719_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1431 VDD a_n4209_39590# a_n4334_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1432 a_18787_45572# a_18341_45572# a_18691_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1433 a_10922_42852# a_10796_42968# a_10518_42984# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1434 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1435 a_3754_39964# a_7754_40130# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1436 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1437 VDD a_526_44458# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1438 a_n1630_35242# a_564_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1439 a_167_45260# a_2202_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1440 VDD a_11967_42832# a_20512_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1441 VDD a_16019_45002# a_15903_45785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1442 a_2896_43646# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1443 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1444 a_n2312_38680# a_n2104_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1445 a_12005_46116# a_10903_43370# a_12005_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1446 a_n2288_47178# a_n2109_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1447 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1448 a_14097_32519# a_22959_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1449 a_6999_46987# a_3877_44458# a_6540_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1450 a_8199_44636# a_10355_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1451 a_3429_45260# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1452 C8_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1453 a_4338_37500# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X1454 a_9293_42558# a_9223_42460# a_8953_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1455 VDD a_n452_47436# a_n815_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1456 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1457 a_14309_45348# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1458 a_13807_45067# a_13556_45296# a_13348_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1459 a_2981_46116# a_2804_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1460 a_1176_45822# a_997_45618# a_1260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X1461 a_4185_45028# a_3877_44458# a_4185_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1462 VDD a_13159_45002# a_n2661_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1463 VSS a_20269_44172# a_19319_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1464 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1465 a_16104_42674# a_15890_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1466 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1467 a_22731_47423# SMPL_ON_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1468 a_n722_46482# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1469 VSS a_n443_42852# a_997_45618# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1470 a_6945_45348# a_5205_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1471 a_21513_45002# a_21363_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1472 a_4791_45118# a_4743_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1473 VSS a_1576_42282# a_1606_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1474 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1475 a_15227_44166# a_22000_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1476 VSS en_comp a_1177_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1477 a_n743_46660# a_n1021_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1478 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1479 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1480 VSS a_5205_44484# a_6756_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1481 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1482 VDD a_327_44734# a_375_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1483 VDD a_19321_45002# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1484 VSS a_3483_46348# a_13829_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1485 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1486 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1487 VDD a_5937_45572# a_6671_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1488 VDD a_n863_45724# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1489 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1490 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1491 VDD a_1756_43548# a_1467_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X1492 VDD a_4791_45118# a_5066_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1493 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1494 a_20269_44172# a_20365_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1495 VDD a_14976_45028# a_15227_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1496 VSS a_13904_45546# a_12594_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1497 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1498 VSS a_8953_45546# a_8568_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1499 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1500 a_16112_44458# a_15227_44166# a_16335_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1501 VSS a_16327_47482# a_17021_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1502 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 VSS a_20974_43370# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1504 a_16388_46812# a_17957_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1505 VSS a_20159_44458# a_19321_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1506 VDD a_9672_43914# a_2107_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1507 a_n4318_37592# a_n1736_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1508 VSS a_6151_47436# a_8189_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1509 VDD a_12549_44172# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1510 a_6229_45572# a_6194_45824# a_5907_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1511 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1512 VDD a_19700_43370# a_n97_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1513 a_6851_47204# a_6491_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1514 VDD a_19615_44636# a_18579_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1515 a_8423_43396# a_n443_42852# a_8317_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1516 VDD a_7499_43078# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1517 a_18799_45938# a_18175_45572# a_18691_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1518 a_1755_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1519 a_n1741_47186# a_12005_46116# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X1520 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1521 VDD a_6765_43638# a_6655_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1522 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1523 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1524 VDD a_22223_47212# a_21588_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1525 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1526 a_685_42968# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1527 a_10467_46802# a_11599_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1528 VDD a_n443_42852# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1529 a_17749_42852# a_17701_42308# a_17665_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1530 a_18599_43230# a_18249_42858# a_18504_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1531 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1532 VDD a_7920_46348# a_7715_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1533 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1534 a_2809_45028# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1535 a_7832_46660# a_7715_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1536 a_3873_46454# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1537 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1538 VSS a_4905_42826# a_4520_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1539 a_6709_45028# a_6431_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1540 VSS a_20202_43084# a_21421_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1541 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1542 a_20623_43914# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1543 a_20193_45348# a_18494_42460# a_20205_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1544 VSS a_9313_45822# a_11459_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1545 a_n4318_39768# a_n2840_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1546 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 VSS a_22469_40625# a_22717_36887# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1548 a_6428_45938# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1549 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1550 a_n2104_46634# a_n1925_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1551 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1552 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1553 EN_VIN_BSTR_N VDD a_19120_35138# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1554 a_2987_42968# a_1847_42826# a_2905_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1555 a_11031_47542# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1556 VSS a_12991_46634# a_12925_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1557 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1558 VDAC_Ni a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1559 VSS a_20894_47436# a_20843_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 a_13076_44458# a_9482_43914# a_13468_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1561 a_10752_42852# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1562 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1563 a_17970_44736# a_18248_44752# a_18204_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1564 a_5663_43940# a_5883_43914# a_5841_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1565 a_n2302_38778# a_n2312_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1566 a_16588_47582# a_15507_47210# a_16241_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1567 VSS a_4099_45572# a_3483_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1568 VSS a_14539_43914# a_16112_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1569 a_16867_43762# a_16243_43396# a_16759_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1570 a_n745_45366# a_n746_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1571 a_10518_42984# a_10835_43094# a_10793_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1572 C2_P_btm a_n3420_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1573 VIN_P EN_VIN_BSTR_P C5_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1574 a_n37_45144# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 a_18287_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1576 a_20159_44458# a_20362_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1577 VSS a_11341_43940# a_22223_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1578 VSS a_8530_39574# a_3754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1579 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1580 a_6969_46634# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1581 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1582 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1583 a_18861_43218# a_18817_42826# a_18695_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1584 a_11322_45546# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1585 a_n3674_37592# a_196_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1586 a_n1809_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1587 a_4419_46090# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1588 VDD a_11189_46129# a_11133_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1589 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1590 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1591 VSS a_7640_43914# a_7584_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1592 VIN_P EN_VIN_BSTR_P a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1593 a_15959_42545# a_15764_42576# a_16269_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1594 a_16375_45002# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1595 VDD a_n1699_44726# a_n1809_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1596 a_4235_43370# a_3935_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1597 a_21177_47436# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1598 a_7418_45394# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1599 a_22000_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1600 VDD a_7542_44172# a_7499_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1601 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1602 a_11309_47204# a_11031_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1603 VDD a_1307_43914# a_3353_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1604 a_3905_42308# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1605 a_8483_43230# a_8037_42858# a_8387_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1606 a_n2104_46634# a_n1925_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1607 a_453_43940# a_175_44278# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1608 a_7281_43914# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1609 a_9028_43914# a_9290_44172# a_9248_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1610 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1611 VDD a_4700_47436# a_3785_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1612 a_18909_45814# a_18691_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1613 a_15521_42308# a_15486_42560# a_15051_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1614 a_11551_42558# a_n97_42460# a_11633_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1615 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1616 VDD a_15227_44166# a_15415_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1617 VSS a_16327_47482# a_20397_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1618 a_n809_44244# a_n984_44318# a_n630_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1619 VDD a_8270_45546# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1620 VDD a_948_46660# a_1123_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1621 VDD a_15009_46634# a_14180_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1622 a_20766_44850# a_20679_44626# a_20362_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1623 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1624 a_13385_45572# a_10903_43370# a_13297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1625 VDD a_13777_45326# a_13807_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1626 VSS a_n755_45592# a_n39_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1627 a_14976_45028# a_14797_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1628 a_6886_37412# VDAC_Pi VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1629 a_6419_46482# a_6165_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X1630 VSS a_768_44030# a_5244_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1631 a_n2302_37690# a_n2810_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1632 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1633 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1634 VDD a_8199_44636# a_8336_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1635 a_20623_45572# a_20273_45572# a_20528_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1636 VSS a_9396_43370# a_5111_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1637 a_n2312_39304# a_n1920_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1638 a_20009_46494# a_18819_46122# a_19900_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1639 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1640 a_7309_42852# a_5891_43370# a_7227_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1641 a_743_42282# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1642 VSS a_n4064_40160# a_n2302_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1643 a_22397_42558# a_n913_45002# a_17303_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1644 a_12991_43230# a_12545_42858# a_12895_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1645 VSS a_3905_42865# a_5013_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1646 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 a_22765_42852# a_15743_43084# a_18184_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1648 a_7705_45326# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1649 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1650 VSS a_10405_44172# a_8016_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1651 a_3065_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1652 a_742_44458# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1653 a_310_45028# a_n37_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1654 VDD a_3232_43370# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1655 VDD a_526_44458# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1656 VSS a_18184_42460# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X1657 VDD a_16241_47178# a_16131_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1658 a_19466_46812# a_13747_46662# a_19929_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1659 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1660 a_20850_46482# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1661 VSS a_768_44030# a_9028_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1662 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1663 a_12089_42308# a_11551_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1664 a_11173_43940# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1665 a_3457_43396# a_1414_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1666 VDD a_5907_46634# a_5894_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1667 a_8034_45724# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1668 a_5841_46660# a_4651_46660# a_5732_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1669 a_22000_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1670 VSS a_3699_46348# a_3160_47472# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1671 VSS a_22223_45036# a_18114_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1672 a_2437_43396# a_1568_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1673 VDD a_n2104_46634# a_n2312_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1674 a_2448_45028# a_2382_45260# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X1675 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1676 a_21167_46155# a_20916_46384# a_20708_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1677 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1678 a_5205_44484# a_5343_44458# a_5289_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1679 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1680 a_948_46660# a_33_46660# a_601_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1681 VSS a_21005_45260# a_19778_44110# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1682 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1683 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X1684 a_9241_46436# a_n237_47217# a_8049_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1685 a_15015_46420# a_14840_46494# a_15194_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1686 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1687 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1688 VDD a_20567_45036# a_12549_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1689 a_21398_44850# a_20640_44752# a_20835_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1690 a_22717_37285# a_22459_39145# a_22609_38406# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1691 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1692 a_1823_45246# a_4704_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1693 a_5527_46155# a_5204_45822# a_5068_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1694 a_1606_42308# a_1576_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1695 VSS a_4235_43370# a_4181_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VDD a_18783_43370# a_18525_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1697 VSS a_18194_35068# a_19120_35138# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1698 a_n881_46662# a_14495_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1699 a_21188_45572# a_20107_45572# a_20841_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1700 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1701 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1702 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1703 VCM a_5534_30871# C7_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1704 VSS a_8270_45546# a_8192_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1705 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1706 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1707 VDD a_n863_45724# a_3059_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1708 VDD a_17609_46634# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1709 VSS a_n755_45592# a_3503_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1710 a_19237_31679# a_22959_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1711 a_12156_46660# a_11813_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1712 a_n4334_38528# a_n4318_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1713 a_n901_43156# a_n1076_43230# a_n722_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1714 a_n2810_45028# a_n2840_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1715 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1716 a_16333_45814# a_16115_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1717 a_16795_42852# a_n97_42460# a_16877_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1718 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1719 VDD a_21188_46660# a_21363_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1720 a_6905_45572# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1721 a_14180_45002# a_13059_46348# a_14403_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1722 a_16405_45348# a_16375_45002# a_16321_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1723 VDD a_5934_30871# a_8515_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1724 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=10.615 ps=76.96 w=3.75 l=15
X1725 VREF a_19963_31679# C3_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1726 VDD a_3422_30871# a_22315_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1727 a_2123_42473# a_n784_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1728 VSS a_n1613_43370# a_n1287_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1729 VSS a_22223_43948# a_14401_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1730 a_19518_43218# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1731 VSS a_20075_46420# a_20009_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1732 VSS a_16922_45042# a_16751_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1733 VDD a_3232_43370# a_11341_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X1734 a_1049_43396# a_458_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1735 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1736 VDD a_n237_47217# a_8270_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1737 a_1848_45724# a_n237_47217# a_1990_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1738 VDD a_14539_43914# a_12465_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1739 VDD a_n881_46662# a_7903_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1740 VDD a_n1423_46090# a_n1533_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1741 VDD a_5111_44636# a_5421_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1742 a_20623_46660# a_20107_46660# a_20528_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1743 a_11778_45572# a_10193_42453# a_11688_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1744 a_6347_46155# a_6165_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1745 a_4700_47436# a_n443_46116# a_4842_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1746 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1747 VDD a_21359_45002# a_21101_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1748 C4_P_btm a_n3565_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1749 a_14113_42308# a_13575_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1750 VDD a_5755_42308# a_5932_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1751 a_10695_43548# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1752 a_4958_30871# a_17124_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1753 a_17333_42852# a_16795_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1754 VSS a_19339_43156# a_19273_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1755 a_8387_43230# a_8037_42858# a_8292_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1756 VDD a_n2840_44458# a_n4318_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1757 VDD a_15004_44636# a_14815_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1758 VSS a_16327_47482# a_18861_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1759 VSS a_1823_45246# a_3602_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1760 VDD a_18780_47178# a_13661_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1761 a_n4334_37440# a_n4318_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1762 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1763 a_2455_43940# a_895_43940# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1764 a_2680_45002# a_3065_45002# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1765 a_13667_43396# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1766 CAL_P a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1767 a_21381_43940# a_21115_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1768 a_380_45546# a_765_45546# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1769 a_15781_43660# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1770 VSS a_22521_39511# a_22469_39537# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1771 a_16019_45002# a_16147_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X1772 VDD a_3537_45260# a_4558_45348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1773 a_12741_44636# a_6755_46942# a_16789_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1774 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1775 a_5534_30871# a_12563_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1776 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1777 VDD a_n473_42460# a_n1761_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1778 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X1779 a_20836_43172# a_20193_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1780 a_12895_43230# a_12545_42858# a_12800_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1781 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1782 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X1783 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1784 a_726_44056# a_626_44172# a_644_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1785 a_6655_43762# a_6031_43396# a_6547_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1786 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1787 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1788 a_2889_44172# a_1414_42308# a_3052_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1789 VDD a_3232_43370# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1790 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1791 a_5343_44458# a_7963_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1792 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1793 a_3483_46348# a_4099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1794 a_9313_44734# a_5883_43914# a_9241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1795 a_2809_45028# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1796 VDD a_6171_45002# a_11827_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1797 VDD a_9625_46129# a_9569_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1798 a_15567_42826# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1799 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1800 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1801 a_7_45899# a_n443_46116# a_n452_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1802 a_n2810_45572# a_n2840_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1803 a_5732_46660# a_4817_46660# a_5385_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1804 a_5708_44484# a_3483_46348# a_5608_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X1805 VDD a_13259_45724# a_22397_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1806 VSS a_22521_40055# a_22459_39145# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1807 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1808 VDD a_13507_46334# a_22765_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1809 a_13678_32519# a_21855_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1810 a_5365_45348# a_5111_44636# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1811 a_17021_43396# a_16977_43638# a_16855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1812 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1813 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1814 a_7989_47542# a_n237_47217# a_7903_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1815 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1816 a_19332_42282# a_19511_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1817 VSS a_6851_47204# a_7227_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1818 a_13607_46688# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1819 a_4880_45572# a_526_44458# a_4808_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1820 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1821 a_20922_43172# a_10193_42453# a_20836_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1822 a_12978_47026# a_11901_46660# a_12816_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1823 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1824 VDD a_13720_44458# a_12607_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1825 VDD a_2952_47436# a_2747_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1826 a_5147_45002# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1827 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1828 VDD a_14513_46634# a_14543_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1829 VDD a_21259_43561# a_16922_45042# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1830 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1831 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1832 VDD a_21137_46414# a_21167_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1833 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1834 a_3905_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1835 VSS a_22959_47212# a_22612_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 a_383_46660# a_33_46660# a_288_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1837 VSS a_6755_46942# a_13556_45296# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1838 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1839 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1840 a_17061_44734# a_11691_44458# a_16979_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1841 a_4149_42891# a_2382_45260# a_3935_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X1842 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1843 VDD a_n755_45592# a_3318_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1844 VDD a_n443_46116# a_1427_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1845 VDD a_5497_46414# a_5527_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1846 a_5937_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1847 a_11323_42473# a_5742_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1848 VSS a_4921_42308# a_5755_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1849 a_21076_30879# a_22959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1850 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1851 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1852 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1853 a_3699_46634# a_3524_46660# a_3878_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1854 VDD a_17583_46090# a_13259_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1855 VSS a_3600_43914# a_3499_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1856 VSS a_n755_45592# a_3318_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1857 a_5111_44636# a_9396_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1858 a_17595_43084# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1859 a_13829_44260# a_13059_46348# a_13483_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1860 a_18341_45572# a_18175_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1861 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 a_12991_46634# a_12816_46660# a_13170_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1863 VSS a_2277_45546# a_2211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1864 a_18429_43548# a_18525_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1865 VSS a_6453_43914# a_n2661_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1866 a_6773_42558# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1867 a_2253_44260# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1868 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1869 a_9885_42558# a_7499_43078# a_9803_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1870 a_16414_43172# a_16137_43396# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1871 a_21811_47423# SINGLE_ENDED VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1872 a_2304_45348# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1873 a_3726_37500# a_6886_37412# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1874 a_13351_46090# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1875 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1876 a_n1435_47204# a_n1605_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1877 a_n935_46688# a_n1151_42308# a_n1021_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1878 VSS a_12549_44172# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X1879 a_6977_45572# a_6598_45938# a_6905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1880 a_11530_34132# EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1881 VSS a_n23_44458# a_n89_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1882 VSS a_n1177_43370# a_n1243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1883 VDD a_13460_43230# a_13635_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1884 VSS a_n913_45002# a_n967_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1885 VDD a_11525_45546# a_11189_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1886 VDD a_n755_45592# a_626_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1887 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1888 VDD a_10227_46804# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1889 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1890 a_895_43940# a_644_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1891 a_n699_43396# a_n1177_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1892 a_11136_42852# a_10922_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1893 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1894 VDD a_8568_45546# a_8162_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1895 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1896 a_11551_42558# a_n97_42460# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1897 a_6293_42852# a_5755_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1898 a_n2840_42826# a_n2661_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1899 a_16131_47204# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1900 a_14033_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1901 a_5289_44734# a_4223_44672# a_5205_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1902 VSS a_n1736_42282# a_n4318_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1903 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1904 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1905 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1906 VDD a_11415_45002# a_22591_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1907 VSS a_5147_45002# a_5708_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X1908 VIN_N EN_VIN_BSTR_N C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1909 VDD a_13259_45724# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1910 VSS a_6886_37412# a_4338_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1911 a_10053_45546# a_10490_45724# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1912 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1913 VDD a_19332_42282# a_4190_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1914 a_n998_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1915 a_3090_45724# a_18911_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X1916 VSS a_18287_44626# a_18248_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1917 a_6671_43940# a_6109_44484# a_6453_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1918 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1919 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1920 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1921 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1922 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1923 a_16131_47204# a_15507_47210# a_16023_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1924 a_n23_44458# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1925 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1926 a_11750_44172# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1927 a_7845_44172# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1928 VIN_N EN_VIN_BSTR_N C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1929 VSS a_6123_31319# a_7963_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1930 a_5907_46634# a_5732_46660# a_6086_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1931 a_8560_45348# a_8746_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1932 a_19095_43396# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1933 a_21363_46634# a_21188_46660# a_21542_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1934 VSS a_n4315_30879# a_n4251_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1935 VSS a_n4064_39616# a_n2302_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1936 a_14180_46482# a_14035_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1937 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1938 a_18315_45260# a_18587_45118# a_18545_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1939 a_8349_46414# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1940 a_2537_44260# a_2479_44172# a_2127_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1941 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1942 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1943 VSS a_3499_42826# a_3445_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1944 VDD a_3815_47204# a_4007_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1945 a_9306_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1946 VDD a_6667_45809# a_6598_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1947 a_7230_45938# a_6511_45714# a_6667_45809# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1948 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1949 a_8685_43396# a_8147_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1950 VDD a_1343_38525# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1951 VSS VSS a_3726_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X1952 a_8270_45546# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1953 a_15765_45572# a_15599_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1954 a_3992_43940# a_768_44030# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1955 a_3815_47204# a_3785_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1956 a_2063_45854# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1957 VSS a_11415_45002# a_22591_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1958 a_6755_46942# a_15015_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1959 VDD a_19431_45546# a_19418_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1960 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1961 VSS a_14021_43940# a_22959_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1962 a_19328_44172# a_19478_44306# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X1963 VSS a_10227_46804# a_14537_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1964 a_21073_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1965 VDD a_768_44030# a_726_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1966 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1967 VDD a_13059_46348# a_15297_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1968 VSS a_12465_44636# a_22223_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1969 VDD a_n1352_43396# a_n1177_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1970 VSS a_n863_45724# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1971 a_19164_43230# a_18083_42858# a_18817_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1972 a_383_46660# a_n133_46660# a_288_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1973 a_3524_46660# a_2443_46660# a_3177_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1974 a_13814_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1975 VSS a_9127_43156# a_9061_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1976 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1977 VDD a_9482_43914# a_10157_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1978 VSS a_12607_44458# a_12553_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1979 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1980 VSS a_10903_43370# a_11963_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1981 VSS a_17499_43370# a_17433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1982 C1_P_btm a_1606_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1983 VDD a_12427_45724# a_10490_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1984 a_13213_44734# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1985 VSS a_14815_43914# a_14761_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1986 a_12513_46660# a_12469_46902# a_12347_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1987 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1988 VSS a_11323_42473# a_10807_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1989 a_18989_43940# a_18451_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1990 VDD a_1209_43370# a_n1557_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1991 VSS a_8667_46634# a_8601_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1992 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1993 a_2889_44172# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1994 VSS a_7281_43914# a_7229_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1995 VSS a_21195_42852# a_21671_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1996 a_n2956_38680# a_n2472_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1997 VSS a_n699_43396# a_4743_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1998 VDD a_n443_46116# a_2437_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1999 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2000 a_10553_43218# a_10518_42984# a_10083_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2001 a_16789_44484# a_14537_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2002 VSS a_13635_43156# a_13569_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2003 a_18834_46812# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2004 a_10405_44172# a_7499_43078# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X2005 a_n1151_42308# a_n1329_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2006 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2007 VSS a_18315_45260# a_18189_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2008 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2009 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2010 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2011 VDD a_17499_43370# a_17486_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2012 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2013 VDD a_22223_42860# a_22400_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2014 VDD a_3524_46660# a_3699_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2015 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2017 VSS a_12861_44030# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2018 a_10765_43646# a_10695_43548# a_10057_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2019 VDD a_12549_44172# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2020 a_15890_42674# a_15803_42450# a_15486_42560# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2021 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2022 a_17433_43396# a_16243_43396# a_17324_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2023 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2024 a_11827_44484# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2025 a_1847_42826# a_2351_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2026 VSS a_6151_47436# a_14955_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2027 a_20205_31679# a_22223_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2028 VSS a_15227_44166# a_15785_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2029 VDD a_1239_47204# a_1431_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2030 VDD a_8667_46634# a_8654_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2031 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2032 a_n452_45724# a_n443_46116# a_n310_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2033 a_700_44734# a_n746_45260# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2034 a_19862_44208# a_13747_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2035 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2036 a_10775_45002# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2037 a_3232_43370# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2038 VDD a_22959_44484# a_19237_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2039 a_1115_44172# a_453_43940# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2040 a_484_44484# a_n863_45724# a_327_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2041 a_n3690_38528# a_n3674_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2042 VDD a_14543_43071# a_13291_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2043 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2044 a_20512_43084# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2045 VSS a_12549_44172# a_21205_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2046 a_20256_43172# a_20202_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X2047 a_6761_42308# a_n913_45002# a_6773_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2048 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2049 VDD a_19864_35138# a_21589_35634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2050 a_n2840_42282# a_n2661_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2051 a_n2661_46098# a_1983_46706# a_2162_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2052 a_5429_46660# a_5385_46902# a_5263_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2053 VSS a_15368_46634# a_15312_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2054 VDD a_8685_43396# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2055 VDD a_16855_45546# a_16842_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2056 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2057 a_11315_46155# a_11133_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2058 a_16522_42674# a_15803_42450# a_15959_42545# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2059 a_1221_42558# a_1184_42692# a_1149_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2060 a_20885_46660# a_20841_46902# a_20719_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2061 a_20719_45572# a_20273_45572# a_20623_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2062 a_1756_43548# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2063 a_n923_35174# EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2064 a_14456_42282# a_14635_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2065 a_n2472_42826# a_n2293_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2066 a_7276_45260# a_6709_45028# a_7418_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2067 VDD a_1823_45246# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2068 VDD a_22400_42852# a_22521_40055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2069 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2070 a_3260_45572# a_3218_45724# a_2957_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2071 a_n2497_47436# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2072 VSS a_3422_30871# a_22315_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2073 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2074 VDD a_10341_42308# a_11554_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2075 a_11280_45822# a_2063_45854# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2076 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2077 a_603_45572# a_310_45028# a_509_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2078 a_15002_46116# a_13925_46122# a_14840_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2079 a_8746_45002# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2080 a_n906_45572# a_n971_45724# a_n1013_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2081 a_11064_45572# a_10903_43370# a_10907_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2082 a_21205_44306# a_20935_43940# a_21115_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2083 a_2479_44172# a_2905_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2084 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2085 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2086 VDD a_n2840_46090# a_n2956_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2087 VDD a_6945_45028# a_22223_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2088 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2089 a_13556_45296# a_6755_46942# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2090 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2091 VCM a_7174_31319# C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2092 VDD a_8199_44636# a_9377_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2093 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2094 a_n4334_39392# a_n4318_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2095 a_12710_44260# a_10903_43370# a_12603_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2096 a_13777_45326# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2097 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2098 a_16522_42674# a_15764_42576# a_15959_42545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2099 a_14205_43396# a_13667_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X2100 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2101 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2102 VDD a_5732_46660# a_5907_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2103 a_6419_46155# a_5807_45002# a_6419_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2104 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2105 a_n2860_39866# a_n2956_39768# a_n2946_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2106 VDD a_13556_45296# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2107 a_18533_44260# a_18326_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2108 a_n901_46420# a_n1076_46494# a_n722_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2109 a_5066_45546# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2110 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X2111 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2112 VSS a_11599_46634# a_18175_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2113 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2114 VSS a_11599_46634# a_18819_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2115 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2116 a_n3690_37440# a_n3674_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2117 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2118 a_n2442_46660# a_n2472_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2119 VSS a_n1435_47204# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2120 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2121 a_8317_43396# a_n755_45592# a_8229_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2122 a_n3674_38216# a_n2104_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2123 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2124 a_n2312_40392# a_n2288_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2125 VDD a_n1079_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2126 VSS a_22591_44484# a_17730_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2127 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2128 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2129 a_n97_42460# a_19700_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2130 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2131 a_3877_44458# a_3699_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2132 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2133 a_15368_46634# a_15143_45578# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2134 a_11206_38545# CAL_N a_4338_37500# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2135 a_4905_42826# a_5379_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2136 VSS a_10467_46802# a_10428_46928# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2137 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2138 a_9313_45822# a_9049_44484# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2139 a_21145_44484# a_20766_44850# a_21073_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2140 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2141 VSS a_22521_40599# a_22717_37285# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2142 VSS a_2680_45002# a_2274_45254# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2143 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2144 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2145 a_10768_47026# a_10554_47026# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2146 VSS a_21671_42860# a_3422_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2147 a_n785_47204# a_n815_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2148 a_5837_45028# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2149 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2150 C0_dummy_P_btm a_7174_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2151 a_14537_43396# a_14358_43442# a_14621_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2152 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2153 a_n1736_43218# a_n1853_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2154 a_6640_46482# a_5257_43370# a_6419_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2155 VDD a_3090_45724# a_17786_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2156 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2157 a_15493_43396# a_14955_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2158 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2159 a_16877_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2160 a_9823_46482# a_9569_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X2161 VDD a_14021_43940# a_22959_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2162 VDD a_n3420_38528# a_n2860_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2163 VSS a_10227_46804# a_12513_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2164 VDD a_3483_46348# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2165 VSS a_17339_46660# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2166 VSS a_n1532_35090# a_n83_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2167 a_3699_46348# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2168 VSS a_10533_42308# a_10723_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2169 VSS a_3537_45260# a_4223_44672# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2170 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2171 a_18214_42558# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2172 VSS a_14537_43396# a_14180_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2173 a_16501_45348# a_10193_42453# a_16405_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2174 VSS a_15743_43084# a_15567_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2175 VSS a_21259_43561# a_16922_45042# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2176 VSS a_n2840_46634# a_n2956_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2177 a_9049_44484# a_8701_44490# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2178 VDD a_22821_38993# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2179 VDD a_2382_45260# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2180 VDD a_n967_45348# a_n961_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2181 a_19615_44636# a_12861_44030# a_19789_44512# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2182 a_9863_46634# a_10150_46912# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2183 VDD a_n881_46662# a_n745_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2184 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2185 VDD a_21496_47436# a_13507_46334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2186 a_n2109_45247# a_n2017_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2187 VSS a_n143_45144# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2188 a_19418_45938# a_18341_45572# a_19256_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2189 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2190 VDD a_n2438_43548# a_n2433_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2191 VDD a_5907_45546# a_5937_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X2192 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2193 C5_P_btm a_n4209_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2194 VSS a_n452_44636# a_n2129_44697# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2195 a_n2472_42282# a_n2293_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2196 a_n4318_38680# a_n2472_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2197 a_5608_44484# a_5111_44636# a_5518_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X2198 VDD a_742_44458# a_700_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2199 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2200 VSS a_768_44030# a_13720_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2201 VSS a_7287_43370# a_7221_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2202 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2203 a_2609_46660# a_2443_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2204 a_n89_44484# a_n467_45028# a_n452_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2205 VDD a_9290_44172# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2206 VSS a_n1613_43370# a_6809_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2207 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2208 a_556_44484# a_526_44458# a_484_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2209 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2210 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2211 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2212 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2213 a_2112_39137# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2214 VSS a_19328_44172# a_19279_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2215 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2216 VDD a_n3420_37440# a_n2860_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2217 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2218 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2219 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2220 a_10554_47026# a_10467_46802# a_10150_46912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2221 a_11387_46155# a_n1151_42308# a_11315_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2222 a_10341_43396# a_9803_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2223 a_13887_32519# a_22223_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2224 VSS a_10227_46804# a_20885_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2225 C0_P_btm a_n3420_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2226 VIN_P EN_VIN_BSTR_P C2_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2227 VSS a_16137_43396# a_18548_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2228 a_n452_45724# a_n743_46660# a_n310_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2229 a_11682_45822# a_11652_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2230 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2231 VDD a_n2472_46090# a_n2956_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2232 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2233 VDD a_11322_45546# a_11280_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2234 VSS a_13747_46662# a_14495_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2235 VDD a_10809_44734# a_n2661_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2236 C0_dummy_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2237 VSS a_n4209_39590# a_n4251_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2238 VSS a_n1329_42308# a_n1151_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2239 a_3381_47502# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2240 VDD a_18479_47436# a_13747_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2241 VSS a_n746_45260# a_261_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2242 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2243 a_5649_42852# a_5111_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2244 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2245 a_11136_45572# a_3483_46348# a_11064_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2246 VSS a_13249_42308# a_13904_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2247 a_17486_43762# a_16409_43396# a_17324_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2248 VSS a_n913_45002# a_8325_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2249 VSS a_1307_43914# a_2675_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2250 VSS a_n1532_35090# a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2251 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2252 a_3699_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2253 VSS a_13259_45724# a_14797_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2254 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2255 a_20841_45814# a_20623_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2256 VIN_N EN_VIN_BSTR_N C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2257 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2258 a_17639_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2259 a_10341_42308# a_9803_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2260 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2261 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2262 a_1260_45572# a_n755_45592# a_1176_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X2263 a_20397_44484# a_20362_44736# a_20159_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2264 a_12991_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2265 a_518_46155# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2266 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2267 VDD a_20841_45814# a_20731_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2268 a_9751_46155# a_9569_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2269 a_1443_43940# a_1414_42308# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2270 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X2271 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2272 VDD a_11823_42460# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2273 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2274 VSS a_n2840_42826# a_n3674_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2275 VSS a_3537_45260# a_5365_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2276 a_21589_35634# a_19864_35138# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2277 a_3065_45002# a_3318_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2278 a_n310_45899# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2279 C8_P_btm a_n3420_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2280 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2281 VDD a_22591_46660# a_20820_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2282 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2283 a_8337_42558# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2284 VDD a_4646_46812# a_7411_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2285 a_11186_47026# a_10428_46928# a_10623_46897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2286 a_20273_46660# a_20107_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2287 VSS a_3877_44458# a_2382_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2288 VDD a_n1331_43914# a_n1441_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2289 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2290 VDD a_10835_43094# a_10796_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2291 VSS a_5066_45546# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2292 VSS a_12883_44458# a_12829_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2293 a_11341_43940# a_10729_43914# a_11257_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2294 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2295 VSS a_564_42282# a_n1630_35242# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2296 a_12549_44172# a_20567_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2297 VDD a_14456_42282# a_5342_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2298 a_645_46660# a_601_46902# a_479_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2299 VDD a_2063_45854# a_10809_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2300 VDD a_2127_44172# a_n2661_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2301 VDD a_10227_46804# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2302 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2303 a_14513_46634# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2304 a_n2840_46090# a_n2661_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2305 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2306 a_21137_46414# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2307 a_1609_45822# a_167_45260# a_1609_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2308 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2309 a_14635_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2310 a_10544_45572# a_10490_45724# a_10053_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X2311 a_10555_44260# a_10949_43914# a_10405_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X2312 C2_P_btm a_n3565_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2313 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2314 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2315 VDD a_1736_39587# a_1239_39587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2316 a_8952_43230# a_7871_42858# a_8605_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2317 a_3067_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2318 a_9377_42558# a_8685_42308# a_9293_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2319 a_4190_30871# a_19332_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2320 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2321 a_15861_45028# a_15595_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2322 a_15194_46482# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2323 a_6469_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2324 a_13720_44458# a_9482_43914# a_14112_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2325 a_15493_43940# a_14955_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2326 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2327 a_16245_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2328 VSS a_n357_42282# a_6101_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2329 a_20692_30879# a_22959_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2330 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2331 a_3177_46902# a_2959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2332 a_5907_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2333 a_5497_46414# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2334 VSS a_104_43370# a_n971_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2335 VREF_GND a_13258_32519# C0_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2336 VDD a_4743_44484# a_4791_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2337 a_19700_43370# a_18579_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2338 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2339 a_21363_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2340 VSS a_n443_42852# a_15940_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X2341 a_12427_45724# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X2342 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2343 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2344 a_n1920_47178# a_n1741_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2345 a_10903_43370# a_13351_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2346 a_n955_45028# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2347 VDD a_n357_42282# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2348 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2349 a_18596_45572# a_18479_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2350 a_4185_45028# a_3065_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2351 a_6575_47204# a_6545_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2352 a_16137_43396# a_15781_43660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2353 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2354 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2355 VSS a_n2472_46634# a_n2442_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2356 a_4649_42852# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2357 VSS a_2711_45572# a_20107_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2358 VSS a_n2104_42282# a_n3674_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2359 VSS a_15015_46420# a_14949_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2360 VIN_N EN_VIN_BSTR_N a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2361 VSS a_5691_45260# a_n2109_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2362 a_17583_46090# a_17715_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2363 a_17730_32519# a_22591_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2364 a_3600_43914# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X2365 a_13925_46122# a_13759_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2366 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2367 VDD a_n901_43156# a_n914_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2368 a_8191_45002# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2369 VDD a_22959_46124# a_20692_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2370 a_n310_44484# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2371 a_21125_42558# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2372 a_5932_42308# a_5755_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2373 VSS a_14543_43071# a_13291_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2374 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2375 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2376 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2377 VDD a_16112_44458# a_14673_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2378 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2379 a_3175_45822# a_3316_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2380 VSS a_16763_47508# a_5807_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2381 VREF a_20447_31679# C5_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2382 a_14226_46660# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2383 VDD a_13348_45260# a_13159_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2384 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2385 VDD a_6491_46660# a_6851_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2386 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2387 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2388 a_6511_45714# a_4646_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2389 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2390 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2391 a_3422_30871# a_21671_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2392 VSS a_16763_47508# a_16697_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2393 VDD a_2889_44172# a_413_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X2394 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2395 VSS a_n443_42852# a_1755_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2396 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2397 a_10405_44172# a_10729_43914# a_10651_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2398 a_n2840_45546# a_n2661_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2399 a_14401_32519# a_22223_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2400 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2401 a_4558_45348# a_4574_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2402 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2403 a_5193_42852# a_3905_42865# a_5111_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2404 a_18143_47464# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2405 a_10533_42308# a_n913_45002# a_10545_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2406 VDD a_16721_46634# a_16751_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2407 a_18909_45814# a_18691_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2408 a_n2840_45002# a_n2661_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2409 a_948_46660# a_n133_46660# a_601_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2410 a_3699_46348# a_3877_44458# a_3873_46454# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2411 a_117_45144# a_n443_42852# a_45_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2412 a_11415_45002# a_13249_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2413 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2414 a_15681_43442# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2415 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2416 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2417 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2418 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X2419 VDD a_n1059_45260# a_18727_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2420 VSS a_5013_44260# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2421 a_9801_43940# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2422 VSS a_10193_42453# a_18797_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2423 a_22521_39511# a_22545_38993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X2424 a_n4251_38304# a_n4318_38216# a_n4334_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2425 a_2779_44458# a_1423_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2426 a_19789_44512# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X2427 VDD a_18057_42282# a_n356_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X2428 a_13113_42826# a_12895_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2429 a_16197_42308# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2430 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2431 VDD a_8034_45724# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2432 VDD a_11691_44458# a_11649_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2433 a_n3690_39392# a_n3674_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2434 a_15761_42308# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2435 a_16680_45572# a_15765_45572# a_16333_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2436 VSS a_1568_43370# a_1512_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2437 VDD a_5066_45546# a_5024_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2438 VSS a_n809_44244# a_n875_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2439 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2440 a_n2267_43396# a_n2433_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2441 a_10518_42984# a_10796_42968# a_10752_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2442 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2443 a_8189_46660# a_8145_46902# a_8023_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2444 VDD a_13661_43548# a_14976_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X2445 a_11691_44458# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2446 VSS a_n4064_39072# a_n2302_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2447 a_20062_46116# a_18985_46122# a_19900_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2448 a_20269_44172# a_20365_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2449 VSS a_5891_43370# a_5837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2450 VSS a_n2472_42826# a_n4318_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2451 VSS a_7754_38470# a_7754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2452 a_18707_42852# a_18083_42858# a_18599_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2453 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2454 a_12638_46436# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2455 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2456 a_n784_42308# a_n961_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2457 a_13157_43218# a_13113_42826# a_12991_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2458 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2459 VDD a_15015_46420# a_15002_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2460 VDD a_16327_47482# a_20159_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2461 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2462 VSS a_n785_47204# a_327_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2463 a_18834_46812# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2464 a_n2840_45546# a_n2661_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2465 VSS a_21177_47436# a_20990_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2466 VSS a_7499_43078# a_11816_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2467 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2468 a_6761_42308# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2469 a_10623_46897# a_10428_46928# a_10933_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2470 a_5263_45724# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2471 VDD a_11823_42460# a_11322_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2472 VSS a_5111_44636# a_8018_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2473 a_7903_47542# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2474 VSS a_8667_46634# a_n237_47217# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2475 a_3357_43084# a_4905_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2476 a_n2472_46090# a_n2293_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2477 VREF a_19237_31679# C0_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2478 VCM a_5742_30871# C6_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2479 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2480 VSS a_22959_46660# a_21076_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2481 a_10249_46116# a_9823_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X2482 VDD a_10775_45002# a_10180_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X2483 a_2684_37794# VDAC_Pi a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2484 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2485 a_8696_44636# a_16855_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2486 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2487 a_13467_32519# a_21487_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2488 a_6633_46155# a_5807_45002# a_6419_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2489 a_n2661_42834# a_8975_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2490 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2491 a_7274_43762# a_6197_43396# a_7112_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2492 a_10922_42852# a_10835_43094# a_10518_42984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2493 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2494 VDD a_5807_45002# a_11691_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2495 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2496 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2497 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2498 VSS RST_Z a_14311_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2499 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2500 a_18285_46348# a_18834_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2501 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2502 a_18597_46090# a_19431_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2503 VSS a_18443_44721# a_18374_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2504 VSS a_8199_44636# a_10951_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2505 a_1176_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2506 a_7735_45067# a_6709_45028# a_7276_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2507 C8_P_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2508 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2509 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2510 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X2511 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2512 VSS a_n2109_45247# en_comp VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2513 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2514 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2515 a_13348_45260# a_13556_45296# a_13490_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2516 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2517 a_n2302_40160# a_n2312_40392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2518 VSS a_21356_42826# a_n357_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2519 VDD a_11453_44696# a_22959_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2520 VSS a_15037_45618# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2521 VSS a_8696_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2522 a_3878_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2523 a_2277_45546# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2524 a_626_44172# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2525 a_18479_45785# a_19268_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2526 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2527 a_20273_45572# a_20107_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2528 a_10555_44260# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2529 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2530 VSS a_n443_42852# a_742_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2531 VSS a_n901_43156# a_n967_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2532 a_20820_30879# a_22591_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2533 VSS a_13076_44458# a_12883_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X2534 a_685_42968# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2535 a_17364_32525# a_22959_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2536 a_13170_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2537 a_11633_42558# a_9290_44172# a_11551_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2538 VDD a_4791_45118# a_6633_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2539 a_20731_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2540 a_19700_43370# a_18579_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2541 VDD a_11599_46634# a_20107_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2542 a_16751_45260# a_17023_45118# a_16981_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2543 a_2382_45260# a_3877_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2544 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2545 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2546 a_12829_44484# a_12741_44636# a_n2293_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2547 a_11257_43940# a_10807_43548# a_11173_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2548 VCM a_6123_31319# C4_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2549 VSS a_14084_46812# a_14035_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2550 VDD a_5937_45572# a_8034_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2551 a_5342_30871# a_14456_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2552 a_17639_46660# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X2553 a_10809_44734# a_10057_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2554 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2555 VDD a_11823_42460# a_14853_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2556 a_20749_43396# a_20974_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2557 VDD a_11967_42832# a_16243_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2558 a_19511_42282# a_n913_45002# a_21125_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2559 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2560 a_1609_45572# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2561 a_17517_44484# a_16979_44734# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2562 a_20075_46420# a_19900_46494# a_20254_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2563 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2564 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2565 a_16020_45572# a_15903_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2566 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2567 a_20731_45938# a_20107_45572# a_20623_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2568 VDD a_n3420_39072# a_n2860_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2569 VSS a_22731_47423# a_13717_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2570 a_16855_45546# a_16680_45572# a_17034_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2571 a_18114_32519# a_22223_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2572 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2573 a_17339_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2574 a_n2472_45546# a_n2293_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2575 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2576 VSS a_18429_43548# a_16823_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2577 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2578 VSS a_8325_42308# a_8791_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2579 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2580 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2581 VSS a_768_44030# a_13076_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2582 VSS a_12861_44030# a_19692_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2583 VDD a_14495_45572# a_n881_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2584 a_18596_45572# a_18479_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2585 a_n2472_45002# a_n2293_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2586 VDD a_n881_46662# a_6431_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2587 a_5326_44056# a_5147_45002# a_5244_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2588 VSS a_22959_42860# a_14097_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2589 a_3445_43172# a_3357_43084# a_n2293_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2590 a_13003_42852# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2591 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2592 a_3503_45724# a_3775_45552# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2593 C6_N_btm a_14401_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2594 a_19929_45028# a_19778_44110# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2595 a_3540_43646# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2596 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2597 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2598 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2599 VDD a_167_45260# a_117_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2600 a_6086_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2601 a_3147_46376# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2602 a_n1533_46116# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2603 VSS a_n3565_38216# a_n3607_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2604 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2605 a_5337_42558# a_5267_42460# a_4905_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2606 a_21542_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2607 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2608 a_10216_45572# a_10180_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2609 a_4699_43561# a_3080_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2610 a_3626_43646# a_3232_43370# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2611 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2612 VDD a_21613_42308# a_22775_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2613 a_16269_42308# a_15890_42674# a_16197_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2614 a_1067_42314# a_1184_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2615 VDD a_5937_45572# a_6945_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2616 a_22545_38993# a_22459_39145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2617 a_21356_42826# a_21381_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2618 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2619 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2620 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2621 VDD a_1307_43914# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2622 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2623 VSS a_19862_44208# a_19808_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2624 VDD a_5891_43370# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2625 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2626 a_20256_43172# a_18494_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2627 a_7927_46660# a_7411_46660# a_7832_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2628 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2629 VREF_GND a_13887_32519# C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2630 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2631 a_n2472_45546# a_n2293_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2632 a_17668_45572# a_n881_46662# a_17568_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X2633 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2634 a_4649_42852# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2635 a_6540_46812# a_3877_44458# a_6682_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2636 VDD a_6511_45714# a_6472_45840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2637 VSS a_15493_43396# a_19478_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2638 a_16664_43396# a_16547_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2639 VDD a_5068_46348# a_4955_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2640 a_9159_44484# a_5883_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2641 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2642 VSS a_10341_43396# a_22591_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2643 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2644 VSS a_17124_42282# a_4958_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2645 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2646 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2647 a_5267_42460# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2648 a_1138_42852# a_791_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2649 a_n4318_40392# a_n2840_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2650 a_n1644_44306# a_n1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2651 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2652 VDD a_1609_45822# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2653 a_5267_42460# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2654 VREF_GND a_17364_32525# C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2655 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2656 a_2127_44172# a_2675_43914# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2657 a_11787_45002# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2658 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2659 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2660 VSS a_19333_46634# a_19123_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2661 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2662 a_n2946_37984# a_n2956_38216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2663 a_3316_45546# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X2664 VSS a_13777_45326# a_13711_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2665 a_20712_42282# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2666 a_19479_31679# a_22223_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2667 a_20573_43172# a_20512_43084# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X2668 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2669 a_n2293_46634# a_14673_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2670 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2671 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2672 VSS a_526_44458# a_5457_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2673 a_33_46660# a_n133_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2674 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2675 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2676 VDD a_10903_43370# a_10849_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2677 VDD a_7754_40130# a_7754_40130# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2678 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2679 a_8495_42852# a_7871_42858# a_8387_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2680 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2681 a_5495_43940# a_5244_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2682 a_16842_45938# a_15765_45572# a_16680_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2683 VDD a_167_45260# a_2521_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2684 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2685 VSS a_n961_42308# a_n784_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2686 a_22780_40945# COMP_P a_22521_40599# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2687 VSS a_13259_45724# a_17303_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2688 VDD a_5937_45572# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2689 a_17538_32519# a_22959_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2690 a_21496_47436# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2691 a_11816_44260# a_11750_44172# a_10729_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2692 a_9801_43940# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2693 a_5742_30871# a_10723_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2694 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2695 a_2123_42473# a_n784_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2696 a_13565_43940# a_12891_46348# a_13483_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2697 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2698 a_7227_42852# a_n97_42460# a_7309_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2699 a_5257_43370# a_5907_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2700 VDD a_13747_46662# a_13607_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2701 a_1667_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2702 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2703 a_n2293_46098# a_5663_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2704 a_13003_42852# a_12379_42858# a_12895_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2705 a_2711_45572# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2706 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2707 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2708 a_16763_47508# a_16588_47582# a_16942_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2709 a_4883_46098# a_21363_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2710 VSS a_16751_45260# a_6171_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2711 VDD a_20835_44721# a_20766_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2712 a_11750_44172# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2713 VSS a_15861_45028# a_17668_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X2714 a_7845_44172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2715 a_15597_42852# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2716 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2717 VSS a_9223_42460# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X2718 VDD a_11967_42832# a_18083_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2719 a_13487_47204# a_13381_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X2720 a_13297_45572# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X2721 a_n923_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2722 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2723 C2_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2724 C10_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2725 VDD a_n3565_38216# a_n3690_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2726 a_6101_43172# a_5891_43370# a_5755_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2727 a_11901_46660# a_11735_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2728 a_16979_44734# a_14539_43914# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2729 VSS a_14955_47212# a_10227_46804# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2730 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2731 a_18443_44721# a_18248_44752# a_18753_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2732 VDD a_18909_45814# a_18799_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2733 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2734 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2735 a_1431_46436# a_1138_42852# a_1337_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2736 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2737 VDD a_n4064_37984# a_n2216_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2738 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2739 VDD a_22521_40599# a_22469_40625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2740 a_18443_44721# a_18287_44626# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2741 VDD a_768_44030# a_5326_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2742 VSS a_n4209_39304# a_n4251_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2743 a_n357_42282# a_21356_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2744 VSS a_n2288_47178# a_n2312_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2745 a_491_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2746 a_n901_46420# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2747 VSS a_3483_46348# a_15301_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2748 VCM a_1606_42308# C1_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2749 VDD a_20712_42282# a_10193_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2750 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 a_5068_46348# a_5204_45822# a_5210_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2752 a_14033_45822# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2753 VSS a_11599_46634# a_20107_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2754 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2755 w_1575_34946# EN_VIN_BSTR_P VDD w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2756 VSS a_6761_42308# a_7227_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2757 VDD a_13661_43548# a_15595_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2758 a_9803_42558# a_n97_42460# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2759 VDD a_10227_46804# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2760 a_n1177_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2761 VREF_GND a_n3420_39616# C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2762 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2763 a_601_46902# a_383_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2764 a_5024_45822# a_n443_46116# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2765 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2766 a_17701_42308# a_17531_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2767 VSS a_12861_44030# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X2768 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X2769 a_4808_45572# a_1823_45246# a_4419_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2770 a_6598_45938# a_6472_45840# a_6194_45824# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2771 a_n229_43646# a_n2497_47436# a_n447_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2772 a_n3607_38304# a_n3674_38216# a_n3690_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2773 VSS a_6969_46634# a_6903_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2774 a_18214_42558# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2775 a_491_47026# a_n133_46660# a_383_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2776 VSS a_4883_46098# a_10355_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2777 VDD a_16327_47482# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2778 VDD a_4646_46812# a_6031_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2779 VSS a_n1613_43370# a_n1655_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2780 a_6812_45938# a_6598_45938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2781 a_8147_43396# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2782 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2783 a_12427_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X2784 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2785 VDD a_19594_46812# a_19551_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2786 VSS a_1736_39043# a_1239_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2787 a_n4318_37592# a_n1736_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2788 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2789 VSS a_2698_46116# a_2804_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2790 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2791 a_1414_42308# a_1067_42314# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2792 VSS a_5649_42852# a_22223_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2793 VDD a_13259_45724# a_14797_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2794 a_n2288_47178# a_n2109_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2795 a_4817_46660# a_4651_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2796 a_8062_46155# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2797 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2798 a_13296_44484# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2799 VDD a_20623_43914# a_20365_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2800 a_11601_46155# a_11309_47204# a_11387_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2801 a_10210_45822# a_8746_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2802 a_18287_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2803 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2804 VSS a_11189_46129# a_11133_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2805 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2806 a_6431_45366# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2807 a_6109_44484# a_5518_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2808 a_14021_43940# a_13483_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2809 a_17499_43370# a_17324_43396# a_17678_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2810 a_3495_45348# a_3429_45260# a_3316_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X2811 VDD a_1115_44172# a_n2293_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2812 VDD a_19787_47423# a_19594_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2813 a_18707_42852# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2814 a_19787_47423# START VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2815 a_8667_46634# a_8492_46660# a_8846_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2816 a_1208_46090# a_n881_46662# a_1431_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2817 a_5431_46482# a_n1151_42308# a_5068_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2818 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2819 a_n2302_39866# a_n2442_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2820 VSS a_n2438_43548# a_2443_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2821 a_18797_44260# a_13661_43548# a_18451_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2822 a_19551_46910# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2823 VDD a_8953_45546# a_8049_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2824 a_8697_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2825 VDD a_10341_43396# a_22591_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2826 a_12005_46116# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2827 VSS a_12861_44030# a_18911_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2828 a_1241_43940# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X2829 VSS a_2123_42473# a_1184_42692# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2830 a_16285_47570# a_16241_47178# a_16119_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2831 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2832 a_1423_45028# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2833 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2834 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2835 a_10617_44484# a_10440_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2836 C7_P_btm a_n4064_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2837 VSS a_961_42354# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2838 VDD a_4704_46090# a_1823_45246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2839 a_18479_47436# a_20075_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2840 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2841 VDD a_9313_45822# a_11459_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2842 a_n1809_44850# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2843 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2844 a_19987_42826# a_10193_42453# a_20573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2845 VSS a_3785_47178# a_3815_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 VDD a_5891_43370# a_8375_44464# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2847 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2848 VSS a_9863_46634# a_2063_45854# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X2849 a_7920_46348# a_n1151_42308# a_8062_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2850 a_19721_31679# a_22959_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2851 a_19808_44306# a_19778_44110# a_19328_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2852 VDD a_10193_42453# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2853 VDD a_15559_46634# a_13059_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2854 VDD a_11189_46129# a_11601_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2855 a_5263_45724# a_5257_43370# a_5437_45600# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2856 a_12495_44260# a_12429_44172# a_10949_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X2857 VSS a_n2840_43370# a_n4318_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2858 a_15037_43396# a_14205_43396# a_14955_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2859 VSS a_4915_47217# a_12891_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2860 a_14084_46812# a_13885_46660# a_14226_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2861 a_6452_43396# a_6293_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2862 a_7705_45326# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2863 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2864 a_16981_45144# a_16922_45042# a_16886_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2865 a_1115_44172# a_1307_43914# a_1241_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2866 a_19478_44306# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2867 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2868 a_4223_44672# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2869 a_7174_31319# a_20107_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2870 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2871 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2872 VDD a_10227_46804# a_15051_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2873 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2874 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2875 a_n2833_47464# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2876 VSS a_8103_44636# a_7640_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2877 a_15146_44811# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2878 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2879 a_2903_45348# a_n971_45724# a_2809_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2880 VSS a_3537_45260# a_8103_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2881 VSS a_21137_46414# a_21071_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2882 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2883 VSS a_1414_42308# a_2889_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2884 VDD a_1848_45724# a_1799_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2885 VSS a_19279_43940# a_21398_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2886 a_1736_39587# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2887 VSS a_n13_43084# a_n1853_43023# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2888 a_18479_45785# a_19268_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2889 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2890 VSS a_22485_44484# a_20974_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2891 VSS a_n3420_37984# a_n2946_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2892 a_5275_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2893 a_5841_44260# a_5495_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2894 C5_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2895 a_n2661_45546# a_4093_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2896 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2897 VSS a_5497_46414# a_5431_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2898 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2899 VDD a_19339_43156# a_19326_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2900 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2901 a_8137_45348# a_8049_45260# a_n2293_42834# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2902 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2903 VDD a_6123_31319# a_7963_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2904 VDD a_12861_44030# a_17339_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2905 a_10849_43646# a_10807_43548# a_10765_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2906 VSS a_13507_46334# a_18997_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2907 a_8560_45348# a_3483_46348# a_8488_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2908 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2909 a_13249_42308# a_13070_42354# a_13333_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2910 a_6969_46634# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2911 a_n2216_37984# a_n2810_45572# a_n2302_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2912 VSS a_22223_46124# a_20205_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2913 a_6194_45824# a_6511_45714# a_6469_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2914 a_17613_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2915 a_n229_43646# a_n97_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2916 VSS a_n1613_43370# a_n1379_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2917 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2918 VSS a_13747_46662# a_19862_44208# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2919 a_22821_38993# a_22400_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2920 a_17303_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2921 a_8649_43218# a_8605_42826# a_8483_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2922 VSS a_n901_46420# a_n967_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2923 a_15004_44636# a_13556_45296# a_15146_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2924 a_11186_47026# a_10467_46802# a_10623_46897# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2925 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2926 VSS a_526_44458# a_4169_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2927 a_n23_45546# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2928 a_3353_43940# a_2998_44172# a_2675_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2929 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2930 a_18326_43940# a_18079_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2931 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2932 a_20922_43172# a_19862_44208# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X2933 a_10334_44484# a_10157_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2934 VSS a_742_44458# a_1756_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2935 C5_P_btm a_5934_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2936 a_n2017_45002# a_19987_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X2937 a_n2956_38216# a_n2472_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2938 VDD a_10193_42453# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2939 a_13885_46660# a_13607_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2940 VDD a_8191_45002# a_n2293_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2941 VSS RST_Z a_7754_39964# VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X2942 VSS a_4223_44672# a_n2497_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2943 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2944 a_4699_43561# a_3080_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2945 a_19511_42282# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2946 a_n1991_46122# a_n2157_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2947 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2948 VSS a_19692_46634# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2949 VDD a_22591_43396# a_14209_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2950 VDD a_7499_43078# a_8746_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2951 a_n971_45724# a_104_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2952 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2953 a_20447_31679# a_22959_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2954 VDD a_15493_43940# a_22959_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2955 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2956 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2957 a_18147_46436# a_17339_46660# a_17957_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2958 a_8336_45822# a_8270_45546# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2959 VDD a_13527_45546# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X2960 a_n4334_39616# a_n4318_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2961 a_n2956_39304# a_n2840_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2962 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2963 VDD a_584_46384# a_766_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2964 a_11361_45348# a_10907_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2965 VDD a_11599_46634# a_11735_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2966 a_19431_45546# a_19256_45572# a_19610_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2967 VSS a_9290_44172# a_12710_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X2968 VDD a_11323_42473# a_10807_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2969 a_2266_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2970 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2971 a_2982_43646# a_2479_44172# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2972 a_18280_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2973 VDD a_8492_46660# a_8667_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2974 C1_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2975 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2976 VDD a_n1076_46494# a_n901_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2977 a_n4251_38528# a_n4318_38680# a_n4334_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2978 a_4361_42308# a_3823_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2979 VDD a_11967_42832# a_12379_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2980 VDD a_21811_47423# a_20916_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2981 VDD a_11599_46634# a_13759_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2982 a_18985_46122# a_18819_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2983 VDD a_n971_45724# a_3775_45552# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2984 VDD a_5649_42852# a_22223_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2985 VSS a_5343_44458# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2986 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2987 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2988 VSS a_3090_45724# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X2989 a_20528_45572# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2990 a_13487_47204# a_13717_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2991 VREF_GND a_13678_32519# C2_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2992 VDD a_20269_44172# a_19319_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2993 a_5807_45002# a_16763_47508# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X2994 VSS a_16327_47482# a_16285_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2995 a_n23_44458# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2996 VDD a_n1059_45260# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2997 a_1847_42826# a_2351_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2998 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2999 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3000 a_19553_46090# a_19335_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3001 VDD a_n2840_45546# a_n2810_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3002 VSS a_3503_45724# a_3218_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X3003 a_15037_45618# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3004 a_14537_43646# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3005 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3006 a_6671_43940# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3007 a_n1699_43638# a_n1917_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3008 C6_P_btm a_n3420_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3009 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3010 VSS a_5111_44636# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3011 VDD a_9313_44734# a_22959_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3012 a_2124_47436# a_2063_45854# a_2266_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3013 VSS a_9625_46129# a_9569_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3014 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3015 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3016 VDD a_19279_43940# a_21398_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3017 VDD a_3483_46348# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3018 a_6171_42473# a_5932_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3019 a_17568_45572# a_8696_44636# a_17478_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3020 a_18588_44850# a_18374_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3021 a_18451_43940# a_18579_44172# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3022 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3023 VSS a_5755_42308# a_5932_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3024 a_2959_46660# a_2609_46660# a_2864_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3025 a_21359_45002# a_21513_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3026 a_7_47243# a_n746_45260# a_n452_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3027 a_15227_46910# a_3090_45724# a_15009_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3028 a_14493_46090# a_14275_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3029 a_19478_44306# a_15493_43396# a_19478_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X3030 a_7287_43370# a_7112_43396# a_7466_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3031 a_12251_46660# a_11901_46660# a_12156_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3032 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3033 a_8495_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3034 a_n4251_37440# a_n4318_37592# a_n4334_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3035 a_11633_42558# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3036 VDD a_7276_45260# a_7227_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3037 VSS a_2479_44172# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3038 a_15279_43071# a_5342_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3039 VREF_GND a_14401_32519# C6_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3040 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3041 VDD a_n815_47178# a_n785_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3042 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3043 a_1239_47204# a_1209_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3044 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3045 VDD a_3877_44458# a_3699_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3046 a_9313_45822# a_5937_45572# a_9241_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3047 a_20841_45814# a_20623_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3048 VDD a_805_46414# a_835_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3049 a_12379_46436# a_12005_46116# a_n1741_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3050 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3051 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3052 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3053 a_961_42354# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3054 a_n2956_39768# a_n2840_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3055 a_n1741_47186# a_12594_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3056 VDD a_5257_43370# a_3905_42865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3057 VSS a_n473_42460# a_n1761_44111# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3058 a_13163_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X3059 VDD a_10227_46804# a_9863_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3060 a_10210_45822# a_10586_45546# a_10053_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3061 VSS a_4185_45028# a_22959_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3062 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3063 VDD a_n2438_43548# a_n2065_43946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3064 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3065 a_5457_43172# a_5111_44636# a_5111_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3066 VDD a_11787_45002# a_11652_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3067 a_10695_43548# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3068 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3069 a_13059_46348# a_15559_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3070 VDD a_n23_44458# a_7_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3071 a_12891_46348# a_4915_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3072 a_8023_46660# a_7577_46660# a_7927_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3073 VSS a_10057_43914# a_9672_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3074 a_n237_47217# a_8667_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X3075 a_n143_45144# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3076 a_20637_44484# a_20159_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3077 a_4520_42826# a_4905_42826# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3078 VSS a_n971_45724# a_8423_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X3079 VSS RST_Z a_8530_39574# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3080 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3081 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3082 a_8697_45822# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3083 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3084 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3085 VSS a_3626_43646# a_19647_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3086 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3087 VDD a_1209_47178# a_1239_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3088 a_3094_47243# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3089 a_15051_42282# a_15486_42560# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3090 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3091 VDD a_13661_43548# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3092 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3093 a_5167_46660# a_4817_46660# a_5072_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3094 VSS a_10835_43094# a_10796_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3095 VDD a_20708_46348# a_20411_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3096 VSS a_16327_47482# a_18005_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3097 VSS a_16292_46812# a_15811_47375# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3098 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3099 a_9482_43914# a_9838_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3100 a_20623_46660# a_20273_46660# a_20528_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3101 VDD a_12594_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3102 a_18374_44850# a_18287_44626# a_17970_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3103 a_16750_47204# a_15673_47210# a_16588_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3104 a_6545_47178# a_6419_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3105 a_8783_44734# a_8696_44636# a_8701_44490# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3106 a_175_44278# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3107 VDD a_22223_43396# a_13887_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3108 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3109 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3110 VDD a_18479_47436# a_20935_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3111 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3112 VSS a_5907_46634# a_5841_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3113 a_5745_43940# a_5883_43914# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3114 a_3754_38470# a_7754_38470# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3115 a_1110_47026# a_33_46660# a_948_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3116 a_16434_46987# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3117 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3118 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3119 a_13381_47204# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3120 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3121 a_2998_44172# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3122 a_20974_43370# a_22485_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3123 VDD a_4921_42308# a_5755_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3124 a_10991_42826# a_10835_43094# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3125 VDD a_6851_47204# a_7227_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3126 a_3052_44056# a_2998_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X3127 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3128 a_3177_46902# a_2959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3129 VSS a_1208_46090# a_472_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3130 a_9241_44734# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3131 a_n1699_43638# a_n1917_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3132 CAL_N a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3133 a_22365_46825# EN_OFFSET_CAL VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3134 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3135 VSS a_13163_45724# a_11962_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3136 a_3055_46660# a_2609_46660# a_2959_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3137 a_19326_42852# a_18249_42858# a_19164_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3138 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3139 a_9885_43646# a_8270_45546# a_9803_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3140 VDD a_18597_46090# a_16375_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3141 a_19431_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3142 VSS a_22959_43396# a_17364_32525# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3143 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3144 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3145 VSS a_n1177_44458# a_n1243_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3146 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3147 VSS a_n23_45546# a_n89_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3148 a_n452_47436# a_n746_45260# a_n310_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3149 a_2952_47436# a_n1151_42308# a_3094_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3150 VDD a_12816_46660# a_12991_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3151 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3152 a_7499_43940# a_7640_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3153 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X3154 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3155 a_4235_43370# a_3935_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X3156 a_5105_45348# a_4558_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3157 a_18051_46116# a_765_45546# a_17957_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X3158 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3159 a_n1441_43940# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3160 a_15301_44260# a_15227_44166# a_14955_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3161 a_n746_45260# a_n1177_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3162 VSS a_n3565_38502# a_n3607_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3163 a_n2840_43914# a_n2661_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3164 a_6809_43396# a_6765_43638# a_6643_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3165 VSS a_376_46348# a_171_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3166 a_19443_46116# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3167 VSS a_13059_46348# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3168 VSS a_8199_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3169 a_7499_43940# a_3090_45724# a_7281_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3170 a_9165_43940# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3171 a_453_43940# a_175_44278# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3172 a_9885_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3173 a_n3674_39304# a_n2840_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3174 a_2959_46660# a_2443_46660# a_2864_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3175 a_14543_46987# a_13885_46660# a_14084_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3176 VDD a_413_45260# a_22959_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3177 a_17969_45144# a_16375_45002# a_17896_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X3178 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3179 a_16292_46812# a_n743_46660# a_16434_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3180 a_21188_46660# a_20107_46660# a_20841_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3181 a_12251_46660# a_11735_46660# a_12156_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3182 a_4365_46436# a_4185_45028# a_n1925_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3183 a_n998_44484# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3184 VDD a_3177_46902# a_3067_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3185 a_7577_46660# a_7411_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3186 VDD a_n2472_45546# a_n2956_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3187 a_14976_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3188 a_10835_43094# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3189 a_12638_46436# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3190 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3191 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3192 VSS a_13661_43548# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3193 a_12839_46116# a_12891_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3194 VSS a_3090_45724# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3195 VSS a_22000_46634# a_15227_44166# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3196 VSS a_n863_45724# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3197 a_14209_32519# a_22591_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3198 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3199 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3200 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3201 a_n2661_43922# a_12465_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3202 a_n2012_43396# a_n2129_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3203 VSS a_11823_42460# a_14635_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3204 a_19692_46634# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3205 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3206 VSS a_4520_42826# a_4093_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3207 a_5013_44260# a_3905_42865# a_5025_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3208 a_8018_44260# a_7499_43078# a_7911_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X3209 VDD a_11823_42460# a_14358_43442# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3210 a_167_45260# a_2202_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3211 a_20254_46482# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3212 VDD a_10405_44172# a_8016_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X3213 VIN_N EN_VIN_BSTR_N C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3214 a_742_44458# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3215 VSS a_19332_42282# a_4190_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3216 a_14840_46494# a_13925_46122# a_14493_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3217 VSS a_1414_42308# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3218 a_20356_42852# a_18184_42460# a_20256_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X3219 a_19006_44850# a_18287_44626# a_18443_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3220 a_9420_43940# a_768_44030# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3221 VDD a_10903_43370# a_12005_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3222 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3223 VSS a_12861_44030# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3224 VSS a_13661_43548# a_15685_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3225 C4_P_btm a_6123_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3226 a_13575_42558# a_n97_42460# a_13657_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3227 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3228 a_8667_46634# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3229 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3230 VDD a_n971_45724# a_n229_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3231 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3232 a_21335_42336# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3233 VSS a_n3565_37414# a_n3607_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3234 a_n2946_38778# a_n2956_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3235 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3236 VSS a_13351_46090# a_10903_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3237 a_14309_45028# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3238 VSS a_413_45260# a_22959_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3239 a_743_42282# a_12549_44172# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3240 VDD a_3877_44458# a_4185_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3241 a_13105_45348# a_13017_45260# a_n2661_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3242 VSS a_6545_47178# a_6575_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3243 a_8229_43396# a_7499_43078# a_8147_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3244 a_19551_46910# a_19466_46812# a_19333_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3245 a_18280_46660# a_12549_44172# a_17609_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3246 VSS a_18285_46348# a_18243_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X3247 a_6945_45028# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3248 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3249 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3250 a_20708_46348# a_20916_46384# a_20850_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3251 a_5167_46660# a_4651_46660# a_5072_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3252 VDD a_n1352_44484# a_n1177_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3253 a_15685_45394# a_15415_45028# a_15595_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3254 VDD a_10193_42453# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3255 a_21350_45938# a_20273_45572# a_21188_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3256 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3257 a_7639_45394# a_n1151_42308# a_7276_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3258 VSS a_526_44458# a_10149_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3259 a_7765_42852# a_7227_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3260 a_501_45348# a_413_45260# a_375_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3261 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3262 a_16547_43609# a_16414_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3263 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3264 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3265 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3266 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3267 a_13857_44734# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3268 a_n2661_46098# a_2107_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3269 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3270 VSS a_16327_47482# a_18953_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3271 VSS a_742_44458# a_1568_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3272 a_19273_43230# a_18083_42858# a_19164_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3273 a_6123_31319# a_7227_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3274 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3275 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3276 VDD a_2711_45572# a_4099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3277 a_12293_43646# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3278 C8_N_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3279 a_8035_47026# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3280 a_10306_45572# a_10193_42453# a_10216_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3281 a_18545_45144# a_13259_45724# a_18450_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X3282 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3283 a_n1423_46090# a_n1641_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3284 a_16977_43638# a_16759_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3285 VDD a_21855_43396# a_13678_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3286 VDD a_6540_46812# a_6491_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3287 VDD a_22223_43948# a_14401_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3288 VDD a_n863_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3289 C10_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3290 a_n2946_37690# a_n2956_37592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3291 a_5111_42852# a_4905_42826# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3292 VDD a_5263_45724# a_5204_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3293 a_n467_45028# a_n745_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3294 VSS a_765_45546# a_1208_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3295 VDD a_15095_43370# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3296 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X3297 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3298 VDD a_2957_45546# a_2905_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3299 a_8855_44734# a_4791_45118# a_8783_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3300 a_11963_45334# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3301 a_n2661_44458# a_11453_44696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X3302 VDD a_4915_47217# a_11415_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3303 a_n1741_47186# a_12005_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3304 a_3600_43914# a_3537_45260# a_3820_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3305 a_21588_30879# a_22223_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3306 a_1848_45724# a_2063_45854# a_1990_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3307 a_14537_46482# a_14493_46090# a_14371_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3308 a_10425_46660# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3309 a_16241_44734# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3310 a_3905_42865# a_5257_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3311 a_21811_47423# SINGLE_ENDED VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3312 a_19365_45572# a_18175_45572# a_19256_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3313 VDD a_22959_45572# a_20447_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3314 a_3090_45724# a_18911_45144# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3315 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3316 a_13777_45326# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3317 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3318 VCM a_5934_30871# C5_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3319 a_n3690_39616# a_n3674_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3320 a_17333_42852# a_16795_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3321 a_11525_45546# a_11962_45724# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3322 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3323 a_17595_43084# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3324 a_n13_43084# a_n755_45592# a_133_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X3325 a_n1838_35608# a_n1386_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3326 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3327 a_n2840_42282# a_n2661_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3328 a_20193_45348# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3329 a_20719_46660# a_20273_46660# a_20623_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3330 a_1756_43548# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3331 VSS a_n1613_43370# a_n1379_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3332 a_n2472_43914# a_n2293_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3333 a_n2302_39072# a_n2312_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3334 a_14456_42282# a_14635_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3335 VDD a_20075_46420# a_20062_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3336 VSS a_2711_45572# a_4099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3337 a_4927_45028# a_5147_45002# a_5105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3338 a_21381_43940# a_21115_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3339 VSS a_10227_46804# a_10185_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3340 a_n3607_38528# a_n3674_38680# a_n3690_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3341 a_4169_42308# a_1823_45246# a_3823_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X3343 VDD a_20894_47436# a_20843_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3344 a_4704_46090# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3345 VSS a_n913_45002# a_6761_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3346 VDD a_12465_44636# a_22223_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3347 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3348 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3349 VDD a_20193_45348# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3350 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3351 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3352 VDD a_5257_43370# a_3357_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3353 VSS a_14113_42308# a_16522_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3354 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3355 a_13460_43230# a_12379_42858# a_13113_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3356 a_19240_46482# a_19123_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3357 a_5829_43940# a_5495_43940# a_5745_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3358 a_22609_37990# a_22521_39511# CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3359 a_10227_46804# a_14955_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3360 VSS a_21487_43396# a_13467_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3361 VDD a_7287_43370# a_7274_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3362 VDD a_12861_44030# a_18911_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X3363 a_14955_43940# a_14537_43396# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3364 a_15953_42852# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3365 a_9114_42852# a_8037_42858# a_8952_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3366 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3367 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3368 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3369 VSS a_8199_44636# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3370 a_18780_47178# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3371 VDD a_15227_44166# a_18285_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3372 a_16375_45002# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3373 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3374 a_15279_43071# a_5342_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3375 a_10193_42453# a_20712_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3376 a_19335_46494# a_18985_46122# a_19240_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3377 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3378 a_5205_44484# a_5111_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3379 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3380 a_4842_47243# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3381 VSS a_685_42968# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3382 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3383 VSS a_22591_45572# a_19963_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3384 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3385 a_509_45572# a_n1099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3386 VSS a_11322_45546# a_12016_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X3387 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3388 a_20753_42852# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3389 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3390 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3391 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3392 a_16789_45572# a_15599_45572# a_16680_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3393 a_20362_44736# a_20640_44752# a_20596_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3394 a_13622_42852# a_12545_42858# a_13460_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3395 a_n1991_42858# a_n2157_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3396 a_15143_45578# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 VSS a_n746_45260# a_556_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3398 a_8701_44490# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3399 a_n3607_37440# a_n3674_37592# a_n3690_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3400 a_10775_45002# a_10951_45334# a_10903_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3401 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3402 VDD a_6151_47436# a_14955_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3403 a_15673_47210# a_15507_47210# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3404 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3405 a_19120_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X3406 a_20679_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3407 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3408 VDD a_10991_42826# a_10922_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X3409 a_5815_47464# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X3410 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X3411 a_n2956_37592# a_n2472_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3412 a_13667_43396# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X3413 VSS a_n1920_47178# a_n2312_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3414 VDD a_n4064_40160# a_n2216_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3415 a_5164_46348# a_4927_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X3416 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3417 a_15940_43402# a_12549_44172# a_15868_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3418 VDD a_4646_46812# a_4651_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3419 a_1427_43646# a_1049_43396# a_1209_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3420 a_19164_43230# a_18249_42858# a_18817_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3421 VDD a_12861_44030# a_21845_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3422 a_2982_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X3423 VDD a_3600_43914# a_3499_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3424 a_648_43396# a_526_44458# a_548_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3425 a_16409_43396# a_16243_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3426 VSS a_2063_45854# a_11136_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3427 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3428 VSS a_1823_45246# a_2202_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3429 a_10903_45394# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X3430 VDD a_n3420_39616# a_n2860_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3431 a_18243_46436# a_18189_46348# a_18147_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X3432 VSS a_n971_45724# a_3775_45552# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3433 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3434 a_4700_47436# a_4915_47217# a_4842_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3435 VDD a_6453_43914# a_n2661_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3436 VSS a_n2438_43548# a_n2433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3437 a_11813_46116# a_11387_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3438 VDD a_380_45546# a_n356_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3439 VDD a_10053_45546# a_9625_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3440 VDD a_12861_44030# a_19615_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3441 a_2253_43940# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X3442 VDD a_13113_42826# a_13003_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3443 a_765_45546# a_17609_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3444 a_3503_45724# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3445 VDD a_3699_46348# a_3160_47472# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3446 VDD a_9625_46129# a_10037_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X3447 VDD a_22223_45036# a_18114_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3448 a_18997_42308# a_18727_42674# a_18907_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3449 a_5755_42852# a_n97_42460# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3450 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3451 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3452 a_12281_43396# a_n913_45002# a_12293_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3453 VDD a_10533_42308# a_10723_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3454 VSS a_9863_47436# a_9804_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3455 a_8049_45260# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3456 a_11387_46482# a_11133_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3457 VDD a_21005_45260# a_19778_44110# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3458 VDD a_8791_42308# a_5934_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3459 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3460 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3461 a_895_43940# a_644_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3462 VSS a_n3420_38528# a_n2946_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3463 VDD a_4646_46812# a_7871_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3464 a_3067_47026# a_2443_46660# a_2959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3465 a_19256_45572# a_18341_45572# a_18909_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3466 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3467 C3_P_btm a_n4064_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3468 VSS a_2713_42308# a_2903_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3469 a_9863_47436# a_2063_45854# a_10037_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3470 a_15037_45618# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3471 a_3726_37500# CAL_P a_11206_38545# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3472 a_10991_42826# a_10796_42968# a_11301_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3473 a_2127_44172# a_1307_43914# a_2253_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3474 a_1823_45246# a_4704_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3475 VDD a_n2438_43548# a_n2433_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3476 a_17678_43396# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3477 a_n452_47436# a_n237_47217# a_n310_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3478 VDD a_10903_43370# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X3479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3480 a_3080_42308# a_2903_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3481 a_18057_42282# a_n1059_45260# a_18310_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3482 VSS a_n452_45724# a_n1853_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3483 a_n3674_39768# a_n2472_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3484 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3485 a_8846_46660# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3486 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3487 a_22365_46825# EN_OFFSET_CAL VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3488 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X3489 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3490 a_n89_45572# a_n743_46660# a_n452_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3491 a_n2472_42282# a_n2293_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3492 VSS a_n2840_45002# a_n2810_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3493 a_15928_47570# a_15811_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3494 a_518_46482# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3495 a_15463_44811# a_11691_44458# a_15004_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3496 VSS a_17767_44458# a_17715_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3497 a_20556_43646# a_19692_46634# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3498 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3499 a_14309_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3500 a_16237_45028# a_16375_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3501 a_8791_43396# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3502 VDD a_n4209_38216# a_n4334_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3503 a_9061_43230# a_7871_42858# a_8952_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3504 a_22780_39857# a_22465_38105# a_22521_39511# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3505 a_1568_43370# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3506 VDD a_n1423_42826# a_n1533_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3507 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3508 a_13575_42558# a_n97_42460# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3509 a_6667_45809# a_6511_45714# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3510 a_3754_39964# a_7754_39964# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3511 VSS a_9290_44172# a_10586_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3512 a_16115_45572# a_15765_45572# a_16020_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3513 VDD a_18911_45144# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X3514 a_2725_42558# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3515 a_18504_43218# a_17333_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3516 VDD a_3499_42826# a_n2293_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3517 a_16979_44734# a_14539_43914# a_17061_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3518 a_2253_43940# a_2479_44172# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3519 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3520 VSS a_1307_43914# a_3681_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3521 a_n310_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3522 a_5025_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3523 VSS a_626_44172# a_648_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3524 VSS a_n3420_37440# a_n2946_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3525 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3526 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3527 a_21356_42826# a_21381_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3528 a_16877_43172# a_16823_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3529 a_20841_46902# a_20623_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3530 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3531 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3532 VSS a_6171_45002# a_6125_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3533 VSS a_17595_43084# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3534 a_21137_46414# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3535 a_5883_43914# a_8333_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3536 a_20766_44850# a_20640_44752# a_20362_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3537 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3538 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3539 a_805_46414# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3540 a_1176_45822# a_997_45618# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3541 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3542 a_21887_42336# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3543 VSS a_11967_42832# a_18083_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3544 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3545 VDD a_1823_45246# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3546 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3547 a_21513_45002# a_21363_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3548 a_8704_45028# a_5937_45572# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3549 a_3232_43370# a_1823_45246# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3550 a_22780_40081# en_comp a_22521_40055# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3551 a_13333_42558# a_13291_42460# a_13249_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3552 a_13661_43548# a_18780_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3553 a_5497_46414# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3554 a_12749_45572# a_12549_44172# a_12649_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X3555 VSS a_n2840_43914# a_n4318_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3556 a_15037_44260# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3557 VSS a_22223_45572# a_19479_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3558 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X3559 VDD a_n2438_43548# a_n133_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3560 VDD a_n984_44318# a_n809_44244# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3561 VDD a_14815_43914# a_n2293_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3562 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3563 VDD a_22521_39511# a_22469_39537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3564 a_11530_34132# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3565 a_8128_46384# a_7903_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3566 VDD a_7281_43914# a_7229_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3567 VDD a_13507_46334# a_18907_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3568 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3569 a_479_46660# a_33_46660# a_383_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3570 VSS a_6667_45809# a_6598_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3571 VDD a_13904_45546# a_12594_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3572 VDD a_n881_46662# a_n1021_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3573 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3574 a_8568_45546# a_8953_45546# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3575 a_17767_44458# a_17970_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3576 VSS a_22400_42852# a_22780_40945# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3577 VREF a_19479_31679# C1_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3578 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3579 VDD a_n755_45592# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3580 a_16241_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3581 a_10867_43940# a_7499_43078# a_10405_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3582 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3583 VDD a_10723_42308# a_5742_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3584 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3585 a_20556_43646# a_20974_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3586 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3587 a_4574_45260# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3588 a_13483_43940# a_13249_42308# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3589 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3590 VDD a_20159_44458# a_19321_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X3591 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3592 a_2583_47243# a_584_46384# a_2124_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3593 a_22612_30879# a_22959_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3594 VDD a_8349_46414# a_8379_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3595 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3596 VSS a_768_44030# a_2711_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3597 a_n2216_40160# a_n2312_40392# a_n2302_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X3598 VSS a_14456_42282# a_5342_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3599 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3600 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3601 a_11608_46482# a_n1151_42308# a_11387_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3602 a_5093_45028# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3603 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3604 a_19862_44208# a_13747_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3605 VDD a_15227_44166# a_15597_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3606 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3607 a_19335_46494# a_18819_46122# a_19240_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3608 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3609 VSS a_1736_39587# a_1239_39587# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3610 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3611 a_8953_45546# a_8685_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3612 a_n4318_38216# a_n2472_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3613 a_18249_42858# a_18083_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3614 a_12816_46660# a_11735_46660# a_12469_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3615 a_19268_43646# a_13661_43548# a_19177_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X3616 a_13258_32519# a_19647_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3617 a_20256_42852# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X3618 VDD a_16680_45572# a_16855_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3619 VSS a_n447_43370# a_n2129_43609# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3620 a_20528_45572# a_19466_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3621 a_11525_45546# a_10586_45546# a_11778_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3622 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3623 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3624 VDD a_2711_45572# a_20107_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3625 a_16147_45260# a_17478_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3626 a_n2109_45247# a_n2017_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3627 a_19610_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3628 a_19963_31679# a_22591_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3629 a_5837_43172# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3630 a_n143_45144# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3631 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3632 VDD a_22959_47212# a_22612_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3633 a_n310_45572# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3634 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3635 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3636 a_15015_46420# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3637 VSS a_7227_45028# a_7230_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3638 a_20596_44850# a_20159_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3639 a_2957_45546# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3640 VSS a_14579_43548# a_14537_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3641 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3642 VDD a_11599_46634# a_15507_47210# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3643 VDD a_6151_47436# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3644 VSS a_5111_44636# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3645 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X3646 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3647 VDD a_20679_44626# a_20640_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3648 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3649 VDD COMP_P a_n1329_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3650 VSS a_19321_45002# a_20567_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3651 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3652 a_14513_46634# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3653 a_10903_43370# a_13351_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3654 VSS a_n2472_45002# a_n2956_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3655 a_10949_43914# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X3656 a_10149_43396# a_5111_44636# a_9803_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3657 VSS a_19431_45546# a_19365_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3658 VSS a_16922_45042# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X3659 a_16112_44458# a_14539_43914# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3660 a_13943_43396# a_11823_42460# a_13837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3661 C8_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3662 VDD a_4099_45572# a_3483_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3663 a_6197_43396# a_6031_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3664 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3665 a_n2840_46634# a_n2661_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3666 a_380_45546# a_n357_42282# a_603_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3667 a_18533_43940# a_18326_43940# a_18451_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3668 a_7309_42852# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3669 VDD a_n863_45724# a_2448_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3670 a_5932_42308# a_5755_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3671 a_16328_43172# a_n97_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3672 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3673 a_17583_46090# a_17715_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3674 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3675 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3676 VDD a_15433_44458# a_15463_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3677 a_n2267_43396# a_n2433_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3678 VDD a_n755_45592# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3679 VSS a_10991_42826# a_10922_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3680 a_5732_46660# a_4651_46660# a_5385_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3681 a_19615_44636# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X3682 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X3683 VDD a_5129_47502# a_5159_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3684 a_n2840_46090# a_n2661_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3685 a_n967_45348# a_n913_45002# a_n955_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3686 a_19006_44850# a_18248_44752# a_18443_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3687 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3688 VDD a_18817_42826# a_18707_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3689 a_15559_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X3690 a_9803_43646# a_8953_45546# a_9885_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3691 VDD a_3232_43370# a_9313_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3692 VDD a_n2840_42282# a_n3674_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3693 a_13460_43230# a_12545_42858# a_13113_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3694 a_20362_44736# a_20679_44626# a_20637_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3695 a_2713_42308# a_n913_45002# a_2725_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3696 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3697 a_16241_47178# a_16023_47582# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3698 a_14955_43396# a_14205_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3699 VSS a_n913_45002# a_10533_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3700 a_7466_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3701 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3702 VDD a_6151_47436# a_5907_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3703 a_16697_47582# a_15507_47210# a_16588_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3704 a_n2267_44484# a_n2433_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3705 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3706 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3707 a_13693_46688# a_6755_46942# a_13607_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3708 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3709 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3710 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3711 VDD a_19778_44110# a_19741_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3712 a_2609_46660# a_2443_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3713 a_5708_44484# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X3714 a_18143_47464# a_18479_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3715 a_5263_46660# a_4817_46660# a_5167_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3716 VSS a_n2472_43914# a_n3674_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3717 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3718 a_12016_45572# a_11962_45724# a_11525_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3719 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3720 VSS a_18057_42282# a_n356_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3721 VDD a_21671_42860# a_3422_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3722 VDD a_8746_45002# a_8704_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3723 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3724 a_3411_47243# a_3160_47472# a_2952_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3725 a_n2840_46634# a_n2661_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3726 VSS a_7705_45326# a_7639_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3727 VSS a_167_45260# a_1423_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3728 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3729 VDD a_9396_43370# a_5111_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3730 a_743_42282# a_13661_43548# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3731 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3732 a_133_43172# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X3733 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3734 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3735 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3736 VDD a_20512_43084# a_19987_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X3737 a_1891_43646# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X3738 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3739 a_14485_44260# a_5807_45002# a_12465_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3740 a_n4318_39304# a_n2840_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3741 VIN_P EN_VIN_BSTR_P C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3742 VSS a_n357_42282# a_17141_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3743 a_11453_44696# a_17719_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X3744 VSS a_n1059_45260# a_8945_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3745 a_17701_42308# a_17531_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3746 a_13657_42558# a_11823_42460# a_13575_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3747 a_10545_42558# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3748 a_8292_43218# a_7765_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3749 a_16751_46987# a_5807_45002# a_16292_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3750 a_10586_45546# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3751 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3752 VSS a_16855_45546# a_16789_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3753 a_45_45144# a_n143_45144# a_n37_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3754 VDD a_3537_45260# a_4223_44672# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3755 a_3626_43646# a_1414_42308# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3756 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3757 VDD a_20107_42308# a_7174_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3758 a_3815_47204# a_3785_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3759 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3760 a_n83_35174# VDD EN_VIN_BSTR_P VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X3761 VCM a_5342_30871# C8_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3762 a_15567_42826# a_15743_43084# a_15953_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3763 VSS a_10341_42308# a_11554_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3764 VSS a_4791_45118# a_6640_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X3765 a_6755_46942# a_15015_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3766 a_2437_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3767 VDAC_Pi a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3768 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3769 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3770 a_9823_46155# a_9804_47204# a_9823_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3771 a_1990_45899# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3772 a_15743_43084# a_19339_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3773 a_5129_47502# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3774 VDD a_5385_46902# a_5275_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3775 a_9145_43396# a_8791_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3776 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3777 VDD a_20841_46902# a_20731_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3778 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3779 VIN_P EN_VIN_BSTR_P C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3780 VDD a_n785_47204# a_327_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3781 a_7276_45260# a_n1151_42308# a_7418_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3782 a_8103_44636# a_8375_44464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3783 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3784 a_4915_47217# a_12991_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3785 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3786 VDD a_8199_44636# a_8855_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3787 VDD a_12549_44172# a_21115_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3788 VDD a_2553_47502# a_2583_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3789 a_n327_42558# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3790 a_19864_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X3791 a_12800_43218# a_12089_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3792 VSS a_20623_43914# a_20365_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3793 VSS a_n743_46660# a_16501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3794 VSS a_22959_45036# a_19721_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3795 VSS a_11967_42832# a_16243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3796 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3797 a_n4318_38680# a_n2472_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3798 a_3363_44484# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3799 a_13483_43940# a_13249_42308# a_13565_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3800 a_7754_40130# RST_Z VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3801 VDD a_4235_43370# a_n2661_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3802 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3803 a_13249_42558# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3804 a_18504_43218# a_17333_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3805 a_n39_42308# a_n97_42460# a_n473_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3806 a_10210_45822# a_10180_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X3807 VSS a_11967_42832# a_20512_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3808 VSS a_n443_46116# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3809 VSS a_4646_46812# a_7411_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3810 a_20273_46660# a_20107_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3811 VDD a_11341_43940# a_22223_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3812 a_n2312_38680# a_n2104_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3813 VDD a_12791_45546# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X3814 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3815 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3816 a_19237_31679# a_22959_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3817 VDD a_19328_44172# a_19279_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X3818 VDD SMPL_ON_P a_n1605_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3819 VSS a_11967_42832# a_12379_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3820 VSS a_15227_44166# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3821 VDD a_18315_45260# a_18189_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X3822 a_10951_45334# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3823 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3824 VDD a_2123_42473# a_1184_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3825 a_4791_45118# a_4743_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3826 a_21195_42852# a_20922_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3827 a_4156_43218# a_3905_42865# a_3935_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3828 a_15227_44166# a_22000_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3829 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3830 a_n1899_43946# a_n2065_43946# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3831 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3832 a_n743_46660# a_n1021_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3833 a_n2293_45546# a_2274_45254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3834 a_11633_42308# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3835 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3836 a_20205_31679# a_22223_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3837 a_n2472_46634# a_n2293_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3838 a_2698_46116# a_2521_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3839 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3840 VDD a_10193_42453# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3841 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3842 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3843 a_22705_37990# a_22521_40055# a_22609_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3844 VDD a_n3565_38502# a_n3690_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3845 a_5342_30871# a_14456_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3846 VDD a_8325_42308# a_8791_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3847 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3848 a_548_43396# a_n863_45724# a_458_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3849 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3850 VSS a_1756_43548# a_1467_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X3851 a_288_46660# a_171_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3852 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3853 VDD a_17517_44484# a_22591_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3854 VSS a_n913_45002# a_19511_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3855 a_20894_47436# a_20990_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3856 a_15312_46660# a_14976_45028# a_15009_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3857 a_n2472_46090# a_n2293_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3858 VDD a_n2438_43548# a_n2157_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3859 VSS a_22959_43948# a_17538_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3860 C9_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3861 VDD a_n4064_38528# a_n2216_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3862 a_8037_42858# a_7871_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3863 a_n1736_43218# a_n1853_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3864 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3865 a_13527_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3866 VDD a_n2472_42282# a_n4318_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3867 a_n2661_43370# a_11415_45002# a_11361_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3868 VSS a_1343_38525# a_2113_38308# VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X3869 VDD a_22165_42308# a_22223_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3870 VDD a_n2840_42826# a_n3674_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3871 VSS a_14180_45002# a_13017_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3872 a_15681_43442# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3873 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3874 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3875 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3876 a_8488_45348# a_8199_44636# a_8191_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X3877 a_16588_47582# a_15673_47210# a_16241_47178# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3878 a_18220_42308# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X3879 a_n1423_46090# a_n1641_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3880 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3881 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3882 a_17609_46634# a_12549_44172# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3883 a_16115_45572# a_15599_45572# a_16020_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3884 VSS a_19700_43370# a_n97_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3885 VSS a_2124_47436# a_1209_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3886 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3887 a_15595_45028# a_15415_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3888 VDD a_6755_46942# a_12741_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3889 VSS a_19615_44636# a_18579_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3890 a_12545_42858# a_12379_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3891 a_16942_47570# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3892 a_8791_45572# a_7499_43078# a_8697_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3893 a_14853_42852# a_n913_45002# a_14635_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3894 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3895 a_8333_44056# a_4223_44672# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3896 VSS a_4958_30871# a_17531_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3897 a_6511_45714# a_4646_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3898 VDD a_10949_43914# a_10867_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X3899 a_17973_43940# a_17737_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X3900 a_18494_42460# a_18907_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3901 a_17061_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3902 a_n2472_46634# a_n2293_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3903 C2_P_btm a_3080_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3904 VSS a_5267_42460# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3905 VSS a_n2438_43548# a_n2065_43946# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3906 VDD a_7754_40130# a_3754_38470# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3907 VDD a_n357_42282# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3908 a_9159_45572# a_5937_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3909 a_3483_46348# a_4099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3910 a_8238_44734# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3911 VSS a_17517_44484# a_22591_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3912 VDD a_n3565_37414# a_n3690_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3913 VDD a_3381_47502# a_3411_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3914 VSS a_21613_42308# a_22775_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3915 a_10150_46912# a_10467_46802# a_10425_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3916 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3917 a_n2810_45572# a_n2840_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3918 a_13675_47204# a_n1435_47204# a_13569_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X3919 VSS a_11827_44484# a_22223_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3920 a_5518_44484# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X3921 VDD a_n4064_37440# a_n2216_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3922 a_22165_42308# a_21887_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3923 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3924 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3925 VDD a_22521_40055# a_22459_39145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3926 a_13678_32519# a_21855_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3927 a_n2312_40392# a_n2288_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3928 VDD a_8605_42826# a_8495_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3929 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3930 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3931 VDD a_20193_45348# a_21887_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3932 a_18691_45572# a_18341_45572# a_18596_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3933 a_13076_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3934 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3935 a_3600_43914# a_1307_43914# a_3992_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3936 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3937 a_4743_43172# a_3537_45260# a_4649_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3938 a_11387_46155# a_11309_47204# a_11387_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3939 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3940 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3941 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3942 a_22609_37990# a_22469_39537# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3943 a_11554_42852# a_10835_43094# a_10991_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3944 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3945 VDD a_2680_45002# a_2274_45254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3946 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3947 VSS a_9313_44734# a_22959_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3948 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3949 VDD a_n1177_43370# a_n1190_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3950 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X3951 VDD a_6755_46942# a_13556_45296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3952 a_n785_47204# a_n815_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3953 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3954 VDD a_n971_45724# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3955 a_n4251_40480# a_n4318_40392# a_n4334_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3956 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3957 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3958 a_19900_46494# a_18819_46122# a_19553_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3959 VSS a_n1386_35608# a_n1838_35608# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3960 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3961 a_12359_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3962 a_12561_45572# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X3963 a_10083_42826# a_10518_42984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3964 VSS a_10355_46116# a_8199_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3965 a_3422_30871# a_21671_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3966 a_5937_45572# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3967 a_21005_45260# a_21101_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X3968 VDD a_16327_47482# a_17767_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3969 a_12649_45572# a_10903_43370# a_12561_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3970 VSS a_19321_45002# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3971 a_5111_44636# a_9396_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3972 a_12469_46902# a_12251_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3973 a_21297_45572# a_20107_45572# a_21188_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3974 a_376_46348# a_584_46384# a_518_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3975 a_15146_44484# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3976 VIN_P EN_VIN_BSTR_P C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3977 VDD a_n971_45724# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3978 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3979 a_14180_45002# a_14537_43396# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3980 VDD a_10193_42453# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3981 a_18681_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3982 VSS a_15009_46634# a_14180_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3983 a_17829_46910# a_12549_44172# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X3984 a_2304_45348# a_2274_45254# a_2232_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3985 a_6598_45938# a_6511_45714# a_6194_45824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3986 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3987 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3988 a_5745_43940# a_5013_44260# a_5663_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3989 VDD a_10193_42453# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3990 a_5742_30871# a_10723_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3991 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3992 a_19478_44056# a_3090_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3993 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3994 a_10185_46660# a_10150_46912# a_9863_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3995 a_8192_45572# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3996 a_15890_42674# a_15764_42576# a_15486_42560# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3997 a_10835_43094# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3998 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3999 a_n699_43396# a_n1177_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4000 a_14033_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4001 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4002 a_6101_44260# a_1307_43914# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4003 a_7927_46660# a_7577_46660# a_7832_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4004 a_21496_47436# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X4005 a_16721_46634# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4006 a_5826_44734# a_5147_45002# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X4007 VDD a_16763_47508# a_16750_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4008 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4009 VDD a_n746_45260# a_175_44278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4010 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4011 a_2813_43396# a_3232_43370# a_2982_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4012 a_6171_42473# a_5932_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4013 VDD a_601_46902# a_491_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4014 VSS a_4646_46812# a_6031_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4015 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4016 VDD a_1123_46634# a_1110_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4017 VSS a_13059_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4018 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4019 a_11787_45002# a_11963_45334# a_11915_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4020 VSS a_584_46384# a_2998_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4021 a_8292_43218# a_7765_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4022 VDD a_n2472_42826# a_n4318_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4023 a_1667_45002# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X4024 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4025 a_20731_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4026 a_8062_46482# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4027 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4028 a_n2216_38778# a_n2312_38680# a_n2302_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4029 VSS a_11599_46634# a_20107_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4030 a_13925_46122# a_13759_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4031 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4032 VSS a_n2104_46634# a_n2312_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4033 a_5385_46902# a_5167_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4034 a_n1177_44458# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4035 VDD a_7499_43078# a_10729_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4036 a_9803_43646# a_8953_45546# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4037 VDD a_19256_45572# a_19431_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4038 a_7911_44260# a_7845_44172# a_7542_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X4039 VDD a_5111_44636# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4040 VDD a_6761_42308# a_7227_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4041 VDD a_19553_46090# a_19443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4042 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4043 a_5205_44484# a_5343_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4044 a_22400_42852# a_22223_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4045 a_12603_44260# a_12549_44172# a_12495_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X4046 VSS a_18194_35068# a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4047 a_3638_45822# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X4048 a_17324_43396# a_16243_43396# a_16977_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4049 a_19452_47524# a_19386_47436# a_13747_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4050 a_5275_47026# a_4651_46660# a_5167_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4051 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4052 a_11915_45394# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X4053 a_14447_46660# a_n1151_42308# a_14084_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4054 a_20731_47026# a_20107_46660# a_20623_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4055 VSS a_n1613_43370# a_n1655_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4056 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4057 a_12800_43218# a_12089_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4058 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4059 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4060 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4061 VSS a_20712_42282# a_10193_42453# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4062 a_15720_42674# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4063 VSS a_n443_42852# a_421_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4064 a_14493_46090# a_14275_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4065 VDD a_11599_46634# a_15599_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4066 a_n659_45366# a_n746_45260# a_n745_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4067 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4068 a_n881_46662# a_14495_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4069 a_8685_43396# a_8147_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4070 C7_P_btm a_n4209_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4071 a_765_45546# a_17609_46634# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4072 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X4073 a_11554_42852# a_10796_42968# a_10991_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4074 a_19386_47436# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4075 a_8492_46660# a_7411_46660# a_8145_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4076 a_2063_45854# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4077 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4078 VDD a_15803_42450# a_15764_42576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4079 a_1337_46436# a_1176_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4080 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4081 VSS a_4419_46090# a_4365_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4082 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4083 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4084 VSS a_6575_47204# a_9067_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4085 a_n1331_43914# a_n1549_44318# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4086 VDD a_3537_45260# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4087 VSS a_11189_46129# a_11608_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4088 a_20835_44721# a_20640_44752# a_21145_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X4089 a_n327_42558# a_n97_42460# a_n473_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X4090 a_8147_43396# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X4091 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4092 a_19431_46494# a_18985_46122# a_19335_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4093 VDD a_12607_44458# a_n2661_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4094 VDD a_17324_43396# a_17499_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4095 a_8685_42308# a_8515_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4096 a_1414_42308# a_1067_42314# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4097 VDD a_4883_46098# a_10355_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4098 a_n2216_37690# a_n2810_45028# a_n2302_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4099 VDD a_10193_42453# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4100 VDD a_21356_42826# a_n357_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4101 a_16977_43638# a_16759_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4102 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4103 VSS a_n237_47217# a_8270_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4104 a_10555_43940# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4105 a_1049_43396# a_458_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4106 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4107 VDD a_n443_42852# a_742_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4108 a_8145_46902# a_7927_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4109 a_21613_42308# a_21335_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4110 VDD a_n23_45546# a_7_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4111 VSS a_16019_45002# a_15903_45785# VSS sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X4112 VCM a_5342_30871# C8_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4113 VDD a_2698_46116# a_2804_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4114 a_20935_43940# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4115 a_2713_42308# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4116 VDD a_n699_43396# a_4743_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4117 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4118 a_17591_47464# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4119 a_9223_42460# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4120 a_12741_44636# a_14537_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4121 a_2684_37794# a_1736_39587# a_1736_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4122 VDD a_20202_43084# a_21335_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4123 a_564_42282# a_743_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4124 a_15367_44484# a_13556_45296# a_15004_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4125 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4126 VSS a_n452_47436# a_n815_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4127 VDD a_2063_45854# a_9863_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4128 a_2981_46116# a_2804_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4129 VSS a_6511_45714# a_6472_45840# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4130 VSS a_13159_45002# a_13105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4131 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4132 a_9223_42460# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4133 VSS a_19987_42826# a_n2017_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X4134 a_20692_30879# a_22959_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4135 a_21188_45572# a_20273_45572# a_20841_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4136 a_9028_43914# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4137 VDD a_17715_44484# a_17737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4138 VSS a_n2840_44458# a_n4318_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4139 VSS a_15004_44636# a_14815_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4140 a_16759_43396# a_16243_43396# a_16664_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4141 a_4574_45260# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4142 a_17829_46910# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4143 VSS a_n443_46116# a_4880_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X4144 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4145 VDD a_1799_45572# a_1983_46706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4146 VDD a_21363_45546# a_21350_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4147 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X4148 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4149 a_13259_45724# a_17583_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4150 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4151 C1_P_btm a_n4064_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4152 VIN_P EN_VIN_BSTR_P C4_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4153 a_6575_47204# a_6545_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4154 VSS a_765_45546# a_380_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4155 VSS a_327_44734# a_501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4156 a_104_43370# a_n699_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4157 VDD a_22959_42860# a_14097_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4158 a_n2293_42282# a_3357_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4159 VSS a_6171_42473# a_5379_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4160 a_3935_42891# a_2382_45260# a_3935_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4161 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD a_8145_46902# a_8035_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4163 VDD a_n863_45724# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4164 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4165 a_17141_43172# a_n1059_45260# a_16795_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4166 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4167 a_15433_44458# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4168 VSS a_10193_42453# a_11897_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4169 VSS a_4791_45118# a_5066_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4170 VDD a_5691_45260# a_n2109_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4171 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4172 VDD a_1983_46706# a_n2661_46098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4173 a_15227_46910# a_15368_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4174 a_18753_44484# a_18374_44850# a_18681_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4175 a_15486_42560# a_15803_42450# a_15761_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X4176 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4177 a_6682_46987# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4178 a_n1079_45724# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4179 a_12429_44172# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X4180 a_1568_43370# a_1847_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4181 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4182 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4183 VDD a_7227_42308# a_6123_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4184 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4185 a_3457_43396# a_3232_43370# a_3626_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4186 a_7174_31319# a_20107_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4187 a_8952_43230# a_8037_42858# a_8605_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4188 VSS a_167_45260# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4189 a_13490_45067# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4190 a_4181_44734# a_3090_45724# a_n2497_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4191 VSS a_6171_45002# a_11909_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4192 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4193 a_33_46660# a_n133_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4194 a_16388_46812# a_17957_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X4195 VDD a_3218_45724# a_3175_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4196 a_8283_46482# a_n1151_42308# a_7920_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4197 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4198 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4199 VDD a_15279_43071# a_14579_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4200 VDD a_16763_47508# a_5807_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4201 VDD a_310_45028# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4202 a_n23_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4203 a_n1099_45572# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X4204 VDD a_10903_43370# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4205 a_3935_43218# a_3681_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4206 a_14949_46494# a_13759_46122# a_14840_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4207 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4208 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4209 a_6851_47204# a_6491_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4210 a_13556_45296# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4211 VDD a_n4315_30879# a_n4334_40480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4212 VSS a_15227_44166# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X4213 a_19987_42826# a_18494_42460# a_20356_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X4214 a_n2833_47464# a_n2497_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4215 a_3524_46660# a_2609_46660# a_3177_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4216 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4217 VSS a_22223_47212# a_21588_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4218 VSS a_6151_47436# a_6229_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X4219 a_18533_43940# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4220 a_14205_43396# a_13667_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4221 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4222 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4223 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4224 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4225 a_16377_45572# a_16333_45814# a_16211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4226 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X4227 a_10044_46482# a_n743_46660# a_9823_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4228 a_19113_45348# a_18911_45144# a_3090_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4229 VSS a_13720_44458# a_12607_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4230 a_n2860_37984# a_n2956_38216# a_n2946_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4231 a_2266_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4232 a_5837_43396# a_5111_44636# a_5147_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4233 a_5934_30871# a_8791_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4234 a_10861_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4235 VSS a_7920_46348# a_7715_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4236 a_14383_46116# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4237 a_2809_45348# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4238 a_2905_42968# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4239 a_6540_46812# a_6755_46942# a_6682_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4240 a_6709_45028# a_6431_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4241 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4242 VSS a_18494_42460# a_20193_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4243 a_n2442_46660# a_n2472_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4244 C7_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4245 a_13249_42308# a_13070_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4246 a_n1991_42858# a_n2157_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4247 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4248 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4249 a_13348_45260# a_12891_46348# a_13490_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4250 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X4251 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4252 a_17061_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4253 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4254 VDD a_18443_44721# a_18374_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4255 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4256 a_1512_43396# a_n443_46116# a_1209_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4257 VDD a_n3565_39304# a_n3690_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4258 VDD a_22591_44484# a_17730_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4259 VSS a_15803_42450# a_15764_42576# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4260 a_11901_46660# a_11735_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4261 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4262 a_21076_30879# a_22959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4263 a_3877_44458# a_3699_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4264 VDD a_n4064_39072# a_n2216_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4265 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4266 a_11691_44458# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4267 a_15368_46634# a_15143_45578# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X4268 VSS a_9028_43914# a_8975_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4269 a_2813_43396# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X4270 C8_N_btm a_17538_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4271 a_5093_45028# a_4558_45348# a_5009_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4272 VSS a_10193_42453# a_13921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4273 a_15597_42852# a_15567_42826# a_15095_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X4274 a_2553_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4275 VDD a_13059_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4276 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4277 a_3823_42558# a_3065_45002# a_3905_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4278 VDD a_526_44458# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4279 VSS a_1667_45002# a_n863_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4280 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4281 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4282 VDD a_21177_47436# a_20990_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4283 a_16855_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4284 a_5495_43940# a_5244_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4285 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4286 VSS a_19787_47423# a_19594_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4287 VDD a_22365_46825# a_20202_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4288 a_5063_47570# a_4915_47217# a_4700_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4289 a_n1736_46482# a_n1853_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4290 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4291 a_11322_45546# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4292 a_19787_47423# START VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4293 a_3754_39466# a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X4294 a_n4251_39616# a_n4318_39768# a_n4334_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4295 VDD a_9127_43156# a_9114_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4296 a_10384_47026# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4297 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4298 VSS a_11525_45546# a_11189_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4299 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4300 a_10729_43914# a_11750_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4301 a_4921_42308# a_n913_45002# a_4933_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4302 VSS a_n23_47502# a_n89_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4303 a_20528_46660# a_20411_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4304 VSS a_8568_45546# a_8162_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4305 a_13657_42558# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4306 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4307 VSS a_4223_44672# a_5205_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4308 a_18005_44484# a_17970_44736# a_17767_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4309 a_13837_43396# a_13259_45724# a_13749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4310 a_19177_43646# a_17339_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X4311 a_196_42282# a_375_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4312 a_791_42968# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4313 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4314 a_11309_47204# a_11031_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4315 VSS a_4646_46812# a_7871_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4316 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4317 a_n23_45546# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4318 a_18691_45572# a_18175_45572# a_18596_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4319 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4320 a_9885_42558# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4321 VSS a_4700_47436# a_3785_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4322 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4323 a_4361_42308# a_3823_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4324 VDD a_n2840_46634# a_n2956_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4325 a_4817_46660# a_4651_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4326 VDD a_13635_43156# a_13622_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4327 VDD a_n2438_43548# a_n2157_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4328 a_8415_44056# a_5343_44458# a_8333_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4329 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4330 VSS a_1307_43914# a_4156_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4331 a_n1699_44726# a_n1917_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4332 a_1525_44260# a_1467_44172# a_1115_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4333 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4334 a_14976_45028# a_14797_45144# a_15060_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X4335 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4336 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4337 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4338 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4339 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4340 VSS a_15959_42545# a_15890_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4341 VDD a_22469_40625# a_22705_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4342 a_n2312_39304# a_n1920_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4343 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4344 VIN_N EN_VIN_BSTR_N C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4345 VDD a_1736_39587# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X4346 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4347 VSS a_21363_45546# a_21297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4348 VDD a_n452_44636# a_n2129_44697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4349 a_19443_46116# a_18819_46122# a_19335_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4350 VDD a_7112_43396# a_7287_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4351 a_310_45028# a_n37_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4352 VDD a_5111_44636# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X4353 VDD EN_VIN_BSTR_N w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4354 a_17719_45144# a_17613_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4355 a_17499_43370# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4356 VDD a_12563_42308# a_5534_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4357 VSS a_13747_46662# a_19466_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4358 a_14112_44734# a_768_44030# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4359 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 a_n357_42282# a_21356_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4361 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4362 VDD a_3483_46348# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4363 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4364 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4365 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4366 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4367 a_14097_32519# a_22959_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4368 a_3094_47570# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4369 a_8270_45546# a_n237_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 a_8781_46436# a_8199_44636# a_8034_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4371 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4372 VSS a_3232_43370# a_11541_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4373 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4374 a_20841_46902# a_20623_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4375 a_13527_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4376 a_10533_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 a_17896_45144# a_16922_45042# a_17801_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X4378 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4379 a_18817_42826# a_18599_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4380 a_104_43370# a_n699_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4381 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4382 a_16211_45572# a_15765_45572# a_16115_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4383 VDD a_4223_44672# a_4181_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4384 VSS a_20835_44721# a_20766_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4385 a_19741_43940# a_19478_44306# a_19328_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4386 VDD a_13747_46662# a_14495_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4387 a_2487_47570# a_2063_45854# a_2124_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4388 VSS a_10809_44734# a_22959_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4389 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4391 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4392 VSS a_20567_45036# a_12549_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4393 a_21359_45002# a_21513_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4394 a_18451_43940# a_18579_44172# a_18533_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4395 a_13904_45546# a_13249_42308# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X4396 VSS a_13661_43548# a_18587_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4397 a_6547_43396# a_6031_43396# a_6452_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
C0 SMPL_ON_N VIN_N 0.587565f
C1 a_2487_47570# DATA[1] 7.79e-21
C2 a_n1853_43023# VDD 0.370563f
C3 a_20107_45572# a_21101_45002# 0.001705f
C4 a_9482_43914# a_13777_45326# 0.206086f
C5 a_10775_45002# a_1307_43914# 2.5e-21
C6 a_13348_45260# a_14180_45002# 5.21e-19
C7 a_7499_43078# a_9313_44734# 0.0624f
C8 a_9049_44484# a_9241_44734# 0.001498f
C9 a_13017_45260# a_14797_45144# 1.84e-19
C10 a_13159_45002# a_14537_43396# 3.64e-20
C11 a_n2109_45247# a_n2661_43370# 0.006863f
C12 a_7276_45260# a_1423_45028# 2.13e-20
C13 a_2274_45254# a_2448_45028# 5.85e-19
C14 a_4558_45348# a_5105_45348# 5.58e-20
C15 a_5147_45002# a_4640_45348# 5.32e-21
C16 a_20273_45572# a_21005_45260# 3.27e-19
C17 a_n4334_40480# a_n2442_46660# 3.24e-19
C18 a_10695_43548# a_n443_42852# 0.042055f
C19 a_133_43172# a_526_44458# 3.34e-20
C20 a_18341_45572# a_12549_44172# 2.55e-20
C21 a_17668_45572# a_n881_46662# 0.005485f
C22 a_413_45260# a_15811_47375# 2.19e-19
C23 a_6709_45028# a_6151_47436# 6.61e-22
C24 a_2232_45348# a_n971_45724# 2.25e-19
C25 a_n863_45724# a_n310_45572# 0.002342f
C26 a_n755_45592# a_509_45822# 2.51e-20
C27 a_n357_42282# a_n443_42852# 0.763015f
C28 a_16137_43396# a_15597_42852# 4.88e-19
C29 a_n13_43084# a_n2293_42282# 7.33e-21
C30 a_10796_42968# a_10341_42308# 0.65943f
C31 a_10991_42826# a_10922_42852# 0.209641f
C32 a_10835_43094# a_12379_42858# 0.001706f
C33 a_3626_43646# a_4921_42308# 0.431551f
C34 a_n97_42460# a_10533_42308# 0.001168f
C35 a_3080_42308# a_6123_31319# 1.45722f
C36 a_n1423_42826# a_n914_42852# 2.6e-19
C37 a_3539_42460# a_4933_42558# 6.41e-19
C38 a_12741_44636# RST_Z 0.004532f
C39 a_3726_37500# a_6886_37412# 0.702909f
C40 a_4338_37500# a_5700_37509# 2.69237f
C41 a_9293_42558# VDD 0.006879f
C42 a_2905_45572# a_n1151_42308# 0.072935f
C43 a_2063_45854# a_3815_47204# 5.54e-20
C44 a_1239_47204# a_n443_46116# 1.76e-21
C45 a_2553_47502# a_3785_47178# 7.79e-20
C46 a_n2833_47464# a_n1435_47204# 2.27e-20
C47 a_n1741_47186# a_9863_47436# 0.006846f
C48 a_n237_47217# a_6545_47178# 0.021104f
C49 a_n971_45724# a_6851_47204# 0.028789f
C50 a_16147_45260# a_15682_43940# 8.35e-19
C51 a_8696_44636# a_15493_43940# 1.53e-19
C52 a_n2661_44458# a_8103_44636# 0.006972f
C53 a_14537_43396# a_11967_42832# 7.01e-19
C54 a_11691_44458# a_16979_44734# 0.12231f
C55 a_11827_44484# a_18287_44626# 0.024541f
C56 a_11823_42460# a_13565_43940# 0.046344f
C57 a_n913_45002# a_895_43940# 3.46e-19
C58 a_n1059_45260# a_2675_43914# 1.32e-21
C59 a_n2017_45002# a_2889_44172# 1.5e-21
C60 a_n3674_37592# a_n2810_45572# 0.025877f
C61 a_6598_45938# VDD 0.204705f
C62 a_12607_44458# a_12891_46348# 0.067773f
C63 a_n2293_42834# a_7577_46660# 1.2e-20
C64 a_5343_44458# a_5807_45002# 4.88e-20
C65 a_n2661_44458# a_n2442_46660# 2.17e-20
C66 a_10057_43914# a_768_44030# 0.041949f
C67 a_13017_45260# a_14976_45028# 2.91e-20
C68 a_20731_45938# a_11415_45002# 0.001207f
C69 a_2711_45572# a_8062_46155# 1.41e-19
C70 a_413_45260# a_13059_46348# 1.63e-20
C71 a_13163_45724# a_10809_44734# 4.78e-21
C72 a_11136_45572# a_10903_43370# 0.002788f
C73 a_11682_45822# a_2324_44458# 1.62e-20
C74 a_n3674_39304# a_n4334_39616# 4.04e-19
C75 a_17701_42308# a_15959_42545# 1.03e-20
C76 a_5534_30871# a_13657_42308# 9.47e-19
C77 a_11599_46634# a_10428_46928# 0.001591f
C78 a_n1435_47204# a_6969_46634# 4e-20
C79 a_13717_47436# a_6755_46942# 9.51e-20
C80 a_6151_47436# a_10384_47026# 2.82e-20
C81 a_4915_47217# a_10768_47026# 4.45e-19
C82 a_6545_47178# a_8270_45546# 4.75e-21
C83 a_n1151_42308# a_12816_46660# 0.008712f
C84 a_4883_46098# a_5385_46902# 6e-21
C85 a_n881_46662# a_491_47026# 3.56e-21
C86 a_768_44030# a_n2438_43548# 6.89e-19
C87 a_20159_44458# a_20640_44752# 0.042415f
C88 a_11967_42832# a_20835_44721# 0.033569f
C89 a_19615_44636# a_20679_44626# 1.02e-20
C90 a_17517_44484# a_21398_44850# 0.01617f
C91 a_n2661_43922# a_175_44278# 0.003068f
C92 a_7640_43914# a_7542_44172# 0.20977f
C93 a_n2293_43922# a_n984_44318# 4.06e-20
C94 a_n2661_42834# a_644_44056# 0.005887f
C95 a_5891_43370# a_6453_43914# 3.53e-20
C96 a_10193_42453# a_18083_42858# 0.037244f
C97 a_n2293_42834# a_n1177_43370# 0.007412f
C98 a_11823_42460# a_5534_30871# 0.511874f
C99 a_1307_43914# a_3539_42460# 1.85e-19
C100 a_13249_42308# a_13113_42826# 0.008586f
C101 a_n356_44636# a_1241_44260# 7.4e-20
C102 en_comp a_12281_43396# 4.34e-21
C103 a_5111_44636# a_7221_43396# 9.51e-19
C104 a_2809_45028# VDD 0.189682f
C105 a_5932_42308# EN_VIN_BSTR_N 0.066129f
C106 a_6123_31319# a_n1532_35090# 1.38e-19
C107 a_4743_44484# a_4185_45028# 0.007252f
C108 a_5518_44484# a_3483_46348# 0.081879f
C109 a_11967_42832# a_3090_45724# 0.12811f
C110 a_14021_43940# a_768_44030# 1.82e-19
C111 a_7845_44172# a_4646_46812# 0.002985f
C112 a_9028_43914# a_2107_46812# 0.110155f
C113 a_14485_44260# a_12549_44172# 2.93e-20
C114 a_14537_43396# a_13259_45724# 0.083218f
C115 a_2382_45260# a_n755_45592# 5.27e-19
C116 a_1667_45002# a_1848_45724# 1.61e-19
C117 a_413_45260# a_3218_45724# 0.016434f
C118 a_n745_45366# a_n443_42852# 4.76e-19
C119 a_3232_43370# a_n2661_45546# 0.038743f
C120 a_11827_44484# a_15682_46116# 6.61e-22
C121 a_11691_44458# a_14275_46494# 1.05e-20
C122 a_19778_44110# a_19553_46090# 4.76e-20
C123 a_n2661_44458# a_8953_45546# 0.019448f
C124 a_n699_43396# a_4419_46090# 1.59e-20
C125 a_11599_46634# VDD 5.64965f
C126 a_17303_42282# a_17531_42308# 0.04615f
C127 a_5932_42308# a_1239_39043# 8.89e-20
C128 a_4958_30871# a_18057_42282# 4.22e-19
C129 a_n2661_46634# a_3483_46348# 0.051915f
C130 a_n2293_46634# a_2698_46116# 3.76e-20
C131 a_n1925_46634# a_2202_46116# 0.00159f
C132 a_n743_46660# a_1138_42852# 0.056829f
C133 a_n2438_43548# a_1176_45822# 0.073092f
C134 a_33_46660# a_472_46348# 0.003485f
C135 a_601_46902# a_376_46348# 8.72e-19
C136 a_n935_46688# a_n2293_46098# 2.46e-19
C137 a_6755_46942# a_14035_46660# 0.040006f
C138 a_12816_46660# a_14084_46812# 6.32e-20
C139 a_12891_46348# a_10903_43370# 0.132903f
C140 a_5807_45002# a_8349_46414# 2.69e-20
C141 a_n881_46662# a_14840_46494# 4.54e-19
C142 a_n1613_43370# a_2324_44458# 0.027159f
C143 a_13717_47436# a_8049_45260# 5.14e-20
C144 SMPL_ON_P a_n2472_45546# 3.24e-19
C145 a_n2497_47436# a_n452_45724# 5.75e-21
C146 a_13483_43940# a_14021_43940# 0.109097f
C147 a_14815_43914# a_14579_43548# 9.4e-21
C148 a_20365_43914# a_15493_43940# 0.048673f
C149 a_20935_43940# a_11341_43940# 0.006081f
C150 a_9313_44734# a_15781_43660# 0.00335f
C151 a_n2661_43922# a_10341_43396# 1.08e-19
C152 a_n2956_37592# a_n2472_42282# 8.96e-21
C153 a_19963_31679# a_n1630_35242# 1.23e-19
C154 a_n2017_45002# a_n4318_37592# 0.043579f
C155 a_n2810_45028# a_n4318_38216# 0.023084f
C156 en_comp a_n3674_38680# 0.014975f
C157 a_n2293_45010# a_n1329_42308# 1.37e-19
C158 a_n1899_43946# VDD 0.475205f
C159 a_10193_42453# a_11688_45572# 0.003765f
C160 a_10490_45724# a_11064_45572# 0.001758f
C161 a_8746_45002# a_11136_45572# 1.91e-20
C162 C0_P_btm VIN_P 0.529671f
C163 C10_N_btm C2_P_btm 3.9e-19
C164 a_9895_44260# a_3483_46348# 1.07e-19
C165 a_2075_43172# a_768_44030# 0.00187f
C166 a_2889_44172# a_526_44458# 2.55e-20
C167 a_n3674_39768# a_n2956_38680# 0.023133f
C168 a_11750_44172# a_10903_43370# 0.135933f
C169 a_8387_43230# a_n1613_43370# 0.163582f
C170 a_5164_46348# a_5497_46414# 0.203417f
C171 a_19636_46660# a_10809_44734# 3.84e-19
C172 a_n2293_46098# a_2324_44458# 0.018455f
C173 a_3483_46348# a_8199_44636# 1.81719f
C174 a_12741_44636# a_18985_46122# 1.17e-19
C175 a_11415_45002# a_20075_46420# 2.53e-20
C176 a_3090_45724# a_13259_45724# 0.261789f
C177 a_14035_46660# a_8049_45260# 0.002246f
C178 a_9028_43914# a_7871_42858# 5.97e-19
C179 a_6031_43396# a_6197_43396# 0.581047f
C180 a_18184_42460# a_17303_42282# 0.027385f
C181 a_14021_43940# a_13678_32519# 0.021333f
C182 a_11967_42832# a_12991_43230# 0.004319f
C183 a_2982_43646# a_2437_43396# 1.82e-20
C184 a_18494_42460# a_4958_30871# 5.63e-20
C185 a_584_46384# DATA[1] 0.007084f
C186 a_14358_43442# VDD 0.170277f
C187 a_11823_42460# a_11691_44458# 0.022559f
C188 a_6511_45714# a_5343_44458# 4.65e-21
C189 a_n467_45028# a_n143_45144# 0.007343f
C190 a_3357_43084# a_7229_43940# 6.23e-21
C191 a_n2017_45002# a_3537_45260# 0.033622f
C192 a_n913_45002# a_3065_45002# 0.225034f
C193 a_15803_42450# a_12549_44172# 1.19e-21
C194 a_1756_43548# a_n863_45724# 9.82e-20
C195 a_4905_42826# a_n2661_45546# 9.27e-20
C196 a_n229_43646# a_n357_42282# 0.00541f
C197 a_4361_42308# a_10903_43370# 0.00974f
C198 a_18997_42308# a_13507_46334# 6.67e-19
C199 a_3422_30871# a_11530_34132# 0.127528f
C200 a_1848_45724# VDD 0.100884f
C201 a_6472_45840# a_n2661_46634# 1.74e-20
C202 a_2711_45572# a_n1925_46634# 0.030736f
C203 a_10193_42453# a_12549_44172# 0.116594f
C204 a_10180_45724# a_768_44030# 7.51e-20
C205 a_10490_45724# a_11309_47204# 2.94e-20
C206 a_13163_45724# a_n881_46662# 2.21e-20
C207 a_3357_43084# a_n237_47217# 0.022871f
C208 a_n2109_45247# a_n2497_47436# 0.001006f
C209 a_2437_43646# a_327_47204# 2.63e-19
C210 a_16115_45572# a_10227_46804# 7.83e-19
C211 a_17478_45572# a_16327_47482# 0.012405f
C212 a_13259_45724# a_15002_46116# 4.39e-20
C213 a_13607_46688# RST_Z 3.83e-19
C214 a_14955_43940# a_15486_42560# 2.71e-19
C215 a_n2433_43396# a_n2104_42282# 1.29e-19
C216 a_8147_43396# a_8495_42852# 4.42e-20
C217 a_16409_43396# a_16795_42852# 0.010927f
C218 a_n2157_42858# a_n1736_43218# 0.089677f
C219 a_n1853_43023# a_n4318_38680# 0.003325f
C220 a_16137_43396# a_18083_42858# 0.005524f
C221 a_15682_43940# a_15051_42282# 2.71e-20
C222 a_3626_43646# a_13291_42460# 0.001564f
C223 a_n4318_39304# a_n3674_38216# 0.023484f
C224 a_n1641_43230# a_n1076_43230# 7.99e-20
C225 a_n1991_42858# a_n3674_39304# 0.002508f
C226 a_17538_32519# COMP_P 1.11e-20
C227 a_7754_39964# VDAC_Pi 0.001576f
C228 a_20273_45572# a_20835_44721# 2.82e-20
C229 a_11322_45546# a_10949_43914# 1.8e-20
C230 a_17023_45118# a_11827_44484# 3.5e-20
C231 a_19778_44110# a_18184_42460# 0.119002f
C232 a_10490_45724# a_10807_43548# 2.96e-21
C233 a_10193_42453# a_12429_44172# 9.75e-19
C234 a_2809_45028# a_n699_43396# 4.51e-19
C235 a_20623_45572# a_20640_44752# 3.53e-20
C236 a_n143_45144# a_n2661_43922# 2.71e-20
C237 a_n37_45144# a_n2661_42834# 3.28e-21
C238 a_6171_45002# a_5891_43370# 9.58e-20
C239 a_22591_45572# a_17517_44484# 3.95e-20
C240 a_3232_43370# a_8238_44734# 2.65e-20
C241 a_5205_44484# a_7640_43914# 2.61e-20
C242 a_n1736_42282# a_n1925_42282# 0.029727f
C243 a_1793_42852# a_n357_42282# 5.15e-19
C244 a_5934_30871# a_9290_44172# 4.13e-20
C245 a_8325_42308# a_8953_45546# 0.002755f
C246 a_8791_42308# a_8199_44636# 6.71e-19
C247 a_9803_42558# a_8016_46348# 1.11e-20
C248 a_17668_45572# a_17609_46634# 1.45e-20
C249 a_18799_45938# a_19466_46812# 2.72e-19
C250 a_7276_45260# a_4646_46812# 0.016809f
C251 a_413_45260# a_7577_46660# 3.89e-21
C252 a_5691_45260# a_5167_46660# 7.13e-20
C253 a_n1059_45260# a_6755_46942# 1.35e-20
C254 a_6194_45824# a_5937_45572# 0.002515f
C255 a_2711_45572# a_10355_46116# 3.59e-20
C256 a_6472_45840# a_8199_44636# 0.001875f
C257 a_7640_43914# a_n971_45724# 5.53e-20
C258 a_5024_45822# a_4419_46090# 8.88e-19
C259 a_5111_42852# a_5932_42308# 0.001025f
C260 a_5755_42852# a_6171_42473# 2.22e-19
C261 a_5649_42852# a_15486_42560# 5.1e-20
C262 a_4361_42308# a_15959_42545# 0.008092f
C263 a_20692_30879# a_18194_35068# 1.16e-19
C264 a_19237_31679# a_22469_40625# 1.24e-20
C265 a_13507_46334# a_768_44030# 0.019457f
C266 a_4883_46098# a_12891_46348# 0.085714f
C267 a_16327_47482# a_19594_46812# 0.004271f
C268 a_10227_46804# a_5807_45002# 0.262866f
C269 a_15673_47210# a_16750_47204# 1.46e-19
C270 a_9863_47436# a_n743_46660# 1.91e-20
C271 a_5815_47464# a_2107_46812# 8.74e-21
C272 a_n237_47217# a_3877_44458# 0.059355f
C273 a_n1741_47186# a_5907_46634# 8.63e-20
C274 a_n971_45724# a_4651_46660# 7.48e-19
C275 a_2952_47436# a_2959_46660# 5.17e-19
C276 a_3160_47472# a_2609_46660# 0.018687f
C277 a_n1151_42308# a_2443_46660# 3.77e-19
C278 a_2905_45572# a_3177_46902# 0.014554f
C279 a_584_46384# a_2864_46660# 2.26e-19
C280 a_n443_46116# a_491_47026# 1.47e-19
C281 a_n2661_43922# a_n2293_43922# 0.05908f
C282 a_n356_44636# a_11967_42832# 0.025796f
C283 a_18248_44752# a_18245_44484# 2.36e-20
C284 a_1307_43914# a_3353_43940# 0.005743f
C285 a_n467_45028# a_n97_42460# 5.34e-19
C286 a_n1059_45260# a_1209_43370# 8.19e-20
C287 a_2437_43646# a_3540_43646# 1.24e-19
C288 a_n2302_39072# a_n2810_45572# 2.61e-19
C289 en_comp VDD 4.26539f
C290 a_22400_42852# a_22821_38993# 0.136515f
C291 a_n2661_43370# a_167_45260# 0.055202f
C292 a_20567_45036# a_11415_45002# 0.011165f
C293 a_19778_44110# a_12741_44636# 0.070586f
C294 a_10903_45394# a_3483_46348# 0.002881f
C295 a_21005_45260# a_20202_43084# 1.88e-19
C296 a_16979_44734# a_15227_44166# 0.181002f
C297 a_18989_43940# a_3090_45724# 0.095784f
C298 a_5013_44260# a_768_44030# 0.064017f
C299 a_3537_45260# a_526_44458# 0.938783f
C300 a_15595_45028# a_15682_46116# 1.03e-20
C301 a_6517_45366# a_5937_45572# 2.26e-19
C302 a_n875_44318# a_n1613_43370# 7.2e-19
C303 a_8953_45002# a_10809_44734# 0.001885f
C304 a_20935_43940# a_16327_47482# 0.004638f
C305 a_10949_43914# a_12465_44636# 3.08e-19
C306 COMP_P a_22465_38105# 0.059345f
C307 a_10545_42558# a_10723_42308# 5.98e-20
C308 a_n3674_38216# a_n4334_40480# 8.37e-20
C309 a_n1630_35242# a_7174_31319# 0.035143f
C310 a_5534_30871# C0_dummy_P_btm 2.22e-20
C311 a_5342_30871# C1_P_btm 9.04e-20
C312 a_18194_35068# VIN_N 0.066301f
C313 a_n1435_47204# a_9625_46129# 2.1e-20
C314 a_6151_47436# a_13925_46122# 5.38e-19
C315 a_4791_45118# a_2324_44458# 0.19212f
C316 a_n2312_39304# a_n2157_46122# 0.00402f
C317 a_1799_45572# a_3090_45724# 1.03e-19
C318 a_8145_46902# a_8492_46660# 0.051162f
C319 a_16131_47204# a_765_45546# 0.005958f
C320 a_5807_45002# a_17339_46660# 0.02927f
C321 a_10440_44484# a_8685_43396# 2.31e-20
C322 a_n2661_43922# a_n97_42460# 6.42e-20
C323 a_n2661_42834# a_104_43370# 0.001459f
C324 a_11691_44458# a_18429_43548# 1.12e-20
C325 a_11827_44484# a_19268_43646# 1.65e-20
C326 a_n2293_42834# a_n1991_42858# 0.02898f
C327 a_7499_43078# a_8515_42308# 1.55e-19
C328 a_2711_45572# a_14113_42308# 5.51e-20
C329 a_n913_45002# a_2987_42968# 1.92e-21
C330 a_413_45260# a_22959_42860# 7.98e-20
C331 a_10617_44484# VDD 0.141193f
C332 a_n4209_38216# C7_P_btm 1.43e-20
C333 a_n3565_38216# C9_P_btm 1.91e-20
C334 a_2711_45572# a_7499_43078# 0.007939f
C335 a_6511_45714# a_4880_45572# 8.15e-21
C336 a_6472_45840# a_6428_45938# 1.46e-19
C337 CAL_N a_n357_42282# 0.001017f
C338 a_3905_42865# a_1823_45246# 0.218008f
C339 a_19478_44306# a_17339_46660# 9.54e-21
C340 a_12281_43396# a_13661_43548# 1.07e-19
C341 a_16137_43396# a_12549_44172# 0.003438f
C342 a_5745_43940# a_3090_45724# 0.003797f
C343 a_2779_44458# a_3218_45724# 3.4e-20
C344 a_n2661_44458# a_1609_45822# 2.15e-19
C345 a_5343_44458# a_n755_45592# 0.349527f
C346 a_n356_44636# a_13259_45724# 0.026337f
C347 a_11967_42832# a_20075_46420# 1.89e-21
C348 a_19615_44636# a_19335_46494# 2.3e-20
C349 a_13678_32519# a_13507_46334# 0.037522f
C350 a_4361_42308# a_4883_46098# 9.17e-20
C351 a_20749_43396# a_18479_47436# 4.66e-19
C352 en_comp a_22469_39537# 0.001226f
C353 a_7411_46660# VDD 0.41059f
C354 a_n4334_38528# a_n4334_38304# 0.052468f
C355 a_n3565_38502# a_n4209_38216# 5.84657f
C356 a_n4209_38502# a_n3565_38216# 0.028468f
C357 a_n2302_38778# a_n2216_38778# 0.011479f
C358 a_n3690_38528# a_n3607_38528# 0.007692f
C359 a_n3420_38528# a_n4251_38528# 0.001487f
C360 a_4958_30871# C10_N_btm 6.95e-19
C361 a_20820_30879# a_12741_44636# 0.103478f
C362 a_22591_46660# a_22959_46660# 7.52e-19
C363 a_11415_45002# a_21076_30879# 8.27e-21
C364 a_20202_43084# a_21297_46660# 4.61e-21
C365 a_765_45546# a_3483_46348# 1.15e-19
C366 a_n2293_46634# a_380_45546# 6.42e-19
C367 a_n1925_46634# a_n1079_45724# 4.37e-19
C368 a_n2438_43548# a_n2472_45546# 0.008798f
C369 a_n1021_46688# a_n2293_45546# 2.36e-21
C370 a_n133_46660# a_n2661_45546# 1.33e-20
C371 a_7715_46873# a_8062_46482# 9.21e-19
C372 a_n2661_46634# a_n357_42282# 3.78e-20
C373 a_11735_46660# a_6945_45028# 1.07e-19
C374 a_3090_45724# a_18189_46348# 0.029136f
C375 a_n4318_37592# a_n3690_37440# 1.65e-19
C376 a_n1761_44111# a_n1736_43218# 3.37e-20
C377 a_n809_44244# a_n1076_43230# 1.8e-20
C378 a_n984_44318# a_n901_43156# 2.43e-19
C379 a_20935_43940# a_10341_43396# 1.76e-20
C380 a_n1352_43396# a_104_43370# 4.33e-20
C381 a_11341_43940# a_14955_43396# 1.96e-20
C382 a_11967_42832# a_12379_42858# 0.492977f
C383 a_5891_43370# a_8292_43218# 0.003655f
C384 a_n1917_43396# a_n1809_43762# 0.057222f
C385 a_n1699_43638# a_n1190_43762# 2.6e-19
C386 a_n2267_43396# a_n1821_43396# 2.28e-19
C387 a_n447_43370# a_n97_42460# 0.00228f
C388 a_n2129_43609# a_n1655_43396# 0.002164f
C389 a_15493_43940# a_14205_43396# 2.04e-19
C390 a_1307_43914# a_16104_42674# 4.76e-21
C391 a_19721_31679# COMP_P 2.4e-20
C392 a_n2956_37592# a_n2216_39866# 1.2e-19
C393 a_n1699_43638# VDD 0.210236f
C394 a_20623_45572# a_21188_45572# 7.99e-20
C395 a_20273_45572# a_20731_45938# 0.034619f
C396 a_7227_45028# a_n2293_42834# 3.08e-20
C397 a_8192_45572# a_8191_45002# 0.001292f
C398 a_12281_43396# a_4185_45028# 1.62e-19
C399 a_10518_42984# a_3090_45724# 0.004978f
C400 a_22400_42852# a_21588_30879# 2.09e-19
C401 a_1049_43396# a_526_44458# 0.121121f
C402 a_8791_43396# a_2324_44458# 3.85e-21
C403 a_9145_43396# a_8953_45546# 0.019849f
C404 a_10053_45546# a_9863_47436# 3.03e-20
C405 a_9159_45572# a_n237_47217# 3.1e-20
C406 a_17715_44484# a_18051_46116# 9.64e-19
C407 a_18985_46122# a_16375_45002# 9.94e-20
C408 a_8199_44636# a_n357_42282# 0.023438f
C409 a_18819_46122# a_19240_46482# 0.089677f
C410 a_5066_45546# a_5210_46155# 0.001301f
C411 a_167_45260# a_2307_45899# 0.005265f
C412 a_104_43370# a_n2293_42282# 6.62e-21
C413 a_16243_43396# a_4361_42308# 7.3e-20
C414 a_17499_43370# a_743_42282# 8.79e-20
C415 a_8791_43396# a_8387_43230# 5.36e-19
C416 a_n2661_42282# a_2123_42473# 8.86e-20
C417 a_18783_43370# a_19177_43646# 2.23e-19
C418 a_18429_43548# a_4190_30871# 0.001307f
C419 a_11967_42832# a_18727_42674# 1.83e-20
C420 a_2982_43646# a_5534_30871# 0.094381f
C421 a_2107_46812# CLK 3e-20
C422 a_22165_42308# VDD 0.336187f
C423 a_16019_45002# a_16922_45042# 7.45e-20
C424 a_3175_45822# a_2998_44172# 1.76e-21
C425 a_8696_44636# a_13468_44734# 0.001421f
C426 a_n143_45144# a_n452_44636# 6.31e-21
C427 a_3065_45002# a_n2661_44458# 0.027917f
C428 a_n1059_45260# a_8103_44636# 8.03e-23
C429 a_12379_42858# a_13259_45724# 0.001312f
C430 a_4649_43172# a_526_44458# 0.005678f
C431 a_421_43172# a_n863_45724# 0.00331f
C432 a_15599_45572# a_6755_46942# 0.024601f
C433 a_6472_45840# a_765_45546# 1.39e-20
C434 a_15143_45578# a_3090_45724# 0.016572f
C435 a_11823_42460# a_15227_44166# 1.79e-19
C436 a_9159_45572# a_8270_45546# 8.13e-20
C437 a_13249_42308# a_15368_46634# 4.76e-21
C438 a_2437_43646# a_1983_46706# 0.01301f
C439 a_n2017_45002# a_n2293_46634# 0.039556f
C440 a_n2810_45028# a_n2956_39768# 0.04304f
C441 a_3232_43370# a_12891_46348# 8.12e-21
C442 a_4927_45028# a_768_44030# 4.62e-21
C443 en_comp a_22612_30879# 5.56e-19
C444 a_6171_45002# a_11309_47204# 3.85e-20
C445 a_n2840_42826# a_n4318_38216# 0.012711f
C446 a_n2472_42826# a_n2472_42282# 0.025171f
C447 a_10835_43094# a_12800_43218# 2.33e-21
C448 a_743_42282# a_1576_42282# 0.007548f
C449 a_2982_43646# a_19647_42308# 0.002685f
C450 a_10922_42852# a_11301_43218# 3.16e-19
C451 a_10991_42826# a_11554_42852# 0.049827f
C452 a_10796_42968# a_10752_42852# 1.46e-19
C453 a_3626_43646# a_18548_42308# 0.001059f
C454 a_n2157_42858# a_n3674_38680# 2.17e-19
C455 a_18819_46122# START 8.36e-19
C456 a_18985_46122# RST_Z 1.22e-21
C457 a_n2216_40160# VDD 0.00515f
C458 a_n237_47217# a_8128_46384# 0.113499f
C459 a_1209_47178# a_n881_46662# 4.08e-21
C460 a_1239_47204# a_n1613_43370# 0.001663f
C461 a_11599_46634# a_16588_47582# 2.07e-20
C462 a_15507_47210# a_16763_47508# 0.043475f
C463 a_7903_47542# a_4883_46098# 3.03e-21
C464 a_14311_47204# a_10227_46804# 2.11e-19
C465 a_15673_47210# a_16327_47482# 0.206019f
C466 a_15811_47375# a_16023_47582# 0.003622f
C467 a_3785_47178# a_2747_46873# 4.9e-20
C468 a_n1151_42308# a_7_47243# 1.92e-19
C469 a_13717_47436# a_18780_47178# 1.64e-19
C470 a_12861_44030# a_18479_47436# 0.065796f
C471 a_18184_42460# a_20159_44458# 0.01449f
C472 a_20567_45036# a_11967_42832# 2.76e-20
C473 a_742_44458# a_n2661_43922# 0.066714f
C474 a_949_44458# a_n2661_42834# 0.009741f
C475 a_4743_44484# a_5708_44484# 1.11e-19
C476 a_9838_44484# a_9313_44734# 0.037628f
C477 a_19778_44110# a_20362_44736# 1.01e-19
C478 a_11691_44458# a_15367_44484# 0.005161f
C479 a_5343_44458# a_5608_44484# 0.004449f
C480 a_7499_43078# a_7466_43396# 1.63e-19
C481 a_2711_45572# a_15781_43660# 1.33e-19
C482 a_11827_44484# a_17061_44484# 0.001186f
C483 a_n2293_42834# a_n1331_43914# 4.35e-19
C484 a_3232_43370# a_11750_44172# 0.020452f
C485 a_6171_45002# a_10807_43548# 3.25e-20
C486 a_n913_45002# a_10555_44260# 3.18e-21
C487 a_8685_42308# a_n443_42852# 6.23e-22
C488 a_13070_42354# a_n357_42282# 1.72e-20
C489 a_18727_42674# a_13259_45724# 8.73e-20
C490 a_n2860_39072# a_n2956_39304# 0.001353f
C491 a_16855_45546# VDD 0.339227f
C492 a_20820_30879# C9_N_btm 3.29e-19
C493 a_9482_43914# a_12741_44636# 0.101234f
C494 a_14180_45002# a_11415_45002# 0.025987f
C495 a_2382_45260# a_3483_46348# 1.72e-21
C496 a_2680_45002# a_3147_46376# 3.68e-20
C497 a_18315_45260# a_3090_45724# 0.061731f
C498 a_4743_44484# a_5257_43370# 7.16e-21
C499 a_5147_45002# a_1823_45246# 0.001658f
C500 a_13296_44484# a_768_44030# 0.001019f
C501 a_15599_45572# a_8049_45260# 0.003996f
C502 a_3733_45822# a_3503_45724# 0.004937f
C503 a_11778_45572# a_10586_45546# 0.006085f
C504 a_3260_45572# a_2957_45546# 0.001377f
C505 a_20273_45572# a_20075_46420# 1.19e-20
C506 a_20107_45572# a_19900_46494# 1.7e-19
C507 a_3357_43084# a_13759_46122# 1.98e-20
C508 a_n1059_45260# a_8953_45546# 0.318691f
C509 a_196_42282# a_6123_31319# 1.36e-20
C510 a_2713_42308# a_2903_42308# 0.23738f
C511 a_n784_42308# a_7227_42308# 3.86e-20
C512 a_15597_42852# a_15764_42576# 9.51e-19
C513 a_13291_42460# a_13921_42308# 2.04e-19
C514 a_n1630_35242# a_5932_42308# 0.033914f
C515 a_4190_30871# C0_dummy_P_btm 1.45e-20
C516 a_22521_40055# a_22521_39511# 0.457858f
C517 a_5807_45002# a_10467_46802# 0.007388f
C518 a_n1925_46634# a_6540_46812# 0.008209f
C519 a_2443_46660# a_3177_46902# 0.053479f
C520 a_2107_46812# a_3055_46660# 0.001203f
C521 a_8128_46384# a_8270_45546# 0.002121f
C522 a_11453_44696# a_19333_46634# 0.026664f
C523 a_16327_47482# a_16388_46812# 0.01513f
C524 a_15811_47375# a_16751_46987# 1.26e-19
C525 a_12861_44030# a_17829_46910# 0.058114f
C526 a_13487_47204# a_765_45546# 0.006318f
C527 a_13717_47436# a_18285_46348# 1.31e-20
C528 a_n2497_47436# a_167_45260# 0.001788f
C529 a_n746_45260# a_n901_46420# 8.55e-20
C530 a_n971_45724# a_n1076_46494# 8.23e-19
C531 a_n2109_47186# a_1823_45246# 7.36e-20
C532 a_1239_47204# a_n2293_46098# 5.76e-21
C533 a_n1741_47186# a_1176_45822# 1.11e-19
C534 a_15433_44458# a_15493_43396# 1.53e-19
C535 a_n809_44244# a_175_44278# 0.001854f
C536 a_n2065_43946# a_453_43940# 2.55e-21
C537 a_n452_44636# a_n97_42460# 4e-21
C538 a_11823_42460# a_14635_42282# 0.087526f
C539 a_n2661_42834# a_11341_43940# 0.007026f
C540 a_14539_43914# a_13565_43940# 4.14e-20
C541 a_n699_43396# a_n1699_43638# 1.54e-20
C542 a_5111_44636# a_5649_42852# 0.121004f
C543 en_comp a_n4318_38680# 0.007648f
C544 a_n2017_45002# a_n1533_42852# 0.004733f
C545 a_n913_45002# a_n967_43230# 8.68e-20
C546 a_n467_45028# a_n901_43156# 4.74e-20
C547 a_3357_43084# a_5755_42852# 8.48e-20
C548 a_n2216_37690# VDD 0.003946f
C549 a_n1699_44726# VDD 0.198612f
C550 a_17303_42282# RST_Z 0.002907f
C551 a_22465_38105# a_22705_37990# 1.35e-19
C552 a_7174_31319# a_11530_34132# 0.001307f
C553 a_15433_44458# a_3483_46348# 4.08e-20
C554 a_20159_44458# a_12741_44636# 0.006194f
C555 a_20679_44626# a_11415_45002# 0.007381f
C556 a_9672_43914# a_8270_45546# 0.003127f
C557 a_4699_43561# a_768_44030# 4.91e-20
C558 a_18326_43940# a_6755_46942# 1.01e-19
C559 a_n2661_43370# a_n863_45724# 0.076347f
C560 a_17719_45144# a_18051_46116# 1.04e-20
C561 a_5891_43370# a_10903_43370# 1.39e-19
C562 a_13667_43396# a_10227_46804# 0.007746f
C563 a_n4334_39616# a_n4064_39616# 0.4504f
C564 a_n3690_39616# a_n3420_39616# 0.431154f
C565 a_n3565_39590# a_n2946_39866# 0.406088f
C566 a_n4209_39590# a_n2302_39866# 0.406459f
C567 a_13661_43548# VDD 3.93017f
C568 SMPL_ON_N a_20205_31679# 0.029367f
C569 a_12861_44030# a_n443_42852# 0.015171f
C570 a_5894_47026# a_5937_45572# 5.36e-21
C571 a_7411_46660# a_7920_46348# 0.004089f
C572 a_n1925_46634# a_1337_46436# 3.83e-19
C573 a_768_44030# a_10586_45546# 3.88e-20
C574 a_n743_46660# a_739_46482# 0.005906f
C575 a_n2442_46660# a_n1925_42282# 8.58e-20
C576 a_n2293_46634# a_526_44458# 0.579444f
C577 a_5807_45002# a_8034_45724# 1.95e-20
C578 a_18834_46812# a_18900_46660# 0.006978f
C579 a_16388_46812# a_16434_46987# 0.006879f
C580 a_15227_44166# a_18280_46660# 0.007923f
C581 a_14513_46634# a_765_45546# 5.52e-20
C582 a_10623_46897# a_3483_46348# 6.27e-20
C583 a_5111_44636# a_7963_42308# 5.33e-19
C584 a_n913_45002# a_13575_42558# 3.5e-19
C585 a_n1059_45260# a_14456_42282# 7.72e-20
C586 en_comp a_11551_42558# 4.34e-21
C587 a_n2017_45002# a_13249_42558# 0.001525f
C588 a_14539_43914# a_5534_30871# 1.4e-20
C589 a_18579_44172# a_18783_43370# 1.04e-19
C590 a_19279_43940# a_19700_43370# 8.74e-21
C591 a_n2661_42834# a_n1076_43230# 5.44e-20
C592 a_n2661_43922# a_n901_43156# 9.27e-21
C593 a_n2293_43922# a_n1641_43230# 9.84e-21
C594 a_n356_44636# a_10518_42984# 1.13e-20
C595 a_15004_44636# a_5342_30871# 5.64e-20
C596 a_19862_44208# VDD 0.588967f
C597 a_4099_45572# a_3537_45260# 5.2e-19
C598 a_2711_45572# a_4558_45348# 0.001943f
C599 a_4093_43548# a_1823_45246# 0.17443f
C600 a_3539_42460# a_n2293_46098# 4.77e-19
C601 a_743_42282# a_8270_45546# 9.44e-21
C602 a_n809_44244# a_n356_45724# 3.24e-21
C603 a_2998_44172# a_n863_45724# 2.34e-19
C604 a_453_43940# a_n755_45592# 0.003942f
C605 a_2127_44172# a_n357_42282# 0.00145f
C606 a_9061_43230# a_n1613_43370# 2.95e-19
C607 a_7754_39964# RST_Z 0.843939f
C608 a_19326_42852# a_16327_47482# 2.94e-19
C609 a_1606_42308# a_4791_45118# 3.68e-20
C610 a_3754_38470# a_n923_35174# 0.002509f
C611 a_4185_45028# VDD 1.65665f
C612 a_n3565_39304# a_n4209_37414# 0.028483f
C613 a_n4209_39304# a_n3565_37414# 0.030571f
C614 a_n3565_38216# a_n3607_38304# 0.001003f
C615 C7_N_btm C10_N_btm 1.39624f
C616 C8_N_btm C9_N_btm 39.4538f
C617 a_765_45546# a_n357_42282# 0.209746f
C618 a_5497_46414# a_5066_45546# 0.05403f
C619 a_5068_46348# a_5210_46155# 0.005572f
C620 a_18819_46122# a_19553_46090# 0.052547f
C621 a_2324_44458# a_6945_45028# 0.183081f
C622 a_15015_46420# a_10809_44734# 6.69e-20
C623 a_n1352_43396# a_n1076_43230# 9.05e-19
C624 a_n447_43370# a_n901_43156# 0.008716f
C625 a_4905_42826# a_4361_42308# 0.005834f
C626 a_14955_43396# a_10341_43396# 0.01411f
C627 a_2982_43646# a_4190_30871# 0.3223f
C628 a_n1809_43762# a_n1853_43023# 4.91e-20
C629 a_14021_43940# a_18083_42858# 1.31e-20
C630 a_9803_43646# a_9885_43396# 0.003935f
C631 a_n97_42460# a_n1641_43230# 3.57e-21
C632 a_n356_44636# a_16197_42308# 1.9e-19
C633 a_n2472_43914# a_n4318_38216# 4.52e-19
C634 a_8685_43396# a_13837_43396# 6.31e-19
C635 a_n1917_43396# a_n3674_39304# 1.1e-19
C636 a_n1699_43638# a_n4318_38680# 1.98e-19
C637 a_11453_44696# CLK 8.57e-19
C638 a_22959_47212# EN_OFFSET_CAL 0.007205f
C639 a_2266_47570# DATA[1] 1.59e-20
C640 a_n2157_42858# VDD 0.424058f
C641 a_n2293_45010# a_n2661_43370# 0.067876f
C642 a_5205_44484# a_1423_45028# 0.821456f
C643 a_8953_45002# a_1307_43914# 1.41e-19
C644 a_n967_45348# a_n2293_42834# 0.038042f
C645 a_4558_45348# a_4640_45348# 0.007001f
C646 a_20273_45572# a_20567_45036# 0.005333f
C647 a_20107_45572# a_21005_45260# 2.5e-19
C648 a_9482_43914# a_13556_45296# 0.726155f
C649 a_8746_45002# a_5891_43370# 1.89e-19
C650 a_13017_45260# a_14537_43396# 0.003458f
C651 a_n2302_40160# a_n2956_39768# 3.63e-19
C652 a_n4315_30879# a_n2442_46660# 0.361271f
C653 a_9803_43646# a_n443_42852# 0.102893f
C654 a_18479_45785# a_12549_44172# 0.105486f
C655 a_17568_45572# a_n881_46662# 0.001221f
C656 a_19479_31679# SMPL_ON_N 0.029207f
C657 a_2437_43646# a_22959_47212# 4.39e-19
C658 a_20447_31679# a_4883_46098# 0.003751f
C659 a_413_45260# a_15507_47210# 3.64e-19
C660 a_n2017_45002# a_18597_46090# 2.49e-21
C661 a_1423_45028# a_n971_45724# 0.021147f
C662 a_13348_45260# a_n1151_42308# 3.18e-22
C663 a_310_45028# a_n443_42852# 0.376934f
C664 a_n357_42282# a_509_45822# 0.039776f
C665 a_10796_42968# a_10922_42852# 0.170059f
C666 a_10835_43094# a_10341_42308# 0.541777f
C667 a_n1076_43230# a_n2293_42282# 3.1e-20
C668 a_14021_43940# a_22775_42308# 1.94e-20
C669 a_n1991_42858# a_n914_42852# 1.46e-19
C670 a_n1853_43023# a_133_42852# 0.001685f
C671 a_5649_42852# a_5837_43172# 1.5e-19
C672 a_3539_42460# a_3905_42558# 0.015463f
C673 a_4905_42826# a_6761_42308# 3.95e-20
C674 a_4338_37500# a_5088_37509# 0.896828f
C675 a_3726_37500# a_5700_37509# 0.574743f
C676 a_20820_30879# RST_Z 0.048737f
C677 a_9803_42558# VDD 0.253745f
C678 a_2905_45572# a_3160_47472# 0.54473f
C679 a_2952_47436# a_n1151_42308# 0.068429f
C680 a_2063_45854# a_3785_47178# 0.001458f
C681 a_n1741_47186# a_9067_47204# 0.012401f
C682 a_n237_47217# a_6151_47436# 0.360224f
C683 a_n971_45724# a_6491_46660# 0.011282f
C684 a_11691_44458# a_14539_43914# 0.268287f
C685 a_n2661_44458# a_6298_44484# 0.025865f
C686 a_11827_44484# a_18248_44752# 0.00953f
C687 a_n2661_43370# a_9313_44734# 3.03e-20
C688 a_1307_43914# a_16335_44484# 8.63e-20
C689 a_15861_45028# a_11341_43940# 3.78e-20
C690 a_n2017_45002# a_2675_43914# 5.66e-22
C691 a_n913_45002# a_2479_44172# 0.003813f
C692 a_n1059_45260# a_895_43940# 2.25e-19
C693 a_6667_45809# VDD 0.195842f
C694 a_10440_44484# a_768_44030# 0.002332f
C695 a_n4318_40392# a_n2442_46660# 0.023735f
C696 a_13017_45260# a_3090_45724# 2.74e-21
C697 a_8975_43940# a_12891_46348# 6.34e-21
C698 a_20623_45572# a_12741_44636# 5.76e-19
C699 a_20731_45938# a_20202_43084# 4.22e-19
C700 a_20528_45572# a_11415_45002# 0.002765f
C701 a_6511_45714# a_8034_45724# 0.001344f
C702 a_12791_45546# a_10809_44734# 3.56e-21
C703 a_5891_43370# a_4883_46098# 0.003161f
C704 a_17701_42308# a_15803_42450# 2.65e-20
C705 a_n3674_39304# a_n4209_39590# 4.47e-20
C706 a_22400_42852# a_22765_42852# 9.38e-19
C707 a_5534_30871# a_11897_42308# 4.24e-20
C708 a_4883_46098# a_4817_46660# 1.29e-19
C709 a_11599_46634# a_10150_46912# 3.38e-21
C710 a_6151_47436# a_8270_45546# 0.142873f
C711 a_n1435_47204# a_6755_46942# 0.006483f
C712 a_6575_47204# a_8035_47026# 3.94e-19
C713 a_2063_45854# a_3090_45724# 0.002495f
C714 a_n1151_42308# a_12991_46634# 0.013856f
C715 a_n1613_43370# a_491_47026# 0.038998f
C716 a_n881_46662# a_288_46660# 0.001197f
C717 a_19594_46812# a_20843_47204# 5.41e-20
C718 a_768_44030# a_n743_46660# 0.028134f
C719 a_8953_45002# a_9396_43370# 6.95e-20
C720 a_5111_44636# a_8685_43396# 0.078598f
C721 a_3537_45260# a_8317_43396# 7.25e-21
C722 a_20159_44458# a_20362_44736# 0.233657f
C723 a_11967_42832# a_20679_44626# 0.863531f
C724 a_n2661_43922# a_n984_44318# 0.004148f
C725 a_n2661_42834# a_175_44278# 0.010875f
C726 a_8975_43940# a_11750_44172# 1.78e-19
C727 a_5891_43370# a_5663_43940# 1.27e-19
C728 a_13249_42308# a_12545_42858# 0.030353f
C729 a_n2293_42834# a_n1917_43396# 0.006976f
C730 a_1307_43914# a_3626_43646# 0.012223f
C731 a_10193_42453# a_17701_42308# 5.98e-19
C732 a_11823_42460# a_14543_43071# 0.028488f
C733 a_17517_44484# a_20980_44850# 0.026284f
C734 a_7640_43914# a_7281_43914# 0.003713f
C735 a_n2293_43922# a_n809_44244# 4.38e-21
C736 a_6109_44484# a_7542_44172# 2.12e-20
C737 a_2448_45028# VDD 0.004293f
C738 a_5932_42308# a_11530_34132# 0.001408f
C739 a_n2946_37984# a_n2956_38680# 0.004795f
C740 a_n699_43396# a_4185_45028# 0.027874f
C741 a_5343_44458# a_3483_46348# 0.046505f
C742 a_17517_44484# a_19692_46634# 0.023737f
C743 a_11341_43940# a_19321_45002# 0.009893f
C744 a_15493_43940# a_13747_46662# 0.049242f
C745 a_14021_43940# a_12549_44172# 0.150377f
C746 a_7542_44172# a_4646_46812# 0.012612f
C747 a_19006_44850# a_3090_45724# 0.001921f
C748 a_14180_45002# a_13259_45724# 0.04353f
C749 a_413_45260# a_2957_45546# 0.012841f
C750 a_2274_45254# a_n755_45592# 1.63e-19
C751 a_n913_45002# a_n443_42852# 0.796158f
C752 a_2382_45260# a_n357_42282# 0.025504f
C753 a_11827_44484# a_2324_44458# 0.03555f
C754 a_19778_44110# a_18985_46122# 3.49e-19
C755 a_n2661_44458# a_5937_45572# 0.061693f
C756 a_3539_42460# a_4791_45118# 6.9e-19
C757 a_4223_44672# a_4419_46090# 1.94e-20
C758 a_14955_47212# VDD 0.301751f
C759 a_4958_30871# a_17531_42308# 0.192941f
C760 a_5742_30871# a_n4209_39590# 1.2e-21
C761 a_5934_30871# a_n3565_39304# 5.05e-21
C762 a_5342_30871# a_n3420_37984# 0.028488f
C763 a_5534_30871# a_n4064_37984# 0.047233f
C764 a_171_46873# a_472_46348# 0.008963f
C765 a_n2661_46634# a_3147_46376# 8.89e-20
C766 a_n1925_46634# a_1823_45246# 0.001679f
C767 a_n743_46660# a_1176_45822# 0.08607f
C768 a_n2438_43548# a_1208_46090# 0.005695f
C769 a_n133_46660# a_805_46414# 0.001959f
C770 a_33_46660# a_376_46348# 5.66e-19
C771 a_22612_30879# a_4185_45028# 2.99e-19
C772 a_6755_46942# a_13885_46660# 0.078788f
C773 a_12816_46660# a_13607_46688# 3.63e-19
C774 a_5807_45002# a_8016_46348# 3.22e-19
C775 a_12891_46348# a_11387_46155# 1.97e-20
C776 a_11309_47204# a_10903_43370# 1.95e-19
C777 a_n881_46662# a_15015_46420# 2.18e-20
C778 SMPL_ON_P a_n2661_45546# 0.002242f
C779 a_n2497_47436# a_n863_45724# 0.337007f
C780 a_n2109_47186# a_n2293_45546# 4.56e-21
C781 a_n452_44636# a_n901_43156# 6.5e-20
C782 a_18287_44626# a_16823_43084# 9.2e-20
C783 a_n1899_43946# a_n1809_43762# 8.11e-19
C784 a_n809_44244# a_n97_42460# 3.09e-19
C785 a_20269_44172# a_15493_43940# 0.051355f
C786 a_20935_43940# a_21115_43940# 0.185422f
C787 a_20623_43914# a_11341_43940# 0.007271f
C788 a_9313_44734# a_15681_43442# 0.001424f
C789 a_13483_43940# a_13829_44260# 0.013377f
C790 a_14539_43914# a_4190_30871# 8.06e-21
C791 a_10193_42453# a_21613_42308# 1.95e-19
C792 a_n2661_42834# a_10341_43396# 2.59e-19
C793 a_n2017_45002# a_n1736_42282# 0.017988f
C794 a_n2810_45028# a_n2472_42282# 9.69e-21
C795 a_n2956_37592# a_n3674_38680# 0.02294f
C796 en_comp a_n2840_42282# 0.001493f
C797 a_n1761_44111# VDD 0.620042f
C798 a_10490_45724# a_10544_45572# 0.004398f
C799 a_8746_45002# a_11064_45572# 9.37e-21
C800 a_2711_45572# a_16377_45572# 4.3e-19
C801 C1_P_btm VIN_P 0.39234f
C802 C10_N_btm C3_P_btm 0.001117f
C803 C9_N_btm C2_P_btm 2.13e-19
C804 a_22959_43948# a_4185_45028# 0.014665f
C805 a_9801_44260# a_3483_46348# 0.002837f
C806 a_1847_42826# a_768_44030# 4.92e-19
C807 a_2982_43646# a_15227_44166# 8.62e-20
C808 a_556_44484# a_n443_42852# 4.78e-20
C809 a_n2661_43922# a_3503_45724# 5.64e-21
C810 a_2675_43914# a_526_44458# 0.03283f
C811 a_n3674_39768# a_n2956_39304# 0.02324f
C812 a_n4318_39768# a_n2956_38680# 0.023254f
C813 a_22959_44484# a_8049_45260# 5.34e-19
C814 a_10807_43548# a_10903_43370# 0.193971f
C815 a_8605_42826# a_n1613_43370# 0.159791f
C816 a_19164_43230# a_18597_46090# 2.45e-21
C817 a_20922_43172# a_18479_47436# 9.43e-20
C818 a_18083_42858# a_13507_46334# 1.81e-19
C819 a_14543_46987# VDD 8.63e-19
C820 a_5164_46348# a_5204_45822# 0.132894f
C821 a_18900_46660# a_10809_44734# 8.2e-19
C822 a_21350_47026# a_6945_45028# 1.62e-19
C823 a_3483_46348# a_8349_46414# 4.04e-20
C824 a_12741_44636# a_18819_46122# 2.26e-20
C825 a_11415_45002# a_19335_46494# 3.95e-20
C826 a_14976_45028# a_15194_46482# 5.51e-19
C827 a_13885_46660# a_8049_45260# 5.7e-22
C828 a_15009_46634# a_13259_45724# 9.93e-20
C829 a_8333_44056# a_7871_42858# 5.27e-20
C830 a_6031_43396# a_6293_42852# 0.163953f
C831 a_3626_43646# a_9396_43370# 2.73e-20
C832 a_n97_42460# a_14955_43396# 2e-20
C833 a_14021_43940# a_21855_43396# 0.025748f
C834 a_11967_42832# a_12800_43218# 0.025258f
C835 a_5343_44458# a_8791_42308# 3.69e-19
C836 a_18184_42460# a_4958_30871# 0.004748f
C837 a_584_46384# DATA[0] 3.21e-20
C838 a_2124_47436# DATA[1] 0.00138f
C839 a_14579_43548# VDD 0.278225f
C840 a_12427_45724# a_11691_44458# 3.08e-21
C841 a_n1059_45260# a_3065_45002# 0.023485f
C842 a_n967_45348# a_413_45260# 9.61e-20
C843 a_791_42968# a_1138_42852# 0.100783f
C844 a_15764_42576# a_12549_44172# 7.49e-20
C845 a_10793_43218# a_3090_45724# 9.54e-20
C846 a_1568_43370# a_n863_45724# 0.202455f
C847 a_3080_42308# a_n2661_45546# 0.155045f
C848 a_5649_42852# a_9290_44172# 3.77e-19
C849 a_13258_32519# SMPL_ON_N 0.030848f
C850 a_22775_42308# a_13507_46334# 0.022177f
C851 a_997_45618# VDD 0.12359f
C852 a_6194_45824# a_n2661_46634# 1.76e-20
C853 a_10193_42453# a_12891_46348# 1.13e-20
C854 a_n2293_45010# a_n2497_47436# 0.233882f
C855 a_16333_45814# a_10227_46804# 3.14e-19
C856 a_15861_45028# a_16327_47482# 0.030602f
C857 a_526_44458# a_2277_45546# 5.37e-21
C858 a_14955_43940# a_15051_42282# 1.74e-20
C859 a_15682_43940# a_14113_42308# 2.3e-19
C860 a_n2157_42858# a_n4318_38680# 9.64e-19
C861 a_n1853_43023# a_n3674_39304# 1.5e-19
C862 a_16409_43396# a_16414_43172# 4.62e-21
C863 a_743_42282# a_5755_42852# 2.61e-20
C864 a_16137_43396# a_17701_42308# 0.025497f
C865 a_2982_43646# a_14635_42282# 3.39e-19
C866 a_n1423_42826# a_n1076_43230# 0.051162f
C867 a_16547_43609# a_16795_42852# 0.081093f
C868 a_n2433_43396# a_n4318_38216# 0.002497f
C869 a_10384_47026# CLK 9.6e-20
C870 a_3357_43084# a_17517_44484# 0.001645f
C871 a_n143_45144# a_n2661_42834# 2.16e-21
C872 a_n467_45028# a_n2661_43922# 0.024697f
C873 a_6171_45002# a_8375_44464# 4.23e-20
C874 a_3232_43370# a_5891_43370# 0.137859f
C875 a_2382_45260# a_3363_44484# 9.62e-20
C876 a_5205_44484# a_6109_44484# 0.029986f
C877 a_20273_45572# a_20679_44626# 3.84e-19
C878 a_10193_42453# a_11750_44172# 0.01114f
C879 a_11322_45546# a_10729_43914# 3.04e-19
C880 a_20107_45572# a_20835_44721# 6.77e-20
C881 a_16922_45042# a_11827_44484# 0.032223f
C882 a_11551_42558# a_4185_45028# 8.71e-20
C883 a_n3674_38216# a_n1925_42282# 0.004354f
C884 a_1709_42852# a_n357_42282# 5.74e-19
C885 a_8685_42308# a_8199_44636# 0.114007f
C886 a_8337_42558# a_8953_45546# 1.56e-19
C887 a_4880_45572# a_3483_46348# 4.49e-19
C888 a_19256_45572# a_19692_46634# 2.88e-19
C889 a_626_44172# a_1123_46634# 7.29e-21
C890 a_18596_45572# a_19466_46812# 7.53e-21
C891 a_13490_45394# a_768_44030# 1.56e-19
C892 a_413_45260# a_7715_46873# 5.62e-20
C893 a_3537_45260# a_5275_47026# 7.68e-22
C894 a_5205_44484# a_4646_46812# 0.094488f
C895 a_5691_45260# a_5385_46902# 3.11e-22
C896 a_5147_45002# a_5732_46660# 5.29e-20
C897 a_n2017_45002# a_6755_46942# 1.28e-20
C898 a_5907_45546# a_5937_45572# 0.104991f
C899 a_2711_45572# a_9823_46155# 5.98e-20
C900 a_6598_45938# a_6419_46155# 1.5e-19
C901 a_11691_44458# a_11453_44696# 0.035893f
C902 a_n2012_44484# a_n1151_42308# 9.03e-20
C903 a_5755_42852# a_5755_42308# 3.59e-19
C904 a_5649_42852# a_15051_42282# 3.72e-19
C905 a_16823_43084# a_17124_42282# 6.14e-21
C906 a_4361_42308# a_15803_42450# 0.055869f
C907 a_11301_43218# a_11554_42852# 4.61e-19
C908 a_20205_31679# a_18194_35068# 1.48e-19
C909 a_20692_30879# EN_VIN_BSTR_N 2.04e-19
C910 a_19237_31679# a_22521_40599# 1.41e-20
C911 a_13507_46334# a_12549_44172# 0.363125f
C912 a_4883_46098# a_11309_47204# 0.012799f
C913 a_16327_47482# a_19321_45002# 0.925259f
C914 a_17591_47464# a_5807_45002# 0.001206f
C915 a_12861_44030# a_n2661_46634# 0.03828f
C916 a_n1741_47186# a_5167_46660# 2.91e-20
C917 a_n971_45724# a_4646_46812# 0.303249f
C918 a_2063_45854# a_3699_46634# 7.49e-20
C919 a_2952_47436# a_3177_46902# 1.43e-19
C920 a_n1151_42308# a_n2661_46098# 0.024549f
C921 a_3160_47472# a_2443_46660# 0.019074f
C922 a_2905_45572# a_2609_46660# 0.027251f
C923 a_n2109_47186# a_5732_46660# 0.009505f
C924 a_584_46384# a_3524_46660# 4.24e-20
C925 a_18287_44626# a_19279_43940# 4.65e-20
C926 a_18989_43940# a_20679_44626# 4.34e-21
C927 a_n2661_42834# a_n2293_43922# 0.034793f
C928 a_n699_43396# a_n1761_44111# 0.018554f
C929 a_10193_42453# a_4361_42308# 0.274131f
C930 a_17970_44736# a_18245_44484# 0.007416f
C931 a_1307_43914# a_3052_44056# 0.001611f
C932 a_n2661_44458# a_2479_44172# 1.07e-19
C933 a_15861_45028# a_10341_43396# 2.08e-20
C934 a_n467_45028# a_n447_43370# 6.82e-20
C935 a_n1059_45260# a_458_43396# 3e-19
C936 a_n2017_45002# a_1209_43370# 4.18e-21
C937 a_2437_43646# a_2982_43646# 0.0016f
C938 a_n2956_37592# VDD 1.25966f
C939 a_14097_32519# a_22521_39511# 7.51e-21
C940 a_22400_42852# a_22545_38993# 0.038805f
C941 a_8560_45348# a_3483_46348# 0.021507f
C942 a_18494_42460# a_11415_45002# 0.006745f
C943 a_18911_45144# a_12741_44636# 0.013476f
C944 a_14539_43914# a_15227_44166# 0.520312f
C945 a_18374_44850# a_3090_45724# 3.45e-19
C946 a_5244_44056# a_768_44030# 0.167173f
C947 a_3429_45260# a_526_44458# 0.010386f
C948 a_3065_45002# a_n1925_42282# 0.04956f
C949 a_15595_45028# a_2324_44458# 0.04743f
C950 a_n1287_44306# a_n1613_43370# 0.003155f
C951 a_15493_43396# a_10227_46804# 0.003705f
C952 a_20623_43914# a_16327_47482# 0.009946f
C953 a_10807_43548# a_4883_46098# 2.5e-20
C954 a_564_42282# a_7174_31319# 9.76e-21
C955 a_n4318_38216# a_n4064_40160# 0.052465f
C956 a_10545_42558# a_10533_42308# 0.011812f
C957 a_5534_30871# C0_P_btm 8.49e-20
C958 EN_VIN_BSTR_N VIN_N 1.41696f
C959 EN_VIN_BSTR_P VCM 0.929333f
C960 a_4190_30871# a_n4064_37984# 0.032018f
C961 a_10227_46804# a_3483_46348# 0.057984f
C962 a_9313_45822# a_9823_46155# 6.69e-21
C963 a_6151_47436# a_13759_46122# 3.56e-19
C964 a_4915_47217# a_14275_46494# 0.01257f
C965 a_n1435_47204# a_8953_45546# 5.89e-20
C966 a_n2312_39304# a_n2293_46098# 0.027561f
C967 a_5807_45002# a_15312_46660# 3.46e-19
C968 a_13747_46662# a_14226_46660# 0.001089f
C969 a_3877_44458# a_8189_46660# 9.93e-21
C970 a_6540_46812# a_6999_46987# 6.64e-19
C971 a_5907_46634# a_6086_46660# 0.007399f
C972 a_5732_46660# a_5841_46660# 0.007416f
C973 a_7577_46660# a_8492_46660# 0.118423f
C974 a_n913_45002# a_1793_42852# 0.00284f
C975 a_n967_45348# a_n914_42852# 1.98e-19
C976 a_10334_44484# a_8685_43396# 1.89e-20
C977 a_n2661_42834# a_n97_42460# 9.39e-19
C978 a_11691_44458# a_17324_43396# 1.34e-21
C979 a_11827_44484# a_15743_43084# 3.38e-21
C980 a_n2293_42834# a_n1853_43023# 0.053782f
C981 a_9482_43914# a_10991_42826# 8.72e-21
C982 a_1307_43914# a_8037_42858# 2.06e-21
C983 a_7499_43078# a_5934_30871# 0.00463f
C984 a_5708_44484# VDD 9.68e-19
C985 a_n3565_38216# C10_P_btm 2.25e-20
C986 a_n4209_38216# C8_P_btm 1.65e-20
C987 a_2711_45572# a_8568_45546# 0.011004f
C988 a_6194_45824# a_6428_45938# 0.006453f
C989 a_3600_43914# a_1823_45246# 0.016141f
C990 a_11341_43940# a_13059_46348# 0.025185f
C991 a_10341_43396# a_19321_45002# 1.67e-19
C992 a_15493_43396# a_17339_46660# 0.075223f
C993 a_12293_43646# a_13661_43548# 8.56e-20
C994 a_5326_44056# a_3090_45724# 2.02e-19
C995 a_8317_43396# a_n2293_46634# 3.08e-19
C996 a_2779_44458# a_2957_45546# 6.96e-19
C997 a_n2661_44458# a_n443_42852# 0.045408f
C998 a_5343_44458# a_n357_42282# 0.022768f
C999 a_11967_42832# a_19335_46494# 4.62e-21
C1000 a_21855_43396# a_13507_46334# 0.003121f
C1001 a_8605_42826# a_4791_45118# 1.13e-21
C1002 en_comp a_22821_38993# 1.42e-19
C1003 a_19479_31679# a_18194_35068# 8.48e-20
C1004 a_5257_43370# VDD 0.922495f
C1005 a_n4209_38502# a_n4334_38304# 3.3e-19
C1006 a_n4334_38528# a_n4209_38216# 3.3e-19
C1007 a_n3565_38502# a_n3607_38528# 0.001003f
C1008 a_n4064_38528# a_n2216_38778# 0.005567f
C1009 a_4958_30871# C9_N_btm 0.209166f
C1010 a_22591_46660# a_12741_44636# 0.0686f
C1011 a_11415_45002# a_22959_46660# 3.29e-19
C1012 a_20202_43084# a_21076_30879# 6.04e-20
C1013 a_765_45546# a_3147_46376# 2.61e-20
C1014 a_17339_46660# a_3483_46348# 7.08e-22
C1015 a_n2293_46634# a_n452_45724# 0.002803f
C1016 a_n2661_46634# a_310_45028# 4.45e-20
C1017 a_8667_46634# a_5066_45546# 4.03e-20
C1018 a_n2438_43548# a_n2661_45546# 0.065227f
C1019 a_n1925_46634# a_n2293_45546# 7.25e-20
C1020 a_3090_45724# a_17715_44484# 0.108364f
C1021 a_12156_46660# a_10903_43370# 8.13e-19
C1022 a_15559_46634# a_2324_44458# 0.012623f
C1023 a_n4318_37592# a_n3565_37414# 4.06e-19
C1024 a_n809_44244# a_n901_43156# 0.001977f
C1025 a_n1549_44318# a_n1076_43230# 2.38e-20
C1026 a_15682_43940# a_15781_43660# 0.005099f
C1027 a_20623_43914# a_10341_43396# 7.45e-20
C1028 a_n1699_43638# a_n1809_43762# 0.097745f
C1029 a_11341_43940# a_15095_43370# 4.91e-20
C1030 a_n2293_43922# a_n2293_42282# 0.19201f
C1031 a_n4318_40392# a_n3674_38216# 0.023361f
C1032 a_n1917_43396# a_n2012_43396# 0.049827f
C1033 a_n2267_43396# a_n1190_43762# 1.46e-19
C1034 a_3905_42865# a_5649_42852# 3.85e-20
C1035 a_n2129_43609# a_n1821_43396# 0.004509f
C1036 a_5891_43370# a_7573_43172# 5.51e-21
C1037 a_11967_42832# a_10341_42308# 0.001434f
C1038 a_14539_43914# a_14635_42282# 1.26e-19
C1039 a_18114_32519# COMP_P 1.46e-20
C1040 en_comp a_n2302_39866# 4.43e-20
C1041 a_n2956_37592# a_n2860_39866# 3.22e-20
C1042 a_n2267_43396# VDD 0.570924f
C1043 a_20107_45572# a_20731_45938# 9.73e-19
C1044 a_20841_45814# a_21188_45572# 0.051162f
C1045 a_20273_45572# a_20528_45572# 0.064178f
C1046 a_14495_45572# a_14537_43396# 2.49e-19
C1047 a_10907_45822# a_10951_45334# 0.002454f
C1048 a_2711_45572# a_n2661_43370# 0.112998f
C1049 a_10083_42826# a_3090_45724# 0.005497f
C1050 a_1209_43370# a_526_44458# 0.057216f
C1051 a_13070_42354# a_12861_44030# 2.94e-20
C1052 a_9803_43646# a_8199_44636# 0.009804f
C1053 a_8685_43396# a_9290_44172# 0.207262f
C1054 a_1337_46116# VDD 0.20087f
C1055 a_11823_42460# a_4915_47217# 0.016758f
C1056 a_8568_45546# a_9313_45822# 0.002981f
C1057 a_11652_45724# a_6151_47436# 9.87e-21
C1058 a_17583_46090# a_18051_46116# 3.98e-20
C1059 a_18819_46122# a_16375_45002# 0.002016f
C1060 a_167_45260# a_1990_45899# 0.006879f
C1061 a_n97_42460# a_n2293_42282# 5.22e-19
C1062 a_8147_43396# a_8387_43230# 1.33e-19
C1063 a_16759_43396# a_743_42282# 1.02e-20
C1064 a_3626_43646# a_13635_43156# 1.89e-19
C1065 a_2982_43646# a_14543_43071# 2.24e-21
C1066 a_16137_43396# a_4361_42308# 0.019831f
C1067 a_11967_42832# a_18057_42282# 0.002498f
C1068 a_n2661_42282# a_1755_42282# 0.145244f
C1069 a_3422_30871# a_15890_42674# 2.49e-20
C1070 a_16664_43396# a_16855_43396# 4.61e-19
C1071 a_17324_43396# a_4190_30871# 2.14e-20
C1072 a_21671_42860# VDD 0.229963f
C1073 a_n913_45002# CAL_N 0.002966f
C1074 en_comp VDAC_N 7.58e-19
C1075 a_15595_45028# a_16922_45042# 1.97e-20
C1076 a_2711_45572# a_2998_44172# 1.79e-21
C1077 a_16019_45002# a_16501_45348# 2.93e-19
C1078 a_8696_44636# a_13213_44734# 0.004648f
C1079 a_4640_45348# a_n2661_43370# 4.5e-19
C1080 a_2680_45002# a_n2661_44458# 7.59e-20
C1081 a_n467_45028# a_n452_44636# 0.092885f
C1082 a_n1059_45260# a_6298_44484# 2.2e-22
C1083 a_133_43172# a_n863_45724# 7.15e-19
C1084 a_n3420_37440# w_1575_34946# 2.64e-19
C1085 a_6194_45824# a_765_45546# 9.06e-22
C1086 a_13904_45546# a_15368_46634# 8.27e-21
C1087 a_8791_45572# a_8270_45546# 9.56e-20
C1088 a_413_45260# a_13747_46662# 3.67e-20
C1089 a_2437_43646# a_2107_46812# 0.185914f
C1090 a_n2109_45247# a_n2293_46634# 0.016559f
C1091 a_n913_45002# a_n2661_46634# 8.11e-21
C1092 a_5111_44636# a_768_44030# 0.154519f
C1093 a_n2017_45002# a_n2442_46660# 1.18e-21
C1094 en_comp a_21588_30879# 4.44e-19
C1095 a_3232_43370# a_11309_47204# 9.11e-20
C1096 a_n2661_43370# a_9313_45822# 8.9e-20
C1097 a_8191_45002# a_n881_46662# 2.82e-21
C1098 a_8685_43396# a_15051_42282# 7.21e-19
C1099 a_10796_42968# a_11554_42852# 0.056391f
C1100 a_743_42282# a_1067_42314# 0.010185f
C1101 a_2982_43646# a_19511_42282# 0.014171f
C1102 a_10991_42826# a_11301_43218# 0.013793f
C1103 a_10922_42852# a_11229_43218# 3.69e-19
C1104 a_n2472_42826# a_n3674_38680# 0.004228f
C1105 a_4361_42308# a_n784_42308# 2.34e-20
C1106 a_9145_43396# a_13575_42558# 4.11e-19
C1107 a_13887_32519# COMP_P 6.33e-21
C1108 a_3626_43646# a_18310_42308# 0.00142f
C1109 a_13925_46122# CLK 1.2e-20
C1110 a_18819_46122# RST_Z 7.83e-21
C1111 a_n4251_40480# VDD 3.95e-19
C1112 a_n1741_47186# a_12549_44172# 9.64e-19
C1113 a_n971_45724# a_9804_47204# 1.23e-20
C1114 a_327_47204# a_n881_46662# 3.68e-20
C1115 a_1209_47178# a_n1613_43370# 0.006245f
C1116 a_15673_47210# a_16241_47178# 0.183195f
C1117 a_15507_47210# a_16023_47582# 0.109156f
C1118 a_11599_46634# a_16763_47508# 4.36e-20
C1119 a_15811_47375# a_16327_47482# 0.038827f
C1120 a_3381_47502# a_2747_46873# 2.58e-20
C1121 a_2063_45854# a_2583_47243# 2.21e-19
C1122 a_n1151_42308# a_n310_47243# 3.07e-19
C1123 a_13717_47436# a_18479_47436# 2.23e-19
C1124 a_13487_47204# a_10227_46804# 2.54e-19
C1125 a_12861_44030# a_18143_47464# 0.394543f
C1126 a_6171_45002# a_10949_43914# 9.46e-21
C1127 a_3232_43370# a_10807_43548# 0.001324f
C1128 a_2437_43646# a_2253_43940# 0.003306f
C1129 a_18494_42460# a_11967_42832# 0.025796f
C1130 a_n452_44636# a_n2661_43922# 0.009547f
C1131 a_5883_43914# a_9313_44734# 0.124999f
C1132 a_8975_43940# a_5891_43370# 0.021307f
C1133 a_742_44458# a_n2661_42834# 0.034578f
C1134 a_19778_44110# a_20159_44458# 2.12e-20
C1135 a_n2293_42834# a_n1899_43946# 0.001698f
C1136 a_n2012_44484# a_n1821_44484# 4.61e-19
C1137 a_7499_43078# a_7221_43396# 4.61e-20
C1138 a_1423_45028# a_7281_43914# 0.001025f
C1139 a_18479_45785# a_19478_44056# 3.95e-19
C1140 a_11827_44484# a_16789_44484# 2.76e-19
C1141 a_12563_42308# a_n357_42282# 9.02e-20
C1142 a_18057_42282# a_13259_45724# 4.22e-19
C1143 a_8325_42308# a_n443_42852# 0.001008f
C1144 a_16115_45572# VDD 0.194492f
C1145 a_20820_30879# C8_N_btm 9.97e-19
C1146 a_21076_30879# C5_N_btm 1.31e-19
C1147 a_5342_30871# EN_VIN_BSTR_N 0.010795f
C1148 a_13348_45260# a_12741_44636# 5.41e-21
C1149 a_13777_45326# a_11415_45002# 0.021087f
C1150 a_4558_45348# a_1823_45246# 1.95e-19
C1151 a_2382_45260# a_3147_46376# 1.77e-20
C1152 a_2680_45002# a_2804_46116# 1.03e-20
C1153 a_17719_45144# a_3090_45724# 0.001738f
C1154 a_14309_45028# a_15227_44166# 8.19e-20
C1155 a_13857_44734# a_13661_43548# 0.012574f
C1156 a_12829_44484# a_768_44030# 3.4e-20
C1157 a_3638_45822# a_3503_45724# 0.008535f
C1158 a_11688_45572# a_10586_45546# 7.93e-19
C1159 a_15297_45822# a_8049_45260# 1.34e-19
C1160 a_20107_45572# a_20075_46420# 0.001614f
C1161 a_3357_43084# a_13351_46090# 3.73e-21
C1162 a_n913_45002# a_8199_44636# 0.018004f
C1163 a_n1059_45260# a_5937_45572# 2.49e-20
C1164 a_n2017_45002# a_8953_45546# 0.080521f
C1165 a_413_45260# a_4419_46090# 7.46e-21
C1166 a_564_42282# a_5932_42308# 8.68e-21
C1167 a_n784_42308# a_6761_42308# 2.26e-20
C1168 a_2725_42558# a_2903_42308# 5.98e-20
C1169 a_13291_42460# a_13657_42308# 0.001043f
C1170 a_4190_30871# C0_P_btm 6.53e-20
C1171 a_22521_40055# a_22780_40081# 0.010228f
C1172 a_5807_45002# a_10428_46928# 0.002901f
C1173 a_n1925_46634# a_5732_46660# 0.006885f
C1174 a_n743_46660# a_5167_46660# 2.34e-20
C1175 a_1799_45572# a_2959_46660# 3.87e-20
C1176 a_2443_46660# a_2609_46660# 0.579196f
C1177 a_1983_46706# a_2162_46660# 0.006978f
C1178 a_n2661_46634# a_5894_47026# 1.44e-19
C1179 a_8128_46384# a_8189_46660# 6.01e-19
C1180 a_11453_44696# a_15227_44166# 0.979188f
C1181 a_3080_42308# a_3754_38470# 3.23e-19
C1182 a_10227_46804# a_14513_46634# 0.004612f
C1183 a_16241_47178# a_16388_46812# 1.22e-19
C1184 a_15673_47210# a_16721_46634# 2.97e-19
C1185 a_15811_47375# a_16434_46987# 8.78e-19
C1186 a_16327_47482# a_13059_46348# 5.25e-20
C1187 a_12861_44030# a_765_45546# 0.190301f
C1188 a_n2109_47186# a_1138_42852# 1.13e-20
C1189 a_n971_45724# a_n901_46420# 0.021388f
C1190 a_n1151_42308# a_11415_45002# 2.84e-20
C1191 a_n785_47204# a_n1853_46287# 2.37e-20
C1192 a_n452_44636# a_n447_43370# 0.001136f
C1193 a_15004_44636# a_15037_43940# 1.72e-20
C1194 a_n809_44244# a_n984_44318# 0.234322f
C1195 a_11823_42460# a_13291_42460# 0.257506f
C1196 a_n699_43396# a_n2267_43396# 1.05e-19
C1197 a_n2661_45010# a_685_42968# 5.86e-22
C1198 a_3357_43084# a_5111_42852# 5.76e-19
C1199 a_n2956_37592# a_n4318_38680# 0.023187f
C1200 en_comp a_n3674_39304# 3.39e-19
C1201 a_5147_45002# a_5649_42852# 2.35e-21
C1202 a_n2860_37690# VDD 0.004184f
C1203 a_n2267_44484# VDD 0.289888f
C1204 a_4958_30871# RST_Z 0.087554f
C1205 a_22465_38105# a_22609_37990# 3.5e-19
C1206 a_19615_44636# a_12741_44636# 0.001298f
C1207 a_20640_44752# a_11415_45002# 0.0058f
C1208 a_20679_44626# a_20202_43084# 0.035147f
C1209 a_14815_43914# a_3483_46348# 0.036548f
C1210 a_9028_43914# a_8270_45546# 0.233359f
C1211 a_18079_43940# a_6755_46942# 2.17e-19
C1212 a_n2661_43370# a_n1079_45724# 2.43e-20
C1213 a_8103_44636# a_526_44458# 3.01e-21
C1214 a_18494_42460# a_13259_45724# 1.69e-19
C1215 a_14209_32519# w_11334_34010# 7.84e-19
C1216 a_10695_43548# a_10227_46804# 2.31e-19
C1217 a_3626_43646# a_n1613_43370# 1.21e-19
C1218 a_n356_44636# a_17715_44484# 1.89e-21
C1219 a_n2661_43922# a_5164_46348# 8.9e-20
C1220 a_n4209_39590# a_n4064_39616# 0.269818f
C1221 a_n3565_39590# a_n3420_39616# 0.281955f
C1222 a_5807_45002# VDD 1.75047f
C1223 a_10227_46804# a_n357_42282# 0.103631f
C1224 a_11309_47204# a_11608_46482# 6.71e-19
C1225 a_n1925_46634# a_n914_46116# 5.09e-20
C1226 a_12549_44172# a_10586_45546# 0.003919f
C1227 a_n743_46660# a_518_46482# 7.72e-19
C1228 a_14180_46812# a_765_45546# 4.49e-21
C1229 a_16388_46812# a_16721_46634# 0.222024f
C1230 a_19692_46634# a_20731_47026# 9.71e-20
C1231 a_10467_46802# a_3483_46348# 9.89e-19
C1232 a_14539_43914# a_14543_43071# 8.67e-19
C1233 a_18579_44172# a_18525_43370# 0.012789f
C1234 a_742_44458# a_n2293_42282# 0.006579f
C1235 a_19279_43940# a_19268_43646# 5.83e-21
C1236 a_n2661_42834# a_n901_43156# 0.001144f
C1237 a_n2293_43922# a_n1423_42826# 1.71e-20
C1238 a_n356_44636# a_10083_42826# 4.56e-20
C1239 a_375_42282# a_1184_42692# 1.26e-19
C1240 a_5111_44636# a_6123_31319# 1.17e-19
C1241 a_n913_45002# a_13070_42354# 4.84e-20
C1242 a_n1059_45260# a_13575_42558# 8.82e-21
C1243 a_n2017_45002# a_14456_42282# 0.003727f
C1244 en_comp a_5742_30871# 0.092238f
C1245 a_19478_44306# VDD 0.127794f
C1246 a_2711_45572# a_4574_45260# 8.29e-19
C1247 a_1756_43548# a_1823_45246# 5.06e-21
C1248 a_10341_43396# a_13059_46348# 0.014853f
C1249 a_17324_43396# a_15227_44166# 0.010717f
C1250 a_16664_43396# a_3090_45724# 1.05e-21
C1251 a_453_43940# a_n357_42282# 0.027908f
C1252 a_2889_44172# a_n863_45724# 4.42e-22
C1253 a_1414_42308# a_n755_45592# 0.013035f
C1254 a_5013_44260# a_n2661_45546# 1.73e-19
C1255 a_8649_43218# a_n1613_43370# 0.001903f
C1256 a_n3420_37984# VIN_P 0.06991f
C1257 a_n39_42308# a_n1151_42308# 9.43e-20
C1258 a_19721_31679# a_22609_37990# 7.56e-21
C1259 a_3699_46348# VDD 0.208984f
C1260 C6_N_btm C10_N_btm 0.895671f
C1261 C7_N_btm C9_N_btm 0.22201f
C1262 a_n4209_39304# a_n4334_37440# 4.61e-19
C1263 a_1736_39043# a_3754_38802# 7.66e-20
C1264 a_3483_46348# a_8034_45724# 1.49e-19
C1265 a_765_45546# a_310_45028# 0.012232f
C1266 a_17339_46660# a_n357_42282# 1.31e-19
C1267 a_5204_45822# a_5066_45546# 0.402457f
C1268 a_8953_45546# a_526_44458# 0.037032f
C1269 a_18819_46122# a_18985_46122# 0.749955f
C1270 a_14275_46494# a_10809_44734# 6.38e-20
C1271 a_18189_46348# a_19335_46494# 1.11e-21
C1272 a_n2840_43914# a_n4318_38216# 8.56e-19
C1273 a_n1177_43370# a_n1076_43230# 9.51e-21
C1274 a_15095_43370# a_10341_43396# 0.013375f
C1275 a_3080_42308# a_4361_42308# 8.53e-19
C1276 a_2982_43646# a_21259_43561# 0.034927f
C1277 a_n1809_43762# a_n2157_42858# 2.44e-20
C1278 a_n1352_43396# a_n901_43156# 1.07e-20
C1279 a_9801_43940# a_9127_43156# 5.84e-20
C1280 a_14021_43940# a_17701_42308# 9.5e-20
C1281 a_n2661_42834# a_10533_42308# 4.35e-22
C1282 a_13667_43396# a_12281_43396# 1.88e-20
C1283 a_n97_42460# a_n1423_42826# 6.33e-21
C1284 a_8685_43396# a_13749_43396# 6.06e-19
C1285 a_n1699_43638# a_n3674_39304# 2.54e-19
C1286 a_n2267_43396# a_n4318_38680# 3e-19
C1287 a_11453_44696# EN_OFFSET_CAL 7.26e-19
C1288 a_n2472_42826# VDD 0.229608f
C1289 a_10193_42453# a_5891_43370# 0.001973f
C1290 a_20107_45572# a_20567_45036# 9.82e-19
C1291 a_13348_45260# a_13556_45296# 0.189446f
C1292 a_13017_45260# a_14180_45002# 0.079928f
C1293 a_13159_45002# a_13777_45326# 8.25e-20
C1294 a_18799_45938# a_11691_44458# 7.04e-20
C1295 a_n2472_45002# a_n2661_43370# 0.017331f
C1296 a_6431_45366# a_1423_45028# 1.36e-20
C1297 en_comp a_n2293_42834# 0.103485f
C1298 a_4574_45260# a_4640_45348# 0.006978f
C1299 a_413_45260# a_2809_45028# 0.005798f
C1300 a_4558_45348# a_4185_45348# 1.34e-19
C1301 a_3537_45260# a_5105_45348# 3.16e-19
C1302 a_20273_45572# a_18494_42460# 0.002243f
C1303 a_n4064_40160# a_n2956_39768# 0.002282f
C1304 a_9145_43396# a_n443_42852# 2.32123f
C1305 a_18175_45572# a_12549_44172# 1.35e-20
C1306 a_5024_45822# a_5257_43370# 1.25e-19
C1307 a_2437_43646# a_11453_44696# 0.189184f
C1308 a_413_45260# a_11599_46634# 3.55e-19
C1309 a_5205_44484# a_6545_47178# 1.89e-20
C1310 a_626_44172# a_n746_45260# 0.011647f
C1311 a_n2661_45546# a_603_45572# 8.65e-19
C1312 a_3316_45546# a_3503_45724# 0.024901f
C1313 a_n1099_45572# a_n443_42852# 0.026572f
C1314 a_310_45028# a_509_45822# 0.039722f
C1315 a_n901_43156# a_n2293_42282# 7.23e-20
C1316 a_10796_42968# a_10991_42826# 0.206455f
C1317 a_10518_42984# a_10341_42308# 0.00245f
C1318 a_10835_43094# a_10922_42852# 0.053385f
C1319 a_2982_43646# a_4921_42308# 0.001781f
C1320 a_n97_42460# a_9885_42558# 0.011255f
C1321 a_3539_42460# a_3581_42558# 0.002471f
C1322 a_5649_42852# a_5457_43172# 1.97e-19
C1323 a_3626_43646# a_3905_42558# 0.004928f
C1324 a_4905_42826# a_6773_42558# 8.37e-21
C1325 a_20202_43084# SINGLE_ENDED 1.07e-19
C1326 a_22591_46660# RST_Z 4.25e-19
C1327 a_3726_37500# a_5088_37509# 0.189392f
C1328 a_9223_42460# VDD 0.205797f
C1329 a_327_47204# a_n443_46116# 1.72e-19
C1330 a_2553_47502# a_n1151_42308# 0.007448f
C1331 a_2952_47436# a_3160_47472# 0.192116f
C1332 a_2063_45854# a_3381_47502# 1.06e-19
C1333 a_584_46384# a_3785_47178# 1.58e-20
C1334 a_n1741_47186# a_6575_47204# 0.075265f
C1335 a_n971_45724# a_6545_47178# 0.295443f
C1336 a_16855_45546# a_15493_43940# 1.91e-22
C1337 a_8696_44636# a_11341_43940# 1.44e-19
C1338 a_n2661_44458# a_5518_44484# 0.01193f
C1339 a_11827_44484# a_17970_44736# 0.012326f
C1340 a_11691_44458# a_16112_44458# 0.012386f
C1341 a_18494_42460# a_18989_43940# 1.47e-20
C1342 a_10193_42453# a_18533_43940# 0.007041f
C1343 a_1307_43914# a_16241_44484# 0.001942f
C1344 a_n467_45028# a_n809_44244# 0.010788f
C1345 a_n1059_45260# a_2479_44172# 0.004979f
C1346 a_n2017_45002# a_895_43940# 2.49e-20
C1347 a_n1630_35242# a_20692_30879# 2.27e-19
C1348 a_6511_45714# VDD 0.405279f
C1349 a_21188_45572# a_11415_45002# 0.009324f
C1350 a_10334_44484# a_768_44030# 0.001784f
C1351 a_7639_45394# a_7715_46873# 2.05e-20
C1352 a_6472_45840# a_8034_45724# 1.02e-19
C1353 a_8975_43940# a_11309_47204# 4.06e-22
C1354 a_3357_43084# a_20731_47026# 0.00277f
C1355 a_17730_32519# w_11334_34010# 0.027505f
C1356 a_15433_44458# a_12861_44030# 0.002244f
C1357 a_10907_45822# a_2324_44458# 0.025622f
C1358 a_11136_45572# a_11133_46155# 5.62e-20
C1359 a_11823_42460# a_10809_44734# 0.215753f
C1360 a_13163_45724# a_6945_45028# 3.09e-21
C1361 a_22400_42852# a_20753_42852# 6.01e-21
C1362 a_17701_42308# a_15764_42576# 1.32e-20
C1363 a_4883_46098# a_4955_46873# 0.09516f
C1364 a_11599_46634# a_9863_46634# 3.12e-21
C1365 a_n1435_47204# a_10249_46116# 7.87e-20
C1366 a_7903_47542# a_8035_47026# 9.4e-20
C1367 a_13381_47204# a_6755_46942# 9.89e-20
C1368 a_6151_47436# a_8189_46660# 0.001903f
C1369 a_n1151_42308# a_12251_46660# 0.00985f
C1370 a_584_46384# a_3090_45724# 0.001068f
C1371 a_2747_46873# a_2959_46660# 0.010672f
C1372 a_n1613_43370# a_288_46660# 0.01808f
C1373 a_19321_45002# a_20843_47204# 1.68e-20
C1374 a_12549_44172# a_n743_46660# 0.03191f
C1375 a_13747_46662# a_20916_46384# 2.31e-20
C1376 a_12607_44458# a_10949_43914# 7.79e-20
C1377 a_19615_44636# a_20362_44736# 2.51e-19
C1378 a_11967_42832# a_20640_44752# 0.588649f
C1379 a_19006_44850# a_20679_44626# 6.41e-22
C1380 a_n2661_43922# a_n809_44244# 0.010689f
C1381 a_n2293_43922# a_n1549_44318# 1.15e-19
C1382 a_n2661_42834# a_n984_44318# 0.012148f
C1383 a_8975_43940# a_10807_43548# 2.16e-19
C1384 a_n2293_42834# a_n1699_43638# 0.005603f
C1385 a_11823_42460# a_13460_43230# 0.00394f
C1386 a_1307_43914# a_3540_43646# 0.005727f
C1387 a_10193_42453# a_17595_43084# 2.47e-19
C1388 a_13249_42308# a_12089_42308# 0.002934f
C1389 a_18479_45785# a_4361_42308# 5.55e-20
C1390 a_8953_45002# a_8791_43396# 4.51e-19
C1391 a_5111_44636# a_6809_43396# 0.002123f
C1392 a_3537_45260# a_8229_43396# 1.13e-20
C1393 a_117_45144# VDD 2.04e-19
C1394 a_n1630_35242# VIN_N 0.040646f
C1395 a_n3420_37984# a_n2956_38680# 8.07e-19
C1396 a_4223_44672# a_4185_45028# 0.031094f
C1397 a_n699_43396# a_3699_46348# 1.2e-21
C1398 a_4743_44484# a_3483_46348# 6.71e-19
C1399 a_17517_44484# a_19466_46812# 1.01e-19
C1400 a_15493_43940# a_13661_43548# 1.28948f
C1401 a_7281_43914# a_4646_46812# 0.021965f
C1402 a_14021_43940# a_12891_46348# 3.26e-20
C1403 a_n2293_43922# a_13059_46348# 5.13e-21
C1404 a_13565_44260# a_768_44030# 7.87e-20
C1405 a_13829_44260# a_12549_44172# 4.49e-19
C1406 a_13777_45326# a_13259_45724# 0.043567f
C1407 a_413_45260# a_1848_45724# 2.84e-21
C1408 a_1667_45002# a_n755_45592# 0.002f
C1409 a_n1059_45260# a_n443_42852# 0.130036f
C1410 a_3537_45260# a_n863_45724# 1.54e-20
C1411 a_4927_45028# a_n2661_45546# 0.001509f
C1412 a_19778_44110# a_18819_46122# 5.3e-21
C1413 a_11691_44458# a_13925_46122# 3.94e-21
C1414 a_n2661_44458# a_8199_44636# 0.069807f
C1415 a_18911_45144# a_18985_46122# 7.42e-22
C1416 a_3626_43646# a_4791_45118# 0.006599f
C1417 a_14311_47204# VDD 0.241476f
C1418 a_15890_42674# a_7174_31319# 2.06e-20
C1419 a_4958_30871# a_17303_42282# 0.168656f
C1420 a_n2293_46634# a_167_45260# 0.087596f
C1421 a_171_46873# a_376_46348# 0.080253f
C1422 a_n1925_46634# a_1138_42852# 5.27e-19
C1423 a_n743_46660# a_1208_46090# 0.045297f
C1424 a_n133_46660# a_472_46348# 6.87e-19
C1425 a_21588_30879# a_4185_45028# 2.74e-19
C1426 a_n2438_43548# a_805_46414# 2.09e-19
C1427 a_12991_46634# a_13607_46688# 0.002207f
C1428 a_5894_47026# a_765_45546# 1.39e-19
C1429 a_5807_45002# a_7920_46348# 3.4e-20
C1430 a_768_44030# a_9290_44172# 0.189655f
C1431 a_12549_44172# a_11189_46129# 3.08e-20
C1432 a_11309_47204# a_11387_46155# 0.061891f
C1433 a_n881_46662# a_14275_46494# 0.004854f
C1434 a_22959_47212# a_10809_44734# 0.005622f
C1435 a_4915_47217# a_14371_46494# 0.001038f
C1436 a_n1151_42308# a_13259_45724# 5.41e-19
C1437 a_n2288_47178# a_n2293_45546# 5.3e-21
C1438 SMPL_ON_P a_n2810_45572# 0.039568f
C1439 a_n2497_47436# a_n1079_45724# 5.93e-19
C1440 a_18248_44752# a_16823_43084# 1.7e-19
C1441 a_n1761_44111# a_n1809_43762# 4.8e-19
C1442 a_n809_44244# a_n447_43370# 0.003582f
C1443 a_19862_44208# a_15493_43940# 0.534481f
C1444 a_20365_43914# a_11341_43940# 0.010232f
C1445 a_10057_43914# a_4361_42308# 3.62e-20
C1446 a_n984_44318# a_n1352_43396# 5.83e-20
C1447 a_13483_43940# a_13565_44260# 0.003935f
C1448 a_10193_42453# a_21887_42336# 3.37e-21
C1449 a_n2956_37592# a_n2840_42282# 8.96e-21
C1450 a_n2017_45002# a_n3674_38216# 0.004889f
C1451 a_n2810_45028# a_n3674_38680# 0.022953f
C1452 a_n2065_43946# VDD 0.4213f
C1453 a_10490_45724# a_10306_45572# 8.03e-20
C1454 a_8746_45002# a_10544_45572# 4.52e-20
C1455 a_2711_45572# a_16211_45572# 0.001012f
C1456 C9_N_btm C3_P_btm 6.09e-19
C1457 C8_N_btm C2_P_btm 1.77e-19
C1458 a_15493_43940# a_4185_45028# 0.039364f
C1459 a_791_42968# a_768_44030# 1.22e-19
C1460 a_484_44484# a_n443_42852# 3.87e-19
C1461 a_n2661_42834# a_3503_45724# 2.21e-21
C1462 a_n2661_43922# a_3316_45546# 3.15e-20
C1463 a_895_43940# a_526_44458# 0.018069f
C1464 a_14815_43914# a_n357_42282# 1.18e-20
C1465 a_n4318_39768# a_n2956_39304# 0.023377f
C1466 a_2479_44172# a_n1925_42282# 3.15e-21
C1467 a_17730_32519# a_8049_45260# 3.56e-20
C1468 a_17701_42308# a_13507_46334# 7.88e-21
C1469 a_8037_42858# a_n1613_43370# 0.047354f
C1470 a_13483_43940# a_9290_44172# 0.005971f
C1471 a_n2661_42282# a_2324_44458# 0.001316f
C1472 a_10949_43914# a_10903_43370# 0.451961f
C1473 a_14226_46987# VDD 6.34e-20
C1474 a_5068_46348# a_5204_45822# 0.20685f
C1475 a_18280_46660# a_10809_44734# 0.002977f
C1476 a_3483_46348# a_8016_46348# 0.019798f
C1477 a_12741_44636# a_17957_46116# 9.01e-21
C1478 a_n97_42460# a_15095_43370# 0.002411f
C1479 a_3626_43646# a_8791_43396# 1.23e-21
C1480 a_14021_43940# a_4361_42308# 0.003147f
C1481 a_5891_43370# a_n784_42308# 6.43e-20
C1482 a_n356_44636# a_2351_42308# 1.17e-19
C1483 a_5883_43914# a_8515_42308# 5.6e-22
C1484 a_5343_44458# a_8685_42308# 5.14e-19
C1485 a_18533_43940# a_16137_43396# 4.77e-20
C1486 a_1431_47204# DATA[1] 0.334099f
C1487 a_2124_47436# DATA[0] 2.79e-21
C1488 a_13667_43396# VDD 0.402378f
C1489 a_5907_45546# a_5518_44484# 2.57e-19
C1490 a_2711_45572# a_5883_43914# 2.93e-21
C1491 a_n913_45002# a_2382_45260# 0.021705f
C1492 a_n2017_45002# a_3065_45002# 0.043491f
C1493 a_3357_43084# a_5205_44484# 0.020505f
C1494 a_685_42968# a_1138_42852# 6.59e-20
C1495 a_15486_42560# a_12549_44172# 1.17e-21
C1496 a_10553_43218# a_3090_45724# 8.81e-20
C1497 a_5934_30871# a_n2312_38680# 4.54e-21
C1498 a_4699_43561# a_n2661_45546# 0.013733f
C1499 a_1049_43396# a_n863_45724# 1.03e-19
C1500 a_10149_43396# a_526_44458# 0.003062f
C1501 a_n1190_43762# a_n755_45592# 2.34e-20
C1502 a_21613_42308# a_13507_46334# 0.035917f
C1503 a_3422_30871# EN_VIN_BSTR_P 0.182769f
C1504 a_n755_45592# VDD 2.41485f
C1505 a_3357_43084# a_n971_45724# 0.565799f
C1506 a_5907_45546# a_n2661_46634# 7.09e-21
C1507 a_9049_44484# a_768_44030# 0.006069f
C1508 a_3175_45822# a_n2293_46634# 1.98e-19
C1509 a_10193_42453# a_11309_47204# 0.006435f
C1510 a_11823_42460# a_n881_46662# 0.036994f
C1511 a_15765_45572# a_10227_46804# 4.04e-19
C1512 a_8696_44636# a_16327_47482# 0.087584f
C1513 a_n1925_42282# a_n443_42852# 0.02261f
C1514 a_526_44458# a_1609_45822# 3.1e-20
C1515 a_n2433_43396# a_n2472_42282# 2.98e-20
C1516 a_16547_43609# a_16414_43172# 0.143695f
C1517 a_16243_43396# a_16795_42852# 8.18e-20
C1518 a_n2472_42826# a_n4318_38680# 0.158196f
C1519 a_n2157_42858# a_n3674_39304# 2.93e-19
C1520 a_n1991_42858# a_n1076_43230# 0.123255f
C1521 a_n1853_43023# a_n13_43084# 0.109925f
C1522 a_743_42282# a_5111_42852# 8.1e-20
C1523 a_16137_43396# a_17595_43084# 0.001749f
C1524 a_2982_43646# a_13291_42460# 2.6e-19
C1525 a_n4318_39304# a_n4318_38216# 0.023477f
C1526 a_14401_32519# COMP_P 8.68e-21
C1527 a_8270_45546# CLK 7.07e-21
C1528 a_20256_43172# VDD 7.47e-19
C1529 a_20107_45572# a_20679_44626# 0.001176f
C1530 a_16751_45260# a_14539_43914# 3.77e-20
C1531 a_2809_45028# a_2779_44458# 0.001617f
C1532 a_8746_45002# a_10949_43914# 4.6e-20
C1533 a_10490_45724# a_10729_43914# 2.89e-21
C1534 a_10193_42453# a_10807_43548# 0.060211f
C1535 a_21188_45572# a_11967_42832# 2.72e-22
C1536 a_3232_43370# a_8375_44464# 0.022129f
C1537 a_n467_45028# a_n2661_42834# 0.001028f
C1538 a_19479_31679# a_17517_44484# 0.002614f
C1539 a_6431_45366# a_6109_44484# 2.93e-19
C1540 a_5691_45260# a_5891_43370# 3.67e-21
C1541 a_3537_45260# a_9313_44734# 6.69e-20
C1542 a_5205_44484# a_5826_44734# 0.003766f
C1543 a_6171_45002# a_7640_43914# 8.9e-20
C1544 a_20273_45572# a_20640_44752# 7.28e-19
C1545 a_5742_30871# a_4185_45028# 0.062132f
C1546 a_n2104_42282# a_n1925_42282# 0.166917f
C1547 a_945_42968# a_n357_42282# 4.86e-19
C1548 a_8325_42308# a_8199_44636# 0.004591f
C1549 a_4808_45572# a_3483_46348# 3.56e-19
C1550 a_17478_45572# a_16388_46812# 5.42e-21
C1551 a_16020_45572# a_13059_46348# 2.07e-20
C1552 a_19431_45546# a_19692_46634# 5.98e-20
C1553 a_19256_45572# a_19466_46812# 0.041135f
C1554 a_18799_45938# a_15227_44166# 7.44e-21
C1555 a_13711_45394# a_12891_46348# 0.003687f
C1556 a_15903_45785# a_765_45546# 2.27e-20
C1557 a_5111_44636# a_5167_46660# 1.66e-20
C1558 a_413_45260# a_7411_46660# 2.01e-20
C1559 a_5691_45260# a_4817_46660# 8.09e-19
C1560 a_5205_44484# a_3877_44458# 5.39e-21
C1561 a_6431_45366# a_4646_46812# 8.39e-19
C1562 a_3775_45552# a_5204_45822# 9.09e-22
C1563 a_2711_45572# a_9569_46155# 6.07e-20
C1564 a_6667_45809# a_6419_46155# 6.84e-19
C1565 a_5263_45724# a_5937_45572# 0.002746f
C1566 a_14539_43914# a_4915_47217# 1.6e-19
C1567 a_n356_44636# a_584_46384# 0.268036f
C1568 a_19268_43646# a_19332_42282# 2.41e-19
C1569 a_4361_42308# a_15764_42576# 0.009129f
C1570 a_5649_42852# a_14113_42308# 9.77e-20
C1571 a_5342_30871# a_n1630_35242# 0.035143f
C1572 a_20205_31679# EN_VIN_BSTR_N 0.003421f
C1573 a_13507_46334# a_12891_46348# 0.076674f
C1574 a_16588_47582# a_5807_45002# 0.040789f
C1575 a_n2312_40392# a_n1613_43370# 4.82e-21
C1576 a_10227_46804# a_16942_47570# 0.00186f
C1577 a_4915_47217# a_2107_46812# 6.45e-20
C1578 a_6575_47204# a_n743_46660# 5.55e-20
C1579 a_n971_45724# a_3877_44458# 0.927248f
C1580 a_n1741_47186# a_5385_46902# 1.59e-20
C1581 a_2063_45854# a_2959_46660# 2.88e-19
C1582 a_n1151_42308# a_1799_45572# 2.59e-19
C1583 a_2952_47436# a_2609_46660# 0.006778f
C1584 a_2905_45572# a_2443_46660# 0.026052f
C1585 a_n2109_47186# a_5907_46634# 0.001384f
C1586 a_8696_44636# a_10341_43396# 6.7e-21
C1587 a_n1352_44484# a_n984_44318# 7.43e-19
C1588 a_n452_44636# a_n809_44244# 0.002409f
C1589 a_n2661_42834# a_n2661_43922# 0.841361f
C1590 a_1307_43914# a_2455_43940# 0.047238f
C1591 a_7499_43078# a_5649_42852# 2.19e-19
C1592 a_18989_43940# a_20640_44752# 1.37e-21
C1593 a_10193_42453# a_13467_32519# 0.005873f
C1594 a_626_44172# a_726_44056# 7.66e-19
C1595 a_n2661_45010# a_1756_43548# 2.49e-21
C1596 en_comp a_n2012_43396# 4.42e-20
C1597 a_2437_43646# a_2896_43646# 5.48e-19
C1598 a_n1059_45260# a_n229_43646# 3.39e-19
C1599 a_n3565_39304# a_n2956_38216# 0.02162f
C1600 a_n2810_45028# VDD 0.526631f
C1601 a_22400_42852# a_22521_39511# 0.031206f
C1602 a_2455_43940# a_n443_46116# 0.010179f
C1603 a_17538_32519# w_11334_34010# 0.036508f
C1604 a_n2661_43370# a_1823_45246# 0.112095f
C1605 a_18184_42460# a_11415_45002# 0.006818f
C1606 a_18587_45118# a_12741_44636# 0.005591f
C1607 a_18494_42460# a_20202_43084# 0.166633f
C1608 a_8488_45348# a_3483_46348# 0.003238f
C1609 a_n2293_42834# a_4185_45028# 0.022725f
C1610 a_n2661_44458# a_765_45546# 1.25e-21
C1611 a_18443_44721# a_3090_45724# 3.2e-20
C1612 a_16112_44458# a_15227_44166# 0.073746f
C1613 a_3905_42865# a_768_44030# 0.011432f
C1614 a_3065_45002# a_526_44458# 0.138202f
C1615 a_20365_43914# a_16327_47482# 0.007136f
C1616 a_10949_43914# a_4883_46098# 3.15e-21
C1617 a_n1453_44318# a_n1613_43370# 9.54e-19
C1618 a_5837_45348# a_5937_45572# 2.99e-19
C1619 a_15415_45028# a_2324_44458# 0.03757f
C1620 a_9885_42558# a_10533_42308# 5.68e-21
C1621 a_9803_42558# a_5742_30871# 0.002197f
C1622 a_n4318_38216# a_n4334_40480# 9.74e-20
C1623 a_5534_30871# C1_P_btm 1.06e-19
C1624 EN_VIN_BSTR_P VREF_GND 0.85739f
C1625 a_11530_34132# VIN_N 1.547f
C1626 a_4915_47217# a_14493_46090# 1.95e-19
C1627 a_6151_47436# a_13351_46090# 4.87e-21
C1628 a_9313_45822# a_9569_46155# 0.019679f
C1629 a_n1435_47204# a_5937_45572# 1.19e-20
C1630 a_n2312_40392# a_n2293_46098# 7.25e-19
C1631 a_n2312_39304# a_n2472_46090# 0.006797f
C1632 a_5807_45002# a_14447_46660# 8.93e-19
C1633 a_7715_46873# a_8492_46660# 5.47e-21
C1634 a_3877_44458# a_8023_46660# 1.47e-20
C1635 a_6540_46812# a_6682_46987# 0.005572f
C1636 a_7577_46660# a_8667_46634# 0.041879f
C1637 a_8145_46902# a_7927_46660# 0.209641f
C1638 a_7411_46660# a_9863_46634# 2.84e-21
C1639 a_n2661_42834# a_n447_43370# 0.006056f
C1640 a_n2293_43922# a_n1177_43370# 1.47e-22
C1641 a_11691_44458# a_17499_43370# 3.7e-20
C1642 a_11827_44484# a_18783_43370# 1.47e-20
C1643 a_n2293_42834# a_n2157_42858# 0.058852f
C1644 a_1423_45028# a_3935_42891# 2.7e-22
C1645 a_7499_43078# a_7963_42308# 5.61e-19
C1646 a_n913_45002# a_1709_42852# 0.0021f
C1647 a_3357_43084# a_3863_42891# 5.79e-19
C1648 a_n1059_45260# a_1793_42852# 4.52e-19
C1649 a_n4209_38216# C9_P_btm 1.91e-20
C1650 a_n4064_39072# VCM 0.035838f
C1651 a_2711_45572# a_8162_45546# 0.019489f
C1652 a_6194_45824# a_4880_45572# 4.69e-20
C1653 a_5263_45724# a_5437_45600# 0.006584f
C1654 a_3775_45552# a_3733_45822# 7.47e-21
C1655 a_2998_44172# a_1823_45246# 0.062531f
C1656 a_5025_43940# a_3090_45724# 4.03e-19
C1657 a_8229_43396# a_n2293_46634# 2.24e-19
C1658 a_n2661_43922# a_5066_45546# 4.26e-20
C1659 a_n699_43396# a_n755_45592# 0.185444f
C1660 a_4743_44484# a_n357_42282# 5.15e-21
C1661 a_4361_42308# a_13507_46334# 0.040714f
C1662 a_10341_42308# a_2063_45854# 6.99e-21
C1663 en_comp a_22545_38993# 7.26e-21
C1664 a_19479_31679# EN_VIN_BSTR_N 0.007584f
C1665 a_n4209_38502# a_n4209_38216# 0.041706f
C1666 a_n4064_38528# a_n2860_38778# 0.003766f
C1667 a_4958_30871# C8_N_btm 0.001147f
C1668 a_n4318_37592# a_n4334_37440# 0.083644f
C1669 a_22591_46660# a_20820_30879# 0.166885f
C1670 a_11415_45002# a_12741_44636# 1.07921f
C1671 a_20202_43084# a_22959_46660# 2.07e-19
C1672 a_765_45546# a_2804_46116# 1.28e-20
C1673 a_n2661_46634# a_n1099_45572# 5.05e-20
C1674 a_n2293_46634# a_n863_45724# 0.157683f
C1675 a_n743_46660# a_n2661_45546# 0.013544f
C1676 a_n2438_43548# a_n2810_45572# 4.17e-19
C1677 a_3090_45724# a_17583_46090# 0.003153f
C1678 a_15368_46634# a_2324_44458# 0.00404f
C1679 a_10933_46660# a_9290_44172# 2.81e-19
C1680 a_7542_44172# a_743_42282# 2.49e-21
C1681 a_20365_43914# a_10341_43396# 1.17e-20
C1682 a_5013_44260# a_4361_42308# 1.27e-20
C1683 a_14539_43914# a_13291_42460# 2.89e-21
C1684 a_n1352_43396# a_n447_43370# 4.88e-19
C1685 a_15682_43940# a_15681_43442# 1.6e-19
C1686 a_11341_43940# a_14205_43396# 0.001925f
C1687 a_n2267_43396# a_n1809_43762# 0.034619f
C1688 a_5891_43370# a_7309_43172# 0.002083f
C1689 a_n2433_43396# a_n1821_43396# 3.82e-19
C1690 a_11967_42832# a_10922_42852# 4.37e-20
C1691 a_n2956_37592# a_n2302_39866# 0.006499f
C1692 a_n2129_43609# VDD 0.400674f
C1693 a_20273_45572# a_21188_45572# 0.125324f
C1694 a_14495_45572# a_14180_45002# 9.07e-19
C1695 a_11823_42460# a_1307_43914# 0.049611f
C1696 a_13249_42308# a_14537_43396# 0.020089f
C1697 a_7227_45028# a_7418_45394# 2.88e-19
C1698 a_10907_45822# a_10775_45002# 1.92e-19
C1699 a_20107_45572# a_20528_45572# 0.086377f
C1700 a_8952_43230# a_3090_45724# 1.36e-19
C1701 a_458_43396# a_526_44458# 0.085782f
C1702 a_9145_43396# a_8199_44636# 0.020485f
C1703 a_835_46155# VDD 7.28e-19
C1704 a_9049_44484# a_9067_47204# 3.2e-20
C1705 a_17957_46116# a_16375_45002# 0.017118f
C1706 a_18189_46348# a_19240_46482# 1.71e-21
C1707 a_8016_46348# a_n357_42282# 3.18e-20
C1708 a_167_45260# a_2277_45546# 0.214157f
C1709 a_8147_43396# a_8605_42826# 0.003157f
C1710 a_8791_43396# a_8037_42858# 0.001631f
C1711 a_16977_43638# a_743_42282# 1.08e-20
C1712 a_17499_43370# a_4190_30871# 2.22e-19
C1713 a_15781_43660# a_5649_42852# 4.06e-21
C1714 a_15743_43084# a_16823_43084# 0.031733f
C1715 a_n2661_42282# a_1606_42308# 0.082268f
C1716 a_3422_30871# a_15959_42545# 5.29e-20
C1717 a_11967_42832# a_17531_42308# 0.003854f
C1718 a_21195_42852# VDD 0.285496f
C1719 a_n1059_45260# CAL_N 0.001614f
C1720 a_15415_45028# a_16922_45042# 9.08e-21
C1721 a_16019_45002# a_16405_45348# 5.59e-19
C1722 a_1307_43914# a_16321_45348# 8.2e-20
C1723 a_8696_44636# a_n2293_43922# 0.002811f
C1724 a_4185_45348# a_n2661_43370# 1.42e-19
C1725 a_2382_45260# a_n2661_44458# 0.032484f
C1726 a_n467_45028# a_n1352_44484# 1.49e-19
C1727 a_n913_45002# a_5343_44458# 0.020508f
C1728 a_5907_45546# a_765_45546# 6.13e-21
C1729 a_13249_42308# a_3090_45724# 0.032019f
C1730 a_413_45260# a_13661_43548# 2.4e-20
C1731 a_2437_43646# a_948_46660# 2.21e-20
C1732 a_n2661_45010# a_n2312_38680# 1.97e-21
C1733 a_n2293_45010# a_n2293_46634# 0.036081f
C1734 a_5147_45002# a_768_44030# 0.191082f
C1735 a_14309_45028# a_4915_47217# 0.004859f
C1736 a_16751_45260# a_11453_44696# 0.002984f
C1737 a_8191_45002# a_n1613_43370# 2.41e-21
C1738 a_7705_45326# a_n881_46662# 3.83e-20
C1739 a_8685_43396# a_14113_42308# 5.76e-20
C1740 a_n2840_42826# a_n3674_38680# 0.019613f
C1741 a_10835_43094# a_11554_42852# 0.086334f
C1742 a_743_42282# a_n1630_35242# 0.004023f
C1743 a_n2293_42282# a_3445_43172# 0.009537f
C1744 a_10518_42984# a_10752_42852# 0.006453f
C1745 a_10991_42826# a_11229_43218# 0.001705f
C1746 a_10796_42968# a_11301_43218# 2.28e-19
C1747 a_13467_32519# a_n784_42308# 0.014901f
C1748 a_3626_43646# a_18220_42308# 9.35e-19
C1749 a_13759_46122# CLK 2.17e-20
C1750 a_n2302_40160# VDD 0.428934f
C1751 a_n2109_47186# a_768_44030# 2.81e-21
C1752 a_n1741_47186# a_12891_46348# 0.107238f
C1753 a_n971_45724# a_8128_46384# 0.041637f
C1754 a_n785_47204# a_n881_46662# 6.65e-20
C1755 a_4915_47217# a_11453_44696# 0.026396f
C1756 a_327_47204# a_n1613_43370# 0.002699f
C1757 a_15507_47210# a_16327_47482# 0.425757f
C1758 a_15811_47375# a_16241_47178# 0.003645f
C1759 a_11599_46634# a_16023_47582# 1.42e-20
C1760 a_n1151_42308# a_2747_46873# 0.009962f
C1761 a_2952_47436# a_3094_47570# 0.007833f
C1762 a_2063_45854# a_2266_47243# 4.14e-19
C1763 a_13717_47436# a_18143_47464# 3.4e-19
C1764 a_12861_44030# a_10227_46804# 0.291378f
C1765 a_19778_44110# a_19615_44636# 0.012379f
C1766 a_18184_42460# a_11967_42832# 0.024012f
C1767 a_n1352_44484# a_n2661_43922# 0.007747f
C1768 a_n452_44636# a_n2661_42834# 0.002825f
C1769 a_7499_43078# a_8685_43396# 0.153217f
C1770 a_n2293_42834# a_n1761_44111# 0.03111f
C1771 a_10057_43914# a_5891_43370# 0.197199f
C1772 a_5883_43914# a_9241_44734# 0.010354f
C1773 a_8975_43940# a_8375_44464# 2.42e-20
C1774 a_20193_45348# a_17517_44484# 0.015762f
C1775 a_8701_44490# a_9313_44734# 5.25e-19
C1776 a_16922_45042# a_19279_43940# 0.018289f
C1777 a_8696_44636# a_n97_42460# 9.12e-22
C1778 a_11827_44484# a_16335_44484# 7.13e-19
C1779 a_3232_43370# a_10949_43914# 0.093316f
C1780 a_6171_45002# a_10729_43914# 2.56e-21
C1781 a_20447_31679# a_14021_43940# 1.09e-20
C1782 a_17531_42308# a_13259_45724# 0.009212f
C1783 a_16333_45814# VDD 0.201203f
C1784 a_20820_30879# C7_N_btm 0.184297f
C1785 a_5342_30871# a_11530_34132# 0.012973f
C1786 a_13159_45002# a_12741_44636# 7.19e-20
C1787 a_13556_45296# a_11415_45002# 0.16025f
C1788 a_4574_45260# a_1823_45246# 3.32e-19
C1789 a_2382_45260# a_2804_46116# 1.18e-21
C1790 a_2680_45002# a_2698_46116# 2.37e-20
C1791 a_17613_45144# a_3090_45724# 1.41e-19
C1792 a_413_45260# a_4185_45028# 0.191095f
C1793 a_4223_44672# a_5257_43370# 0.016657f
C1794 a_9313_44734# a_n2293_46634# 0.022598f
C1795 a_12829_44484# a_12549_44172# 3.48e-20
C1796 a_13296_44484# a_12891_46348# 3.98e-19
C1797 a_3775_45552# a_3503_45724# 0.13675f
C1798 a_11136_45572# a_10586_45546# 0.006861f
C1799 a_5024_45822# a_n755_45592# 1.65e-20
C1800 a_15225_45822# a_8049_45260# 7.33e-20
C1801 a_2437_43646# a_13925_46122# 1.99e-20
C1802 a_n1059_45260# a_8199_44636# 0.019728f
C1803 a_n2017_45002# a_5937_45572# 2.08e-20
C1804 a_3357_43084# a_12594_46348# 9.87e-21
C1805 a_n822_43940# a_n1151_42308# 3.16e-20
C1806 a_1755_42282# a_5379_42460# 0.045501f
C1807 a_15597_42852# a_15051_42282# 3.4e-19
C1808 a_2725_42558# a_2713_42308# 0.01129f
C1809 COMP_P a_5934_30871# 0.028728f
C1810 a_4190_30871# C1_P_btm 7.67e-20
C1811 a_22521_40055# a_22459_39145# 0.129251f
C1812 a_5807_45002# a_10150_46912# 0.007534f
C1813 a_n1925_46634# a_5907_46634# 0.010645f
C1814 a_n743_46660# a_5385_46902# 5.02e-22
C1815 a_1799_45572# a_3177_46902# 7.67e-21
C1816 a_n2661_46098# a_2609_46660# 6e-19
C1817 a_2107_46812# a_2162_46660# 0.002508f
C1818 a_8128_46384# a_8023_46660# 8e-19
C1819 a_11453_44696# a_18834_46812# 0.010577f
C1820 a_12465_44636# a_19692_46634# 6.79e-20
C1821 a_4883_46098# a_10425_46660# 2.44e-19
C1822 a_10227_46804# a_14180_46812# 0.008201f
C1823 a_15673_47210# a_16388_46812# 4.51e-19
C1824 a_15811_47375# a_16721_46634# 2.3e-19
C1825 a_12861_44030# a_17339_46660# 1.25428f
C1826 a_13717_47436# a_765_45546# 0.009975f
C1827 a_n2497_47436# a_1823_45246# 0.025359f
C1828 a_n2109_47186# a_1176_45822# 1.41e-19
C1829 a_n815_47178# a_n1076_46494# 6.69e-19
C1830 a_327_47204# a_n2293_46098# 8.71e-21
C1831 a_n699_43396# a_n2129_43609# 0.062898f
C1832 a_n1549_44318# a_n984_44318# 7.99e-20
C1833 a_n1899_43946# a_644_44056# 2.13e-20
C1834 a_11823_42460# a_13003_42852# 0.002475f
C1835 a_3357_43084# a_4520_42826# 5.54e-19
C1836 a_n967_45348# a_n1076_43230# 0.019022f
C1837 a_n2956_37592# a_n3674_39304# 0.023366f
C1838 a_n2810_45028# a_n4318_38680# 0.023185f
C1839 a_n2017_45002# a_n967_43230# 3.36e-21
C1840 a_5205_44484# a_743_42282# 2.08e-20
C1841 a_n2302_37690# VDD 0.350133f
C1842 a_n2129_44697# VDD 1.4165f
C1843 a_7174_31319# EN_VIN_BSTR_P 0.053205f
C1844 a_22465_38105# a_22705_38406# 0.003319f
C1845 a_13258_32519# EN_VIN_BSTR_N 0.040234f
C1846 a_4958_30871# C2_P_btm 9.53e-20
C1847 a_743_42282# a_n971_45724# 2.96e-19
C1848 a_11967_42832# a_12741_44636# 0.004783f
C1849 a_20362_44736# a_11415_45002# 0.001672f
C1850 a_20640_44752# a_20202_43084# 0.027593f
C1851 a_14112_44734# a_3483_46348# 2.1e-20
C1852 a_8333_44056# a_8270_45546# 0.001906f
C1853 a_4093_43548# a_768_44030# 1.82e-19
C1854 a_n4318_39304# a_n2956_39768# 0.02353f
C1855 a_17973_43940# a_6755_46942# 6e-19
C1856 a_18587_45118# a_16375_45002# 2.59e-20
C1857 a_18184_42460# a_13259_45724# 0.001266f
C1858 a_6298_44484# a_526_44458# 8.53e-21
C1859 a_n2661_43370# a_n2293_45546# 0.131199f
C1860 a_19721_31679# a_8049_45260# 7.57e-19
C1861 a_9803_43646# a_10227_46804# 0.003261f
C1862 a_16131_47204# VDD 0.142103f
C1863 a_n3565_39590# a_n3690_39616# 0.246863f
C1864 a_n4334_39616# a_n3420_39616# 0.015897f
C1865 a_n4209_39590# a_n2946_39866# 0.022704f
C1866 a_22223_47212# a_20205_31679# 8.22e-20
C1867 a_4883_46098# a_21167_46155# 3.61e-19
C1868 a_5257_43370# a_6419_46155# 0.186651f
C1869 a_2107_46812# a_10809_44734# 1.51e-20
C1870 a_11309_47204# a_11387_46482# 0.006175f
C1871 a_n2661_46634# a_n1925_42282# 8.9e-20
C1872 a_171_46873# a_n1379_46482# 8.94e-21
C1873 a_19692_46634# a_20528_46660# 0.021985f
C1874 a_17609_46634# a_18280_46660# 0.094543f
C1875 a_14035_46660# a_765_45546# 9.28e-19
C1876 a_10428_46928# a_3483_46348# 3.44e-19
C1877 a_19279_43940# a_15743_43084# 6.64e-19
C1878 a_18579_44172# a_18429_43548# 6.43e-20
C1879 a_n2661_42834# a_n1641_43230# 9.58e-19
C1880 a_n2293_43922# a_n1991_42858# 0.007113f
C1881 a_n356_44636# a_8952_43230# 4.57e-21
C1882 a_n2661_42282# a_3539_42460# 1.44e-19
C1883 a_16789_44484# a_16823_43084# 4.65e-20
C1884 a_5111_44636# a_7227_42308# 1.41e-20
C1885 a_3537_45260# a_8515_42308# 3.86e-22
C1886 a_n913_45002# a_12563_42308# 1.51e-19
C1887 a_n1059_45260# a_13070_42354# 2.07e-20
C1888 a_n2017_45002# a_13575_42558# 0.006408f
C1889 en_comp a_11323_42473# 4.34e-21
C1890 a_15493_43396# VDD 2.34659f
C1891 a_15861_45028# a_17478_45572# 0.080824f
C1892 a_8696_44636# a_16020_45572# 1.4e-20
C1893 a_2711_45572# a_3537_45260# 0.0026f
C1894 a_4099_45572# a_3065_45002# 3.74e-19
C1895 a_17499_43370# a_15227_44166# 0.021724f
C1896 a_1414_42308# a_n357_42282# 0.027118f
C1897 a_2675_43914# a_n863_45724# 2e-20
C1898 a_7309_42852# a_n1613_43370# 8.11e-20
C1899 a_7754_40130# RST_Z 0.022036f
C1900 a_22400_42852# a_16327_47482# 1.22e-21
C1901 a_3823_42558# a_584_46384# 3.7e-20
C1902 a_n327_42308# a_n1151_42308# 1.59e-19
C1903 VDAC_Ni a_n923_35174# 7.46e-19
C1904 a_3483_46348# VDD 2.29096f
C1905 C5_N_btm C10_N_btm 0.51798f
C1906 C6_N_btm C9_N_btm 0.165353f
C1907 C7_N_btm C8_N_btm 31.072699f
C1908 a_22465_38105# a_22469_40625# 0.072192f
C1909 a_n4064_40160# VDAC_P 0.003375f
C1910 a_12741_44636# a_13259_45724# 0.113445f
C1911 a_11415_45002# a_16375_45002# 0.080382f
C1912 a_765_45546# a_n1099_45572# 7.06e-19
C1913 a_5164_46348# a_5066_45546# 0.096188f
C1914 a_5204_45822# a_5431_46482# 0.004982f
C1915 a_5937_45572# a_526_44458# 7.57e-20
C1916 a_15015_46420# a_6945_45028# 4.64e-20
C1917 a_n3565_38216# a_n2302_37984# 0.067194f
C1918 a_n4209_39304# a_n4209_37414# 0.029637f
C1919 a_n4334_38304# a_n4251_38304# 0.007692f
C1920 a_n4209_38216# a_n3607_38304# 0.002352f
C1921 a_n1177_43370# a_n901_43156# 0.002573f
C1922 a_4699_43561# a_4361_42308# 1.18e-20
C1923 a_14205_43396# a_10341_43396# 0.033299f
C1924 a_8685_43396# a_15781_43660# 0.001931f
C1925 a_n2012_43396# a_n2157_42858# 4.38e-19
C1926 a_n1352_43396# a_n1641_43230# 0.001129f
C1927 a_9165_43940# a_8952_43230# 7.02e-20
C1928 a_14021_43940# a_17595_43084# 2.59e-21
C1929 a_15493_43940# a_21671_42860# 2.52e-21
C1930 a_3080_42308# a_13467_32519# 1.61e-19
C1931 a_n2267_43396# a_n3674_39304# 0.001257f
C1932 a_n2129_43609# a_n4318_38680# 7.92e-19
C1933 a_10695_43548# a_12281_43396# 5.09e-20
C1934 a_n97_42460# a_n1991_42858# 7.96e-21
C1935 a_11341_43940# a_22223_42860# 4.04e-19
C1936 SMPL_ON_N EN_OFFSET_CAL 0.066251f
C1937 a_n89_47570# DATA[0] 2.46e-19
C1938 a_n2840_42826# VDD 0.302305f
C1939 a_3775_45552# a_n2661_43922# 1.64e-20
C1940 a_20107_45572# a_18494_42460# 0.010062f
C1941 a_13348_45260# a_9482_43914# 0.352976f
C1942 a_13017_45260# a_13777_45326# 0.195607f
C1943 a_10180_45724# a_5891_43370# 2.51e-20
C1944 a_13159_45002# a_13556_45296# 0.006136f
C1945 a_7499_43078# a_8783_44734# 1.04e-19
C1946 a_13249_42308# a_n356_44636# 6.2e-20
C1947 a_20841_45814# a_19778_44110# 7.65e-21
C1948 a_n2661_45010# a_n2661_43370# 0.077441f
C1949 a_6171_45002# a_1423_45028# 3.32e-19
C1950 a_413_45260# a_2448_45028# 5.27e-19
C1951 a_4743_43172# a_1823_45246# 1.5e-19
C1952 a_n4334_40480# a_n2956_39768# 4.08e-19
C1953 a_12281_43396# a_n357_42282# 0.022975f
C1954 a_8423_43396# a_n443_42852# 0.007509f
C1955 a_16147_45260# a_12549_44172# 9.2e-20
C1956 a_2711_45572# a_6969_46634# 5.57e-20
C1957 a_16223_45938# a_13747_46662# 0.02646f
C1958 a_3357_43084# a_12465_44636# 1.30897f
C1959 a_2437_43646# SMPL_ON_N 2.94e-19
C1960 a_20447_31679# a_13507_46334# 8.21e-20
C1961 a_413_45260# a_14955_47212# 2.11e-19
C1962 a_n913_45002# a_10227_46804# 0.344574f
C1963 a_5205_44484# a_6151_47436# 0.010575f
C1964 a_8191_45002# a_4791_45118# 5e-20
C1965 a_n2661_45546# a_509_45572# 4.21e-19
C1966 a_380_45546# a_n443_42852# 0.030032f
C1967 a_n1099_45572# a_509_45822# 0.026885f
C1968 a_n863_45724# a_2277_45546# 0.00198f
C1969 a_3218_45724# a_3503_45724# 0.099872f
C1970 a_10341_43396# a_22400_42852# 0.004171f
C1971 a_n1641_43230# a_n2293_42282# 1.64e-20
C1972 a_10083_42826# a_10341_42308# 0.001156f
C1973 a_10835_43094# a_10991_42826# 0.105839f
C1974 a_14021_43940# a_21887_42336# 5.15e-21
C1975 a_3539_42460# a_3497_42558# 0.002673f
C1976 a_10518_42984# a_10922_42852# 0.051162f
C1977 a_16547_43609# a_17141_43172# 5.08e-20
C1978 a_4905_42826# a_6481_42558# 1.25e-20
C1979 a_11415_45002# RST_Z 4.24e-19
C1980 a_n4064_37440# VDAC_P 3.73e-19
C1981 a_3726_37500# a_4338_37500# 0.212154f
C1982 a_8791_42308# VDD 0.226318f
C1983 a_2952_47436# a_2905_45572# 0.318161f
C1984 a_2063_45854# a_n1151_42308# 0.425035f
C1985 a_2553_47502# a_3160_47472# 2.08e-19
C1986 a_n785_47204# a_n443_46116# 2.37e-20
C1987 a_19721_31679# a_22469_40625# 1.46e-20
C1988 a_n1741_47186# a_7903_47542# 0.00805f
C1989 a_n971_45724# a_6151_47436# 0.29974f
C1990 a_n1352_44484# a_n452_44636# 1.85e-19
C1991 a_n2661_44458# a_5343_44458# 0.003787f
C1992 a_13556_45296# a_11967_42832# 1.65e-21
C1993 a_11691_44458# a_15004_44636# 0.221929f
C1994 a_11827_44484# a_17767_44458# 0.014019f
C1995 a_18184_42460# a_18989_43940# 2.27e-20
C1996 a_10193_42453# a_19319_43548# 1.94e-20
C1997 a_16115_45572# a_15493_43940# 3.81e-20
C1998 a_n913_45002# a_453_43940# 2.62e-21
C1999 a_n2661_45010# a_2998_44172# 5.85e-20
C2000 a_n2017_45002# a_2479_44172# 1.51e-20
C2001 a_n1630_35242# a_20205_31679# 1.48e-19
C2002 a_7174_31319# a_10903_43370# 4.88e-21
C2003 a_6472_45840# VDD 0.257073f
C2004 a_20273_45572# a_12741_44636# 0.028616f
C2005 a_n2661_43370# a_5732_46660# 6.03e-21
C2006 a_21188_45572# a_20202_43084# 0.013137f
C2007 a_21363_45546# a_11415_45002# 0.011178f
C2008 a_4223_44672# a_5807_45002# 4.42e-21
C2009 a_n2661_44458# a_n2956_39768# 1.99e-20
C2010 a_n2293_42834# a_5257_43370# 5.57e-19
C2011 a_10157_44484# a_768_44030# 0.00283f
C2012 a_5437_45600# a_526_44458# 2.03e-20
C2013 a_3357_43084# a_20528_46660# 0.002704f
C2014 a_n913_45002# a_17339_46660# 4.56e-21
C2015 a_9313_44734# a_18597_46090# 0.029282f
C2016 a_10210_45822# a_2324_44458# 3.44e-20
C2017 a_11136_45572# a_11189_46129# 0.042798f
C2018 a_12427_45724# a_10809_44734# 0.01284f
C2019 a_14539_43914# a_n881_46662# 1.15e-20
C2020 a_16795_42852# a_15803_42450# 6.31e-20
C2021 a_20836_43172# a_20753_42852# 1.48e-19
C2022 a_5342_30871# a_15720_42674# 9.9e-20
C2023 a_4883_46098# a_4651_46660# 2e-19
C2024 a_n1435_47204# a_10554_47026# 3.08e-20
C2025 a_11459_47204# a_6755_46942# 1.05e-19
C2026 a_6151_47436# a_8023_46660# 1.79e-19
C2027 a_n1151_42308# a_12469_46902# 0.007465f
C2028 a_n1741_47186# a_12359_47026# 8.57e-21
C2029 a_n1613_43370# a_1983_46706# 0.020434f
C2030 a_2747_46873# a_3177_46902# 3.64e-20
C2031 a_n881_46662# a_2107_46812# 0.138703f
C2032 a_19321_45002# a_19594_46812# 0.267862f
C2033 a_12891_46348# a_n743_46660# 0.044305f
C2034 a_768_44030# a_n1925_46634# 5.22e-20
C2035 a_8975_43940# a_10949_43914# 2.76e-19
C2036 a_11967_42832# a_20362_44736# 0.052989f
C2037 a_19615_44636# a_20159_44458# 0.001766f
C2038 a_10057_43914# a_10807_43548# 0.039192f
C2039 a_6109_44484# a_6453_43914# 0.165572f
C2040 a_n2293_43922# a_n1331_43914# 1.37e-19
C2041 a_n2661_42834# a_n809_44244# 0.021917f
C2042 a_n2661_43922# a_n1549_44318# 0.004791f
C2043 a_1307_43914# a_2982_43646# 0.028987f
C2044 a_n2293_42834# a_n2267_43396# 0.010565f
C2045 a_3363_44484# a_1414_42308# 1.44e-20
C2046 a_11823_42460# a_13635_43156# 0.040348f
C2047 a_13249_42308# a_12379_42858# 0.029761f
C2048 a_10193_42453# a_16795_42852# 1.71e-19
C2049 a_17517_44484# a_20596_44850# 3.5e-19
C2050 a_n1059_45260# a_8945_43396# 0.002485f
C2051 a_5111_44636# a_6643_43396# 0.004357f
C2052 a_3537_45260# a_7466_43396# 1.01e-19
C2053 a_45_45144# VDD 3.5e-19
C2054 a_n1630_35242# VIN_P 0.049047f
C2055 a_5932_42308# EN_VIN_BSTR_P 0.067144f
C2056 a_n784_42308# VCM 0.195503f
C2057 a_n699_43396# a_3483_46348# 2.82e-19
C2058 a_18989_43940# a_12741_44636# 0.002238f
C2059 a_5883_43914# a_1823_45246# 3.03e-19
C2060 a_15493_43940# a_5807_45002# 1.03e-20
C2061 a_11341_43940# a_13747_46662# 0.008288f
C2062 a_6453_43914# a_4646_46812# 8.23e-20
C2063 a_20935_43940# a_19321_45002# 9.4e-19
C2064 a_13565_44260# a_12549_44172# 4.96e-19
C2065 a_13829_44260# a_12891_46348# 1.39e-19
C2066 a_12710_44260# a_768_44030# 6.85e-19
C2067 a_13556_45296# a_13259_45724# 0.019616f
C2068 a_327_44734# a_n755_45592# 0.00429f
C2069 a_n2017_45002# a_n443_42852# 0.033337f
C2070 a_5111_44636# a_n2661_45546# 0.001037f
C2071 a_n913_45002# a_n906_45572# 1.9e-19
C2072 a_11691_44458# a_13759_46122# 7.99e-21
C2073 a_18911_45144# a_18819_46122# 4e-21
C2074 a_20974_43370# a_18597_46090# 0.025672f
C2075 a_2982_43646# a_n443_46116# 0.140614f
C2076 a_15959_42545# a_7174_31319# 4.42e-20
C2077 a_5934_30871# a_n4209_39304# 5.64e-21
C2078 a_6123_31319# a_n3565_39304# 4.63e-21
C2079 a_13487_47204# VDD 0.273369f
C2080 a_5534_30871# a_n3420_37984# 0.043974f
C2081 a_171_46873# a_n1076_46494# 9.82e-20
C2082 a_n2661_46634# a_2698_46116# 1.4e-20
C2083 a_n1925_46634# a_1176_45822# 0.001268f
C2084 a_n743_46660# a_805_46414# 0.064413f
C2085 a_n2438_43548# a_472_46348# 4.71e-19
C2086 a_n133_46660# a_376_46348# 0.004089f
C2087 a_12991_46634# a_12816_46660# 0.233657f
C2088 a_12891_46348# a_11189_46129# 3.11e-20
C2089 a_5807_45002# a_6419_46155# 0.072498f
C2090 a_12549_44172# a_9290_44172# 0.053193f
C2091 a_11309_47204# a_11133_46155# 0.040357f
C2092 a_n881_46662# a_14493_46090# 0.011925f
C2093 a_11453_44696# a_10809_44734# 0.274367f
C2094 a_11459_47204# a_8049_45260# 2.62e-22
C2095 a_4915_47217# a_14180_46482# 4.16e-19
C2096 a_9313_45822# a_9241_46436# 1.86e-19
C2097 a_n2497_47436# a_n2293_45546# 0.307373f
C2098 a_n1151_42308# a_14383_46116# 1.15e-19
C2099 SMPL_ON_P a_n2840_45546# 8.99e-19
C2100 a_19478_44306# a_15493_43940# 0.025498f
C2101 a_20269_44172# a_11341_43940# 0.006087f
C2102 a_n984_44318# a_n1177_43370# 1.43e-19
C2103 a_18579_44172# a_2982_43646# 1.56e-20
C2104 a_n1352_44484# a_n1641_43230# 4.5e-21
C2105 a_n1177_44458# a_n901_43156# 7.62e-22
C2106 a_1307_43914# a_5837_42852# 4.88e-20
C2107 a_20623_43914# a_20935_43940# 0.040559f
C2108 a_10193_42453# a_21335_42336# 3.27e-20
C2109 a_n2017_45002# a_n2104_42282# 0.010745f
C2110 a_n2810_45028# a_n2840_42282# 9.69e-21
C2111 a_19479_31679# a_n1630_35242# 8.9e-20
C2112 a_n2472_43914# VDD 0.236691f
C2113 a_11823_42460# a_11682_45822# 4.41e-19
C2114 a_8746_45002# a_10306_45572# 0.007074f
C2115 a_10490_45724# a_10216_45572# 4.26e-20
C2116 C8_N_btm C3_P_btm 5.08e-19
C2117 C7_N_btm C2_P_btm 1.06e-19
C2118 a_22223_43948# a_4185_45028# 9.96e-19
C2119 a_685_42968# a_768_44030# 5.63e-19
C2120 a_n2661_42834# a_3316_45546# 6.51e-21
C2121 a_n2661_43922# a_3218_45724# 3.16e-20
C2122 a_2479_44172# a_526_44458# 0.08343f
C2123 a_11967_42832# a_16375_45002# 9.56e-20
C2124 a_7765_42852# a_n1613_43370# 0.081834f
C2125 a_12429_44172# a_9290_44172# 0.040422f
C2126 a_10729_43914# a_10903_43370# 0.082892f
C2127 a_14513_46634# VDD 0.223375f
C2128 a_5068_46348# a_5164_46348# 0.31819f
C2129 a_4704_46090# a_5204_45822# 1.24e-19
C2130 a_17639_46660# a_10809_44734# 3.03e-19
C2131 a_12741_44636# a_18189_46348# 0.00488f
C2132 a_3483_46348# a_7920_46348# 4.08e-21
C2133 a_11415_45002# a_18985_46122# 9.02e-21
C2134 a_765_45546# a_n1925_42282# 4.84e-20
C2135 a_3626_43646# a_8147_43396# 1.64e-21
C2136 a_2982_43646# a_9396_43370# 2.9e-20
C2137 a_n97_42460# a_14205_43396# 4.02e-21
C2138 a_n356_44636# a_2123_42473# 1.17e-19
C2139 a_5883_43914# a_5934_30871# 1.2e-20
C2140 a_5343_44458# a_8325_42308# 0.014133f
C2141 a_14021_43940# a_13467_32519# 0.016437f
C2142 a_11967_42832# a_11554_42852# 9.86e-20
C2143 a_1239_47204# DATA[1] 0.01925f
C2144 a_1431_47204# DATA[0] 3.79e-20
C2145 a_10695_43548# VDD 0.201247f
C2146 a_6511_45714# a_4223_44672# 1.22e-21
C2147 a_11652_45724# a_11691_44458# 8.35e-19
C2148 a_5907_45546# a_5343_44458# 1.37e-20
C2149 a_n967_45348# a_n143_45144# 1.34e-20
C2150 a_n1059_45260# a_2382_45260# 0.025598f
C2151 a_n659_45366# a_n467_45028# 5.76e-19
C2152 a_421_43172# a_1138_42852# 3.71e-20
C2153 a_8515_42308# a_n2293_46634# 1.72e-21
C2154 a_15051_42282# a_12549_44172# 1.32e-20
C2155 a_4235_43370# a_n2661_45546# 0.088313f
C2156 a_1209_43370# a_n863_45724# 8.74e-19
C2157 a_n1809_43762# a_n755_45592# 1.04e-19
C2158 a_21887_42336# a_13507_46334# 0.002462f
C2159 a_11967_42832# RST_Z 4.49e-20
C2160 a_3422_30871# a_n923_35174# 0.036845f
C2161 a_n357_42282# VDD 1.90108f
C2162 a_2437_43646# a_n237_47217# 0.076344f
C2163 a_n2661_45010# a_n2497_47436# 0.281004f
C2164 a_2711_45572# a_n2293_46634# 0.003426f
C2165 a_7499_43078# a_768_44030# 0.101779f
C2166 a_13297_45572# a_12861_44030# 8.01e-20
C2167 a_16680_45572# a_16327_47482# 0.223571f
C2168 a_15903_45785# a_10227_46804# 0.00138f
C2169 a_10306_45572# a_4883_46098# 1.7e-19
C2170 a_13259_45724# a_16375_45002# 0.60955f
C2171 a_526_44458# a_n443_42852# 2.06448f
C2172 a_n2840_43370# a_n4318_38216# 0.003324f
C2173 a_n2840_42826# a_n4318_38680# 0.044261f
C2174 a_n1423_42826# a_n1641_43230# 0.209641f
C2175 a_n2157_42858# a_n13_43084# 9.69e-21
C2176 a_n1991_42858# a_n901_43156# 0.041762f
C2177 a_n1853_43023# a_n1076_43230# 0.040291f
C2178 a_16243_43396# a_16414_43172# 9.71e-20
C2179 a_743_42282# a_4520_42826# 5.99e-20
C2180 a_16137_43396# a_16795_42852# 0.010001f
C2181 a_10341_43396# a_22223_42860# 2.12e-20
C2182 a_n2472_42826# a_n3674_39304# 7.06e-19
C2183 a_3422_30871# a_n4064_39072# 0.007014f
C2184 a_7754_40130# a_7754_39964# 0.301877f
C2185 a_18707_42852# VDD 0.132317f
C2186 a_20273_45572# a_20362_44736# 1.1e-20
C2187 a_20107_45572# a_20640_44752# 3.77e-19
C2188 a_18587_45118# a_19778_44110# 1.74e-20
C2189 a_16922_45042# a_21101_45002# 2.6e-19
C2190 a_1307_43914# a_14539_43914# 0.131617f
C2191 a_10193_42453# a_10949_43914# 0.032349f
C2192 a_21363_45546# a_11967_42832# 3.52e-22
C2193 a_6171_45002# a_6109_44484# 1.77e-19
C2194 a_3232_43370# a_7640_43914# 1.47e-19
C2195 a_n967_45348# a_n2293_43922# 0.001623f
C2196 a_n913_45002# a_14815_43914# 9.21e-19
C2197 a_5205_44484# a_5289_44734# 0.011388f
C2198 a_3537_45260# a_9241_44734# 1.1e-21
C2199 a_11323_42473# a_4185_45028# 6.87e-20
C2200 a_133_42852# a_n755_45592# 0.020885f
C2201 a_3059_42968# a_n863_45724# 0.003162f
C2202 a_n4318_38216# a_n1925_42282# 1.9e-19
C2203 a_n1630_35242# a_n2956_38680# 6.62e-19
C2204 a_873_42968# a_n357_42282# 5.83e-19
C2205 a_3080_42308# VCM 0.148824f
C2206 a_19431_45546# a_19466_46812# 0.038922f
C2207 a_2304_45348# a_n2438_43548# 2.8e-21
C2208 a_15861_45028# a_16388_46812# 1.87e-21
C2209 a_1307_43914# a_2107_46812# 0.015866f
C2210 a_13490_45394# a_12891_46348# 5.25e-19
C2211 a_8696_44636# a_16721_46634# 2.23e-19
C2212 a_6171_45002# a_4646_46812# 0.032849f
C2213 a_2437_43646# a_8270_45546# 5.82e-21
C2214 a_5147_45002# a_5167_46660# 4.02e-21
C2215 a_4927_45028# a_4817_46660# 1.88e-20
C2216 a_413_45260# a_5257_43370# 1.46e-20
C2217 a_2711_45572# a_9625_46129# 0.019316f
C2218 a_6511_45714# a_6419_46155# 3.42e-19
C2219 a_n2661_44458# a_10227_46804# 0.034728f
C2220 a_18114_32519# a_18597_46090# 4.06e-20
C2221 a_16112_44458# a_4915_47217# 7.03e-21
C2222 a_743_42282# a_15720_42674# 1.14e-19
C2223 a_4361_42308# a_15486_42560# 0.005067f
C2224 a_15743_43084# a_19332_42282# 1.97e-20
C2225 a_13259_45724# RST_Z 0.003467f
C2226 a_17730_32519# a_22521_40599# 1.2e-20
C2227 a_16327_47482# a_13747_46662# 0.128159f
C2228 a_16763_47508# a_5807_45002# 0.127783f
C2229 a_11453_44696# a_n881_46662# 4.06e-20
C2230 a_10227_46804# a_16697_47582# 8.41e-19
C2231 a_7903_47542# a_n743_46660# 8.42e-22
C2232 a_n1435_47204# a_n2661_46634# 0.002772f
C2233 a_n2109_47186# a_5167_46660# 0.004784f
C2234 a_n1741_47186# a_4817_46660# 8.55e-20
C2235 a_3160_47472# a_1799_45572# 1.08e-20
C2236 a_2553_47502# a_2609_46660# 0.001405f
C2237 a_2952_47436# a_2443_46660# 5.83e-19
C2238 a_n443_46116# a_2107_46812# 0.075963f
C2239 a_584_46384# a_2959_46660# 1.91e-19
C2240 a_n1177_44458# a_n984_44318# 1.7e-20
C2241 a_18989_43940# a_20362_44736# 5.76e-19
C2242 a_1307_43914# a_2253_43940# 0.056967f
C2243 a_17767_44458# a_18005_44484# 0.007399f
C2244 a_9313_44734# a_10809_44484# 1.08e-19
C2245 a_14539_43914# a_18579_44172# 3.18e-21
C2246 a_11649_44734# a_n2661_43922# 1.92e-19
C2247 a_n2661_45010# a_1568_43370# 5.03e-22
C2248 a_n967_45348# a_n97_42460# 3.72e-20
C2249 a_2437_43646# a_1987_43646# 2.32e-21
C2250 a_n745_45366# VDD 0.20887f
C2251 a_22400_42852# a_22780_40081# 1.96e-20
C2252 a_2253_43940# a_n443_46116# 0.011444f
C2253 a_19778_44110# a_11415_45002# 0.030651f
C2254 a_18315_45260# a_12741_44636# 0.011294f
C2255 a_18184_42460# a_20202_43084# 0.299795f
C2256 a_n2661_43370# a_1138_42852# 0.023497f
C2257 a_15004_44636# a_15227_44166# 7.56e-19
C2258 a_18287_44626# a_3090_45724# 0.037072f
C2259 a_9313_44734# a_6755_46942# 3.88e-20
C2260 a_3600_43914# a_768_44030# 0.182408f
C2261 a_20269_44172# a_16327_47482# 8.13e-19
C2262 a_n2661_42282# a_n2312_39304# 6.22e-20
C2263 a_8191_45002# a_6945_45028# 8.52e-21
C2264 a_n1644_44306# a_n1613_43370# 0.001113f
C2265 a_14797_45144# a_2324_44458# 0.048583f
C2266 a_5093_45028# a_5164_46348# 0.003673f
C2267 a_14537_43396# a_15682_46116# 2.16e-21
C2268 a_2382_45260# a_n1925_42282# 4.45e-19
C2269 a_2680_45002# a_526_44458# 0.119733f
C2270 a_9223_42460# a_5742_30871# 8.72e-20
C2271 a_n3674_38680# a_n4064_40160# 0.022279f
C2272 C3_P_btm C2_P_btm 5.99608f
C2273 a_4190_30871# a_n3420_37984# 0.032285f
C2274 a_4915_47217# a_13925_46122# 0.029041f
C2275 a_9313_45822# a_9625_46129# 0.018694f
C2276 a_n1435_47204# a_8199_44636# 1.19e-20
C2277 a_6151_47436# a_12594_46348# 2.73e-20
C2278 a_n2312_39304# a_n2840_46090# 0.007641f
C2279 a_5807_45002# a_14226_46660# 2.03e-19
C2280 a_7715_46873# a_8667_46634# 1.39e-20
C2281 a_7411_46660# a_8492_46660# 0.102325f
C2282 a_7577_46660# a_7927_46660# 0.206455f
C2283 a_22315_44484# a_14021_43940# 2.03e-21
C2284 a_n2661_42834# a_n1352_43396# 0.005746f
C2285 a_n2293_43922# a_n1917_43396# 3.53e-21
C2286 a_11827_44484# a_18525_43370# 8.62e-21
C2287 a_n2293_42834# a_n2472_42826# 0.199703f
C2288 a_1307_43914# a_7871_42858# 9.1e-21
C2289 a_7499_43078# a_6123_31319# 0.002947f
C2290 a_9482_43914# a_10835_43094# 1.01e-21
C2291 a_7845_44172# a_8333_44056# 0.065494f
C2292 a_11691_44458# a_16759_43396# 3.94e-20
C2293 a_n913_45002# a_945_42968# 0.001032f
C2294 a_n1059_45260# a_1709_42852# 4.99e-19
C2295 a_3363_44484# VDD 1.62e-19
C2296 a_n4209_38216# C10_P_btm 2.25e-20
C2297 a_n4064_39072# VREF_GND 0.048253f
C2298 a_2711_45572# a_7230_45938# 0.004731f
C2299 a_2889_44172# a_1823_45246# 3.93e-19
C2300 a_10341_43396# a_13747_46662# 4.28e-20
C2301 a_18451_43940# a_17339_46660# 0.012866f
C2302 a_9396_43370# a_2107_46812# 0.001284f
C2303 a_7466_43396# a_n2293_46634# 2.46e-19
C2304 a_n2661_42834# a_5066_45546# 1.32e-20
C2305 a_949_44458# a_1848_45724# 4.69e-19
C2306 a_18248_44752# a_18051_46116# 4.95e-21
C2307 a_n699_43396# a_n357_42282# 0.055761f
C2308 a_4223_44672# a_n755_45592# 3.55e-19
C2309 a_9313_44734# a_8049_45260# 5.74e-21
C2310 a_11967_42832# a_18985_46122# 1.38e-21
C2311 a_13467_32519# a_13507_46334# 0.043891f
C2312 a_10922_42852# a_2063_45854# 1.31e-20
C2313 en_comp a_22521_39511# 0.008551f
C2314 a_n4064_38528# a_n2302_38778# 0.239588f
C2315 a_n4334_38528# a_n4251_38528# 0.007692f
C2316 a_n2946_38778# a_n2860_38778# 0.011479f
C2317 a_n4209_38502# a_n3607_38528# 0.002294f
C2318 a_4958_30871# C7_N_btm 1.47e-19
C2319 a_n4318_37592# a_n4209_37414# 0.105251f
C2320 a_n3674_38216# a_n3565_37414# 3.9e-20
C2321 COMP_P a_8530_39574# 2.33e-19
C2322 a_11415_45002# a_20820_30879# 0.056772f
C2323 a_20202_43084# a_12741_44636# 0.22243f
C2324 a_765_45546# a_2698_46116# 4.07e-20
C2325 a_n2293_46634# a_n1079_45724# 0.002861f
C2326 a_n1021_46688# a_n2661_45546# 5.88e-21
C2327 a_n2312_38680# a_n2956_38216# 0.044798f
C2328 a_n2438_43548# a_n2840_45546# 9.23e-19
C2329 a_8145_46902# a_5066_45546# 6.07e-19
C2330 a_3090_45724# a_15682_46116# 6.43e-19
C2331 a_15368_46634# a_14840_46494# 2.19e-19
C2332 a_14976_45028# a_2324_44458# 0.086305f
C2333 a_n2472_43914# a_n4318_38680# 5.56e-21
C2334 a_n1899_43946# a_n1076_43230# 5.62e-21
C2335 a_20269_44172# a_10341_43396# 3.22e-20
C2336 a_5244_44056# a_4361_42308# 2.42e-21
C2337 a_n1177_43370# a_n447_43370# 0.010921f
C2338 a_n2267_43396# a_n2012_43396# 0.064178f
C2339 a_5829_43940# a_6031_43396# 3.18e-19
C2340 a_11341_43940# a_14358_43442# 1.43e-20
C2341 a_n1549_44318# a_n1641_43230# 1.17e-21
C2342 a_14673_44172# a_15567_42826# 4.79e-22
C2343 a_n4318_40392# a_n4318_38216# 0.023287f
C2344 a_5891_43370# a_6101_43172# 0.003606f
C2345 a_11967_42832# a_10991_42826# 7.44e-20
C2346 a_n2810_45028# a_n2302_39866# 4.97e-19
C2347 a_n2956_37592# a_n4064_39616# 0.015429f
C2348 a_n2433_43396# VDD 0.416276f
C2349 a_20273_45572# a_21363_45546# 0.042415f
C2350 a_13249_42308# a_14180_45002# 0.014749f
C2351 a_8746_45002# a_1423_45028# 2.1e-19
C2352 a_15143_45578# a_13556_45296# 9.68e-20
C2353 a_20107_45572# a_21188_45572# 0.102355f
C2354 a_10907_45822# a_8953_45002# 1.29e-20
C2355 a_20841_45814# a_20623_45572# 0.209641f
C2356 a_9127_43156# a_3090_45724# 8.78e-19
C2357 a_8292_43218# a_4646_46812# 2.63e-20
C2358 a_9803_43646# a_8016_46348# 7.46e-19
C2359 a_518_46155# VDD 0.00166f
C2360 a_2711_45572# a_18597_46090# 2.61e-20
C2361 a_8791_45572# a_n971_45724# 1.43e-20
C2362 a_18189_46348# a_16375_45002# 0.165328f
C2363 a_17957_46116# a_18243_46436# 0.010132f
C2364 a_1823_45246# a_1990_45899# 0.001705f
C2365 a_2202_46116# a_2277_45546# 0.006767f
C2366 a_167_45260# a_1609_45822# 0.141505f
C2367 a_8147_43396# a_8037_42858# 3.54e-19
C2368 a_16409_43396# a_743_42282# 8.5e-21
C2369 a_2982_43646# a_13635_43156# 1.77e-19
C2370 a_3626_43646# a_13113_42826# 5.26e-21
C2371 a_11967_42832# a_17303_42282# 0.058225f
C2372 a_3422_30871# a_15803_42450# 1.13e-19
C2373 a_19862_44208# a_20753_42852# 0.008633f
C2374 a_18783_43370# a_16823_43084# 5.12e-19
C2375 a_2107_46812# DATA[4] 2.5e-21
C2376 a_21356_42826# VDD 0.225688f
C2377 a_8696_44636# a_n2661_43922# 0.257466f
C2378 a_2711_45572# a_2675_43914# 1.32e-20
C2379 a_10193_42453# a_3422_30871# 0.404849f
C2380 a_16019_45002# a_16321_45348# 0.002468f
C2381 a_n745_45366# a_n699_43396# 2.06e-22
C2382 a_2274_45254# a_n2661_44458# 8.17e-20
C2383 a_327_44734# a_n2129_44697# 0.00201f
C2384 a_n467_45028# a_n1177_44458# 0.001271f
C2385 a_n1059_45260# a_5343_44458# 0.019826f
C2386 a_n722_43218# a_n863_45724# 6.21e-21
C2387 a_18114_32519# w_11334_34010# 9.7e-19
C2388 a_15037_45618# a_6755_46942# 1.85e-20
C2389 a_8192_45572# a_8270_45546# 0.048422f
C2390 a_1423_45028# a_4883_46098# 0.022493f
C2391 a_1307_43914# a_11453_44696# 0.037741f
C2392 a_6709_45028# a_n881_46662# 0.011804f
C2393 a_6171_45002# a_9804_47204# 7.74e-21
C2394 a_n2472_45002# a_n2293_46634# 0.001349f
C2395 a_4558_45348# a_768_44030# 5.74e-21
C2396 a_413_45260# a_5807_45002# 1.49e-19
C2397 a_n2840_42826# a_n2840_42282# 0.025171f
C2398 a_743_42282# a_564_42282# 0.169821f
C2399 a_10922_42852# a_10793_43218# 4.2e-19
C2400 a_3626_43646# a_18214_42558# 5.05e-20
C2401 a_10835_43094# a_11301_43218# 3.82e-19
C2402 a_13351_46090# CLK 4.09e-21
C2403 a_n1741_47186# a_11309_47204# 0.01734f
C2404 a_n237_47217# a_7989_47542# 5.29e-20
C2405 a_6151_47436# a_12465_44636# 0.025929f
C2406 a_n785_47204# a_n1613_43370# 3.89e-19
C2407 a_6491_46660# a_4883_46098# 5.95e-21
C2408 a_15811_47375# a_15673_47210# 0.281607f
C2409 a_15507_47210# a_16241_47178# 0.06628f
C2410 a_11599_46634# a_16327_47482# 0.526398f
C2411 a_2124_47436# a_2583_47243# 6.64e-19
C2412 a_3160_47472# a_2747_46873# 2.93e-19
C2413 a_13717_47436# a_10227_46804# 3.27e-19
C2414 a_12861_44030# a_17591_47464# 0.079093f
C2415 a_n4064_40160# VDD 2.37253f
C2416 a_18175_45572# a_18533_43940# 1.04e-21
C2417 a_19778_44110# a_11967_42832# 0.024799f
C2418 a_n1177_44458# a_n2661_43922# 0.010791f
C2419 a_n1352_44484# a_n2661_42834# 0.002886f
C2420 a_n699_43396# a_3363_44484# 0.07346f
C2421 a_10440_44484# a_5891_43370# 0.001688f
C2422 a_n2293_42834# a_n2065_43946# 9.75e-19
C2423 a_18479_45785# a_19319_43548# 0.102555f
C2424 a_11691_44458# a_17517_44484# 0.058911f
C2425 a_8975_43940# a_7640_43914# 1.34e-20
C2426 a_8103_44636# a_9313_44734# 1.28e-19
C2427 a_7499_43078# a_6809_43396# 1.07e-19
C2428 a_11827_44484# a_16241_44484# 6.75e-19
C2429 a_3232_43370# a_10729_43914# 0.090148f
C2430 a_11551_42558# a_n357_42282# 1.33e-19
C2431 a_5742_30871# a_n755_45592# 5.83e-20
C2432 a_17303_42282# a_13259_45724# 0.460497f
C2433 a_15765_45572# VDD 0.249471f
C2434 a_20820_30879# C6_N_btm 0.001067f
C2435 a_5534_30871# EN_VIN_BSTR_N 0.007335f
C2436 a_9482_43914# a_11415_45002# 0.309633f
C2437 a_13017_45260# a_12741_44636# 9.29e-21
C2438 a_3537_45260# a_1823_45246# 0.482502f
C2439 a_2382_45260# a_2698_46116# 4.99e-21
C2440 a_17023_45118# a_3090_45724# 1.26e-20
C2441 a_12553_44484# a_12549_44172# 4.66e-19
C2442 a_15037_45618# a_8049_45260# 0.001405f
C2443 a_2711_45572# a_2277_45546# 0.01233f
C2444 a_1990_45572# a_1848_45724# 0.007833f
C2445 a_11064_45572# a_10586_45546# 6.98e-19
C2446 a_3357_43084# a_12005_46116# 8.11e-21
C2447 a_2437_43646# a_13759_46122# 5.19e-20
C2448 a_n2017_45002# a_8199_44636# 0.020035f
C2449 a_n913_45002# a_8016_46348# 1.22e-20
C2450 a_22315_44484# a_13507_46334# 1.46e-19
C2451 a_3499_42826# a_584_46384# 0.036739f
C2452 a_1755_42282# a_5267_42460# 2.48e-19
C2453 a_1606_42308# a_5379_42460# 9.76e-20
C2454 a_17538_32519# a_22521_40599# 4.64e-21
C2455 a_3080_42308# VDAC_Ni 6.28e-19
C2456 a_5807_45002# a_9863_46634# 0.009219f
C2457 a_n1925_46634# a_5167_46660# 0.008646f
C2458 a_n743_46660# a_4817_46660# 7.71e-20
C2459 a_n2661_46098# a_2443_46660# 0.063999f
C2460 a_1799_45572# a_2609_46660# 9.48e-20
C2461 a_8128_46384# a_8654_47026# 1.16e-19
C2462 a_11453_44696# a_17609_46634# 0.079593f
C2463 a_12465_44636# a_19466_46812# 3.79e-20
C2464 a_10227_46804# a_14035_46660# 0.035412f
C2465 a_15811_47375# a_16388_46812# 0.010369f
C2466 a_11599_46634# a_16434_46987# 8.38e-20
C2467 a_n1435_47204# a_765_45546# 0.00799f
C2468 a_n815_47178# a_n901_46420# 3.99e-19
C2469 a_n2497_47436# a_1138_42852# 0.144386f
C2470 a_n971_45724# a_n1423_46090# 5.47e-19
C2471 a_n1352_44484# a_n1352_43396# 1.58e-19
C2472 a_13720_44458# a_13565_43940# 6.18e-20
C2473 a_n699_43396# a_n2433_43396# 1.5e-20
C2474 a_n1331_43914# a_n984_44318# 0.051162f
C2475 a_10193_42453# a_18504_43218# 0.003216f
C2476 a_n1899_43946# a_175_44278# 6.25e-20
C2477 a_5111_44636# a_4361_42308# 0.009091f
C2478 a_n967_45348# a_n901_43156# 0.002872f
C2479 a_3357_43084# a_3935_42891# 0.025181f
C2480 en_comp a_n1076_43230# 4.2e-20
C2481 a_n2810_45028# a_n3674_39304# 0.023324f
C2482 a_n913_45002# a_n1736_43218# 7.53e-21
C2483 a_n2017_45002# a_n1379_43218# 2.45e-19
C2484 a_n4064_37440# VDD 1.65981f
C2485 a_n2433_44484# VDD 0.40658f
C2486 a_7174_31319# a_n923_35174# 0.007133f
C2487 a_22465_38105# a_22609_38406# 0.20695f
C2488 a_13258_32519# a_11530_34132# 0.002091f
C2489 a_4958_30871# C3_P_btm 1.05e-19
C2490 a_13887_32519# w_11334_34010# 3.17e-19
C2491 a_13857_44734# a_3483_46348# 0.005876f
C2492 a_20159_44458# a_11415_45002# 5.37e-19
C2493 a_19006_44850# a_12741_44636# 0.001054f
C2494 a_1756_43548# a_768_44030# 0.093469f
C2495 a_17737_43940# a_6755_46942# 5.46e-19
C2496 a_9145_43396# a_10227_46804# 0.066362f
C2497 a_2982_43646# a_n1613_43370# 8.34e-20
C2498 a_18989_43940# a_18985_46122# 5.94e-20
C2499 a_9313_44734# a_8953_45546# 3.9e-19
C2500 a_18114_32519# a_8049_45260# 5.83e-20
C2501 a_n2661_43370# a_n2956_38216# 0.028301f
C2502 a_5343_44458# a_n1925_42282# 5.11e-21
C2503 a_n2293_42834# a_n755_45592# 0.059468f
C2504 a_19778_44110# a_13259_45724# 1.81e-20
C2505 a_18315_45260# a_16375_45002# 4.03e-21
C2506 a_n2661_44458# a_8034_45724# 7.74e-21
C2507 a_n2302_40160# a_n2302_39866# 0.050477f
C2508 a_n4209_39590# a_n3420_39616# 0.234699f
C2509 a_4958_30871# a_n4064_38528# 0.030901f
C2510 a_n4334_39616# a_n3690_39616# 8.67e-19
C2511 a_4883_46098# a_20850_46155# 3.81e-19
C2512 a_11309_47204# a_10586_45546# 1.36e-19
C2513 a_5257_43370# a_6165_46155# 0.11382f
C2514 a_n1925_46634# a_518_46482# 5.09e-19
C2515 a_171_46873# a_n1545_46494# 1.06e-20
C2516 a_n2956_39768# a_n1925_42282# 7.32e-20
C2517 a_n2661_46634# a_526_44458# 9.72e-20
C2518 a_19466_46812# a_20528_46660# 9.92e-21
C2519 a_13885_46660# a_765_45546# 1.88e-20
C2520 a_13059_46348# a_16388_46812# 8.68e-20
C2521 a_17609_46634# a_17639_46660# 0.094289f
C2522 a_12816_46660# a_11415_45002# 5.41e-22
C2523 a_13720_44458# a_5534_30871# 6.17e-22
C2524 a_626_44172# a_564_42282# 2.14e-19
C2525 a_1307_43914# a_1184_42692# 2.31e-21
C2526 a_14021_43940# a_19319_43548# 0.026713f
C2527 a_n2293_43922# a_n1853_43023# 0.001113f
C2528 a_n356_44636# a_9127_43156# 1.19e-19
C2529 a_3422_30871# a_16137_43396# 2.61e-20
C2530 a_n2661_42282# a_3626_43646# 0.02843f
C2531 a_n2661_42834# a_n1423_42826# 7.48e-19
C2532 a_3537_45260# a_5934_30871# 9.2e-20
C2533 a_5111_44636# a_6761_42308# 2.87e-20
C2534 a_n1059_45260# a_12563_42308# 5.81e-20
C2535 a_n2017_45002# a_13070_42354# 0.002239f
C2536 en_comp a_10723_42308# 8.68e-21
C2537 a_3065_45002# a_3905_42308# 0.001599f
C2538 a_n913_45002# a_11633_42558# 1.3e-20
C2539 a_19328_44172# VDD 0.263964f
C2540 a_8696_44636# a_17478_45572# 0.185985f
C2541 a_2711_45572# a_3429_45260# 9.02e-20
C2542 a_1568_43370# a_1138_42852# 9.74e-20
C2543 a_19268_43646# a_3090_45724# 0.003095f
C2544 a_16759_43396# a_15227_44166# 8.01e-19
C2545 a_453_43940# a_n1099_45572# 2.55e-20
C2546 a_10807_43548# a_10586_45546# 1.23e-21
C2547 a_1467_44172# a_n357_42282# 0.002404f
C2548 a_895_43940# a_n863_45724# 0.015488f
C2549 a_3905_42865# a_n2661_45546# 0.001705f
C2550 a_1115_44172# a_n755_45592# 2.69e-21
C2551 a_20836_43172# a_16327_47482# 0.001598f
C2552 a_1184_42692# a_n443_46116# 3.57e-21
C2553 a_3318_42354# a_584_46384# 1.04e-20
C2554 a_3147_46376# VDD 0.341038f
C2555 C5_N_btm C9_N_btm 0.150576f
C2556 C4_N_btm C10_N_btm 0.703336f
C2557 C6_N_btm C8_N_btm 0.163943f
C2558 a_22465_38105# a_22521_40599# 0.132396f
C2559 a_765_45546# a_380_45546# 0.141908f
C2560 a_22000_46634# a_20692_30879# 4.17e-19
C2561 a_5068_46348# a_5066_45546# 0.04842f
C2562 a_8199_44636# a_526_44458# 0.019697f
C2563 a_5204_45822# a_5210_46482# 6.82e-19
C2564 a_17957_46116# a_18819_46122# 4.51e-21
C2565 a_13925_46122# a_10809_44734# 6.72e-20
C2566 a_18189_46348# a_18985_46122# 3.95e-21
C2567 a_n3565_38216# a_n4064_37984# 0.342209f
C2568 a_n4209_38216# a_n4251_38304# 0.00226f
C2569 a_n2129_43609# a_n3674_39304# 4.16e-19
C2570 a_n2433_43396# a_n4318_38680# 0.001035f
C2571 a_n1177_43370# a_n1641_43230# 0.003712f
C2572 a_n97_42460# a_n1853_43023# 0.151542f
C2573 a_15095_43370# a_14955_43396# 0.130374f
C2574 a_14358_43442# a_10341_43396# 0.00838f
C2575 a_8685_43396# a_15681_43442# 0.002304f
C2576 a_15493_43940# a_21195_42852# 2.39e-21
C2577 a_9165_43940# a_9127_43156# 8.16e-20
C2578 a_3626_43646# a_16823_43084# 1.31e-20
C2579 a_n1557_42282# a_743_42282# 2.06e-19
C2580 a_9313_44734# a_14456_42282# 6.48e-20
C2581 a_n356_44636# a_17124_42282# 0.025455f
C2582 a_3422_30871# a_n784_42308# 0.022792f
C2583 a_n2840_43914# a_n3674_38680# 0.001131f
C2584 a_4235_43370# a_4361_42308# 0.006227f
C2585 a_11341_43940# a_22165_42308# 0.003146f
C2586 a_22731_47423# EN_OFFSET_CAL 1.57e-20
C2587 a_n310_47570# DATA[0] 6.14e-19
C2588 a_20749_43396# VDD 7.57e-19
C2589 a_20273_45572# a_19778_44110# 3.15e-20
C2590 a_3775_45552# a_n2661_42834# 3.12e-21
C2591 a_19256_45572# a_11691_44458# 0.001053f
C2592 a_20107_45572# a_18184_42460# 0.001559f
C2593 a_13159_45002# a_9482_43914# 0.020865f
C2594 a_13017_45260# a_13556_45296# 0.049621f
C2595 a_10053_45546# a_5891_43370# 3.54e-20
C2596 a_n2840_45002# a_n2661_43370# 0.005868f
C2597 a_3232_43370# a_1423_45028# 0.396815f
C2598 a_4649_43172# a_1823_45246# 3.11e-19
C2599 a_n4315_30879# a_n2956_39768# 0.056491f
C2600 a_8317_43396# a_n443_42852# 0.00203f
C2601 a_2711_45572# a_6755_46942# 0.612305f
C2602 a_16020_45572# a_13747_46662# 0.016423f
C2603 a_16223_45938# a_13661_43548# 3.77e-20
C2604 a_2437_43646# a_22731_47423# 3.67e-19
C2605 a_3357_43084# a_21811_47423# 9.16e-21
C2606 a_413_45260# a_14311_47204# 8.86e-20
C2607 a_n1059_45260# a_10227_46804# 0.036978f
C2608 en_comp a_16327_47482# 3.13e-20
C2609 a_6431_45366# a_6151_47436# 8.2e-20
C2610 a_6171_45002# a_6545_47178# 3.78e-20
C2611 a_375_42282# a_n746_45260# 0.41439f
C2612 a_7705_45326# a_4791_45118# 9.46e-20
C2613 a_n452_45724# a_n443_42852# 0.005182f
C2614 a_3218_45724# a_3316_45546# 0.162813f
C2615 a_n863_45724# a_1609_45822# 0.117311f
C2616 a_n1099_45572# a_n906_45572# 0.001923f
C2617 a_380_45546# a_509_45822# 0.062574f
C2618 a_n755_45592# a_n310_45899# 6.91e-19
C2619 a_n2661_45546# a_n89_45572# 4.62e-19
C2620 a_4905_42826# a_5932_42308# 0.058059f
C2621 a_n1423_42826# a_n2293_42282# 3.12e-20
C2622 a_10835_43094# a_10796_42968# 0.671797f
C2623 a_10518_42984# a_10991_42826# 7.99e-20
C2624 a_16547_43609# a_16877_43172# 9.85e-19
C2625 a_16137_43396# a_18504_43218# 0.002301f
C2626 a_2982_43646# a_3905_42558# 4.96e-19
C2627 a_20885_46660# SINGLE_ENDED 2.32e-21
C2628 a_20202_43084# RST_Z 7.21e-20
C2629 a_8685_42308# VDD 0.286875f
C2630 a_584_46384# a_n1151_42308# 0.047349f
C2631 a_2553_47502# a_2905_45572# 8.68e-19
C2632 a_2063_45854# a_3160_47472# 0.005303f
C2633 a_18114_32519# a_22469_40625# 9.95e-21
C2634 a_19721_31679# a_22521_40599# 1.69e-20
C2635 a_n237_47217# a_4915_47217# 0.071869f
C2636 a_n1741_47186# a_7227_47204# 0.016018f
C2637 a_n971_45724# a_5815_47464# 7.7e-19
C2638 a_n1177_44458# a_n452_44636# 0.011059f
C2639 a_n2661_44458# a_4743_44484# 0.006148f
C2640 a_9482_43914# a_11967_42832# 3.07e-21
C2641 a_11691_44458# a_13720_44458# 0.029855f
C2642 a_11827_44484# a_16979_44734# 0.012885f
C2643 a_19778_44110# a_18989_43940# 6.83e-20
C2644 a_n913_45002# a_1414_42308# 0.021774f
C2645 a_n1059_45260# a_453_43940# 2.04e-20
C2646 a_n967_45348# a_n984_44318# 0.00756f
C2647 a_n2293_45010# a_895_43940# 0.283316f
C2648 a_n2661_45010# a_2889_44172# 1.48e-20
C2649 a_3357_43084# a_6453_43914# 4.6e-20
C2650 COMP_P a_n2956_38216# 1.9e-21
C2651 a_6194_45824# VDD 0.274689f
C2652 a_4190_30871# EN_VIN_BSTR_N 0.043599f
C2653 a_20107_45572# a_12741_44636# 0.029025f
C2654 a_13159_45002# a_12816_46660# 3.88e-19
C2655 a_21363_45546# a_20202_43084# 0.029873f
C2656 a_20623_45572# a_11415_45002# 0.006621f
C2657 a_13348_45260# a_12991_46634# 7.26e-22
C2658 a_9838_44484# a_768_44030# 0.00219f
C2659 a_n4318_40392# a_n2956_39768# 0.023582f
C2660 a_11064_45572# a_11189_46129# 7.76e-20
C2661 a_11136_45572# a_9290_44172# 0.008811f
C2662 a_11962_45724# a_10809_44734# 0.033571f
C2663 a_11823_42460# a_6945_45028# 9.85e-22
C2664 a_n1059_45260# a_17339_46660# 2.95e-19
C2665 a_2711_45572# a_8049_45260# 2.31131f
C2666 a_15567_42826# a_15959_42545# 8.04e-19
C2667 a_16414_43172# a_15803_42450# 1.98e-19
C2668 a_n4318_38680# a_n4064_40160# 0.079598f
C2669 a_5342_30871# a_15890_42674# 0.001531f
C2670 a_4883_46098# a_4646_46812# 0.028054f
C2671 a_4915_47217# a_8270_45546# 1.62e-19
C2672 a_9313_45822# a_6755_46942# 0.031706f
C2673 a_6491_46660# a_6682_46660# 2.88e-19
C2674 a_6151_47436# a_8654_47026# 7.05e-19
C2675 a_6545_47178# a_6903_46660# 5.61e-19
C2676 a_n1151_42308# a_11901_46660# 0.020194f
C2677 a_n1741_47186# a_12156_46660# 0.005703f
C2678 a_n881_46662# a_948_46660# 0.002487f
C2679 a_n1613_43370# a_2107_46812# 0.05377f
C2680 a_2747_46873# a_2609_46660# 0.347674f
C2681 a_11309_47204# a_n743_46660# 0.001744f
C2682 a_5807_45002# a_20916_46384# 3.09e-20
C2683 a_11967_42832# a_20159_44458# 0.056889f
C2684 a_19006_44850# a_20362_44736# 3.32e-21
C2685 a_n2661_43922# a_n1331_43914# 0.002577f
C2686 a_6109_44484# a_5663_43940# 1.88e-19
C2687 a_n2293_43922# a_n1899_43946# 0.013114f
C2688 a_n2661_42834# a_n1549_44318# 0.011433f
C2689 a_626_44172# a_n1557_42282# 0.003837f
C2690 a_8975_43940# a_10729_43914# 2.43e-19
C2691 a_n2293_42834# a_n2129_43609# 0.017516f
C2692 a_11823_42460# a_12895_43230# 0.0142f
C2693 a_10057_43914# a_10949_43914# 5.37e-19
C2694 a_18479_45785# a_19095_43396# 0.001675f
C2695 a_8191_45002# a_8147_43396# 1.42e-20
C2696 a_n913_45002# a_12281_43396# 0.28203f
C2697 a_n1059_45260# a_8873_43396# 6.35e-19
C2698 a_3537_45260# a_7221_43396# 9.66e-20
C2699 a_5932_42308# a_n923_35174# 0.006295f
C2700 a_n784_42308# VREF_GND 0.068593f
C2701 a_4223_44672# a_3483_46348# 4.16e-19
C2702 a_18374_44850# a_12741_44636# 0.002579f
C2703 a_17517_44484# a_15227_44166# 0.104904f
C2704 a_11341_43940# a_13661_43548# 0.15891f
C2705 a_20623_43914# a_19321_45002# 0.294126f
C2706 a_21115_43940# a_13747_46662# 0.02491f
C2707 a_5663_43940# a_4646_46812# 2.23e-19
C2708 a_13565_44260# a_12891_46348# 9.26e-19
C2709 a_n2661_42834# a_13059_46348# 2.13e-21
C2710 a_12710_44260# a_12549_44172# 7.8e-19
C2711 a_12603_44260# a_768_44030# 0.00112f
C2712 a_9482_43914# a_13259_45724# 0.321549f
C2713 a_5093_45028# a_5066_45546# 5.33e-19
C2714 a_413_45260# a_n755_45592# 0.032345f
C2715 a_327_44734# a_n357_42282# 0.078335f
C2716 a_1667_45002# a_310_45028# 6.44e-21
C2717 a_5147_45002# a_n2661_45546# 6.41e-20
C2718 a_3065_45002# a_n863_45724# 2.64e-21
C2719 a_3537_45260# a_n2293_45546# 8.32e-21
C2720 a_16922_45042# a_19900_46494# 3.54e-21
C2721 a_11827_44484# a_14275_46494# 2.75e-21
C2722 a_n2661_44458# a_8016_46348# 0.030129f
C2723 a_19778_44110# a_18189_46348# 1.37e-20
C2724 a_14401_32519# a_18597_46090# 3e-20
C2725 a_2896_43646# a_n443_46116# 0.039985f
C2726 a_2982_43646# a_4791_45118# 0.002472f
C2727 a_15803_42450# a_7174_31319# 9.34e-20
C2728 a_5934_30871# a_1343_38525# 1.69e-19
C2729 a_16269_42308# a_4958_30871# 0.001757f
C2730 a_12861_44030# VDD 3.56689f
C2731 a_n2293_46634# a_1823_45246# 0.230429f
C2732 a_n2661_46634# a_2521_46116# 4.54e-20
C2733 a_n1925_46634# a_1208_46090# 0.005309f
C2734 a_n743_46660# a_472_46348# 0.076758f
C2735 a_2107_46812# a_n2293_46098# 1.3e-19
C2736 a_171_46873# a_n901_46420# 2.27e-19
C2737 a_12251_46660# a_12816_46660# 7.99e-20
C2738 a_5807_45002# a_6165_46155# 0.039202f
C2739 a_12891_46348# a_9290_44172# 1.02e-19
C2740 a_11309_47204# a_11189_46129# 0.03753f
C2741 a_n881_46662# a_13925_46122# 0.019683f
C2742 a_11453_44696# a_22223_46124# 1.39e-21
C2743 SMPL_ON_N a_10809_44734# 0.002895f
C2744 a_4915_47217# a_12638_46436# 2.75e-20
C2745 a_9313_45822# a_8049_45260# 0.086184f
C2746 a_n2497_47436# a_n2956_38216# 8.23e-20
C2747 a_n2109_47186# a_n2661_45546# 4.99e-20
C2748 a_17767_44458# a_16823_43084# 7.97e-22
C2749 a_n2065_43946# a_n2012_43396# 8.21e-20
C2750 a_n809_44244# a_n1177_43370# 0.002467f
C2751 a_n1549_44318# a_n1352_43396# 2.22e-19
C2752 a_14815_43914# a_9145_43396# 2.41e-19
C2753 a_15493_43396# a_15493_43940# 0.188034f
C2754 a_19862_44208# a_11341_43940# 0.07932f
C2755 a_1307_43914# a_5193_42852# 2.47e-20
C2756 a_10193_42453# a_7174_31319# 0.020527f
C2757 a_12429_44172# a_12710_44260# 0.008628f
C2758 a_3422_30871# a_3080_42308# 0.022126f
C2759 a_14539_43914# a_17678_43396# 1.74e-19
C2760 a_n2017_45002# a_n4318_38216# 7.46e-19
C2761 a_n2840_43914# VDD 0.304745f
C2762 a_10193_42453# a_10306_45572# 0.002653f
C2763 a_8746_45002# a_10216_45572# 0.001575f
C2764 a_2711_45572# a_14127_45572# 0.001525f
C2765 C7_N_btm C3_P_btm 3.05e-19
C2766 C6_N_btm C2_P_btm 7.09e-20
C2767 a_15493_43940# a_3483_46348# 0.026486f
C2768 a_11341_43940# a_4185_45028# 1.23e-19
C2769 a_7871_42858# a_n1613_43370# 0.659491f
C2770 a_11750_44172# a_9290_44172# 0.001116f
C2771 a_10405_44172# a_10903_43370# 0.026421f
C2772 a_22485_44484# a_8049_45260# 2.49e-20
C2773 a_2127_44172# a_526_44458# 0.001334f
C2774 a_n2661_42834# a_3218_45724# 1.7e-20
C2775 a_14180_46812# VDD 0.755623f
C2776 a_4958_30871# a_7754_40130# 5.49e-20
C2777 a_4704_46090# a_5164_46348# 5.86e-19
C2778 a_4419_46090# a_5204_45822# 0.001858f
C2779 a_11415_45002# a_18819_46122# 1.5e-20
C2780 a_12741_44636# a_17715_44484# 0.029877f
C2781 a_3483_46348# a_6419_46155# 2.02e-21
C2782 a_12816_46660# a_13259_45724# 1.31e-19
C2783 a_765_45546# a_526_44458# 5.75e-20
C2784 a_n97_42460# a_14358_43442# 1.05e-20
C2785 a_2982_43646# a_8791_43396# 1.3e-21
C2786 a_n356_44636# a_1755_42282# 0.00959f
C2787 a_5883_43914# a_7963_42308# 1.91e-21
C2788 a_14021_43940# a_19095_43396# 1.04e-19
C2789 a_11967_42832# a_11301_43218# 8.99e-21
C2790 a_5343_44458# a_8337_42558# 9.56e-19
C2791 a_1239_47204# DATA[0] 2.02e-19
C2792 a_1209_47178# DATA[1] 0.076054f
C2793 a_9803_43646# VDD 0.261557f
C2794 a_11823_42460# a_11827_44484# 0.024482f
C2795 a_5263_45724# a_5343_44458# 1.81e-20
C2796 a_2711_45572# a_8103_44636# 5.76e-21
C2797 a_11525_45546# a_11691_44458# 4.12e-20
C2798 a_10193_42453# a_16981_45144# 0.001232f
C2799 a_n2017_45002# a_2382_45260# 0.032443f
C2800 a_3357_43084# a_6171_45002# 0.003278f
C2801 a_n967_45348# a_n467_45028# 0.005391f
C2802 a_5934_30871# a_n2293_46634# 2.22e-19
C2803 a_16877_42852# a_6755_46942# 1.98e-19
C2804 a_6123_31319# a_n2312_38680# 4.19e-21
C2805 a_9306_43218# a_3090_45724# 2.03e-20
C2806 a_458_43396# a_n863_45724# 0.122956f
C2807 a_4093_43548# a_n2661_45546# 0.343267f
C2808 a_4361_42308# a_9290_44172# 0.1126f
C2809 a_21335_42336# a_13507_46334# 2.39e-19
C2810 a_310_45028# VDD 0.360949f
C2811 a_4099_45572# a_n2661_46634# 2.95e-20
C2812 a_7499_43078# a_12549_44172# 1.93e-19
C2813 a_1609_45572# a_n2293_46634# 1.5e-19
C2814 a_16020_45572# a_11599_46634# 2.63e-20
C2815 a_16855_45546# a_16327_47482# 0.305145f
C2816 a_15599_45572# a_10227_46804# 0.001084f
C2817 a_10216_45572# a_4883_46098# 5.19e-19
C2818 a_526_44458# a_509_45822# 1.55e-20
C2819 a_13483_43940# a_13657_42558# 8.24e-21
C2820 a_n1991_42858# a_n1641_43230# 0.229804f
C2821 a_n2840_42826# a_n3674_39304# 0.16082f
C2822 a_n2157_42858# a_n1076_43230# 0.102325f
C2823 a_n1853_43023# a_n901_43156# 0.081949f
C2824 a_16137_43396# a_16414_43172# 0.179708f
C2825 a_743_42282# a_3935_42891# 1.46e-20
C2826 a_16547_43609# a_5342_30871# 1.72e-20
C2827 a_10341_43396# a_22165_42308# 3.24e-19
C2828 a_n4318_39304# a_n3674_38680# 0.031218f
C2829 a_3754_39964# VDAC_Pi 0.296508f
C2830 a_20273_45572# a_20159_44458# 1.49e-21
C2831 a_10193_42453# a_10729_43914# 0.010339f
C2832 a_20107_45572# a_20362_44736# 1.08e-21
C2833 a_1307_43914# a_16112_44458# 0.012033f
C2834 a_18587_45118# a_18911_45144# 0.010993f
C2835 a_1423_45028# a_8975_43940# 0.331942f
C2836 a_7499_43078# a_12429_44172# 0.001488f
C2837 a_8746_45002# a_10405_44172# 1.94e-20
C2838 a_20623_45572# a_11967_42832# 7.43e-21
C2839 a_3232_43370# a_6109_44484# 0.072011f
C2840 a_5111_44636# a_5891_43370# 0.702087f
C2841 en_comp a_n2293_43922# 0.412872f
C2842 a_n1059_45260# a_14815_43914# 2.69e-20
C2843 a_5205_44484# a_5205_44734# 0.015405f
C2844 a_n967_45348# a_n2661_43922# 0.024232f
C2845 a_2437_43646# a_17517_44484# 3.17e-20
C2846 a_17303_42282# a_20202_43084# 0.00102f
C2847 a_10723_42308# a_4185_45028# 1.64e-19
C2848 a_8515_42308# a_8953_45546# 6.71e-19
C2849 a_n1630_35242# a_n2956_39304# 0.001241f
C2850 a_2987_42968# a_n863_45724# 0.002594f
C2851 a_n2472_42282# a_n1925_42282# 2.81e-19
C2852 a_133_42852# a_n357_42282# 0.011275f
C2853 a_3080_42308# VREF_GND 0.001083f
C2854 a_14495_45572# a_12741_44636# 3.7e-20
C2855 a_8696_44636# a_16388_46812# 2.13e-19
C2856 a_n2661_43370# a_768_44030# 0.024666f
C2857 a_626_44172# a_33_46660# 1.58e-20
C2858 a_19431_45546# a_19333_46634# 4.38e-20
C2859 a_19256_45572# a_15227_44166# 2.59e-20
C2860 a_18691_45572# a_19466_46812# 2.36e-19
C2861 a_15861_45028# a_13059_46348# 2.15e-21
C2862 a_3232_43370# a_4646_46812# 0.305673f
C2863 a_5111_44636# a_4817_46660# 2.19e-22
C2864 a_5691_45260# a_4651_46660# 1.21e-20
C2865 a_4927_45028# a_4955_46873# 7.8e-21
C2866 a_6171_45002# a_3877_44458# 1.79e-21
C2867 a_5147_45002# a_5385_46902# 9.06e-21
C2868 a_2711_45572# a_8953_45546# 0.032277f
C2869 a_6472_45840# a_6419_46155# 6.52e-19
C2870 a_15004_44636# a_4915_47217# 0.008914f
C2871 a_18525_43370# a_18214_42558# 8.42e-21
C2872 a_15743_43084# a_18907_42674# 1.64e-20
C2873 a_5755_42852# a_4921_42308# 0.002018f
C2874 a_4361_42308# a_15051_42282# 0.016131f
C2875 a_743_42282# a_15890_42674# 0.010042f
C2876 a_16137_43396# a_7174_31319# 2.14e-20
C2877 a_5534_30871# a_n1630_35242# 0.033914f
C2878 a_2747_46873# a_3094_47570# 2.88e-19
C2879 a_4883_46098# a_9804_47204# 0.020011f
C2880 a_16327_47482# a_13661_43548# 0.132061f
C2881 a_16023_47582# a_5807_45002# 0.00104f
C2882 a_10227_46804# a_16285_47570# 0.002099f
C2883 a_6575_47204# a_n1925_46634# 3.37e-19
C2884 a_n1435_47204# a_n2956_39768# 1.18e-19
C2885 a_n2109_47186# a_5385_46902# 0.013334f
C2886 a_n1741_47186# a_4955_46873# 2.85e-19
C2887 a_2063_45854# a_2609_46660# 0.005947f
C2888 a_2905_45572# a_1799_45572# 0.002025f
C2889 a_2553_47502# a_2443_46660# 0.001147f
C2890 a_4791_45118# a_2107_46812# 0.078338f
C2891 a_584_46384# a_3177_46902# 9.68e-20
C2892 a_n1177_44458# a_n809_44244# 0.00369f
C2893 a_18989_43940# a_20159_44458# 1.23e-19
C2894 a_18287_44626# a_20679_44626# 5.48e-21
C2895 a_n2661_44458# a_1414_42308# 6.41e-20
C2896 a_n1352_44484# a_n1549_44318# 3.11e-20
C2897 a_8696_44636# a_14955_43396# 2.57e-23
C2898 a_9159_44484# a_n2661_43922# 0.004106f
C2899 a_1307_43914# a_1443_43940# 0.042476f
C2900 a_8953_45002# a_9801_43940# 4.55e-20
C2901 a_n2293_45010# a_458_43396# 1.65e-19
C2902 a_n2661_45010# a_1049_43396# 1.29e-21
C2903 en_comp a_n97_42460# 5.85e-20
C2904 a_n2017_45002# a_n1655_43396# 4.3e-19
C2905 a_n4209_39304# a_n2956_38216# 0.020992f
C2906 a_n913_45002# VDD 9.190901f
C2907 a_22400_42852# a_22459_39145# 0.242947f
C2908 a_1443_43940# a_n443_46116# 2.66e-19
C2909 a_14401_32519# w_11334_34010# 0.023412f
C2910 a_n2661_43370# a_1176_45822# 4.9e-20
C2911 a_18911_45144# a_11415_45002# 0.006861f
C2912 a_17719_45144# a_12741_44636# 0.011019f
C2913 a_n2293_42834# a_3483_46348# 0.033766f
C2914 a_19778_44110# a_20202_43084# 2.92e-20
C2915 a_18248_44752# a_3090_45724# 0.027743f
C2916 a_2998_44172# a_768_44030# 0.571981f
C2917 a_22959_43948# a_12861_44030# 1.04e-19
C2918 a_19862_44208# a_16327_47482# 0.209324f
C2919 a_n2661_42282# a_n2312_40392# 3.67e-19
C2920 a_n3674_39768# a_n1613_43370# 5.31e-19
C2921 a_5009_45028# a_5164_46348# 4.03e-19
C2922 a_14537_43396# a_2324_44458# 0.341957f
C2923 a_2382_45260# a_526_44458# 0.072916f
C2924 a_n784_42308# a_7174_31319# 1.93626f
C2925 a_8791_42308# a_5742_30871# 4.57e-20
C2926 a_n3674_38680# a_n4334_40480# 1.51e-19
C2927 a_n83_35174# VIN_P 0.001664f
C2928 C4_P_btm C2_P_btm 7.72909f
C2929 a_16327_47482# a_4185_45028# 1.37e-19
C2930 a_4915_47217# a_13759_46122# 0.024639f
C2931 a_9313_45822# a_8953_45546# 0.038855f
C2932 a_13759_47204# a_765_45546# 5.9e-19
C2933 a_12549_44172# a_20411_46873# 1.31e-20
C2934 a_5807_45002# a_16751_46987# 0.001109f
C2935 a_7715_46873# a_7927_46660# 3.12e-19
C2936 a_5385_46902# a_5841_46660# 4.2e-19
C2937 a_3877_44458# a_6903_46660# 0.007019f
C2938 a_5732_46660# a_6969_46634# 3.02e-20
C2939 a_6540_46812# a_6755_46942# 0.057503f
C2940 a_7577_46660# a_8145_46902# 0.170059f
C2941 a_7411_46660# a_8667_46634# 0.043475f
C2942 a_5883_43914# a_8685_43396# 3.79e-19
C2943 a_3422_30871# a_14021_43940# 0.018792f
C2944 a_n2661_43922# a_n1917_43396# 1.76e-20
C2945 a_n2661_42834# a_n1177_43370# 8.78e-19
C2946 a_11827_44484# a_18429_43548# 4.78e-21
C2947 a_18494_42460# a_19700_43370# 3.28e-20
C2948 a_n2293_42834# a_n2840_42826# 9.62e-19
C2949 a_1423_45028# a_2905_42968# 6.76e-22
C2950 a_7845_44172# a_8018_44260# 0.007688f
C2951 a_7542_44172# a_8333_44056# 7.67e-20
C2952 a_11691_44458# a_16977_43638# 3.52e-19
C2953 a_16237_45028# a_16547_43609# 3.95e-21
C2954 a_n913_45002# a_873_42968# 7.48e-19
C2955 a_556_44484# VDD 0.004463f
C2956 a_n3420_39072# VCM 0.007907f
C2957 a_2711_45572# a_6812_45938# 0.003338f
C2958 a_2675_43914# a_1823_45246# 8.17e-19
C2959 a_10341_43396# a_13661_43548# 0.053085f
C2960 a_18326_43940# a_17339_46660# 0.006409f
C2961 a_4905_42826# a_4646_46812# 5.08e-20
C2962 a_15781_43660# a_12549_44172# 0.062935f
C2963 a_7221_43396# a_n2293_46634# 1.49e-19
C2964 a_742_44458# a_1848_45724# 1.5e-20
C2965 a_949_44458# a_997_45618# 5.82e-20
C2966 a_2779_44458# a_n755_45592# 1.49e-20
C2967 a_n699_43396# a_310_45028# 9.49e-22
C2968 a_4223_44672# a_n357_42282# 7.15e-20
C2969 a_11967_42832# a_18819_46122# 5.34e-22
C2970 a_19095_43396# a_13507_46334# 3.23e-19
C2971 a_10991_42826# a_2063_45854# 8.1e-19
C2972 a_7871_42858# a_4791_45118# 2.66e-21
C2973 en_comp a_22780_40081# 4.3e-20
C2974 a_n4209_38502# a_n4251_38528# 0.00226f
C2975 a_n2946_38778# a_n2302_38778# 6.68e-19
C2976 a_n3420_38528# a_n2860_38778# 0.002301f
C2977 a_5894_47026# VDD 4.6e-19
C2978 a_4958_30871# C6_N_btm 0.005441f
C2979 a_n3674_38216# a_n4334_37440# 6.7e-20
C2980 COMP_P a_7754_38470# 1.8e-19
C2981 a_11415_45002# a_22591_46660# 0.172844f
C2982 a_20202_43084# a_20820_30879# 0.005846f
C2983 a_765_45546# a_2521_46116# 3.87e-20
C2984 a_22365_46825# a_12741_44636# 0.062216f
C2985 a_n2293_46634# a_n2293_45546# 0.065405f
C2986 a_7577_46660# a_5066_45546# 1.32e-19
C2987 a_n1925_46634# a_n2661_45546# 5.29e-20
C2988 a_3090_45724# a_2324_44458# 0.684819f
C2989 a_15368_46634# a_15015_46420# 0.012546f
C2990 a_14976_45028# a_14840_46494# 0.010576f
C2991 a_n1899_43946# a_n901_43156# 0.001167f
C2992 a_n984_44318# a_n1853_43023# 1.28e-20
C2993 a_19862_44208# a_10341_43396# 0.028065f
C2994 a_n1177_43370# a_n1352_43396# 0.233657f
C2995 a_n2129_43609# a_n2012_43396# 0.183186f
C2996 a_n2433_43396# a_n1809_43762# 9.73e-19
C2997 a_n1331_43914# a_n1641_43230# 1.38e-21
C2998 a_n1761_44111# a_n1076_43230# 2.91e-19
C2999 a_3905_42865# a_4361_42308# 3.2e-19
C3000 a_11967_42832# a_10796_42968# 0.001301f
C3001 a_n4318_39304# a_n1190_43762# 3.5e-21
C3002 a_5891_43370# a_5837_43172# 4.79e-20
C3003 a_n2956_37592# a_n2946_39866# 3.12e-19
C3004 a_n4318_39304# VDD 0.643395f
C3005 a_20273_45572# a_20623_45572# 0.219856f
C3006 a_14495_45572# a_13556_45296# 1.1e-20
C3007 a_13904_45546# a_14180_45002# 1.92e-19
C3008 a_13249_42308# a_13777_45326# 2.35e-21
C3009 a_15143_45578# a_9482_43914# 7.52e-21
C3010 a_20107_45572# a_21363_45546# 0.043567f
C3011 a_10210_45822# a_8953_45002# 1.45e-19
C3012 a_9159_45572# a_6171_45002# 0.00193f
C3013 a_10341_43396# a_4185_45028# 0.019539f
C3014 a_9145_43396# a_8016_46348# 2.69e-19
C3015 a_15493_43940# a_n357_42282# 2.07e-19
C3016 a_n1557_42282# a_n2956_38680# 1.47e-20
C3017 a_8387_43230# a_3090_45724# 2.71e-20
C3018 a_13249_42308# a_n1151_42308# 2.6e-20
C3019 a_8697_45572# a_n971_45724# 2.34e-19
C3020 a_4419_46090# a_3503_45724# 3.27e-21
C3021 a_17715_44484# a_16375_45002# 0.026655f
C3022 a_17957_46116# a_18147_46436# 0.011458f
C3023 a_10809_44734# a_12638_46436# 0.003187f
C3024 a_167_45260# a_n443_42852# 0.246952f
C3025 a_1823_45246# a_2277_45546# 3.97e-20
C3026 a_5663_43940# a_6171_42473# 3.37e-21
C3027 a_n1177_43370# a_n2293_42282# 2.19e-22
C3028 a_16547_43609# a_743_42282# 1.93e-20
C3029 a_11967_42832# a_4958_30871# 0.239255f
C3030 a_18525_43370# a_16823_43084# 0.009621f
C3031 a_3457_43396# a_3681_42891# 0.001119f
C3032 a_8147_43396# a_7765_42852# 7.06e-19
C3033 a_8791_43396# a_7871_42858# 1.26e-19
C3034 a_3626_43646# a_12545_42858# 8.41e-20
C3035 a_2982_43646# a_12895_43230# 2.86e-20
C3036 a_3422_30871# a_15764_42576# 7.68e-20
C3037 a_2107_46812# DATA[3] 2.5e-21
C3038 a_20922_43172# VDD 0.192467f
C3039 a_8696_44636# a_n2661_42834# 0.004739f
C3040 a_1667_45002# a_n2661_44458# 1.72e-20
C3041 a_327_44734# a_n2433_44484# 1.63e-21
C3042 a_n1059_45260# a_4743_44484# 6.94e-22
C3043 a_n913_45002# a_n699_43396# 2.01e-19
C3044 a_6171_45002# a_16237_45028# 0.05704f
C3045 a_n2017_45002# a_5343_44458# 0.027073f
C3046 a_n467_45028# a_n1917_44484# 1.34e-20
C3047 a_n13_43084# a_n755_45592# 0.113444f
C3048 a_n967_43230# a_n863_45724# 3.46e-21
C3049 a_1709_42852# a_526_44458# 3.71e-19
C3050 a_16019_45002# a_11453_44696# 0.006638f
C3051 a_6709_45028# a_n1613_43370# 0.037165f
C3052 a_7229_43940# a_n881_46662# 0.002123f
C3053 a_6171_45002# a_8128_46384# 4.91e-20
C3054 a_n2017_45002# a_n2956_39768# 1.08e-21
C3055 a_n2661_45010# a_n2293_46634# 0.003275f
C3056 a_4574_45260# a_768_44030# 6.09e-21
C3057 a_4099_45572# a_765_45546# 1.94e-21
C3058 a_3626_43646# a_19332_42282# 0.013212f
C3059 a_13678_32519# COMP_P 2.06e-19
C3060 a_3080_42308# a_7174_31319# 0.22305f
C3061 a_4190_30871# a_n1630_35242# 0.039258f
C3062 a_743_42282# a_n3674_37592# 2.16e-19
C3063 a_10341_43396# a_9803_42558# 6.46e-20
C3064 a_10695_43548# a_5742_30871# 3.57e-19
C3065 a_12594_46348# CLK 1.08e-20
C3066 a_n4334_40480# VDD 0.390668f
C3067 a_n2497_47436# a_768_44030# 0.023758f
C3068 a_n1741_47186# a_11117_47542# 2.77e-19
C3069 a_n237_47217# a_n881_46662# 0.958566f
C3070 a_n23_47502# a_n1613_43370# 5.76e-20
C3071 a_15507_47210# a_15673_47210# 0.81159f
C3072 a_6545_47178# a_4883_46098# 0.008688f
C3073 a_11599_46634# a_16241_47178# 2.85e-20
C3074 a_14955_47212# a_16327_47482# 1.03e-19
C3075 a_2905_45572# a_2747_46873# 0.010677f
C3076 a_2124_47436# a_2266_47243# 0.005572f
C3077 a_n1435_47204# a_10227_46804# 0.004624f
C3078 a_13717_47436# a_17591_47464# 3.4e-19
C3079 a_12861_44030# a_16588_47582# 9.72e-20
C3080 a_18911_45144# a_11967_42832# 5.48e-20
C3081 a_n1917_44484# a_n2661_43922# 0.010578f
C3082 a_6298_44484# a_9313_44734# 7.5e-22
C3083 a_10334_44484# a_5891_43370# 7.17e-19
C3084 a_n1177_44458# a_n2661_42834# 0.002427f
C3085 a_16922_45042# a_20835_44721# 2.59e-21
C3086 a_1423_45028# a_5495_43940# 1.89e-20
C3087 a_n2293_42834# a_n2472_43914# 4.12e-19
C3088 a_8701_44490# a_8855_44734# 0.008678f
C3089 a_11691_44458# a_17061_44734# 0.001749f
C3090 a_7499_43078# a_6643_43396# 1.32e-19
C3091 a_11827_44484# a_15367_44484# 6.14e-19
C3092 a_3232_43370# a_10405_44172# 2.4e-20
C3093 a_5111_44636# a_10807_43548# 1.74e-20
C3094 a_4958_30871# a_13259_45724# 0.054732f
C3095 a_5742_30871# a_n357_42282# 0.001298f
C3096 a_15903_45785# VDD 0.291109f
C3097 a_20820_30879# C5_N_btm 1.83e-19
C3098 a_5534_30871# a_11530_34132# 0.010307f
C3099 a_5342_30871# EN_VIN_BSTR_P 0.010795f
C3100 a_13348_45260# a_11415_45002# 0.036052f
C3101 a_3429_45260# a_1823_45246# 0.047931f
C3102 a_16922_45042# a_3090_45724# 0.206138f
C3103 a_n2293_43922# a_13661_43548# 7.4e-20
C3104 a_413_45260# a_3483_46348# 5.51e-19
C3105 a_16501_45348# a_14976_45028# 7.45e-21
C3106 a_12189_44484# a_12549_44172# 6.62e-21
C3107 a_8696_44636# a_5066_45546# 1.84e-20
C3108 a_14033_45822# a_8049_45260# 0.004947f
C3109 a_10544_45572# a_10586_45546# 3.58e-19
C3110 a_2437_43646# a_13351_46090# 1.08e-20
C3111 a_n1059_45260# a_8016_46348# 2.52e-20
C3112 a_3357_43084# a_10903_43370# 9.87e-21
C3113 a_18245_44484# a_11453_44696# 1.9e-19
C3114 a_3422_30871# a_13507_46334# 0.074924f
C3115 a_20512_43084# a_18597_46090# 0.023158f
C3116 a_8333_44056# a_n971_45724# 0.017284f
C3117 a_2351_42308# a_2903_42308# 8.7e-20
C3118 a_1755_42282# a_3823_42558# 2.57e-19
C3119 a_1606_42308# a_5267_42460# 1.69e-20
C3120 a_n784_42308# a_5932_42308# 0.151611f
C3121 COMP_P a_6123_31319# 0.02889f
C3122 a_5807_45002# a_8492_46660# 0.005311f
C3123 a_n743_46660# a_4955_46873# 0.0023f
C3124 a_n1925_46634# a_5385_46902# 0.003429f
C3125 a_1799_45572# a_2443_46660# 1.77e-19
C3126 a_n2661_46634# a_5275_47026# 0.003477f
C3127 a_n881_46662# a_8270_45546# 9.01e-20
C3128 a_12465_44636# a_19333_46634# 2.86e-20
C3129 a_4883_46098# a_19692_46634# 0.058277f
C3130 a_11599_46634# a_16721_46634# 0.00139f
C3131 a_10227_46804# a_13885_46660# 6.78e-19
C3132 a_15507_47210# a_16388_46812# 5.7e-19
C3133 a_15811_47375# a_13059_46348# 0.001466f
C3134 a_13381_47204# a_765_45546# 0.002617f
C3135 a_n971_45724# a_n1991_46122# 0.010501f
C3136 a_n746_45260# a_n1853_46287# 3.3e-21
C3137 a_n2497_47436# a_1176_45822# 2.85e-20
C3138 a_n1352_44484# a_n1177_43370# 8.8e-22
C3139 a_n1177_44458# a_n1352_43396# 7.26e-20
C3140 a_n1899_43946# a_n984_44318# 0.118759f
C3141 a_n2065_43946# a_644_44056# 6.01e-22
C3142 a_9313_44734# a_10555_44260# 0.005264f
C3143 a_11823_42460# a_13569_43230# 7.84e-20
C3144 a_n467_45028# a_n1853_43023# 5.11e-21
C3145 a_3357_43084# a_3681_42891# 0.052403f
C3146 a_3537_45260# a_5649_42852# 0.048691f
C3147 en_comp a_n901_43156# 4.8e-21
C3148 a_n913_45002# a_n4318_38680# 4.18e-21
C3149 a_n1059_45260# a_n1736_43218# 5.17e-20
C3150 a_n2017_45002# a_n1545_43230# 6.01e-19
C3151 a_n967_45348# a_n1641_43230# 0.00611f
C3152 a_n2946_37690# VDD 0.38221f
C3153 a_n2661_44458# VDD 1.06317f
C3154 a_15761_42308# RST_Z 2.8e-20
C3155 a_22465_38105# CAL_P 0.026947f
C3156 a_7174_31319# a_n1532_35090# 1.2e-19
C3157 a_4958_30871# C4_P_btm 1.18e-19
C3158 a_n2661_43922# a_4419_46090# 4.13e-20
C3159 a_20159_44458# a_20202_43084# 1.9e-19
C3160 a_n2293_43922# a_4185_45028# 0.093999f
C3161 a_18588_44850# a_12741_44636# 0.002114f
C3162 a_n356_44636# a_2324_44458# 0.00124f
C3163 a_9313_44734# a_5937_45572# 0.006008f
C3164 a_5891_43370# a_9290_44172# 0.302383f
C3165 a_n2661_43370# a_n2472_45546# 0.002286f
C3166 a_18911_45144# a_13259_45724# 9.82e-20
C3167 a_4743_44484# a_n1925_42282# 1.27e-19
C3168 a_n2293_42834# a_n357_42282# 4.06139f
C3169 a_5343_44458# a_526_44458# 0.015378f
C3170 a_17719_45144# a_16375_45002# 0.201099f
C3171 a_1568_43370# a_768_44030# 0.077231f
C3172 a_n97_42460# a_13661_43548# 0.02781f
C3173 a_15682_43940# a_6755_46942# 0.028635f
C3174 a_11322_45546# CLK 0.003637f
C3175 a_11652_45724# DATA[5] 1.16e-19
C3176 a_n4064_40160# a_n2302_39866# 2.59e-20
C3177 a_n4209_39590# a_n3690_39616# 0.045251f
C3178 a_n2302_40160# a_n4064_39616# 2.59e-20
C3179 a_n4334_39616# a_n3565_39590# 2e-19
C3180 a_4883_46098# a_20692_30879# 9.38e-20
C3181 a_n1925_46634# a_n1533_46116# 0.001581f
C3182 a_5257_43370# a_5497_46414# 0.002158f
C3183 a_2107_46812# a_6945_45028# 0.028356f
C3184 a_15227_46910# a_16388_46812# 1e-19
C3185 a_19692_46634# a_21188_46660# 0.022017f
C3186 a_15227_44166# a_20731_47026# 1.96e-20
C3187 a_9863_46634# a_3483_46348# 3.53e-22
C3188 a_20835_44721# a_15743_43084# 1.25e-21
C3189 a_14673_44172# a_743_42282# 6.85e-21
C3190 a_n2293_43922# a_n2157_42858# 0.040551f
C3191 a_n2661_43922# a_n1853_43023# 1.11e-20
C3192 a_n2661_42834# a_n1991_42858# 8.85e-19
C3193 a_n356_44636# a_8387_43230# 1.68e-20
C3194 a_375_42282# a_n1630_35242# 0.036312f
C3195 a_3232_43370# a_6171_42473# 5.89e-23
C3196 a_3537_45260# a_7963_42308# 4.5e-20
C3197 a_n913_45002# a_11551_42558# 3.95e-19
C3198 a_n2017_45002# a_12563_42308# 0.003288f
C3199 en_comp a_10533_42308# 4.34e-21
C3200 a_18451_43940# VDD 0.172318f
C3201 a_16680_45572# a_17478_45572# 0.001111f
C3202 a_8696_44636# a_15861_45028# 0.26484f
C3203 a_16115_45572# a_16223_45938# 0.057222f
C3204 a_14033_45822# a_14127_45572# 1.26e-19
C3205 a_2711_45572# a_3065_45002# 0.012727f
C3206 a_1049_43396# a_1138_42852# 0.022078f
C3207 a_n97_42460# a_4185_45028# 0.022167f
C3208 a_16977_43638# a_15227_44166# 0.002041f
C3209 a_15743_43084# a_3090_45724# 0.005519f
C3210 a_3681_42891# a_3877_44458# 1.24e-20
C3211 a_1115_44172# a_n357_42282# 0.011627f
C3212 a_15682_43940# a_8049_45260# 6.17e-21
C3213 a_644_44056# a_n755_45592# 1.74e-20
C3214 a_2479_44172# a_n863_45724# 0.047943f
C3215 a_9165_43940# a_2324_44458# 1.24e-20
C3216 a_20573_43172# a_16327_47482# 0.001116f
C3217 a_1576_42282# a_n443_46116# 2.01e-21
C3218 a_2903_42308# a_584_46384# 1.37e-20
C3219 a_5934_30871# w_11334_34010# 2.35e-19
C3220 a_2804_46116# VDD 0.159351f
C3221 a_22465_38105# CAL_N 0.072253f
C3222 a_n4315_30879# VDAC_P 0.011363f
C3223 a_n4334_38304# a_n4064_37984# 0.410244f
C3224 a_n3565_38216# a_n2946_37984# 0.411006f
C3225 a_n4209_38216# a_n2302_37984# 0.407312f
C3226 a_2684_37794# a_2113_38308# 0.468006f
C3227 C6_N_btm C7_N_btm 26.0771f
C3228 C5_N_btm C8_N_btm 0.145019f
C3229 C3_N_btm C10_N_btm 0.321945f
C3230 C4_N_btm C9_N_btm 0.154834f
C3231 a_21188_46660# a_20692_30879# 3.94e-20
C3232 a_4704_46090# a_5066_45546# 0.002532f
C3233 a_13759_46122# a_10809_44734# 6.06e-20
C3234 a_18189_46348# a_18819_46122# 1.04e-20
C3235 a_n2433_43396# a_n3674_39304# 9.78e-19
C3236 a_n1917_43396# a_n1641_43230# 0.00125f
C3237 a_n1352_43396# a_n1991_42858# 0.00171f
C3238 a_n1177_43370# a_n1423_42826# 0.0016f
C3239 a_14205_43396# a_14955_43396# 0.157423f
C3240 a_14579_43548# a_10341_43396# 0.029139f
C3241 a_n97_42460# a_n2157_42858# 9.01e-21
C3242 a_14021_43940# a_16414_43172# 9.19e-22
C3243 a_15493_43940# a_21356_42826# 1.97e-20
C3244 a_11341_43940# a_21671_42860# 6.71e-21
C3245 a_n2293_43922# a_9803_42558# 4.58e-20
C3246 a_n4318_39304# a_n4318_38680# 0.059432f
C3247 a_10695_43548# a_10849_43646# 0.010303f
C3248 a_9145_43396# a_12281_43396# 0.032945f
C3249 a_n356_44636# a_16522_42674# 0.001524f
C3250 a_4093_43548# a_4361_42308# 1.72e-21
C3251 a_12465_44636# CLK 0.795478f
C3252 a_22223_47212# EN_OFFSET_CAL 0.011048f
C3253 a_n2312_39304# DATA[0] 0.001796f
C3254 a_17364_32525# VDD 0.511443f
C3255 a_19431_45546# a_11691_44458# 1.76e-20
C3256 a_20107_45572# a_19778_44110# 1.5e-19
C3257 a_13159_45002# a_13348_45260# 0.105274f
C3258 a_13017_45260# a_9482_43914# 0.048717f
C3259 a_9049_44484# a_5891_43370# 1.84e-20
C3260 a_5691_45260# a_1423_45028# 1.19e-19
C3261 a_n37_45144# a_117_45144# 0.008535f
C3262 a_3537_45260# a_3602_45348# 2.49e-19
C3263 a_7229_43940# a_1307_43914# 0.004598f
C3264 a_5342_30871# a_10903_43370# 2.1e-21
C3265 a_8229_43396# a_n443_42852# 2.56e-19
C3266 a_2711_45572# a_10249_46116# 9.85e-22
C3267 a_17478_45572# a_13747_46662# 0.073886f
C3268 a_18596_45572# a_n881_46662# 1.26e-20
C3269 a_2437_43646# a_22223_47212# 0.001377f
C3270 a_3357_43084# a_4883_46098# 0.060164f
C3271 a_19963_31679# a_13507_46334# 1.83e-19
C3272 a_n2017_45002# a_10227_46804# 0.030377f
C3273 a_6171_45002# a_6151_47436# 0.006279f
C3274 a_413_45260# a_13487_47204# 4.31e-19
C3275 a_9482_43914# a_2063_45854# 0.018952f
C3276 a_11787_45002# a_n1151_42308# 2.96e-21
C3277 a_375_42282# a_n971_45724# 1.02e-19
C3278 a_6709_45028# a_4791_45118# 0.017539f
C3279 a_n2293_45546# a_2277_45546# 1.67e-19
C3280 a_n863_45724# a_n443_42852# 0.556081f
C3281 a_997_45618# a_n356_45724# 2.02e-19
C3282 a_n755_45592# a_n23_45546# 0.001003f
C3283 a_n1099_45572# a_n1013_45572# 0.00411f
C3284 a_2957_45546# a_3316_45546# 0.001625f
C3285 a_n2661_45546# a_n310_45572# 1.2e-19
C3286 a_15681_43442# a_15597_42852# 1.25e-19
C3287 a_n1991_42858# a_n2293_42282# 9.15e-21
C3288 a_10518_42984# a_10796_42968# 0.118759f
C3289 a_3626_43646# a_5379_42460# 0.057009f
C3290 a_n97_42460# a_9803_42558# 0.099148f
C3291 a_3080_42308# a_5932_42308# 14.0282f
C3292 a_16547_43609# a_16328_43172# 1.96e-19
C3293 a_4905_42826# a_6171_42473# 2.44e-20
C3294 a_14021_43940# a_7174_31319# 9.94e-21
C3295 a_22365_46825# RST_Z 1.22e-19
C3296 a_n3420_37440# VDAC_P 4.18e-19
C3297 a_8325_42308# VDD 0.313956f
C3298 a_18114_32519# a_22521_40599# 1.3e-20
C3299 a_n237_47217# a_n443_46116# 0.110841f
C3300 a_2124_47436# a_n1151_42308# 0.006002f
C3301 a_2553_47502# a_2952_47436# 0.002785f
C3302 a_2063_45854# a_2905_45572# 0.037943f
C3303 a_584_46384# a_3160_47472# 2.16e-20
C3304 a_n971_45724# a_5129_47502# 3.14e-19
C3305 a_n1741_47186# a_6851_47204# 0.030234f
C3306 a_18911_45144# a_18989_43940# 0.016276f
C3307 a_n1177_44458# a_n1352_44484# 0.233657f
C3308 a_n2661_44458# a_n699_43396# 0.002525f
C3309 a_11691_44458# a_13076_44458# 0.03093f
C3310 a_11827_44484# a_14539_43914# 0.044058f
C3311 a_10193_42453# a_18797_44260# 0.003033f
C3312 a_14537_43396# a_16789_44484# 2.77e-19
C3313 a_15765_45572# a_15493_43940# 2.68e-20
C3314 a_n1059_45260# a_1414_42308# 0.031011f
C3315 a_n2017_45002# a_453_43940# 8.57e-22
C3316 a_n2661_45010# a_2675_43914# 1.7e-19
C3317 a_3357_43084# a_5663_43940# 0.015908f
C3318 a_n2293_45010# a_2479_44172# 1.92e-20
C3319 a_n4318_37592# a_n2956_38216# 0.023126f
C3320 a_17303_42282# a_17715_44484# 3.11e-21
C3321 a_5907_45546# VDD 0.390381f
C3322 a_17364_32525# a_22469_39537# 1.61e-20
C3323 a_4190_30871# a_11530_34132# 0.031248f
C3324 a_9313_44734# a_18479_47436# 4.54e-21
C3325 a_11652_45724# a_10809_44734# 0.073342f
C3326 a_15004_44636# a_n881_46662# 9.62e-22
C3327 a_n2017_45002# a_17339_46660# 4.48e-20
C3328 a_413_45260# a_14513_46634# 1.94e-20
C3329 a_4880_45572# a_526_44458# 0.02064f
C3330 a_7227_45028# a_5066_45546# 8.68e-20
C3331 a_20623_45572# a_20202_43084# 9.54e-19
C3332 a_1307_43914# a_8270_45546# 0.050297f
C3333 a_5883_43914# a_768_44030# 0.087568f
C3334 a_13159_45002# a_12991_46634# 2.16e-21
C3335 a_20841_45814# a_11415_45002# 0.004448f
C3336 a_13017_45260# a_12816_46660# 2.41e-21
C3337 a_n2661_43370# a_5167_46660# 2.93e-21
C3338 a_16414_43172# a_15764_42576# 0.001182f
C3339 a_15567_42826# a_15803_42450# 1.29e-20
C3340 a_17701_42308# a_14113_42308# 4.89e-20
C3341 a_n4318_38680# a_n4334_40480# 1.45e-19
C3342 a_5342_30871# a_15959_42545# 7.85e-19
C3343 a_n3674_39304# a_n4064_40160# 0.024923f
C3344 a_2747_46873# a_2443_46660# 0.129886f
C3345 a_4883_46098# a_3877_44458# 0.002191f
C3346 a_n1435_47204# a_10467_46802# 1.8e-20
C3347 a_9313_45822# a_10249_46116# 1.36e-19
C3348 a_11031_47542# a_6755_46942# 0.001571f
C3349 a_6151_47436# a_6903_46660# 4.55e-19
C3350 a_n1151_42308# a_11813_46116# 0.019835f
C3351 a_n881_46662# a_1123_46634# 0.004455f
C3352 a_n1613_43370# a_948_46660# 0.281392f
C3353 a_5807_45002# a_16750_47204# 5.29e-19
C3354 a_13747_46662# a_19594_46812# 0.03826f
C3355 a_10057_43914# a_10729_43914# 0.063518f
C3356 a_11967_42832# a_19615_44636# 0.065767f
C3357 a_n2661_43922# a_n1899_43946# 0.00455f
C3358 a_n2293_43922# a_n1761_44111# 0.005057f
C3359 a_n2661_42834# a_n1331_43914# 0.01077f
C3360 a_8975_43940# a_10405_44172# 1.35e-19
C3361 a_n2293_42834# a_n2433_43396# 0.025997f
C3362 a_11823_42460# a_13113_42826# 0.003218f
C3363 a_10193_42453# a_15567_42826# 1.05e-20
C3364 a_1307_43914# a_1987_43646# 0.002379f
C3365 a_6109_44484# a_5495_43940# 2.63e-20
C3366 a_626_44172# a_766_43646# 9.22e-19
C3367 a_5205_44484# a_6655_43762# 5.14e-19
C3368 a_3232_43370# a_3457_43396# 0.131408f
C3369 a_3537_45260# a_8685_43396# 0.023888f
C3370 a_n1059_45260# a_12281_43396# 0.025081f
C3371 a_5111_44636# a_5837_43396# 7.68e-19
C3372 a_5932_42308# a_n1532_35090# 1.05e-19
C3373 a_18443_44721# a_12741_44636# 0.002904f
C3374 a_11341_43940# a_5807_45002# 0.002004f
C3375 a_17061_44734# a_15227_44166# 0.07208f
C3376 a_20365_43914# a_19321_45002# 0.006039f
C3377 a_20935_43940# a_13747_46662# 2.52e-19
C3378 a_12603_44260# a_12549_44172# 0.00397f
C3379 a_14955_43940# a_n2293_46634# 0.004724f
C3380 a_12495_44260# a_768_44030# 0.001355f
C3381 a_5009_45028# a_5066_45546# 1.52e-19
C3382 a_13348_45260# a_13259_45724# 0.016055f
C3383 a_413_45260# a_n357_42282# 0.032207f
C3384 a_327_44734# a_310_45028# 0.006962f
C3385 a_n37_45144# a_n755_45592# 0.050738f
C3386 a_2680_45002# a_n863_45724# 0.024737f
C3387 a_n2293_45010# a_n443_42852# 0.003134f
C3388 a_4558_45348# a_n2661_45546# 0.050441f
C3389 a_3429_45260# a_n2293_45546# 3.77e-21
C3390 a_16922_45042# a_20075_46420# 9.42e-20
C3391 a_n2661_44458# a_7920_46348# 4.63e-21
C3392 a_18911_45144# a_18189_46348# 1.91e-19
C3393 a_11691_44458# a_12594_46348# 4.78e-21
C3394 a_20974_43370# a_18479_47436# 0.008175f
C3395 a_21381_43940# a_18597_46090# 0.080234f
C3396 a_15764_42576# a_7174_31319# 6.35e-20
C3397 a_16197_42308# a_4958_30871# 9.31e-19
C3398 a_6123_31319# a_n4209_39304# 5.16e-21
C3399 a_13717_47436# VDD 0.314317f
C3400 a_n2661_46634# a_167_45260# 2.09e-19
C3401 a_n2293_46634# a_1138_42852# 0.023262f
C3402 a_n1925_46634# a_805_46414# 9.66e-19
C3403 a_n743_46660# a_376_46348# 0.076781f
C3404 a_n2438_43548# a_n1076_46494# 2.06e-20
C3405 a_171_46873# a_n1641_46494# 5.78e-21
C3406 a_12469_46902# a_12816_46660# 0.051162f
C3407 a_5275_47026# a_765_45546# 0.002883f
C3408 a_11309_47204# a_9290_44172# 4.41e-19
C3409 a_n881_46662# a_13759_46122# 0.01582f
C3410 a_10227_46804# a_526_44458# 5.93e-20
C3411 a_11453_44696# a_6945_45028# 0.022389f
C3412 a_22731_47423# a_10809_44734# 0.005082f
C3413 a_n2288_47178# a_n2661_45546# 1.03e-20
C3414 a_n2833_47464# a_n2956_38216# 1e-20
C3415 a_n1549_44318# a_n1177_43370# 0.003012f
C3416 a_20365_43914# a_20623_43914# 0.22264f
C3417 a_19328_44172# a_15493_43940# 0.062184f
C3418 a_19478_44306# a_11341_43940# 6.59e-19
C3419 a_19862_44208# a_21115_43940# 0.064973f
C3420 a_n1331_43914# a_n1352_43396# 1.74e-20
C3421 a_1307_43914# a_4649_42852# 1.56e-19
C3422 a_n356_44636# a_15743_43084# 2.51e-20
C3423 a_10193_42453# a_20712_42282# 0.157661f
C3424 a_12429_44172# a_12603_44260# 0.011572f
C3425 a_3499_42826# a_3992_43940# 2.6e-19
C3426 a_n1761_44111# a_n97_42460# 0.001173f
C3427 a_14539_43914# a_17433_43396# 1.68e-19
C3428 a_n2017_45002# a_n2472_42282# 0.001176f
C3429 a_19237_31679# VDD 0.746512f
C3430 a_11962_45724# a_11682_45822# 0.014813f
C3431 a_11823_42460# a_10907_45822# 1.3e-19
C3432 a_7499_43078# a_11136_45572# 1.89e-21
C3433 a_10193_42453# a_10216_45572# 0.003165f
C3434 a_10053_45546# a_10544_45572# 0.00278f
C3435 a_10180_45724# a_10306_45572# 9.37e-19
C3436 a_2711_45572# a_14033_45572# 6.82e-19
C3437 C6_N_btm C3_P_btm 2.03e-19
C3438 C5_N_btm C2_P_btm 3.54e-20
C3439 a_5193_42852# a_4791_45118# 0.004916f
C3440 a_5534_30871# a_12465_44636# 1.02e-21
C3441 a_7227_42852# a_n1613_43370# 0.007002f
C3442 a_10807_43548# a_9290_44172# 0.364112f
C3443 a_20512_43084# a_8049_45260# 5.74e-21
C3444 a_9313_44734# a_n443_42852# 0.02484f
C3445 a_1414_42308# a_n1925_42282# 5.84e-21
C3446 a_453_43940# a_526_44458# 0.028123f
C3447 a_17364_32525# a_22612_30879# 0.062457f
C3448 a_9396_43370# a_8270_45546# 8.62e-19
C3449 a_14035_46660# VDD 0.363878f
C3450 a_5742_30871# a_n4064_37440# 0.004687f
C3451 a_4704_46090# a_5068_46348# 5.06e-19
C3452 a_12991_46634# a_13259_45724# 6.17e-19
C3453 a_765_45546# a_2981_46116# 3.97e-21
C3454 a_12741_44636# a_17583_46090# 2.35e-20
C3455 a_11415_45002# a_17957_46116# 4.92e-22
C3456 a_3483_46348# a_6165_46155# 1.15e-21
C3457 a_22959_43948# a_17364_32525# 0.005227f
C3458 a_3626_43646# a_7287_43370# 2.15e-20
C3459 a_2982_43646# a_8147_43396# 1.75e-21
C3460 a_n97_42460# a_14579_43548# 0.001021f
C3461 a_14021_43940# a_21487_43396# 0.023941f
C3462 a_n356_44636# a_1606_42308# 0.282657f
C3463 a_11967_42832# a_11229_43218# 3.74e-21
C3464 a_18494_42460# a_17124_42282# 4.91e-20
C3465 a_3080_42308# a_4181_43396# 2.84e-19
C3466 a_n237_47217# DATA[4] 0.001087f
C3467 a_1209_47178# DATA[0] 3.05e-20
C3468 a_327_47204# DATA[1] 2.2e-19
C3469 a_9145_43396# VDD 2.43736f
C3470 a_12427_45724# a_11827_44484# 3.2e-21
C3471 a_11322_45546# a_11691_44458# 1.74e-19
C3472 a_2711_45572# a_6298_44484# 6.39e-20
C3473 a_10193_42453# a_16886_45144# 0.001731f
C3474 a_3357_43084# a_3232_43370# 0.118744f
C3475 a_n967_45348# a_n955_45028# 0.014419f
C3476 a_n745_45366# a_413_45260# 4.33e-20
C3477 a_19164_43230# a_17339_46660# 9.04e-20
C3478 a_n784_42308# a_4646_46812# 4.29e-21
C3479 a_7963_42308# a_n2293_46634# 2.47e-20
C3480 a_5934_30871# a_n2442_46660# 7.2e-21
C3481 a_9061_43230# a_3090_45724# 3.86e-21
C3482 a_104_43370# a_n755_45592# 0.029812f
C3483 a_n229_43646# a_n863_45724# 4.39e-19
C3484 a_743_42282# a_10903_43370# 0.029178f
C3485 a_7174_31319# a_13507_46334# 0.041342f
C3486 a_21125_42558# a_18597_46090# 0.002227f
C3487 a_19237_31679# a_22469_39537# 2.75e-20
C3488 a_n1099_45572# VDD 0.89411f
C3489 a_2437_43646# a_n971_45724# 0.204278f
C3490 a_17478_45572# a_11599_46634# 0.025658f
C3491 a_16115_45572# a_16327_47482# 0.163022f
C3492 a_9159_45572# a_4883_46098# 6.4e-19
C3493 a_11652_45724# a_n881_46662# 4.56e-21
C3494 a_1260_45572# a_n2293_46634# 6.07e-19
C3495 a_8162_45546# a_768_44030# 2.17e-21
C3496 a_n2840_43370# a_n3674_38680# 0.003987f
C3497 a_n1991_42858# a_n1423_42826# 0.186387f
C3498 a_n2157_42858# a_n901_43156# 0.043475f
C3499 a_n1853_43023# a_n1641_43230# 0.036072f
C3500 a_10341_43396# a_21671_42860# 1.14e-19
C3501 a_743_42282# a_3681_42891# 1.37e-20
C3502 a_3422_30871# a_n3420_39072# 0.096346f
C3503 a_16137_43396# a_15567_42826# 6.67e-19
C3504 a_8270_45546# DATA[4] 0.003852f
C3505 a_20107_45572# a_20159_44458# 2.4e-19
C3506 a_18315_45260# a_18911_45144# 7.05e-19
C3507 a_16922_45042# a_20567_45036# 0.002083f
C3508 a_16019_45002# a_16112_44458# 3.78e-19
C3509 a_1307_43914# a_15004_44636# 1.02e-20
C3510 a_7499_43078# a_11750_44172# 0.195997f
C3511 a_n2293_42834# a_n2433_44484# 4.65e-21
C3512 a_327_44734# a_556_44484# 0.033015f
C3513 a_21513_45002# a_17517_44484# 2.37e-19
C3514 a_5111_44636# a_8375_44464# 0.001962f
C3515 a_5147_45002# a_5891_43370# 0.049542f
C3516 a_n967_45348# a_n2661_42834# 0.027185f
C3517 en_comp a_n2661_43922# 0.237031f
C3518 a_n2956_37592# a_n2293_43922# 2.05e-20
C3519 a_10533_42308# a_4185_45028# 9.41e-20
C3520 a_5934_30871# a_8953_45546# 0.113715f
C3521 a_1793_42852# a_n863_45724# 5.96e-19
C3522 a_n3674_37592# a_n2956_38680# 0.026013f
C3523 a_13249_42308# a_12741_44636# 0.028381f
C3524 a_8696_44636# a_13059_46348# 0.020156f
C3525 a_19431_45546# a_15227_44166# 2.07e-20
C3526 a_17668_45572# a_3090_45724# 0.071363f
C3527 a_18909_45814# a_19466_46812# 0.001786f
C3528 a_1423_45028# a_n2438_43548# 0.242599f
C3529 a_n2661_43370# a_12549_44172# 3e-20
C3530 a_4927_45028# a_4651_46660# 5.26e-21
C3531 a_5147_45002# a_4817_46660# 6.83e-20
C3532 a_3232_43370# a_3877_44458# 0.016642f
C3533 a_5691_45260# a_4646_46812# 1.06e-21
C3534 a_2711_45572# a_5937_45572# 0.063757f
C3535 a_11827_44484# a_11453_44696# 0.170003f
C3536 a_11691_44458# a_12465_44636# 0.15589f
C3537 a_18114_32519# a_18479_47436# 3.09e-20
C3538 a_13720_44458# a_4915_47217# 0.006519f
C3539 a_700_44734# a_n746_45260# 0.009437f
C3540 a_15743_43084# a_18727_42674# 1.5e-19
C3541 a_5111_42852# a_4921_42308# 3.76e-20
C3542 a_22959_42860# a_14097_32519# 0.166017f
C3543 a_743_42282# a_15959_42545# 0.006675f
C3544 a_4361_42308# a_14113_42308# 0.075467f
C3545 a_21195_42852# a_20753_42852# 7.65e-19
C3546 a_16867_43762# a_4958_30871# 4.18e-20
C3547 a_11599_46634# a_19594_46812# 0.001035f
C3548 a_16327_47482# a_5807_45002# 0.451783f
C3549 a_16588_47582# a_16697_47582# 0.007416f
C3550 a_16763_47508# a_16942_47570# 0.007399f
C3551 a_16023_47582# a_16131_47204# 0.057222f
C3552 a_4883_46098# a_8128_46384# 0.010382f
C3553 a_7903_47542# a_n1925_46634# 8.56e-21
C3554 a_11459_47204# a_n2661_46634# 1.65e-19
C3555 a_13717_47436# a_22612_30879# 0.00542f
C3556 a_n1151_42308# a_1110_47026# 1.25e-19
C3557 a_n971_45724# a_3686_47026# 1.68e-19
C3558 a_584_46384# a_2609_46660# 3.91e-19
C3559 a_4700_47436# a_2107_46812# 3.8e-22
C3560 a_2063_45854# a_2443_46660# 0.017518f
C3561 a_n443_46116# a_1123_46634# 8.72e-19
C3562 a_n1741_47186# a_4651_46660# 4.72e-20
C3563 a_n2109_47186# a_4817_46660# 0.028101f
C3564 a_18989_43940# a_19615_44636# 8.51e-19
C3565 a_n1177_44458# a_n1549_44318# 0.004943f
C3566 a_18248_44752# a_20679_44626# 1.77e-21
C3567 a_n1352_44484# a_n1331_43914# 7.59e-19
C3568 a_1307_43914# a_1241_43940# 0.038832f
C3569 a_7499_43078# a_4361_42308# 0.04291f
C3570 a_10193_42453# a_20556_43646# 1.67e-19
C3571 a_10617_44484# a_n2661_43922# 0.004461f
C3572 a_n967_45348# a_n1352_43396# 0.010028f
C3573 a_3357_43084# a_4905_42826# 0.062628f
C3574 a_n2661_45010# a_1209_43370# 9.39e-22
C3575 a_n2017_45002# a_n1821_43396# 0.001012f
C3576 a_n3565_39304# a_n2810_45572# 0.030572f
C3577 a_n1059_45260# VDD 4.75361f
C3578 a_22400_42852# a_22521_40055# 0.681186f
C3579 a_1241_43940# a_n443_46116# 1.44e-19
C3580 a_17613_45144# a_12741_44636# 0.006096f
C3581 a_18587_45118# a_11415_45002# 0.005313f
C3582 a_19478_44306# a_16327_47482# 3.2e-19
C3583 a_15493_43940# a_12861_44030# 0.370814f
C3584 a_9672_43914# a_4883_46098# 0.009886f
C3585 a_6709_45028# a_6945_45028# 0.060282f
C3586 a_n4318_39768# a_n1613_43370# 1.98e-19
C3587 a_14180_45002# a_2324_44458# 0.026932f
C3588 a_14797_45144# a_15015_46420# 2.32e-20
C3589 a_413_45260# a_518_46155# 3.64e-20
C3590 a_2274_45254# a_526_44458# 0.019853f
C3591 a_19237_31679# a_22612_30879# 0.062542f
C3592 a_2889_44172# a_768_44030# 0.011283f
C3593 a_17970_44736# a_3090_45724# 1.26e-19
C3594 a_9803_42558# a_10533_42308# 5.35e-19
C3595 a_8685_42308# a_5742_30871# 4.1e-20
C3596 COMP_P a_22775_42308# 4.23e-19
C3597 EN_VIN_BSTR_P VIN_P 1.41696f
C3598 C5_P_btm C2_P_btm 0.13795f
C3599 C4_P_btm C3_P_btm 9.61674f
C3600 a_9313_45822# a_5937_45572# 0.137696f
C3601 a_6151_47436# a_10903_43370# 6.84e-20
C3602 a_4915_47217# a_13351_46090# 3.17e-21
C3603 a_n1435_47204# a_8016_46348# 1.14e-20
C3604 a_13675_47204# a_765_45546# 7.69e-19
C3605 a_7715_46873# a_8145_46902# 2.33e-20
C3606 a_5732_46660# a_6755_46942# 1.39e-20
C3607 a_3877_44458# a_6682_46660# 0.002161f
C3608 a_4817_46660# a_5841_46660# 2.36e-20
C3609 a_7411_46660# a_7927_46660# 0.105839f
C3610 a_9482_43914# a_10083_42826# 4.71e-19
C3611 a_n2293_43922# a_n2267_43396# 0.020404f
C3612 a_19237_31679# a_22959_43948# 5.09e-19
C3613 a_n2661_42834# a_n1917_43396# 0.007372f
C3614 a_11691_44458# a_16409_43396# 6.27e-20
C3615 a_11827_44484# a_17324_43396# 2.91e-21
C3616 a_18184_42460# a_19700_43370# 0.003845f
C3617 a_18494_42460# a_19268_43646# 5.16e-21
C3618 a_1307_43914# a_5755_42852# 2.6e-19
C3619 a_n356_44636# a_3539_42460# 1.86e-19
C3620 a_7845_44172# a_7911_44260# 0.010598f
C3621 a_7542_44172# a_8018_44260# 0.001923f
C3622 a_5708_44484# a_n97_42460# 4.19e-21
C3623 a_5343_44458# a_8317_43396# 1.12e-19
C3624 a_8701_44490# a_8685_43396# 1.11e-20
C3625 a_n967_45348# a_n2293_42282# 5.08e-19
C3626 a_n913_45002# a_133_42852# 0.046777f
C3627 a_n3420_39072# VREF_GND 0.066097f
C3628 a_2711_45572# a_5437_45600# 5.64e-19
C3629 a_895_43940# a_1823_45246# 1.63e-20
C3630 a_2127_44172# a_167_45260# 3.83e-20
C3631 a_10341_43396# a_5807_45002# 1.82e-19
C3632 a_n97_42460# a_5257_43370# 0.167676f
C3633 a_3080_42308# a_4646_46812# 2.88e-19
C3634 a_15681_43442# a_12549_44172# 0.080982f
C3635 a_15301_44260# a_15227_44166# 0.003263f
C3636 a_8685_43396# a_n2293_46634# 0.335608f
C3637 a_949_44458# a_n755_45592# 0.011024f
C3638 a_2779_44458# a_n357_42282# 8.49e-21
C3639 a_17767_44458# a_18051_46116# 5.87e-22
C3640 a_21487_43396# a_13507_46334# 4.46e-21
C3641 a_743_42282# a_4883_46098# 1.38e-19
C3642 a_5649_42852# a_18597_46090# 9.18e-20
C3643 a_10796_42968# a_2063_45854# 7.47e-21
C3644 en_comp a_22459_39145# 0.415926f
C3645 a_n2946_38778# a_n4064_38528# 0.053228f
C3646 a_n3420_38528# a_n2302_38778# 1.28e-19
C3647 a_4958_30871# C5_N_btm 1.35e-19
C3648 a_20202_43084# a_22591_46660# 0.001634f
C3649 a_765_45546# a_167_45260# 0.276049f
C3650 a_22365_46825# a_20820_30879# 0.00309f
C3651 a_n2661_46634# a_n863_45724# 3.34e-20
C3652 a_n2312_38680# a_n2661_45546# 5.53e-19
C3653 a_7715_46873# a_5066_45546# 0.020181f
C3654 a_n2293_46634# a_n2956_38216# 5.44e-19
C3655 a_14976_45028# a_15015_46420# 0.012921f
C3656 a_3090_45724# a_14840_46494# 0.002524f
C3657 a_n3674_38216# a_n4209_37414# 1.61e-20
C3658 a_n4318_38216# a_n3565_37414# 2.51e-20
C3659 a_n1899_43946# a_n1641_43230# 3.58e-20
C3660 a_n809_44244# a_n1853_43023# 4.45e-20
C3661 a_n2065_43946# a_n1076_43230# 2.53e-21
C3662 a_n1549_44318# a_n1991_42858# 6.41e-19
C3663 a_5663_43940# a_743_42282# 7.52e-22
C3664 a_19478_44306# a_10341_43396# 5.01e-20
C3665 a_n2433_43396# a_n2012_43396# 0.089677f
C3666 a_11341_43940# a_13667_43396# 9.28e-19
C3667 a_n1761_44111# a_n901_43156# 0.013702f
C3668 a_11967_42832# a_10835_43094# 0.263495f
C3669 a_n4318_40392# a_n3674_38680# 0.023225f
C3670 a_n1917_43396# a_n1352_43396# 7.99e-20
C3671 a_n4318_39304# a_n1809_43762# 1.53e-19
C3672 a_n2129_43609# a_104_43370# 3.36e-19
C3673 a_n2810_45028# a_n2946_39866# 5.51e-20
C3674 a_n2956_37592# a_n3420_39616# 3.18e-19
C3675 a_n2840_43370# VDD 0.246858f
C3676 a_20273_45572# a_20841_45814# 0.175891f
C3677 a_14495_45572# a_9482_43914# 2.35e-20
C3678 a_13249_42308# a_13556_45296# 0.059719f
C3679 a_13904_45546# a_13777_45326# 1.68e-19
C3680 a_20107_45572# a_20623_45572# 0.103168f
C3681 a_8791_45572# a_6171_45002# 6.13e-19
C3682 a_n1557_42282# a_n2956_39304# 1.75e-20
C3683 a_n1925_42282# VDD 0.728242f
C3684 a_2711_45572# a_18479_47436# 1.11e-19
C3685 a_8746_45002# a_6151_47436# 8.1e-20
C3686 a_13904_45546# a_n1151_42308# 1.84e-19
C3687 a_8192_45572# a_n971_45724# 0.005205f
C3688 a_17583_46090# a_16375_45002# 4.13e-20
C3689 a_17957_46116# a_13259_45724# 0.011559f
C3690 a_14840_46494# a_15002_46116# 0.006453f
C3691 a_10809_44734# a_12379_46436# 0.011204f
C3692 a_18189_46348# a_18147_46436# 9.33e-19
C3693 a_167_45260# a_509_45822# 2.36e-20
C3694 a_1823_45246# a_1609_45822# 0.35471f
C3695 a_5013_44260# a_5932_42308# 4.06e-21
C3696 a_n1917_43396# a_n2293_42282# 9.44e-21
C3697 a_8147_43396# a_7871_42858# 1.53e-19
C3698 a_15781_43660# a_4361_42308# 1.85e-20
C3699 a_16243_43396# a_743_42282# 7.51e-20
C3700 a_18429_43548# a_16823_43084# 0.130506f
C3701 a_3499_42826# a_1755_42282# 2.38e-20
C3702 a_3626_43646# a_12089_42308# 0.002196f
C3703 a_2982_43646# a_13113_42826# 1.09e-20
C3704 a_n2661_42282# a_961_42354# 1.35e-19
C3705 a_5663_43940# a_5755_42308# 1e-20
C3706 a_17324_43396# a_17433_43396# 0.007416f
C3707 a_17499_43370# a_17678_43396# 0.007399f
C3708 a_15743_43084# a_17486_43762# 2.49e-19
C3709 a_16409_43396# a_4190_30871# 4.44e-21
C3710 a_11967_42832# a_16269_42308# 6.4e-20
C3711 a_2107_46812# DATA[2] 5.18e-20
C3712 a_19987_42826# VDD 0.588466f
C3713 a_5009_45028# a_5093_45028# 0.092725f
C3714 a_2711_45572# a_2479_44172# 9.28e-20
C3715 a_8696_44636# a_11649_44734# 5.17e-19
C3716 a_327_44734# a_n2661_44458# 0.027103f
C3717 a_n967_45348# a_n1352_44484# 0.007805f
C3718 a_n1059_45260# a_n699_43396# 0.021143f
C3719 a_n467_45028# a_n1699_44726# 1.68e-21
C3720 a_n913_45002# a_4223_44672# 6.25e-20
C3721 a_n13_43084# a_n357_42282# 0.194173f
C3722 a_n1076_43230# a_n755_45592# 2.49e-20
C3723 a_n1379_43218# a_n863_45724# 3.89e-21
C3724 a_8530_39574# w_11334_34010# 2.13e-19
C3725 a_15595_45028# a_11453_44696# 0.007267f
C3726 a_7229_43940# a_n1613_43370# 0.059621f
C3727 a_7276_45260# a_n881_46662# 4.09e-20
C3728 a_3232_43370# a_8128_46384# 1.19e-20
C3729 a_n2840_45002# a_n2293_46634# 7.08e-19
C3730 a_3537_45260# a_768_44030# 0.341201f
C3731 a_n2661_45010# a_n2442_46660# 1.33e-20
C3732 a_10180_45724# a_10185_46660# 7.92e-20
C3733 a_10193_42453# a_19692_46634# 0.010323f
C3734 a_11823_42460# a_15368_46634# 0.014491f
C3735 a_3626_43646# a_18907_42674# 0.003037f
C3736 a_10796_42968# a_10793_43218# 2.36e-20
C3737 a_12005_46116# CLK 8.86e-21
C3738 a_17583_46090# RST_Z 1.08e-21
C3739 a_n4315_30879# VDD 4.0486f
C3740 a_n1741_47186# a_10037_47542# 4.61e-19
C3741 a_n746_45260# a_n881_46662# 0.190303f
C3742 a_n971_45724# a_7989_47542# 1.99e-19
C3743 a_n237_47217# a_n1613_43370# 0.034341f
C3744 a_15507_47210# a_15811_47375# 0.170975f
C3745 a_6151_47436# a_4883_46098# 0.032223f
C3746 a_11599_46634# a_15673_47210# 0.012504f
C3747 a_2952_47436# a_2747_46873# 0.078913f
C3748 a_13717_47436# a_16588_47582# 6.43e-20
C3749 a_13381_47204# a_10227_46804# 7.94e-20
C3750 a_12861_44030# a_16763_47508# 0.008377f
C3751 a_18587_45118# a_11967_42832# 4.11e-20
C3752 a_18911_45144# a_19006_44850# 3.38e-19
C3753 a_n1699_44726# a_n2661_43922# 0.006002f
C3754 a_n1917_44484# a_n2661_42834# 0.002676f
C3755 a_10157_44484# a_5891_43370# 0.001885f
C3756 a_16922_45042# a_20679_44626# 5.14e-20
C3757 a_n2267_44484# a_n2293_43922# 6.94e-19
C3758 a_1423_45028# a_5013_44260# 3.14e-20
C3759 a_1307_43914# a_7845_44172# 0.002954f
C3760 a_8701_44490# a_8783_44734# 0.004999f
C3761 a_2779_44458# a_3363_44484# 0.020864f
C3762 a_11691_44458# a_16241_44734# 4.13e-19
C3763 a_n699_43396# a_484_44484# 1.33e-19
C3764 a_11827_44484# a_15146_44484# 1.1e-19
C3765 a_3232_43370# a_9672_43914# 4.68e-20
C3766 a_n913_45002# a_15493_43940# 1.64e-20
C3767 a_7229_43940# a_7584_44260# 0.001386f
C3768 a_n2302_39072# a_n2956_38680# 2.87e-19
C3769 a_11323_42473# a_n357_42282# 7.85e-20
C3770 a_8515_42308# a_n443_42852# 2.59e-21
C3771 a_15599_45572# VDD 0.390565f
C3772 a_5342_30871# a_n923_35174# 0.00897f
C3773 a_13159_45002# a_11415_45002# 0.141106f
C3774 a_3065_45002# a_1823_45246# 0.607468f
C3775 a_2382_45260# a_167_45260# 0.002522f
C3776 a_413_45260# a_3147_46376# 0.015235f
C3777 a_16405_45348# a_14976_45028# 1.42e-20
C3778 a_5891_43370# a_n1925_46634# 1.42e-20
C3779 a_11541_44484# a_768_44030# 0.003356f
C3780 a_2711_45572# a_n443_42852# 9.23e-22
C3781 a_1609_45572# a_1609_45822# 0.009518f
C3782 a_10306_45572# a_10586_45546# 1.95e-19
C3783 a_17517_44484# a_n881_46662# 2.63e-20
C3784 a_n2017_45002# a_8016_46348# 2.05e-20
C3785 a_2437_43646# a_12594_46348# 3.38e-20
C3786 a_18005_44484# a_11453_44696# 1e-19
C3787 a_21398_44850# a_13507_46334# 2.03e-20
C3788 a_21145_44484# a_18597_46090# 0.001307f
C3789 a_n630_44306# a_n1151_42308# 0.001084f
C3790 a_2351_42308# a_2713_42308# 0.00357f
C3791 a_1755_42282# a_3318_42354# 2.48e-19
C3792 a_1606_42308# a_3823_42558# 1.77e-20
C3793 a_n784_42308# a_6171_42473# 1.56e-20
C3794 a_5807_45002# a_8667_46634# 0.008461f
C3795 a_n743_46660# a_4651_46660# 9.85e-20
C3796 a_n1925_46634# a_4817_46660# 0.008055f
C3797 a_1799_45572# a_n2661_46098# 0.003478f
C3798 a_948_46660# a_1057_46660# 0.007416f
C3799 a_1123_46634# a_1302_46660# 0.007399f
C3800 a_n2661_46634# a_5072_46660# 0.002463f
C3801 a_15928_47570# a_6755_46942# 3.42e-19
C3802 a_n881_46662# a_8189_46660# 5.68e-19
C3803 a_n1613_43370# a_8270_45546# 9.43e-20
C3804 a_11453_44696# a_15559_46634# 1.71e-21
C3805 a_12465_44636# a_15227_44166# 1.22e-19
C3806 a_4883_46098# a_19466_46812# 0.028345f
C3807 a_21496_47436# a_19692_46634# 2.68e-21
C3808 a_11599_46634# a_16388_46812# 0.24092f
C3809 a_15507_47210# a_13059_46348# 2.35e-19
C3810 a_10227_46804# a_13170_46660# 0.003988f
C3811 a_15811_47375# a_15227_46910# 6.58e-19
C3812 a_11459_47204# a_765_45546# 0.005723f
C3813 a_n971_45724# a_n1853_46287# 0.08556f
C3814 a_n1741_47186# a_n1076_46494# 9.46e-21
C3815 a_n237_47217# a_n2293_46098# 0.044593f
C3816 a_21359_45002# a_2982_43646# 3.84e-21
C3817 a_n1177_44458# a_n1177_43370# 7.08e-19
C3818 a_n1331_43914# a_n1549_44318# 0.209641f
C3819 a_n2065_43946# a_175_44278# 5.71e-21
C3820 a_n1899_43946# a_n809_44244# 0.042737f
C3821 a_n1761_44111# a_n984_44318# 0.056404f
C3822 a_8704_45028# a_8685_43396# 1.1e-21
C3823 a_3232_43370# a_743_42282# 2.67e-20
C3824 en_comp a_n1641_43230# 6.37e-21
C3825 a_3357_43084# a_2905_42968# 0.025927f
C3826 a_n2017_45002# a_n1736_43218# 0.0083f
C3827 a_n967_45348# a_n1423_42826# 0.010397f
C3828 a_n3420_37440# VDD 2.26579f
C3829 a_n4318_40392# VDD 0.573389f
C3830 a_15521_42308# RST_Z 4.66e-20
C3831 a_4958_30871# C5_P_btm 1.35e-19
C3832 a_9241_44734# a_5937_45572# 9.79e-19
C3833 a_9313_44734# a_8199_44636# 0.016063f
C3834 a_n2661_43370# a_n2661_45546# 0.145941f
C3835 a_2809_45028# a_3316_45546# 9.97e-20
C3836 a_n699_43396# a_n1925_42282# 0.024581f
C3837 a_18587_45118# a_13259_45724# 0.099974f
C3838 a_17613_45144# a_16375_45002# 0.040514f
C3839 a_4743_44484# a_526_44458# 5.55e-19
C3840 a_14955_43940# a_6755_46942# 0.00126f
C3841 a_1049_43396# a_768_44030# 5.52e-20
C3842 a_n97_42460# a_5807_45002# 1.62e-22
C3843 a_11967_42832# a_11415_45002# 0.007699f
C3844 a_n2661_43922# a_4185_45028# 0.022579f
C3845 a_10490_45724# CLK 0.029352f
C3846 a_n4064_40160# a_n4064_39616# 5.80394f
C3847 a_n4209_39590# a_n3565_39590# 6.15218f
C3848 a_4958_30871# a_n3420_38528# 0.030871f
C3849 a_5257_43370# a_5204_45822# 0.005904f
C3850 a_4883_46098# a_20205_31679# 3.29e-19
C3851 a_15227_46910# a_13059_46348# 0.043664f
C3852 a_19692_46634# a_21363_46634# 0.00151f
C3853 a_15227_44166# a_20528_46660# 4.16e-21
C3854 a_5807_45002# a_6640_46482# 9.8e-19
C3855 a_n1925_46634# a_n722_46482# 2.37e-19
C3856 a_8492_46660# a_3483_46348# 1.74e-20
C3857 a_20679_44626# a_15743_43084# 9.47e-21
C3858 a_13720_44458# a_13460_43230# 1.78e-21
C3859 a_n2293_43922# a_n2472_42826# 1.92e-19
C3860 a_19478_44306# a_n97_42460# 6.27e-19
C3861 a_1307_43914# a_1067_42314# 3.75e-21
C3862 a_n2661_42834# a_n1853_43023# 0.002855f
C3863 a_n2661_43922# a_n2157_42858# 2.6e-21
C3864 a_n356_44636# a_8605_42826# 1.43e-20
C3865 a_375_42282# a_564_42282# 0.022891f
C3866 a_5745_43940# a_5829_43940# 0.092725f
C3867 a_n2661_42282# a_2982_43646# 0.076578f
C3868 a_3232_43370# a_5755_42308# 2.19e-21
C3869 a_n913_45002# a_5742_30871# 0.028271f
C3870 a_3065_45002# a_5934_30871# 1.09e-20
C3871 a_3537_45260# a_6123_31319# 9.93e-19
C3872 a_n1059_45260# a_11551_42558# 9.25e-20
C3873 a_2382_45260# a_3905_42308# 4.58e-19
C3874 a_n2017_45002# a_11633_42558# 0.005942f
C3875 a_18326_43940# VDD 0.129408f
C3876 a_16333_45814# a_16223_45938# 0.097745f
C3877 a_16680_45572# a_15861_45028# 1.57e-19
C3878 a_16855_45546# a_17478_45572# 3.95e-19
C3879 a_14033_45822# a_14033_45572# 6.96e-20
C3880 a_16115_45572# a_16020_45572# 0.049827f
C3881 a_2711_45572# a_2680_45002# 2.69e-19
C3882 a_1209_43370# a_1138_42852# 0.01435f
C3883 a_14205_43396# a_13059_46348# 0.049915f
C3884 a_16409_43396# a_15227_44166# 0.003488f
C3885 a_644_44056# a_n357_42282# 0.007544f
C3886 a_2998_44172# a_n2661_45546# 0.060624f
C3887 a_10729_43914# a_10586_45546# 2.76e-22
C3888 a_175_44278# a_n755_45592# 0.01086f
C3889 a_20256_43172# a_16327_47482# 0.054992f
C3890 a_5934_30871# w_1575_34946# 0.002787f
C3891 a_2698_46116# VDD 0.195879f
C3892 C5_N_btm C7_N_btm 0.151416f
C3893 C2_N_btm C10_N_btm 0.327137f
C3894 C3_N_btm C9_N_btm 0.137552f
C3895 C4_N_btm C8_N_btm 0.145646f
C3896 a_1177_38525# a_2113_38308# 1.21e-19
C3897 a_n4209_38216# a_n4064_37984# 0.19304f
C3898 a_n3565_38216# a_n3420_37984# 0.238595f
C3899 a_n4064_39616# a_n4064_37440# 0.050913f
C3900 a_11415_45002# a_13259_45724# 0.505354f
C3901 a_765_45546# a_n863_45724# 0.00497f
C3902 a_21363_46634# a_20692_30879# 2.83e-19
C3903 a_8016_46348# a_526_44458# 0.005011f
C3904 a_5068_46348# a_5210_46482# 0.007833f
C3905 a_18189_46348# a_17957_46116# 0.038851f
C3906 a_17715_44484# a_18819_46122# 1.03e-20
C3907 a_13925_46122# a_6945_45028# 3.29e-20
C3908 a_13351_46090# a_10809_44734# 5.63e-20
C3909 a_4419_46090# a_5066_45546# 8.55e-19
C3910 a_n2840_43370# a_n4318_38680# 0.001904f
C3911 a_n1917_43396# a_n1423_42826# 0.001812f
C3912 a_n1352_43396# a_n1853_43023# 5.05e-20
C3913 a_n1177_43370# a_n1991_42858# 0.003015f
C3914 a_4905_42826# a_743_42282# 0.0175f
C3915 a_14205_43396# a_15095_43370# 0.086245f
C3916 a_13667_43396# a_10341_43396# 0.007486f
C3917 a_n2129_43609# a_n1076_43230# 3.31e-20
C3918 a_14021_43940# a_15567_42826# 4.16e-20
C3919 a_15493_43940# a_20922_43172# 1.71e-21
C3920 a_11341_43940# a_21195_42852# 4.62e-21
C3921 a_2982_43646# a_16823_43084# 1.31e-20
C3922 a_n2293_43922# a_9223_42460# 4.38e-20
C3923 a_9313_44734# a_13070_42354# 3.27e-21
C3924 a_n4318_39304# a_n3674_39304# 2.9537f
C3925 a_10695_43548# a_10765_43646# 0.011552f
C3926 a_9145_43396# a_12293_43646# 0.003544f
C3927 a_n2661_42282# a_5837_42852# 0.002566f
C3928 a_12465_44636# EN_OFFSET_CAL 2.39e-20
C3929 a_n2312_39304# CLK_DATA 0.003547f
C3930 a_22959_43396# VDD 0.303237f
C3931 a_19431_45546# a_19113_45348# 0.001195f
C3932 a_13017_45260# a_13348_45260# 0.044101f
C3933 a_11963_45334# a_9482_43914# 2.68e-20
C3934 a_7499_43078# a_5891_43370# 1.00892f
C3935 a_18691_45572# a_11691_44458# 7.43e-20
C3936 a_4927_45028# a_1423_45028# 1.19e-20
C3937 a_n913_45002# a_n2293_42834# 0.055202f
C3938 a_n37_45144# a_45_45144# 0.004937f
C3939 a_3429_45260# a_3602_45348# 0.007688f
C3940 a_3537_45260# a_3495_45348# 7.3e-19
C3941 a_20528_45572# a_16922_45042# 7.24e-19
C3942 a_7466_43396# a_n443_42852# 2.62e-19
C3943 a_15861_45028# a_13747_46662# 0.021551f
C3944 a_2437_43646# a_12465_44636# 0.18195f
C3945 a_3357_43084# a_21496_47436# 2.47e-20
C3946 a_22591_45572# a_13507_46334# 9.32e-20
C3947 a_3232_43370# a_6151_47436# 7.33e-19
C3948 a_413_45260# a_12861_44030# 2.92e-19
C3949 a_10951_45334# a_n1151_42308# 1.15e-20
C3950 a_1307_43914# a_n746_45260# 1.91e-20
C3951 a_7229_43940# a_4791_45118# 0.026326f
C3952 a_2957_45546# a_3218_45724# 0.063846f
C3953 a_n755_45592# a_n356_45724# 0.016853f
C3954 a_n2293_45546# a_1609_45822# 0.159696f
C3955 a_n1099_45572# a_7_45899# 5.1e-20
C3956 a_n1853_43023# a_n2293_42282# 4.92e-20
C3957 a_10083_42826# a_10796_42968# 0.042737f
C3958 a_10518_42984# a_10835_43094# 0.102355f
C3959 a_3539_42460# a_3823_42558# 0.07742f
C3960 a_3626_43646# a_5267_42460# 1.19e-19
C3961 a_n97_42460# a_9223_42460# 0.004352f
C3962 a_14021_43940# a_20712_42282# 1.2e-20
C3963 a_4905_42826# a_5755_42308# 0.001861f
C3964 a_8337_42558# VDD 0.006426f
C3965 a_n746_45260# a_n443_46116# 0.060788f
C3966 a_1431_47204# a_n1151_42308# 0.013895f
C3967 a_n237_47217# a_4791_45118# 0.10712f
C3968 a_2063_45854# a_2952_47436# 2.96e-19
C3969 a_584_46384# a_2905_45572# 1.24e-20
C3970 a_n971_45724# a_4915_47217# 0.017974f
C3971 a_n1741_47186# a_6491_46660# 0.023524f
C3972 a_n2661_44458# a_4223_44672# 0.019953f
C3973 a_11691_44458# a_12883_44458# 0.058264f
C3974 a_11827_44484# a_16112_44458# 0.00849f
C3975 a_n1917_44484# a_n1352_44484# 7.99e-20
C3976 a_14537_43396# a_16335_44484# 0.003972f
C3977 a_10193_42453# a_18533_44260# 0.003163f
C3978 a_n967_45348# a_n1549_44318# 5.66e-19
C3979 a_n913_45002# a_1115_44172# 1.07e-21
C3980 a_n2017_45002# a_1414_42308# 0.015426f
C3981 a_3357_43084# a_5495_43940# 0.004364f
C3982 a_n2661_45010# a_895_43940# 0.020382f
C3983 a_n1736_42282# a_n2956_38216# 2.12e-20
C3984 a_20753_42852# a_n357_42282# 0.013117f
C3985 a_5263_45724# VDD 0.202719f
C3986 a_20273_45572# a_11415_45002# 0.01364f
C3987 a_11525_45546# a_10809_44734# 2.29e-19
C3988 a_8953_45002# a_3090_45724# 8.01e-20
C3989 a_413_45260# a_14180_46812# 1.15e-20
C3990 a_3357_43084# a_21363_46634# 2.28e-20
C3991 a_2711_45572# a_6633_46155# 1.05e-19
C3992 a_4808_45572# a_526_44458# 0.005047f
C3993 a_6598_45938# a_5066_45546# 1.62e-19
C3994 a_20841_45814# a_20202_43084# 0.001988f
C3995 a_8701_44490# a_768_44030# 0.00464f
C3996 a_15567_42826# a_15764_42576# 2.66e-20
C3997 a_5342_30871# a_15803_42450# 0.001339f
C3998 a_20256_43172# a_20356_42852# 0.001534f
C3999 a_n3674_39304# a_n4334_40480# 1.8e-19
C4000 a_22400_42852# a_14097_32519# 3.83e-19
C4001 a_n1613_43370# a_1123_46634# 0.358475f
C4002 a_2747_46873# a_n2661_46098# 0.004275f
C4003 a_n1435_47204# a_10428_46928# 1.94e-20
C4004 a_9313_45822# a_10554_47026# 3.34e-20
C4005 a_11031_47542# a_10249_46116# 0.003514f
C4006 a_n1151_42308# a_11735_46660# 0.050593f
C4007 a_4791_45118# a_8270_45546# 0.001618f
C4008 a_768_44030# a_n2293_46634# 0.26984f
C4009 a_13661_43548# a_19594_46812# 0.003227f
C4010 a_13747_46662# a_19321_45002# 0.080725f
C4011 a_n881_46662# a_383_46660# 0.001801f
C4012 a_10057_43914# a_10405_44172# 0.028414f
C4013 a_n2661_43922# a_n1761_44111# 0.006596f
C4014 a_n2293_43922# a_n2065_43946# 0.02752f
C4015 a_n2661_42834# a_n1899_43946# 0.049432f
C4016 a_8975_43940# a_9672_43914# 4.08e-19
C4017 a_17517_44484# a_18579_44172# 0.031747f
C4018 a_1423_45028# a_4699_43561# 1.02e-20
C4019 a_11823_42460# a_12545_42858# 0.039145f
C4020 a_10193_42453# a_5342_30871# 0.151919f
C4021 a_375_42282# a_n1557_42282# 0.450989f
C4022 a_1307_43914# a_1891_43646# 0.00299f
C4023 a_n1243_44484# a_n4318_39768# 6.55e-21
C4024 a_3232_43370# a_2813_43396# 0.05929f
C4025 a_n2017_45002# a_12281_43396# 0.028019f
C4026 a_5147_45002# a_5837_43396# 0.009374f
C4027 a_5111_44636# a_5565_43396# 3.27e-19
C4028 a_3537_45260# a_6809_43396# 5.68e-19
C4029 a_n784_42308# VIN_N 0.004358f
C4030 a_2779_44458# a_3147_46376# 2.99e-20
C4031 a_18287_44626# a_12741_44636# 0.004901f
C4032 a_18989_43940# a_11415_45002# 2.61e-19
C4033 a_13857_44734# a_14035_46660# 9.44e-21
C4034 a_16241_44734# a_15227_44166# 0.105126f
C4035 a_20269_44172# a_19321_45002# 6.92e-19
C4036 a_13483_43940# a_n2293_46634# 8.18e-21
C4037 a_12495_44260# a_12549_44172# 0.002899f
C4038 a_11816_44260# a_768_44030# 5.23e-19
C4039 a_13159_45002# a_13259_45724# 0.047761f
C4040 a_327_44734# a_n1099_45572# 3.5e-20
C4041 a_n143_45144# a_n755_45592# 0.07862f
C4042 a_413_45260# a_310_45028# 0.025313f
C4043 a_2382_45260# a_n863_45724# 0.119625f
C4044 a_4574_45260# a_n2661_45546# 0.014727f
C4045 a_n37_45144# a_n357_42282# 1.32e-21
C4046 a_3065_45002# a_n2293_45546# 9.28e-21
C4047 a_n2661_45010# a_1609_45822# 0.003846f
C4048 a_11827_44484# a_13925_46122# 5.41e-21
C4049 a_16922_45042# a_19335_46494# 1.17e-20
C4050 a_18315_45260# a_17957_46116# 3.37e-20
C4051 a_11691_44458# a_12005_46116# 8.12e-21
C4052 a_n2661_44458# a_6419_46155# 1.98e-22
C4053 a_18587_45118# a_18189_46348# 5.47e-19
C4054 a_14401_32519# a_18479_47436# 3.18e-21
C4055 a_15486_42560# a_7174_31319# 1.69e-21
C4056 a_6123_31319# a_1343_38525# 1.91e-19
C4057 a_17124_42282# a_17531_42308# 0.003716f
C4058 a_15761_42308# a_4958_30871# 1.41e-19
C4059 a_n1435_47204# VDD 0.267875f
C4060 a_17364_32525# VDAC_N 0.002958f
C4061 a_n2293_46634# a_1176_45822# 0.001481f
C4062 a_n1925_46634# a_472_46348# 0.002778f
C4063 a_n743_46660# a_n1076_46494# 0.001766f
C4064 a_n2438_43548# a_n901_46420# 5.58e-20
C4065 a_1123_46634# a_n2293_46098# 4.36e-20
C4066 a_171_46873# a_n1423_46090# 1.51e-20
C4067 a_11735_46660# a_14084_46812# 3.45e-21
C4068 a_11901_46660# a_12816_46660# 0.125324f
C4069 a_6755_46942# a_12978_47026# 3.05e-19
C4070 a_5072_46660# a_765_45546# 0.001239f
C4071 a_n881_46662# a_13351_46090# 5.07e-21
C4072 a_11453_44696# a_21137_46414# 7.06e-21
C4073 a_22223_47212# a_10809_44734# 0.009267f
C4074 a_n2497_47436# a_n2661_45546# 0.030609f
C4075 a_19279_43940# a_2982_43646# 9.07e-21
C4076 a_n1899_43946# a_n1352_43396# 4.29e-19
C4077 a_18451_43940# a_15493_43940# 0.051906f
C4078 a_15493_43396# a_11341_43940# 0.020569f
C4079 a_20269_44172# a_20623_43914# 0.001885f
C4080 a_19862_44208# a_20935_43940# 0.03846f
C4081 a_n1549_44318# a_n1917_43396# 9.82e-19
C4082 a_n1331_43914# a_n1177_43370# 1.74e-19
C4083 a_n1761_44111# a_n447_43370# 0.004447f
C4084 a_10193_42453# a_20107_42308# 0.007306f
C4085 a_n4318_40392# a_n4318_38680# 0.023692f
C4086 a_12429_44172# a_12495_44260# 0.012714f
C4087 a_1307_43914# a_4149_42891# 0.006879f
C4088 a_3499_42826# a_3737_43940# 0.002888f
C4089 a_14539_43914# a_16823_43084# 0.058282f
C4090 a_3357_43084# a_n784_42308# 4.03e-21
C4091 a_n2017_45002# a_n3674_38680# 2.15e-19
C4092 a_22959_44484# VDD 0.303517f
C4093 a_11652_45724# a_11682_45822# 0.006313f
C4094 a_10053_45546# a_10306_45572# 0.011897f
C4095 a_10180_45724# a_10216_45572# 0.002048f
C4096 a_12427_45724# a_10907_45822# 1.82e-21
C4097 a_2711_45572# a_13485_45572# 1.99e-20
C4098 C5_N_btm C3_P_btm 1.02e-19
C4099 C4_N_btm C2_P_btm 3.54e-20
C4100 a_4649_42852# a_4791_45118# 3.78e-19
C4101 a_21195_42852# a_16327_47482# 5.9e-20
C4102 a_14543_43071# a_12465_44636# 2.17e-22
C4103 a_3499_42826# a_2324_44458# 1.36e-21
C4104 a_10949_43914# a_9290_44172# 0.113864f
C4105 a_n2293_43922# a_n755_45592# 4.58e-19
C4106 a_11967_42832# a_13259_45724# 0.141918f
C4107 a_1414_42308# a_526_44458# 0.097596f
C4108 a_3626_43646# a_3090_45724# 4.54e-20
C4109 a_17364_32525# a_21588_30879# 0.05857f
C4110 a_8791_43396# a_8270_45546# 6.22e-19
C4111 a_11341_43940# a_3483_46348# 0.017129f
C4112 a_6171_45002# CLK 0.032376f
C4113 a_13885_46660# VDD 0.499249f
C4114 a_20731_47026# a_10809_44734# 0.003685f
C4115 a_4419_46090# a_5068_46348# 5.78e-21
C4116 a_765_45546# a_1431_46436# 4.27e-19
C4117 a_12741_44636# a_15682_46116# 3.17e-20
C4118 a_4185_45028# a_5164_46348# 1.41e-19
C4119 a_3483_46348# a_5497_46414# 8.7e-21
C4120 a_11415_45002# a_18189_46348# 0.028334f
C4121 a_1823_45246# a_5937_45572# 3.25e-20
C4122 a_22959_43948# a_22959_43396# 0.025171f
C4123 a_15493_43940# a_17364_32525# 9.31e-19
C4124 a_3626_43646# a_6547_43396# 1.95e-20
C4125 a_n97_42460# a_13667_43396# 2.99e-20
C4126 a_14021_43940# a_20556_43646# 0.085306f
C4127 a_18184_42460# a_17124_42282# 9.36e-20
C4128 a_n356_44636# a_1221_42558# 3.42e-19
C4129 a_3080_42308# a_3457_43396# 1.33e-19
C4130 a_n237_47217# DATA[3] 0.0265f
C4131 a_327_47204# DATA[0] 0.353891f
C4132 a_n785_47204# DATA[1] 2.65e-19
C4133 a_2711_45572# CAL_N 6.22e-19
C4134 a_5907_45546# a_4223_44672# 3.43e-21
C4135 a_10193_42453# a_16237_45028# 0.049386f
C4136 a_10490_45724# a_11691_44458# 2.02e-20
C4137 a_11136_45572# a_n2661_43370# 5.37e-20
C4138 a_n745_45366# a_n37_45144# 6.85e-19
C4139 a_3357_43084# a_5691_45260# 0.011637f
C4140 a_n1059_45260# a_327_44734# 1.06e-21
C4141 a_n913_45002# a_413_45260# 9.09e-20
C4142 a_5755_42852# a_n2293_46098# 4.28e-20
C4143 a_6123_31319# a_n2293_46634# 4.66e-20
C4144 a_n97_42460# a_n755_45592# 1.02989f
C4145 a_104_43370# a_n357_42282# 0.026213f
C4146 a_20712_42282# a_13507_46334# 4.89e-19
C4147 a_380_45546# VDD 0.154763f
C4148 a_15861_45028# a_11599_46634# 4.02e-19
C4149 a_16333_45814# a_16327_47482# 0.168559f
C4150 a_15225_45822# a_10227_46804# 7.94e-20
C4151 a_10907_45822# a_11453_44696# 3.71e-19
C4152 a_7499_43078# a_11309_47204# 3.32e-22
C4153 a_1176_45572# a_n2293_46634# 4.47e-19
C4154 a_2711_45572# a_n2661_46634# 0.032616f
C4155 a_7287_43370# a_7309_42852# 6.34e-20
C4156 a_n2157_42858# a_n1641_43230# 0.110532f
C4157 a_n1853_43023# a_n1423_42826# 0.022091f
C4158 a_10341_43396# a_21195_42852# 1.4e-20
C4159 a_743_42282# a_2905_42968# 8.11e-20
C4160 a_16137_43396# a_5342_30871# 1.45e-19
C4161 a_20273_45572# a_11967_42832# 1.95e-21
C4162 a_18315_45260# a_18587_45118# 0.13675f
C4163 a_16922_45042# a_18494_42460# 0.242236f
C4164 a_15415_45028# a_14539_43914# 4.93e-21
C4165 a_7499_43078# a_10807_43548# 0.119721f
C4166 a_1307_43914# a_13720_44458# 1.84e-20
C4167 a_10180_45724# a_10405_44172# 1.31e-21
C4168 a_n2293_42834# a_n2661_44458# 0.0289f
C4169 a_5111_44636# a_7640_43914# 0.001351f
C4170 a_327_44734# a_484_44484# 0.004093f
C4171 en_comp a_n2661_42834# 0.080292f
C4172 a_413_45260# a_556_44484# 2.84e-19
C4173 a_n2810_45028# a_n2293_43922# 2.3e-20
C4174 a_3537_45260# a_8333_44734# 1.47e-20
C4175 a_1709_42852# a_n863_45724# 7.55e-19
C4176 a_n3674_37592# a_n2956_39304# 0.026377f
C4177 a_3080_42308# VIN_N 0.025929f
C4178 a_13904_45546# a_12741_44636# 2.6e-21
C4179 a_15143_45578# a_11415_45002# 0.003102f
C4180 a_16680_45572# a_13059_46348# 1.67e-21
C4181 a_15037_45618# a_765_45546# 3e-21
C4182 a_16855_45546# a_16388_46812# 4.77e-21
C4183 a_18691_45572# a_15227_44166# 5.63e-21
C4184 a_626_44172# a_n133_46660# 1.1e-21
C4185 a_375_42282# a_33_46660# 2.38e-20
C4186 a_18341_45572# a_19466_46812# 0.02497f
C4187 a_17568_45572# a_3090_45724# 4.36e-20
C4188 a_6945_45348# a_5807_45002# 2.54e-21
C4189 a_18479_45785# a_19692_46634# 5.23e-20
C4190 a_1423_45028# a_n743_46660# 4.79e-20
C4191 a_5111_44636# a_4651_46660# 7.15e-21
C4192 a_3537_45260# a_5167_46660# 9.28e-22
C4193 a_5691_45260# a_3877_44458# 4.47e-21
C4194 a_6511_45714# a_5204_45822# 2.92e-21
C4195 a_5907_45546# a_6419_46155# 2.91e-20
C4196 a_2711_45572# a_8199_44636# 0.098064f
C4197 a_6194_45824# a_6165_46155# 5.54e-19
C4198 a_20193_45348# a_4883_46098# 3.03e-20
C4199 a_3775_45552# a_4419_46090# 2.91e-21
C4200 a_19700_43370# a_17303_42282# 4.48e-21
C4201 a_18783_43370# a_18727_42674# 1.92e-19
C4202 a_22959_42860# a_22400_42852# 8.07e-19
C4203 a_5649_42852# a_14456_42282# 1.31e-19
C4204 a_743_42282# a_15803_42450# 0.037845f
C4205 a_4190_30871# a_15890_42674# 2.93e-20
C4206 a_22223_42860# a_14097_32519# 5.42e-19
C4207 a_5342_30871# a_n784_42308# 0.049079f
C4208 a_4520_42826# a_4921_42308# 4.91e-19
C4209 a_16664_43396# a_4958_30871# 1.61e-19
C4210 a_11599_46634# a_19321_45002# 0.091019f
C4211 a_16327_47482# a_16131_47204# 0.016621f
C4212 a_16241_47178# a_5807_45002# 0.002482f
C4213 a_10227_46804# a_13675_47204# 1.49e-19
C4214 a_7227_47204# a_n1925_46634# 1.2e-19
C4215 a_9313_45822# a_n2661_46634# 0.032598f
C4216 a_6491_46660# a_n743_46660# 4.83e-21
C4217 a_13717_47436# a_21588_30879# 0.052863f
C4218 a_n443_46116# a_383_46660# 0.001079f
C4219 a_n1151_42308# a_n935_46688# 0.001606f
C4220 a_4007_47204# a_2107_46812# 7.24e-20
C4221 a_584_46384# a_2443_46660# 0.004099f
C4222 a_2063_45854# a_n2661_46098# 0.021195f
C4223 a_n2109_47186# a_4955_46873# 0.001032f
C4224 a_n1741_47186# a_4646_46812# 1.57e-19
C4225 a_n1917_44484# a_n1549_44318# 6.05e-19
C4226 a_n1352_44484# a_n1899_43946# 3.68e-19
C4227 a_n1177_44458# a_n1331_43914# 1.54e-19
C4228 a_n452_44636# a_n1761_44111# 4.05e-21
C4229 a_9313_44734# a_15433_44458# 1.54e-20
C4230 a_18989_43940# a_11967_42832# 0.039137f
C4231 a_18287_44626# a_20362_44736# 5.63e-20
C4232 a_8696_44636# a_14205_43396# 8.74e-22
C4233 a_10193_42453# a_743_42282# 1.1645f
C4234 a_5708_44484# a_n2661_43922# 0.004801f
C4235 a_8953_45002# a_9165_43940# 4.13e-20
C4236 a_3357_43084# a_3080_42308# 0.233522f
C4237 a_n967_45348# a_n1177_43370# 0.013627f
C4238 a_n2017_45002# VDD 3.8321f
C4239 a_22400_42852# a_22780_40945# 2e-19
C4240 a_9028_43914# a_4883_46098# 0.002203f
C4241 a_15493_43396# a_16327_47482# 0.025969f
C4242 a_22223_43948# a_12861_44030# 0.001164f
C4243 a_7229_43940# a_6945_45028# 0.001224f
C4244 a_7845_44172# a_n1613_43370# 5.96e-21
C4245 a_13777_45326# a_2324_44458# 0.002856f
C4246 a_14537_43396# a_15015_46420# 1.61e-20
C4247 a_14797_45144# a_14275_46494# 1.37e-19
C4248 a_1667_45002# a_526_44458# 2.21e-19
C4249 a_19256_45572# a_19443_46116# 2.91e-19
C4250 a_19237_31679# a_21588_30879# 0.055917f
C4251 a_n2661_43922# a_5257_43370# 0.030003f
C4252 a_17767_44458# a_3090_45724# 1.66e-19
C4253 a_2675_43914# a_768_44030# 0.026212f
C4254 a_5837_45028# a_4185_45028# 1.38e-19
C4255 a_17023_45118# a_12741_44636# 0.005061f
C4256 a_18315_45260# a_11415_45002# 0.00724f
C4257 a_8325_42308# a_5742_30871# 1.69e-20
C4258 a_9223_42460# a_10533_42308# 4.9e-20
C4259 COMP_P a_21613_42308# 1.34e-20
C4260 a_n923_35174# VIN_P 1.547f
C4261 C5_P_btm C3_P_btm 0.135528f
C4262 C6_P_btm C2_P_btm 0.137206f
C4263 a_16327_47482# a_3483_46348# 0.003076f
C4264 a_4915_47217# a_12594_46348# 3.27e-20
C4265 a_9313_45822# a_8199_44636# 0.015956f
C4266 a_n2497_47436# a_n1533_46116# 0.006317f
C4267 a_n1151_42308# a_2324_44458# 0.075066f
C4268 a_n237_47217# a_6945_45028# 0.072758f
C4269 a_5807_45002# a_16721_46634# 0.112018f
C4270 a_13747_46662# a_13059_46348# 0.273684f
C4271 a_7715_46873# a_7577_46660# 0.205227f
C4272 a_7411_46660# a_8145_46902# 0.053385f
C4273 a_4817_46660# a_6999_46987# 1.63e-20
C4274 a_4646_46812# a_7832_46660# 3.69e-20
C4275 a_5907_46634# a_6755_46942# 5.62e-20
C4276 a_5257_43370# a_7927_46660# 7.79e-22
C4277 a_13661_43548# a_16388_46812# 2.4e-20
C4278 a_13569_47204# a_765_45546# 7.71e-19
C4279 a_12549_44172# a_19551_46910# 1.88e-19
C4280 a_19778_44110# a_19700_43370# 0.009715f
C4281 a_22959_44484# a_22959_43948# 0.026152f
C4282 a_n2293_43922# a_n2129_43609# 0.028035f
C4283 a_n2661_42834# a_n1699_43638# 0.00613f
C4284 a_n2661_43922# a_n2267_43396# 1.14e-20
C4285 a_11827_44484# a_17499_43370# 3.5e-20
C4286 a_18494_42460# a_15743_43084# 0.027791f
C4287 a_18184_42460# a_19268_43646# 1.21e-21
C4288 a_1307_43914# a_5111_42852# 2.66e-19
C4289 a_7542_44172# a_7911_44260# 0.00411f
C4290 a_n356_44636# a_3626_43646# 0.073377f
C4291 a_5343_44458# a_8229_43396# 0.00134f
C4292 a_11691_44458# a_16547_43609# 4.26e-20
C4293 a_16237_45028# a_16137_43396# 5.13e-20
C4294 a_n1059_45260# a_133_42852# 0.045134f
C4295 en_comp a_n2293_42282# 0.026f
C4296 a_n913_45002# a_n914_42852# 9.04e-20
C4297 a_n89_44484# VDD 6.07e-19
C4298 a_n4064_39072# VIN_P 0.039352f
C4299 a_n4064_38528# C5_P_btm 0.042017f
C4300 a_n3565_39304# VCM 0.035438f
C4301 a_2711_45572# a_6428_45938# 1.42e-19
C4302 a_895_43940# a_1138_42852# 0.017458f
C4303 a_2479_44172# a_1823_45246# 7.38e-19
C4304 a_14955_43396# a_13661_43548# 3.87e-20
C4305 a_17973_43940# a_17339_46660# 8.68e-20
C4306 a_4699_43561# a_4646_46812# 2.54e-20
C4307 a_14021_43940# a_19692_46634# 0.775991f
C4308 a_15037_44260# a_15227_44166# 6.14e-19
C4309 a_6809_43396# a_n2293_46634# 3.99e-19
C4310 a_949_44458# a_n357_42282# 0.016511f
C4311 a_742_44458# a_n755_45592# 3e-20
C4312 a_5883_43914# a_n2661_45546# 3.15e-21
C4313 a_11967_42832# a_18189_46348# 2.07e-20
C4314 a_16823_43084# a_11453_44696# 7.31e-22
C4315 a_10835_43094# a_2063_45854# 8.1e-21
C4316 en_comp a_22521_40055# 0.260972f
C4317 a_n3420_38528# a_n4064_38528# 8.203589f
C4318 a_n3565_38502# a_n2860_38778# 2.96e-19
C4319 a_2112_39137# a_2684_37794# 0.091415f
C4320 a_4958_30871# C4_N_btm 1.18e-19
C4321 a_20202_43084# a_11415_45002# 0.041726f
C4322 a_765_45546# a_2202_46116# 4.62e-20
C4323 a_22365_46825# a_22591_46660# 0.08571f
C4324 a_768_44030# a_2277_45546# 0.027945f
C4325 a_n2661_46634# a_n1079_45724# 4.39e-21
C4326 a_7411_46660# a_5066_45546# 7.26e-20
C4327 a_n2312_38680# a_n2810_45572# 0.062154f
C4328 a_5257_43370# a_6419_46482# 0.006417f
C4329 a_n2293_46634# a_n2472_45546# 1.2e-19
C4330 a_n2442_46660# a_n2956_38216# 0.048086f
C4331 a_8270_45546# a_6945_45028# 3.18e-19
C4332 a_15009_46634# a_14840_46494# 0.001393f
C4333 a_3090_45724# a_15015_46420# 0.019425f
C4334 COMP_P a_3754_38470# 4.61e-19
C4335 a_n2065_43946# a_n901_43156# 6.54e-19
C4336 a_n1549_44318# a_n1853_43023# 7.93e-21
C4337 a_5495_43940# a_743_42282# 7.52e-22
C4338 a_14673_44172# a_5534_30871# 1.22e-19
C4339 a_15493_43396# a_10341_43396# 0.039468f
C4340 a_n1761_44111# a_n1641_43230# 2.7e-21
C4341 a_n2433_43396# a_104_43370# 2.99e-21
C4342 a_n1331_43914# a_n1991_42858# 3.18e-20
C4343 a_n1699_43638# a_n1352_43396# 0.051162f
C4344 a_n4318_39304# a_n2012_43396# 1.24e-19
C4345 a_n2129_43609# a_n97_42460# 3.26e-19
C4346 a_11967_42832# a_10518_42984# 5.09e-21
C4347 a_2998_44172# a_4361_42308# 9.12e-22
C4348 a_15493_43940# a_9145_43396# 3.68e-19
C4349 a_5111_44636# a_7174_31319# 4.88e-21
C4350 a_n2956_37592# a_n3690_39616# 1.91e-20
C4351 a_n2810_45028# a_n3420_39616# 2.09e-19
C4352 en_comp a_n3565_39590# 4.23e-19
C4353 a_21845_43940# VDD 0.00416f
C4354 a_13904_45546# a_13556_45296# 4.14e-19
C4355 a_13249_42308# a_9482_43914# 0.061734f
C4356 a_13527_45546# a_13777_45326# 4.75e-19
C4357 a_20107_45572# a_20841_45814# 0.053479f
C4358 a_8697_45572# a_6171_45002# 3.24e-19
C4359 a_8685_43396# a_8953_45546# 0.062741f
C4360 a_6197_43396# a_2324_44458# 0.001135f
C4361 a_11341_43940# a_n357_42282# 1.86e-19
C4362 a_14021_43940# a_20692_30879# 1.18e-20
C4363 a_15682_43940# a_n443_42852# 0.002992f
C4364 a_8037_42858# a_3090_45724# 1.28e-20
C4365 a_14955_43396# a_4185_45028# 3.39e-21
C4366 a_19268_43646# a_12741_44636# 3.85e-21
C4367 a_10341_43396# a_3483_46348# 2.31e-19
C4368 a_526_44458# VDD 2.35177f
C4369 a_10193_42453# a_6151_47436# 5.26e-20
C4370 a_13527_45546# a_n1151_42308# 1.73e-20
C4371 a_5204_45822# a_n755_45592# 2.71e-20
C4372 a_15682_46116# a_16375_45002# 6.09e-19
C4373 a_18189_46348# a_13259_45724# 0.016675f
C4374 a_4419_46090# a_3218_45724# 4.98e-22
C4375 a_1823_45246# a_n443_42852# 0.125287f
C4376 a_3699_46348# a_3503_45724# 1.91e-19
C4377 a_5495_43940# a_5755_42308# 4.04e-22
C4378 a_5244_44056# a_5932_42308# 1.08e-21
C4379 a_7287_43370# a_7765_42852# 0.002031f
C4380 a_17324_43396# a_16823_43084# 0.038999f
C4381 a_2813_43396# a_2905_42968# 5.2e-19
C4382 a_3626_43646# a_12379_42858# 1.5e-19
C4383 a_2982_43646# a_12545_42858# 9.98e-20
C4384 a_16137_43396# a_743_42282# 0.183525f
C4385 a_n2661_42282# a_1184_42692# 9.09e-20
C4386 a_3422_30871# a_15051_42282# 4.65e-20
C4387 a_n2293_43922# a_n2302_40160# 1.25e-19
C4388 a_3080_42308# a_5342_30871# 0.01896f
C4389 a_15743_43084# a_15940_43402# 0.00103f
C4390 a_11967_42832# a_16197_42308# 1.01e-20
C4391 a_19164_43230# VDD 0.278643f
C4392 a_8696_44636# a_9159_44484# 9.98e-20
C4393 a_413_45260# a_n2661_44458# 0.69469f
C4394 a_6171_45002# a_11691_44458# 0.022104f
C4395 a_n2017_45002# a_n699_43396# 4.86e-20
C4396 a_n967_45348# a_n1177_44458# 0.012502f
C4397 a_n467_45028# a_n2267_44484# 3.24e-21
C4398 a_15890_42674# a_15227_44166# 0.001386f
C4399 a_n901_43156# a_n755_45592# 1.1e-19
C4400 a_n1076_43230# a_n357_42282# 0.001306f
C4401 a_7754_38470# w_11334_34010# 2.62e-19
C4402 a_15415_45028# a_11453_44696# 0.005374f
C4403 a_5205_44484# a_n881_46662# 0.013688f
C4404 a_11823_42460# a_14976_45028# 0.010375f
C4405 a_2711_45572# a_765_45546# 5.89e-20
C4406 a_10903_43370# CLK 0.018377f
C4407 a_743_42282# a_n784_42308# 0.087438f
C4408 a_8685_43396# a_14456_42282# 4.62e-21
C4409 a_3626_43646# a_18727_42674# 0.003134f
C4410 a_2982_43646# a_19332_42282# 2.01e-19
C4411 a_n4318_39304# a_n4064_39616# 0.059009f
C4412 a_10835_43094# a_10793_43218# 2.56e-19
C4413 a_9145_43396# a_5742_30871# 8.14e-20
C4414 a_15682_46116# RST_Z 8.37e-21
C4415 a_n1741_47186# a_9804_47204# 0.010096f
C4416 a_n971_45724# a_n881_46662# 0.236696f
C4417 a_4915_47217# a_12465_44636# 0.07724f
C4418 a_n746_45260# a_n1613_43370# 0.146842f
C4419 a_5815_47464# a_4883_46098# 4.29e-21
C4420 a_11599_46634# a_15811_47375# 0.107881f
C4421 a_14955_47212# a_15673_47210# 3.17e-19
C4422 a_2553_47502# a_2747_46873# 0.14563f
C4423 a_13717_47436# a_16763_47508# 2.89e-19
C4424 a_11459_47204# a_10227_46804# 6.22e-20
C4425 a_12861_44030# a_16023_47582# 2.79e-20
C4426 a_22223_45036# a_17517_44484# 1.7e-20
C4427 a_n2267_44484# a_n2661_43922# 0.010057f
C4428 a_n2129_44697# a_n2293_43922# 3.05e-19
C4429 a_9838_44484# a_5891_43370# 1.24e-20
C4430 a_11691_44458# a_14673_44172# 0.371587f
C4431 a_1423_45028# a_5244_44056# 1.01e-20
C4432 a_1307_43914# a_7542_44172# 0.022371f
C4433 a_5343_44458# a_9313_44734# 6.56e-21
C4434 a_16922_45042# a_20640_44752# 4.09e-19
C4435 a_18315_45260# a_11967_42832# 3.09e-19
C4436 a_11827_44484# a_18204_44850# 1.18e-19
C4437 a_n1699_44726# a_n2661_42834# 0.002084f
C4438 a_3232_43370# a_9028_43914# 1.62e-19
C4439 a_n1059_45260# a_15493_43940# 1.89e-19
C4440 a_n913_45002# a_22223_43948# 3.74e-21
C4441 a_7229_43940# a_6756_44260# 5.36e-21
C4442 a_n4064_39072# a_n2956_38680# 0.001709f
C4443 a_n2302_39072# a_n2956_39304# 0.040755f
C4444 a_10723_42308# a_n357_42282# 7.12e-20
C4445 a_5934_30871# a_n443_42852# 1.89e-19
C4446 a_5534_30871# EN_VIN_BSTR_P 0.007335f
C4447 a_13017_45260# a_11415_45002# 0.100288f
C4448 a_2274_45254# a_167_45260# 8.13e-20
C4449 a_2680_45002# a_1823_45246# 0.073588f
C4450 a_n2661_43922# a_5807_45002# 1.32e-19
C4451 a_8375_44464# a_n1925_46634# 1.53e-21
C4452 a_16321_45348# a_14976_45028# 2.16e-20
C4453 a_10809_44484# a_768_44030# 1.65e-19
C4454 a_15143_45578# a_13259_45724# 0.060775f
C4455 a_3733_45822# a_n755_45592# 4.98e-19
C4456 a_10216_45572# a_10586_45546# 1.7e-19
C4457 a_19431_45546# a_10809_44734# 5.65e-21
C4458 a_3357_43084# a_11133_46155# 1.78e-21
C4459 a_20512_43084# a_18479_47436# 1.2e-19
C4460 a_21073_44484# a_18597_46090# 6.09e-19
C4461 a_n875_44318# a_n1151_42308# 5.38e-21
C4462 a_1755_42282# a_2903_42308# 5e-19
C4463 a_2123_42473# a_2713_42308# 6.03e-20
C4464 a_1606_42308# a_3318_42354# 1.73e-19
C4465 a_n784_42308# a_5755_42308# 3.86e-20
C4466 a_14635_42282# a_15890_42674# 7.2e-22
C4467 a_5807_45002# a_7927_46660# 0.004378f
C4468 a_n2661_46634# a_6540_46812# 0.007418f
C4469 a_n743_46660# a_4646_46812# 0.031686f
C4470 a_n1925_46634# a_4955_46873# 0.033508f
C4471 a_2107_46812# a_2864_46660# 0.002314f
C4472 a_n2438_43548# a_3877_44458# 2.1e-20
C4473 a_768_44030# a_6755_46942# 0.017611f
C4474 a_645_46660# a_n2661_46098# 2.43e-19
C4475 a_8128_46384# a_8035_47026# 0.006018f
C4476 a_n881_46662# a_8023_46660# 0.001443f
C4477 a_11453_44696# a_15368_46634# 6.42e-20
C4478 a_13507_46334# a_19692_46634# 0.823157f
C4479 a_4883_46098# a_19333_46634# 6.67e-20
C4480 a_11599_46634# a_13059_46348# 0.371555f
C4481 a_10227_46804# a_12925_46660# 0.001202f
C4482 a_9313_45822# a_765_45546# 0.034184f
C4483 a_12861_44030# a_16751_46987# 7.13e-19
C4484 a_n746_45260# a_n2293_46098# 0.027821f
C4485 a_n1741_47186# a_n901_46420# 1.81e-20
C4486 a_n971_45724# a_n2157_46122# 0.001149f
C4487 a_2063_45854# a_11415_45002# 5.51e-19
C4488 a_n1899_43946# a_n1549_44318# 0.218775f
C4489 a_n2065_43946# a_n984_44318# 0.102325f
C4490 a_n1761_44111# a_n809_44244# 0.038277f
C4491 a_11823_42460# a_13157_43218# 5.05e-19
C4492 en_comp a_n1423_42826# 1.04e-20
C4493 a_n967_45348# a_n1991_42858# 0.034664f
C4494 a_n913_45002# a_n13_43084# 0.042137f
C4495 a_n2017_45002# a_n4318_38680# 1.48e-19
C4496 a_3357_43084# a_2075_43172# 8.43e-21
C4497 a_n3690_37440# VDD 0.363068f
C4498 a_n2840_44458# VDD 0.247948f
C4499 a_17124_42282# RST_Z 4.07e-20
C4500 a_4958_30871# C6_P_btm 0.005441f
C4501 a_13678_32519# w_11334_34010# 3.98e-19
C4502 a_13076_44458# a_10809_44734# 1.02e-19
C4503 a_18374_44850# a_17957_46116# 8.91e-21
C4504 a_4223_44672# a_n1925_42282# 0.053508f
C4505 a_18315_45260# a_13259_45724# 0.144632f
C4506 a_17023_45118# a_16375_45002# 0.014031f
C4507 a_n699_43396# a_526_44458# 0.285f
C4508 a_9801_43940# a_2107_46812# 3.07e-19
C4509 a_1209_43370# a_768_44030# 1.23e-20
C4510 a_n2661_42834# a_4185_45028# 0.023267f
C4511 a_17061_44484# a_12741_44636# 1.5e-19
C4512 a_11967_42832# a_20202_43084# 0.02752f
C4513 a_8746_45002# CLK 0.018523f
C4514 a_n4334_40480# a_n4064_39616# 7.84e-19
C4515 a_n4209_39590# a_n4334_39616# 0.25243f
C4516 a_n4064_40160# a_n2946_39866# 1.91e-19
C4517 a_n4315_30879# a_n2302_39866# 9.79e-19
C4518 a_13759_47204# VDD 0.004261f
C4519 a_1606_42308# C10_N_btm 1.34e-19
C4520 a_5257_43370# a_5164_46348# 0.02844f
C4521 a_5732_46660# a_5937_45572# 1.49e-19
C4522 a_13507_46334# a_20692_30879# 6.68e-19
C4523 a_4883_46098# a_20062_46116# 9.7e-20
C4524 a_16327_47482# a_n357_42282# 0.49929f
C4525 a_8667_46634# a_3483_46348# 7.36e-19
C4526 a_15227_44166# a_22000_46634# 0.154332f
C4527 a_19692_46634# a_20623_46660# 0.03624f
C4528 a_13885_46660# a_14447_46660# 0.005162f
C4529 a_16292_46812# a_16434_46660# 0.007833f
C4530 a_14035_46660# a_14226_46660# 2.88e-19
C4531 a_13693_46688# a_13059_46348# 1.71e-19
C4532 a_768_44030# a_8049_45260# 0.027975f
C4533 a_5807_45002# a_6419_46482# 0.005524f
C4534 a_n2438_43548# a_n1736_46482# 2.63e-20
C4535 a_n1925_46634# a_n967_46494# 6.65e-20
C4536 a_13720_44458# a_13635_43156# 5.13e-21
C4537 a_15493_43396# a_n97_42460# 0.002057f
C4538 a_n2661_42834# a_n2157_42858# 0.001323f
C4539 a_n2661_43922# a_n2472_42826# 7.7e-20
C4540 a_3499_42826# a_3539_42460# 0.00342f
C4541 a_n356_44636# a_8037_42858# 3.48e-20
C4542 a_375_42282# a_n3674_37592# 0.003119f
C4543 a_5111_44636# a_5932_42308# 0.021257f
C4544 a_n1059_45260# a_5742_30871# 0.002047f
C4545 a_3537_45260# a_7227_42308# 0.001666f
C4546 a_n913_45002# a_11323_42473# 6.5e-19
C4547 a_n2017_45002# a_11551_42558# 0.006777f
C4548 a_18079_43940# VDD 0.162408f
C4549 a_16680_45572# a_8696_44636# 0.004839f
C4550 a_16855_45546# a_15861_45028# 0.001688f
C4551 a_15765_45572# a_16223_45938# 0.027606f
C4552 a_2711_45572# a_2382_45260# 1.81e-20
C4553 a_n97_42460# a_3483_46348# 1.02e-19
C4554 a_14358_43442# a_13059_46348# 0.041731f
C4555 a_16547_43609# a_15227_44166# 1.88e-20
C4556 a_453_43940# a_n863_45724# 0.02533f
C4557 a_n984_44318# a_n755_45592# 0.002789f
C4558 a_175_44278# a_n357_42282# 0.002018f
C4559 a_18707_42852# a_16327_47482# 0.012993f
C4560 a_6123_31319# w_11334_34010# 6.03e-19
C4561 a_2521_46116# VDD 0.163553f
C4562 C4_N_btm C7_N_btm 0.145303f
C4563 C5_N_btm C6_N_btm 22.305399f
C4564 C1_N_btm C10_N_btm 0.31753f
C4565 C2_N_btm C9_N_btm 0.141891f
C4566 C3_N_btm C8_N_btm 0.134581f
C4567 a_20202_43084# a_13259_45724# 2.57e-19
C4568 a_4185_45028# a_5066_45546# 2.04e-20
C4569 a_17583_46090# a_18819_46122# 1.6e-21
C4570 a_17715_44484# a_17957_46116# 0.005313f
C4571 a_13759_46122# a_6945_45028# 7.74e-20
C4572 a_12594_46348# a_10809_44734# 0.082565f
C4573 a_n3565_38216# a_n3690_38304# 0.247167f
C4574 a_n4334_38304# a_n3420_37984# 0.004718f
C4575 a_n4209_38216# a_n2946_37984# 0.022779f
C4576 a_21115_43940# a_21195_42852# 2.21e-21
C4577 a_n2840_43370# a_n3674_39304# 0.008407f
C4578 a_n1917_43396# a_n1991_42858# 1.29e-19
C4579 a_n2267_43396# a_n1641_43230# 0.00175f
C4580 a_n1352_43396# a_n2157_42858# 5.11e-19
C4581 a_n1177_43370# a_n1853_43023# 1.6e-19
C4582 a_3080_42308# a_743_42282# 0.069641f
C4583 a_10695_43548# a_10341_43396# 0.008043f
C4584 a_n1699_43638# a_n1423_42826# 5.89e-19
C4585 a_n2129_43609# a_n901_43156# 0.001317f
C4586 a_14021_43940# a_5342_30871# 0.001922f
C4587 a_15493_43940# a_19987_42826# 7.44e-20
C4588 a_11341_43940# a_21356_42826# 4.25e-20
C4589 a_n2293_43922# a_8791_42308# 8.6e-20
C4590 a_9313_44734# a_12563_42308# 2.09e-20
C4591 a_9145_43396# a_10849_43646# 0.003354f
C4592 a_n2661_42282# a_5193_42852# 2.87e-21
C4593 a_14579_43548# a_14955_43396# 4.82e-20
C4594 a_8685_43396# a_10149_43396# 7.5e-19
C4595 a_n2312_40392# CLK_DATA 0.213071f
C4596 a_4883_46098# CLK 0.032195f
C4597 a_14209_32519# VDD 0.284433f
C4598 a_8568_45546# a_5891_43370# 4.55e-19
C4599 a_6511_45714# a_n2661_43922# 6.22e-21
C4600 a_18909_45814# a_11691_44458# 7.74e-19
C4601 a_18691_45572# a_19113_45348# 0.001513f
C4602 a_13017_45260# a_13159_45002# 0.160415f
C4603 a_11787_45002# a_9482_43914# 8.24e-21
C4604 a_7499_43078# a_8375_44464# 2.35e-19
C4605 a_2711_45572# a_15433_44458# 2.54e-20
C4606 a_9049_44484# a_7640_43914# 7.12e-20
C4607 a_5111_44636# a_1423_45028# 0.028542f
C4608 a_5205_44484# a_1307_43914# 0.006798f
C4609 a_n1059_45260# a_n2293_42834# 0.035031f
C4610 a_3429_45260# a_3495_45348# 0.010598f
C4611 a_n143_45144# a_45_45144# 7.47e-21
C4612 a_3065_45002# a_3602_45348# 5.93e-19
C4613 a_5534_30871# a_10903_43370# 0.134296f
C4614 a_7221_43396# a_n443_42852# 1.62e-19
C4615 a_10341_43396# a_n357_42282# 9.55e-19
C4616 a_8696_44636# a_13747_46662# 0.02273f
C4617 a_17478_45572# a_5807_45002# 1.08e-20
C4618 a_2711_45572# a_10623_46897# 8.62e-20
C4619 a_15861_45028# a_13661_43548# 0.047089f
C4620 a_14127_45572# a_768_44030# 0.002434f
C4621 a_3357_43084# a_13507_46334# 0.050295f
C4622 a_2437_43646# a_21811_47423# 0.025192f
C4623 a_21542_45572# a_18597_46090# 4.51e-19
C4624 a_413_45260# a_13717_47436# 4.36729f
C4625 a_10775_45002# a_n1151_42308# 7.13e-22
C4626 a_1307_43914# a_n971_45724# 0.019541f
C4627 a_7276_45260# a_4791_45118# 0.004255f
C4628 a_n755_45592# a_3503_45724# 0.163919f
C4629 a_n2293_45546# a_n443_42852# 0.084694f
C4630 a_n357_42282# a_n356_45724# 2.1e-19
C4631 a_n863_45724# a_n906_45572# 0.002589f
C4632 a_310_45028# a_n23_45546# 0.022295f
C4633 a_n1099_45572# a_n310_45899# 4.53e-19
C4634 a_6293_42852# a_1755_42282# 1.75e-19
C4635 a_n2157_42858# a_n2293_42282# 5.22e-20
C4636 a_10083_42826# a_10835_43094# 0.043619f
C4637 a_3539_42460# a_3318_42354# 0.161793f
C4638 a_3626_43646# a_3823_42558# 0.017529f
C4639 a_2982_43646# a_5379_42460# 0.068435f
C4640 a_n97_42460# a_8791_42308# 4.89e-19
C4641 a_14021_43940# a_20107_42308# 2.15e-20
C4642 a_4905_42826# a_5421_42558# 0.002476f
C4643 a_8952_43230# a_10796_42968# 2e-20
C4644 a_16137_43396# a_16328_43172# 5.93e-19
C4645 a_22000_46634# EN_OFFSET_CAL 3.46e-20
C4646 a_2063_45854# a_2553_47502# 0.040297f
C4647 a_n971_45724# a_n443_46116# 0.129009f
C4648 a_1239_47204# a_n1151_42308# 0.007713f
C4649 a_1209_47178# a_3381_47502# 7.34e-20
C4650 a_n1741_47186# a_6545_47178# 0.053219f
C4651 a_18587_45118# a_18374_44850# 9.02e-19
C4652 a_n2661_43370# a_5891_43370# 3.67e-19
C4653 a_n2661_44458# a_2779_44458# 0.011596f
C4654 a_11691_44458# a_12607_44458# 0.042423f
C4655 a_11827_44484# a_15004_44636# 0.007895f
C4656 a_19778_44110# a_18287_44626# 5.65e-21
C4657 a_n1699_44726# a_n1352_44484# 0.051162f
C4658 a_14537_43396# a_16241_44484# 0.003767f
C4659 a_413_45260# a_19237_31679# 0.119197f
C4660 a_n1059_45260# a_1115_44172# 2.41e-21
C4661 a_3357_43084# a_5013_44260# 2.89e-19
C4662 a_n967_45348# a_n1331_43914# 0.003919f
C4663 a_n2293_45010# a_453_43940# 0.181603f
C4664 a_n2661_45010# a_2479_44172# 7.5e-19
C4665 a_n3674_38216# a_n2956_38216# 0.028821f
C4666 a_5742_30871# a_n1925_42282# 5.06e-20
C4667 COMP_P a_n2810_45572# 2.2e-21
C4668 a_20356_42852# a_n357_42282# 0.001192f
C4669 a_7174_31319# a_9290_44172# 2.43e-20
C4670 a_4099_45572# VDD 0.296272f
C4671 a_4190_30871# EN_VIN_BSTR_P 0.043599f
C4672 a_14209_32519# a_22469_39537# 1.36e-20
C4673 a_13213_44734# a_12861_44030# 0.002516f
C4674 a_20273_45572# a_20202_43084# 0.003019f
C4675 a_9313_44734# a_10227_46804# 0.875947f
C4676 a_11652_45724# a_6945_45028# 2.08e-20
C4677 a_11322_45546# a_10809_44734# 0.22629f
C4678 a_413_45260# a_14035_46660# 2.37e-20
C4679 a_6171_45002# a_15227_44166# 0.021072f
C4680 a_8191_45002# a_3090_45724# 7.02e-22
C4681 a_2437_43646# a_22000_46634# 0.010034f
C4682 a_3357_43084# a_20623_46660# 0.013905f
C4683 a_2711_45572# a_6347_46155# 1.62e-19
C4684 a_5024_45822# a_526_44458# 1.2e-19
C4685 a_6667_45809# a_5066_45546# 1.76e-19
C4686 a_8103_44636# a_768_44030# 0.004654f
C4687 a_5837_45028# a_5257_43370# 0.008516f
C4688 a_n2661_43370# a_4817_46660# 6.7e-21
C4689 a_20107_45572# a_11415_45002# 0.019157f
C4690 a_15567_42826# a_15486_42560# 1.56e-19
C4691 a_20256_43172# a_20256_42852# 9.31e-19
C4692 a_5342_30871# a_15764_42576# 0.002004f
C4693 a_5837_42852# a_5379_42460# 4.94e-19
C4694 a_5837_43172# a_5932_42308# 3.37e-21
C4695 a_n881_46662# a_601_46902# 4.24e-19
C4696 a_n1613_43370# a_383_46660# 0.182504f
C4697 a_2747_46873# a_1799_45572# 5.65e-19
C4698 a_6151_47436# a_8035_47026# 0.038687f
C4699 a_6575_47204# a_6969_46634# 2.23e-19
C4700 a_n1435_47204# a_10150_46912# 1.49e-20
C4701 a_9067_47204# a_6755_46942# 1.22e-19
C4702 a_11459_47204# a_10467_46802# 4.67e-19
C4703 a_n1151_42308# a_11186_47026# 4.42e-20
C4704 a_2063_45854# a_12251_46660# 2.19e-19
C4705 a_5807_45002# a_19594_46812# 1.59e-19
C4706 a_13661_43548# a_19321_45002# 7.35e-19
C4707 a_12549_44172# a_n2293_46634# 0.005061f
C4708 a_13747_46662# a_19452_47524# 0.003322f
C4709 a_9804_47204# a_n743_46660# 0.295465f
C4710 a_10440_44484# a_10405_44172# 0.001304f
C4711 a_n2293_43922# a_n2472_43914# 0.189122f
C4712 a_n2661_43922# a_n2065_43946# 0.013023f
C4713 a_n2661_42834# a_n1761_44111# 0.073205f
C4714 a_8975_43940# a_9028_43914# 0.184602f
C4715 a_10057_43914# a_9672_43914# 0.143523f
C4716 a_1307_43914# a_1427_43646# 2.4e-19
C4717 a_11823_42460# a_12089_42308# 0.335983f
C4718 a_19006_44850# a_11967_42832# 0.013801f
C4719 a_18479_45785# a_743_42282# 7.51e-20
C4720 a_7705_45326# a_7287_43370# 9.03e-21
C4721 a_3537_45260# a_6643_43396# 0.001481f
C4722 a_5147_45002# a_5565_43396# 2.01e-22
C4723 a_n784_42308# VIN_P 0.004358f
C4724 a_2779_44458# a_2804_46116# 9.85e-20
C4725 a_18248_44752# a_12741_44636# 0.00762f
C4726 a_18374_44850# a_11415_45002# 6.96e-20
C4727 a_5518_44484# a_1823_45246# 4.84e-19
C4728 a_14673_44172# a_15227_44166# 0.357896f
C4729 a_20365_43914# a_13747_46662# 1.31e-20
C4730 a_12429_44172# a_n2293_46634# 9.2e-20
C4731 a_19862_44208# a_19321_45002# 0.090113f
C4732 a_9313_44734# a_17339_46660# 2.43e-19
C4733 a_11173_44260# a_768_44030# 0.005635f
C4734 a_13017_45260# a_13259_45724# 0.078313f
C4735 a_n2293_42834# a_n1925_42282# 0.024873f
C4736 a_413_45260# a_n1099_45572# 0.008675f
C4737 a_327_44734# a_380_45546# 6.27e-19
C4738 a_n37_45144# a_310_45028# 0.112458f
C4739 a_3537_45260# a_n2661_45546# 0.780422f
C4740 a_n467_45028# a_n755_45592# 0.26002f
C4741 a_2274_45254# a_n863_45724# 0.17549f
C4742 a_n2661_45010# a_n443_42852# 0.001666f
C4743 a_2680_45002# a_n2293_45546# 3.47e-20
C4744 a_11827_44484# a_13759_46122# 4.47e-21
C4745 a_11691_44458# a_10903_43370# 0.020718f
C4746 a_n2661_44458# a_6165_46155# 1.3e-22
C4747 a_17719_45144# a_17957_46116# 4.95e-21
C4748 a_18315_45260# a_18189_46348# 0.101775f
C4749 a_21381_43940# a_18479_47436# 8.4e-20
C4750 a_21205_44306# a_18597_46090# 6.68e-19
C4751 a_1427_43646# a_n443_46116# 0.05874f
C4752 a_9396_43370# a_n971_45724# 2.62e-20
C4753 a_1512_43396# a_584_46384# 7.9e-20
C4754 a_17124_42282# a_17303_42282# 0.172579f
C4755 a_15051_42282# a_7174_31319# 6.09e-20
C4756 a_5934_30871# a_1736_39587# 8.81e-20
C4757 a_n1630_35242# a_n3565_38216# 1.42e-19
C4758 a_15521_42308# a_4958_30871# 1.44e-19
C4759 a_5742_30871# a_n4315_30879# 9.24e-21
C4760 a_13381_47204# VDD 0.130765f
C4761 a_n2438_43548# a_n1641_46494# 4.44e-20
C4762 a_n2661_46634# a_1823_45246# 3e-19
C4763 a_n1925_46634# a_376_46348# 0.002206f
C4764 a_n743_46660# a_n901_46420# 0.004763f
C4765 a_n1021_46688# a_n1076_46494# 3.41e-20
C4766 a_171_46873# a_n1991_46122# 7.76e-21
C4767 a_11735_46660# a_13607_46688# 1.3e-20
C4768 a_12469_46902# a_12251_46660# 0.209641f
C4769 a_11901_46660# a_12991_46634# 0.042415f
C4770 a_6540_46812# a_765_45546# 0.00357f
C4771 a_10249_46116# a_12978_47026# 4.67e-21
C4772 a_11813_46116# a_12816_46660# 5.47e-21
C4773 a_6755_46942# a_10933_46660# 5.53e-19
C4774 a_768_44030# a_8953_45546# 0.025581f
C4775 a_5807_45002# a_5164_46348# 5.51e-19
C4776 a_9804_47204# a_11189_46129# 2.45e-20
C4777 a_n881_46662# a_12594_46348# 1.17e-19
C4778 a_22223_47212# a_22223_46124# 8.8e-19
C4779 a_12465_44636# a_10809_44734# 0.099854f
C4780 a_22731_47423# a_6945_45028# 8.58e-20
C4781 a_9067_47204# a_8049_45260# 1.65e-19
C4782 a_n2497_47436# a_n2810_45572# 1.01e-20
C4783 a_n2833_47464# a_n2661_45546# 3.61e-20
C4784 a_n1899_43946# a_n1177_43370# 0.001333f
C4785 a_n984_44318# a_n2129_43609# 5.84e-20
C4786 a_20269_44172# a_20365_43914# 0.419086f
C4787 a_18326_43940# a_15493_43940# 0.075033f
C4788 a_19328_44172# a_11341_43940# 0.004787f
C4789 a_19862_44208# a_20623_43914# 0.023134f
C4790 a_10057_43914# a_743_42282# 4.3e-20
C4791 a_n1761_44111# a_n1352_43396# 1.05e-20
C4792 a_n2267_44484# a_n1641_43230# 7.05e-22
C4793 a_n2129_44697# a_n901_43156# 3.52e-20
C4794 a_10193_42453# a_13258_32519# 0.061618f
C4795 a_n4318_40392# a_n3674_39304# 0.024125f
C4796 a_1307_43914# a_3863_42891# 0.005265f
C4797 a_10949_43914# a_12710_44260# 0.001055f
C4798 a_5883_43914# a_4361_42308# 2.27e-20
C4799 a_14539_43914# a_17021_43396# 5.66e-19
C4800 a_n2017_45002# a_n2840_42282# 7.53e-19
C4801 en_comp a_14097_32519# 5.98e-20
C4802 a_20447_31679# COMP_P 4.66e-20
C4803 a_17730_32519# VDD 0.289738f
C4804 a_11525_45546# a_11682_45822# 0.18824f
C4805 a_10053_45546# a_10216_45572# 0.011381f
C4806 a_11962_45724# a_10907_45822# 2.36e-20
C4807 a_2711_45572# a_13385_45572# 6.27e-20
C4808 C3_N_btm C2_P_btm 1.33e-19
C4809 C4_N_btm C3_P_btm 1.02e-19
C4810 a_21356_42826# a_16327_47482# 0.003181f
C4811 a_10729_43914# a_9290_44172# 0.042243f
C4812 a_n2293_43922# a_n357_42282# 0.02281f
C4813 a_1467_44172# a_526_44458# 0.041836f
C4814 a_n2661_43922# a_n755_45592# 0.037767f
C4815 a_14209_32519# a_22612_30879# 0.059911f
C4816 a_3232_43370# CLK 2.72e-19
C4817 a_11415_45002# a_17715_44484# 0.032854f
C4818 a_12741_44636# a_2324_44458# 0.019655f
C4819 a_3483_46348# a_5204_45822# 2.01e-19
C4820 a_3699_46348# a_5164_46348# 1.23e-21
C4821 a_20528_46660# a_10809_44734# 0.004492f
C4822 a_5742_30871# a_n3420_37440# 0.004591f
C4823 a_4419_46090# a_4704_46090# 0.016592f
C4824 a_15493_43940# a_22959_43396# 3.06e-19
C4825 a_14673_44172# a_14635_42282# 0.002024f
C4826 a_4699_43561# a_3457_43396# 9.15e-20
C4827 a_2982_43646# a_7287_43370# 6.68e-21
C4828 a_548_43396# a_648_43396# 0.005294f
C4829 a_14021_43940# a_743_42282# 0.002697f
C4830 a_3539_42460# a_6197_43396# 4.71e-21
C4831 a_11967_42832# a_10793_43218# 1.94e-21
C4832 a_5343_44458# a_8515_42308# 9e-19
C4833 a_n1761_44111# a_n2293_42282# 8.68e-20
C4834 a_n356_44636# a_1149_42558# 2.72e-19
C4835 a_3080_42308# a_2813_43396# 9.02e-20
C4836 a_22223_43948# a_17364_32525# 6.31e-19
C4837 a_n237_47217# DATA[2] 7.36e-22
C4838 SMPL_ON_P VIN_P 0.587766f
C4839 a_n785_47204# DATA[0] 0.598846f
C4840 a_n23_47502# DATA[1] 1.93e-20
C4841 a_5263_45724# a_4223_44672# 7.35e-19
C4842 a_4099_45572# a_n699_43396# 9.59e-21
C4843 a_2711_45572# a_5343_44458# 3.61e-20
C4844 a_10193_42453# a_20193_45348# 0.305022f
C4845 a_8746_45002# a_11691_44458# 4.34e-20
C4846 a_n745_45366# a_n143_45144# 8.24e-19
C4847 a_n1059_45260# a_413_45260# 1.08e-19
C4848 a_7309_42852# a_3090_45724# 1e-19
C4849 a_18599_43230# a_17339_46660# 0.001489f
C4850 a_7227_42308# a_n2293_46634# 7.23e-22
C4851 a_6123_31319# a_n2442_46660# 6.51e-21
C4852 a_n447_43370# a_n755_45592# 0.017822f
C4853 a_n97_42460# a_n357_42282# 0.900712f
C4854 a_20107_42308# a_13507_46334# 5.01e-19
C4855 a_17730_32519# a_22469_39537# 1.95e-20
C4856 a_n452_45724# VDD 0.112977f
C4857 a_3357_43084# a_n1741_47186# 0.03857f
C4858 a_15765_45572# a_16327_47482# 0.048221f
C4859 a_8696_44636# a_11599_46634# 0.003698f
C4860 a_15037_45618# a_10227_46804# 0.012118f
C4861 a_16137_43396# a_15279_43071# 2.14e-19
C4862 a_n1853_43023# a_n1991_42858# 0.237526f
C4863 a_n2157_42858# a_n1423_42826# 0.07009f
C4864 a_10341_43396# a_21356_42826# 8.92e-20
C4865 a_2113_38308# VDAC_Pi 0.170908f
C4866 a_17749_42852# VDD 0.00742f
C4867 a_19431_45546# a_18579_44172# 2.71e-21
C4868 a_20107_45572# a_11967_42832# 6.49e-21
C4869 a_14797_45144# a_14539_43914# 1.54e-19
C4870 a_16922_45042# a_18184_42460# 0.028064f
C4871 a_7499_43078# a_10949_43914# 0.152939f
C4872 a_10180_45724# a_9672_43914# 9.13e-20
C4873 a_5111_44636# a_6109_44484# 0.003573f
C4874 a_3537_45260# a_8238_44734# 0.001272f
C4875 a_5934_30871# a_8199_44636# 0.159294f
C4876 a_945_42968# a_n863_45724# 0.003329f
C4877 a_3080_42308# VIN_P 0.025929f
C4878 a_13527_45546# a_12741_44636# 1.3e-21
C4879 a_14495_45572# a_11415_45002# 1.03e-19
C4880 a_3775_45552# a_4185_45028# 5.74e-20
C4881 a_18909_45814# a_15227_44166# 6.54e-21
C4882 a_18691_45572# a_18834_46812# 2.2e-20
C4883 a_5837_45028# a_5807_45002# 0.006254f
C4884 a_626_44172# a_n2438_43548# 0.025123f
C4885 a_18479_45785# a_19466_46812# 0.009818f
C4886 a_2903_45348# a_n2293_46634# 5.43e-19
C4887 a_n2661_43370# a_11309_47204# 8.95e-20
C4888 a_5147_45002# a_4651_46660# 3e-19
C4889 a_4558_45348# a_4955_46873# 2.33e-19
C4890 a_3537_45260# a_5385_46902# 8.42e-22
C4891 a_5111_44636# a_4646_46812# 0.078281f
C4892 a_4927_45028# a_3877_44458# 1.65e-20
C4893 a_6511_45714# a_5164_46348# 4.12e-21
C4894 a_2711_45572# a_8349_46414# 8.3e-21
C4895 a_5907_45546# a_6165_46155# 6.1e-19
C4896 a_11691_44458# a_4883_46098# 3.07e-20
C4897 a_n998_44484# a_n971_45724# 5.1e-19
C4898 a_19268_43646# a_17303_42282# 2.14e-21
C4899 a_22223_42860# a_22400_42852# 0.154104f
C4900 a_5649_42852# a_13575_42558# 6.94e-20
C4901 a_743_42282# a_15764_42576# 0.054445f
C4902 a_4190_30871# a_15959_42545# 6.15e-20
C4903 a_15743_43084# a_17531_42308# 2.2e-21
C4904 a_20922_43172# a_20753_42852# 0.08213f
C4905 a_22165_42308# a_14097_32519# 1.3e-19
C4906 a_18597_46090# a_12549_44172# 0.042681f
C4907 a_16241_47178# a_16131_47204# 0.097745f
C4908 a_15673_47210# a_5807_45002# 0.011029f
C4909 a_16327_47482# a_16942_47570# 0.001965f
C4910 a_12465_44636# a_n881_46662# 0.813228f
C4911 a_6545_47178# a_n743_46660# 0.003782f
C4912 a_6851_47204# a_n1925_46634# 6.48e-20
C4913 a_11031_47542# a_n2661_46634# 3.8e-20
C4914 a_13717_47436# a_20916_46384# 1.15e-19
C4915 a_n1151_42308# a_491_47026# 0.002342f
C4916 a_n746_45260# a_1057_46660# 6.69e-20
C4917 a_3815_47204# a_2107_46812# 4.62e-20
C4918 a_584_46384# a_n2661_46098# 0.17431f
C4919 a_2063_45854# a_1799_45572# 5.95e-19
C4920 a_n2109_47186# a_4651_46660# 0.025236f
C4921 a_n1741_47186# a_3877_44458# 1.26e-19
C4922 a_n1352_44484# a_n1761_44111# 1.85e-21
C4923 a_n1177_44458# a_n1899_43946# 7.1e-19
C4924 a_18374_44850# a_11967_42832# 0.053726f
C4925 a_18989_43940# a_19006_44850# 0.168452f
C4926 a_18287_44626# a_20159_44458# 5.37e-21
C4927 a_18248_44752# a_20362_44736# 2.99e-20
C4928 a_n2129_44697# a_n984_44318# 1.03e-20
C4929 a_n2661_44458# a_644_44056# 6.99e-20
C4930 a_n2661_43370# a_10807_43548# 7.36e-20
C4931 a_9313_44734# a_14815_43914# 1.48e-20
C4932 a_10193_42453# a_20301_43646# 2.72e-19
C4933 a_5608_44484# a_n2661_43922# 0.001386f
C4934 a_3357_43084# a_4699_43561# 0.002313f
C4935 a_n913_45002# a_104_43370# 2.19e-20
C4936 a_n2017_45002# a_n1809_43762# 0.003534f
C4937 a_n967_45348# a_n1917_43396# 9.47e-19
C4938 a_n4209_39304# a_n2810_45572# 0.020327f
C4939 a_n2109_45247# VDD 0.266396f
C4940 a_11341_43940# a_12861_44030# 0.064865f
C4941 a_19328_44172# a_16327_47482# 0.0072f
C4942 a_7276_45260# a_6945_45028# 0.00333f
C4943 a_7542_44172# a_n1613_43370# 0.007527f
C4944 a_1423_45028# a_9290_44172# 0.005536f
C4945 a_14537_43396# a_14275_46494# 9.72e-21
C4946 a_13556_45296# a_2324_44458# 0.026317f
C4947 a_413_45260# a_n1925_42282# 4.11e-20
C4948 a_21542_45572# a_8049_45260# 4.32e-19
C4949 a_327_44734# a_526_44458# 0.076983f
C4950 a_19431_45546# a_19443_46116# 1.05e-19
C4951 a_14539_43914# a_14976_45028# 2.57e-19
C4952 a_17730_32519# a_22612_30879# 0.060497f
C4953 a_n2661_42834# a_5257_43370# 0.01982f
C4954 a_895_43940# a_768_44030# 0.06559f
C4955 a_5093_45028# a_4185_45028# 9.16e-19
C4956 a_16922_45042# a_12741_44636# 0.139755f
C4957 a_17719_45144# a_11415_45002# 0.006388f
C4958 a_n784_42308# a_13258_32519# 0.140549f
C4959 a_9803_42558# a_9885_42558# 0.171361f
C4960 a_n1532_35090# VIN_P 0.066301f
C4961 C5_P_btm C4_P_btm 18.6196f
C4962 C7_P_btm C2_P_btm 0.138288f
C4963 C6_P_btm C3_P_btm 0.133742f
C4964 a_9067_47204# a_8953_45546# 0.00218f
C4965 SMPL_ON_P a_n2956_38680# 0.039338f
C4966 a_n1741_47186# a_n1736_46482# 1.99e-19
C4967 a_13661_43548# a_13059_46348# 0.267127f
C4968 a_5807_45002# a_16388_46812# 0.235518f
C4969 a_13747_46662# a_15227_46910# 5.38e-22
C4970 a_7411_46660# a_7577_46660# 0.634781f
C4971 a_4651_46660# a_5841_46660# 2.56e-19
C4972 a_4817_46660# a_6682_46987# 4.3e-20
C4973 a_3877_44458# a_7832_46660# 2.27e-20
C4974 a_12549_44172# a_19123_46287# 1.7e-19
C4975 a_n2293_43922# a_n2433_43396# 0.028793f
C4976 a_1307_43914# a_4520_42826# 6.56e-19
C4977 a_9482_43914# a_9127_43156# 4.2e-19
C4978 a_22959_44484# a_15493_43940# 3.35e-19
C4979 a_17730_32519# a_22959_43948# 0.00961f
C4980 a_n2661_42834# a_n2267_43396# 0.014077f
C4981 a_n2661_43922# a_n2129_43609# 1.04e-20
C4982 a_11691_44458# a_16243_43396# 4.28e-20
C4983 a_18184_42460# a_15743_43084# 0.182123f
C4984 a_18494_42460# a_18783_43370# 4.06e-21
C4985 a_7542_44172# a_7584_44260# 0.009099f
C4986 a_n2017_45002# a_133_42852# 0.001378f
C4987 en_comp a_22959_42860# 1.14e-21
C4988 a_n2956_37592# a_n2293_42282# 1.77e-20
C4989 a_n1059_45260# a_n914_42852# 6.52e-20
C4990 a_n310_44484# VDD 7.01e-20
C4991 a_n3420_38528# C4_P_btm 0.030945f
C4992 a_n4064_38528# C6_P_btm 0.001467f
C4993 a_n3565_39304# VREF_GND 0.010456f
C4994 a_2711_45572# a_4880_45572# 0.006167f
C4995 a_6598_45938# a_7227_45028# 1.78e-20
C4996 a_2479_44172# a_1138_42852# 4.8e-21
C4997 a_7542_44172# a_n2293_46098# 5.6e-21
C4998 a_n4318_39768# a_n2840_46090# 9.97e-22
C4999 a_14761_44260# a_15227_44166# 7.89e-21
C5000 a_15095_43370# a_13661_43548# 1.48e-20
C5001 a_6643_43396# a_n2293_46634# 7e-19
C5002 a_n2661_44458# a_n23_45546# 5.06e-22
C5003 a_n452_44636# a_n755_45592# 0.015469f
C5004 a_18374_44850# a_13259_45724# 0.002311f
C5005 a_18248_44752# a_16375_45002# 1.65e-21
C5006 a_742_44458# a_n357_42282# 0.085409f
C5007 a_11967_42832# a_17715_44484# 0.081495f
C5008 a_743_42282# a_13507_46334# 0.026943f
C5009 a_20749_43396# a_16327_47482# 0.008166f
C5010 a_5111_42852# a_4791_45118# 0.012003f
C5011 a_n3420_38528# a_n2946_38778# 0.236674f
C5012 a_2112_39137# a_1177_38525# 3.38e-19
C5013 a_n3690_38528# a_n4064_38528# 0.085414f
C5014 a_n3565_38502# a_n2302_38778# 0.044367f
C5015 a_n4209_38502# a_n2216_38778# 0.001361f
C5016 a_5275_47026# VDD 0.135766f
C5017 a_4958_30871# C3_N_btm 1.05e-19
C5018 a_n3674_38680# a_n3565_37414# 1.14e-20
C5019 a_765_45546# a_1823_45246# 0.005338f
C5020 a_22365_46825# a_11415_45002# 0.007146f
C5021 a_21350_47026# a_12741_44636# 2.49e-19
C5022 a_5257_43370# a_5066_45546# 0.053231f
C5023 a_n2293_46634# a_n2661_45546# 0.85166f
C5024 a_768_44030# a_1609_45822# 3.5e-21
C5025 a_n2442_46660# a_n2472_45546# 5.69e-20
C5026 a_n2661_46634# a_n2293_45546# 5.66e-20
C5027 a_n2472_46634# a_n2956_38216# 7.81e-20
C5028 a_15009_46634# a_15015_46420# 0.012232f
C5029 a_15368_46634# a_13925_46122# 7.07e-20
C5030 a_n2065_43946# a_n1641_43230# 6.4e-21
C5031 a_n1899_43946# a_n1991_42858# 6.45e-19
C5032 a_n1549_44318# a_n2157_42858# 2.53e-21
C5033 a_5013_44260# a_743_42282# 1.7e-20
C5034 a_14673_44172# a_14543_43071# 2.46e-19
C5035 a_n1331_43914# a_n1853_43023# 6.71e-22
C5036 a_n2267_43396# a_n1352_43396# 0.124988f
C5037 a_n2129_43609# a_n447_43370# 0.119518f
C5038 a_n2956_37592# a_n3565_39590# 0.023811f
C5039 a_17538_32519# VDD 0.352239f
C5040 a_20107_45572# a_20273_45572# 0.667378f
C5041 a_13904_45546# a_9482_43914# 0.002673f
C5042 a_13527_45546# a_13556_45296# 0.006724f
C5043 a_11322_45546# a_1307_43914# 3.56e-20
C5044 a_13249_42308# a_13348_45260# 3.41e-20
C5045 a_11823_42460# a_14537_43396# 0.001649f
C5046 a_9049_44484# a_1423_45028# 0.024539f
C5047 a_2711_45572# a_8560_45348# 0.002436f
C5048 a_8192_45572# a_6171_45002# 0.00429f
C5049 a_n1630_35242# a_n1613_43370# 3.68e-19
C5050 a_6293_42852# a_2324_44458# 0.002463f
C5051 a_8685_43396# a_5937_45572# 7.97e-21
C5052 a_14021_43940# a_20205_31679# 1.01e-20
C5053 a_21115_43940# a_n357_42282# 1.83e-21
C5054 a_14955_43940# a_n443_42852# 5.77e-21
C5055 a_7765_42852# a_3090_45724# 2.34e-20
C5056 a_15743_43084# a_12741_44636# 2.11e-20
C5057 a_8975_43940# CLK 1.38e-19
C5058 a_2981_46116# VDD 0.111597f
C5059 a_2711_45572# a_10227_46804# 0.130695f
C5060 a_10180_45724# a_6151_47436# 9.87e-21
C5061 a_17715_44484# a_13259_45724# 0.391904f
C5062 a_1138_42852# a_n443_42852# 0.14758f
C5063 a_3483_46348# a_3503_45724# 0.009385f
C5064 a_1176_45822# a_1609_45822# 0.010535f
C5065 a_n2267_43396# a_n2293_42282# 6.24e-21
C5066 a_7112_43396# a_7227_42852# 3.34e-19
C5067 a_7287_43370# a_7871_42858# 0.003663f
C5068 a_16243_43396# a_4190_30871# 1.24e-20
C5069 a_17499_43370# a_16823_43084# 0.064861f
C5070 a_3905_42865# a_5932_42308# 0.003844f
C5071 a_3626_43646# a_10341_42308# 0.001954f
C5072 a_2982_43646# a_12089_42308# 1.34e-19
C5073 a_n2661_42282# a_1576_42282# 2.11e-19
C5074 a_3422_30871# a_14113_42308# 5.01e-20
C5075 a_10341_43396# a_20749_43396# 0.003778f
C5076 a_15743_43084# a_15868_43402# 4.12e-21
C5077 a_19339_43156# VDD 0.338297f
C5078 a_3175_45822# a_1414_42308# 7.59e-22
C5079 a_2304_45348# a_n2661_43370# 1.44e-19
C5080 a_8696_44636# a_10617_44484# 0.002097f
C5081 a_n37_45144# a_n2661_44458# 8.09e-19
C5082 a_3232_43370# a_11691_44458# 0.251483f
C5083 a_n913_45002# a_949_44458# 7.6e-21
C5084 a_n1059_45260# a_2779_44458# 8.54e-22
C5085 a_n467_45028# a_n2129_44697# 0.007241f
C5086 a_14097_32519# a_4185_45028# 0.020305f
C5087 a_n901_43156# a_n357_42282# 0.008049f
C5088 a_5649_42852# a_n443_42852# 8.75e-19
C5089 a_14635_42282# a_10903_43370# 1.8e-20
C5090 a_17538_32519# a_22469_39537# 1.77e-20
C5091 a_14797_45144# a_11453_44696# 0.002114f
C5092 a_1307_43914# a_12465_44636# 0.022149f
C5093 a_5205_44484# a_n1613_43370# 0.551795f
C5094 a_6431_45366# a_n881_46662# 0.177591f
C5095 a_3065_45002# a_768_44030# 0.288972f
C5096 a_3357_43084# a_n743_46660# 0.034228f
C5097 a_1609_45572# a_765_45546# 1.84e-19
C5098 a_2711_45572# a_17339_46660# 0.02331f
C5099 a_11823_42460# a_3090_45724# 0.089008f
C5100 a_13527_45546# a_13607_46688# 8.43e-20
C5101 a_22165_42308# a_22959_42860# 6.47e-20
C5102 a_743_42282# a_196_42282# 7.61e-19
C5103 a_10695_43548# a_10533_42308# 9.55e-22
C5104 a_3626_43646# a_18057_42282# 0.01061f
C5105 a_2982_43646# a_18907_42674# 8.43e-20
C5106 a_13467_32519# COMP_P 5.83e-19
C5107 a_3080_42308# a_13258_32519# 7.3e-19
C5108 a_10518_42984# a_10793_43218# 0.007416f
C5109 a_8945_43396# a_5934_30871# 1.73e-20
C5110 a_2324_44458# RST_Z 1.22e-21
C5111 a_22465_38105# VDD 1.3089f
C5112 a_n1741_47186# a_8128_46384# 0.004988f
C5113 a_n971_45724# a_n1613_43370# 0.6298f
C5114 a_11599_46634# a_15507_47210# 0.267808f
C5115 a_6151_47436# a_13507_46334# 7.34e-21
C5116 a_14955_47212# a_15811_47375# 1.55e-19
C5117 a_2063_45854# a_2747_46873# 0.023413f
C5118 a_13717_47436# a_16023_47582# 1.27e-19
C5119 a_9313_45822# a_10227_46804# 1.42e-19
C5120 a_12861_44030# a_16327_47482# 0.120085f
C5121 a_n1151_42308# a_n2312_39304# 2.72e-19
C5122 a_17719_45144# a_11967_42832# 2.77e-21
C5123 a_18587_45118# a_18588_44850# 3.44e-19
C5124 a_11827_44484# a_17517_44484# 0.05115f
C5125 a_n2129_44697# a_n2661_43922# 0.00767f
C5126 a_n2267_44484# a_n2661_42834# 0.002133f
C5127 a_949_44458# a_556_44484# 0.001921f
C5128 a_5883_43914# a_5891_43370# 0.216958f
C5129 a_n2433_44484# a_n2293_43922# 0.010009f
C5130 a_16922_45042# a_20362_44736# 0.00806f
C5131 a_1423_45028# a_3905_42865# 9.59e-20
C5132 a_1307_43914# a_7281_43914# 0.004629f
C5133 a_8103_44636# a_8333_44734# 0.004937f
C5134 a_18374_44850# a_18989_43940# 3.56e-21
C5135 a_3232_43370# a_8333_44056# 2.98e-19
C5136 a_n913_45002# a_11341_43940# 0.001663f
C5137 a_7229_43940# a_n2661_42282# 2.13e-19
C5138 a_n2017_45002# a_15493_43940# 9.45e-20
C5139 a_n2946_39072# a_n2956_38680# 0.004064f
C5140 a_n4064_39072# a_n2956_39304# 0.054199f
C5141 a_10533_42308# a_n357_42282# 7.55e-20
C5142 a_7963_42308# a_n443_42852# 4.91e-20
C5143 a_5534_30871# a_n923_35174# 0.007036f
C5144 a_11963_45334# a_11415_45002# 0.031636f
C5145 a_2382_45260# a_1823_45246# 0.801932f
C5146 a_1667_45002# a_167_45260# 0.05322f
C5147 a_413_45260# a_2698_46116# 9.42e-21
C5148 a_n2661_42834# a_5807_45002# 5.92e-21
C5149 a_5205_44484# a_n2293_46098# 0.001237f
C5150 a_14495_45572# a_13259_45724# 0.020864f
C5151 a_3638_45822# a_n755_45592# 9.05e-19
C5152 a_9159_45572# a_10586_45546# 1.71e-19
C5153 a_3357_43084# a_11189_46129# 3.29e-22
C5154 a_2437_43646# a_10903_43370# 5.87e-20
C5155 a_1241_44260# a_584_46384# 1.06e-19
C5156 a_1755_42282# a_2713_42308# 9.85e-19
C5157 a_1606_42308# a_2903_42308# 0.001317f
C5158 a_5342_30871# a_n3420_39072# 0.062032f
C5159 a_5807_45002# a_8145_46902# 0.003883f
C5160 a_n743_46660# a_3877_44458# 0.034265f
C5161 a_n2661_46634# a_5732_46660# 0.010632f
C5162 a_n1925_46634# a_4651_46660# 0.046762f
C5163 a_2107_46812# a_3524_46660# 0.004383f
C5164 a_948_46660# a_2864_46660# 3.21e-21
C5165 a_12549_44172# a_6755_46942# 0.553062f
C5166 a_479_46660# a_n2661_46098# 3.93e-19
C5167 a_11453_44696# a_14976_45028# 0.014048f
C5168 a_3080_42308# a_3754_38802# 4.08e-21
C5169 a_13507_46334# a_19466_46812# 0.03247f
C5170 a_4883_46098# a_15227_44166# 0.176028f
C5171 a_21177_47436# a_19692_46634# 0.001012f
C5172 a_14955_47212# a_13059_46348# 1.12e-19
C5173 a_10227_46804# a_12513_46660# 0.004052f
C5174 a_15811_47375# a_14543_46987# 2.63e-20
C5175 a_11599_46634# a_15227_46910# 0.006776f
C5176 a_11031_47542# a_765_45546# 0.003176f
C5177 a_12861_44030# a_16434_46987# 0.001423f
C5178 a_n971_45724# a_n2293_46098# 0.110318f
C5179 a_n815_47178# a_n1853_46287# 4.63e-19
C5180 a_n2109_47186# a_n1076_46494# 1.12e-20
C5181 a_n1917_44484# a_n1917_43396# 9.63e-19
C5182 a_n2267_44484# a_n1352_43396# 6.41e-21
C5183 a_n1899_43946# a_n1331_43914# 0.171939f
C5184 a_n2065_43946# a_n809_44244# 0.043475f
C5185 a_n1761_44111# a_n1549_44318# 0.033724f
C5186 a_11541_44484# a_11750_44172# 2.79e-19
C5187 a_n1352_44484# a_n2267_43396# 2.85e-20
C5188 a_n2661_44458# a_104_43370# 8.68e-21
C5189 a_18494_42460# a_3626_43646# 0.066461f
C5190 a_11823_42460# a_12991_43230# 0.001129f
C5191 en_comp a_n1991_42858# 2.41e-19
C5192 a_n1059_45260# a_n13_43084# 0.027848f
C5193 a_n913_45002# a_n1076_43230# 0.05439f
C5194 a_3537_45260# a_4361_42308# 0.017454f
C5195 a_n967_45348# a_n1853_43023# 0.021497f
C5196 a_3357_43084# a_1847_42826# 0.010588f
C5197 a_n2017_45002# a_n3674_39304# 6.29e-20
C5198 a_413_45260# a_22959_43396# 2.15e-19
C5199 a_n3565_37414# VDD 0.783539f
C5200 a_19721_31679# VDD 0.521328f
C5201 a_22465_38105# a_22469_39537# 0.576946f
C5202 a_4958_30871# C7_P_btm 1.47e-19
C5203 a_10341_43396# a_12861_44030# 0.018259f
C5204 a_5608_44484# a_5164_46348# 4.14e-20
C5205 a_18989_43940# a_17715_44484# 1.14e-20
C5206 a_12883_44458# a_10809_44734# 2.59e-19
C5207 a_9313_44734# a_8016_46348# 0.020204f
C5208 a_8855_44734# a_8199_44636# 0.002934f
C5209 a_18287_44626# a_18819_46122# 3.39e-21
C5210 a_18248_44752# a_18985_46122# 4.72e-21
C5211 a_17719_45144# a_13259_45724# 0.039832f
C5212 a_16922_45042# a_16375_45002# 0.170835f
C5213 a_2809_45028# a_2957_45546# 6.81e-20
C5214 a_4223_44672# a_526_44458# 1.22e-19
C5215 a_9420_43940# a_2107_46812# 1.23e-19
C5216 a_17538_32519# a_22612_30879# 0.060018f
C5217 a_458_43396# a_768_44030# 0.001002f
C5218 a_16789_44484# a_12741_44636# 0.009606f
C5219 a_n2661_43922# a_3483_46348# 0.038814f
C5220 a_10193_42453# CLK 0.023289f
C5221 a_n4315_30879# a_n4064_39616# 0.034877f
C5222 a_n4064_40160# a_n3420_39616# 0.05705f
C5223 a_7174_31319# a_n3565_39304# 4.27e-21
C5224 a_13675_47204# VDD 0.004094f
C5225 a_1606_42308# C9_N_btm 9.33e-20
C5226 a_5807_45002# a_5066_45546# 0.027744f
C5227 a_n2438_43548# a_n2956_38680# 0.00293f
C5228 a_12549_44172# a_8049_45260# 0.031115f
C5229 a_n2293_46634# a_n1533_46116# 9.21e-21
C5230 a_n1925_46634# a_n1379_46482# 3.89e-19
C5231 a_5907_46634# a_5937_45572# 1.19e-19
C5232 a_11453_44696# a_18051_46116# 0.00399f
C5233 a_13507_46334# a_20205_31679# 0.023531f
C5234 a_4883_46098# a_21071_46482# 1.62e-19
C5235 a_11901_46660# a_11415_45002# 1.07e-20
C5236 a_15227_44166# a_21188_46660# 3.62e-19
C5237 a_19692_46634# a_20841_46902# 0.025536f
C5238 a_3090_45724# a_18280_46660# 4.52e-21
C5239 a_6453_43914# a_6452_43396# 8.84e-19
C5240 a_19328_44172# a_n97_42460# 9.4e-21
C5241 a_22959_43948# a_17538_32519# 0.168682f
C5242 a_19615_44636# a_19700_43370# 1.17e-20
C5243 a_n2661_42834# a_n2472_42826# 0.03087f
C5244 a_n356_44636# a_7765_42852# 1.83e-20
C5245 a_3499_42826# a_3626_43646# 0.001049f
C5246 a_375_42282# a_n327_42558# 7.38e-21
C5247 a_15493_43940# a_21845_43940# 5.9e-19
C5248 a_11967_42832# a_16664_43396# 1.34e-19
C5249 a_5111_44636# a_6171_42473# 2.14e-20
C5250 a_2382_45260# a_5934_30871# 1.02e-20
C5251 a_3065_45002# a_6123_31319# 9.58e-21
C5252 a_3537_45260# a_6761_42308# 0.057884f
C5253 a_n913_45002# a_10723_42308# 0.006785f
C5254 a_n1059_45260# a_11323_42473# 6.13e-20
C5255 a_n2017_45002# a_5742_30871# 0.007608f
C5256 a_17973_43940# VDD 0.265874f
C5257 a_15765_45572# a_16020_45572# 0.056391f
C5258 a_16855_45546# a_8696_44636# 0.112262f
C5259 a_8530_39574# CAL_P 0.037066f
C5260 a_16243_43396# a_15227_44166# 0.002283f
C5261 a_14579_43548# a_13059_46348# 0.171744f
C5262 a_n809_44244# a_n755_45592# 0.404418f
C5263 a_1414_42308# a_n863_45724# 0.711805f
C5264 a_2675_43914# a_n2661_45546# 1.1e-21
C5265 a_n984_44318# a_n357_42282# 1.05e-19
C5266 a_175_44278# a_310_45028# 1.47e-19
C5267 a_19518_43218# a_16327_47482# 0.002315f
C5268 a_6123_31319# w_1575_34946# 0.002297f
C5269 a_19721_31679# a_22469_39537# 3.67e-20
C5270 a_167_45260# VDD 1.41955f
C5271 C3_N_btm C7_N_btm 0.134911f
C5272 C4_N_btm C6_N_btm 0.143514f
C5273 C0_N_btm C10_N_btm 0.365593f
C5274 C1_N_btm C9_N_btm 0.132506f
C5275 C2_N_btm C8_N_btm 0.138777f
C5276 a_22775_42308# a_22469_40625# 2.08e-20
C5277 a_1823_45246# a_6347_46155# 7.53e-22
C5278 a_3699_46348# a_5066_45546# 1.54e-20
C5279 a_765_45546# a_n2293_45546# 7.13e-22
C5280 a_13351_46090# a_6945_45028# 8.55e-21
C5281 a_12005_46116# a_10809_44734# 0.029593f
C5282 a_17583_46090# a_17957_46116# 0.092344f
C5283 a_17715_44484# a_18189_46348# 0.014348f
C5284 a_n4209_38216# a_n3420_37984# 0.067687f
C5285 a_1343_38525# a_3754_38470# 4.25e-20
C5286 a_n4064_39616# a_n3420_37440# 0.056826f
C5287 a_n3420_39616# a_n4064_37440# 0.047863f
C5288 a_n4334_38304# a_n3690_38304# 8.67e-19
C5289 a_n1699_43638# a_n1991_42858# 4.92e-20
C5290 a_n1917_43396# a_n1853_43023# 0.001737f
C5291 a_n2267_43396# a_n1423_42826# 0.001766f
C5292 a_n1177_43370# a_n2157_42858# 6.59e-19
C5293 a_4699_43561# a_743_42282# 1.35e-20
C5294 a_14358_43442# a_14205_43396# 0.163543f
C5295 a_9803_43646# a_10341_43396# 0.11445f
C5296 a_14579_43548# a_15095_43370# 0.109081f
C5297 a_n2129_43609# a_n1641_43230# 1.1e-19
C5298 a_14021_43940# a_15279_43071# 5.5e-21
C5299 a_15493_43940# a_19164_43230# 3.58e-20
C5300 a_11341_43940# a_20922_43172# 7.6e-21
C5301 a_n2661_42834# a_9223_42460# 8.65e-22
C5302 a_n2293_43922# a_8685_42308# 3.58e-20
C5303 a_9145_43396# a_10765_43646# 0.00303f
C5304 a_n4318_40392# a_n4064_39616# 6.39e-21
C5305 a_8685_43396# a_9885_43396# 4.64e-19
C5306 a_4883_46098# EN_OFFSET_CAL 8.93e-21
C5307 a_22591_43396# VDD 0.280354f
C5308 a_8162_45546# a_5891_43370# 4.81e-19
C5309 a_6511_45714# a_n2661_42834# 6.91e-21
C5310 a_18341_45572# a_11691_44458# 4.3e-20
C5311 a_10951_45334# a_9482_43914# 5.58e-21
C5312 a_7499_43078# a_7640_43914# 0.021219f
C5313 a_2711_45572# a_14815_43914# 9.7e-21
C5314 a_11823_42460# a_n356_44636# 5.09e-19
C5315 a_18479_45785# a_20193_45348# 1.42e-21
C5316 a_6171_45002# a_16751_45260# 0.104212f
C5317 a_5147_45002# a_1423_45028# 0.017515f
C5318 a_n2017_45002# a_n2293_42834# 0.28698f
C5319 a_3065_45002# a_3495_45348# 0.001093f
C5320 a_15743_43084# a_16375_45002# 1.19e-20
C5321 a_n13_43084# a_n1925_42282# 5.01e-21
C5322 a_8685_43396# a_n443_42852# 0.281116f
C5323 a_22465_38105# a_22612_30879# 9.58e-19
C5324 a_22959_42860# a_4185_45028# 0.013205f
C5325 a_15861_45028# a_5807_45002# 3.23e-19
C5326 a_2711_45572# a_10467_46802# 2.47e-20
C5327 a_16680_45572# a_13747_46662# 0.047612f
C5328 a_8696_44636# a_13661_43548# 0.049791f
C5329 a_9241_45822# a_2107_46812# 5.82e-21
C5330 a_12016_45572# a_n2661_46634# 3.65e-19
C5331 a_14033_45572# a_768_44030# 7.13e-19
C5332 a_14127_45572# a_12549_44172# 2.41e-19
C5333 a_18691_45572# a_n881_46662# 3.57e-20
C5334 a_2437_43646# a_4883_46098# 0.458866f
C5335 a_19479_31679# a_13507_46334# 0.061466f
C5336 a_3357_43084# a_21177_47436# 5.54e-20
C5337 a_n913_45002# a_16327_47482# 0.137194f
C5338 a_21297_45572# a_18597_46090# 4.45e-19
C5339 a_413_45260# a_n1435_47204# 0.025027f
C5340 a_6171_45002# a_4915_47217# 0.022258f
C5341 a_5205_44484# a_4791_45118# 0.053467f
C5342 a_8953_45002# a_n1151_42308# 1.04e-19
C5343 a_n755_45592# a_3316_45546# 0.045656f
C5344 a_n2661_45546# a_2277_45546# 0.00928f
C5345 a_n1099_45572# a_n23_45546# 0.042611f
C5346 a_310_45028# a_n356_45724# 0.12349f
C5347 a_n1079_45724# a_n906_45572# 0.007688f
C5348 a_n452_45724# a_7_45899# 6.64e-19
C5349 a_n863_45724# a_n1013_45572# 0.001771f
C5350 a_6031_43396# a_1755_42282# 3.75e-21
C5351 a_10083_42826# a_10518_42984# 0.234322f
C5352 a_n2472_42826# a_n2293_42282# 3.06e-19
C5353 a_2982_43646# a_5267_42460# 1.03e-19
C5354 a_n97_42460# a_8685_42308# 2.19e-19
C5355 a_4905_42826# a_5337_42558# 0.005481f
C5356 a_9127_43156# a_10796_42968# 1.62e-19
C5357 a_3539_42460# a_2903_42308# 6.02e-19
C5358 a_21076_30879# a_21589_35634# 5.95e-20
C5359 a_8530_39574# CAL_N 0.644218f
C5360 a_n1741_47186# a_6151_47436# 0.071065f
C5361 a_n971_45724# a_4791_45118# 0.025426f
C5362 a_1209_47178# a_n1151_42308# 0.024897f
C5363 a_584_46384# a_2553_47502# 0.100103f
C5364 a_n237_47217# a_4007_47204# 2.65e-20
C5365 a_2124_47436# a_2952_47436# 5.21e-19
C5366 a_1307_43914# a_16241_44734# 0.010259f
C5367 a_18587_45118# a_18443_44721# 7.68e-20
C5368 a_18911_45144# a_18287_44626# 3.74e-19
C5369 a_n2267_44484# a_n1352_44484# 0.118759f
C5370 a_n2129_44697# a_n452_44636# 0.079904f
C5371 a_n2661_43370# a_8375_44464# 9.68e-20
C5372 a_n2661_44458# a_949_44458# 0.041721f
C5373 a_11691_44458# a_8975_43940# 0.048259f
C5374 a_11827_44484# a_13720_44458# 0.00996f
C5375 a_14537_43396# a_15367_44484# 0.001966f
C5376 a_413_45260# a_22959_44484# 0.202222f
C5377 a_n967_45348# a_n1899_43946# 0.025102f
C5378 a_n745_45366# a_n984_44318# 1.8e-20
C5379 a_n2661_45010# a_2127_44172# 0.096614f
C5380 a_n1059_45260# a_644_44056# 6.29e-19
C5381 a_n2017_45002# a_1115_44172# 3.58e-21
C5382 a_3357_43084# a_5244_44056# 1.59e-20
C5383 a_n2293_45010# a_1414_42308# 3e-19
C5384 a_n2104_42282# a_n2956_38216# 2.12e-20
C5385 a_5742_30871# a_526_44458# 2.52e-20
C5386 a_n4318_37592# a_n2810_45572# 0.023163f
C5387 a_20256_42852# a_n357_42282# 9.51e-19
C5388 a_3175_45822# VDD 0.193907f
C5389 a_4190_30871# a_n923_35174# 0.025255f
C5390 a_17364_32525# a_22521_39511# 9.72e-21
C5391 a_15743_43084# RST_Z 2.97e-19
C5392 a_14673_44172# a_4915_47217# 0.020025f
C5393 a_n2293_43922# a_12861_44030# 0.008309f
C5394 a_11682_45822# a_12594_46348# 4.71e-19
C5395 a_10490_45724# a_10809_44734# 0.030973f
C5396 a_413_45260# a_13885_46660# 1.99e-20
C5397 a_3357_43084# a_20841_46902# 0.001309f
C5398 a_2437_43646# a_21188_46660# 1.87e-22
C5399 a_3260_45572# a_526_44458# 2.83e-20
C5400 a_6511_45714# a_5066_45546# 2.64e-19
C5401 a_2711_45572# a_8034_45724# 0.035334f
C5402 a_19721_31679# a_22612_30879# 0.068873f
C5403 a_5093_45028# a_5257_43370# 3.11e-21
C5404 a_6298_44484# a_768_44030# 0.015186f
C5405 a_16237_45028# a_n743_46660# 0.038671f
C5406 a_18953_45572# a_11415_45002# 4.28e-19
C5407 a_20107_45572# a_20202_43084# 0.002433f
C5408 a_15567_42826# a_15051_42282# 0.001656f
C5409 a_16414_43172# a_14113_42308# 0.004427f
C5410 a_5193_42852# a_5379_42460# 3.15e-19
C5411 a_5342_30871# a_15486_42560# 0.006845f
C5412 a_12089_42308# a_11897_42308# 1.97e-19
C5413 a_4190_30871# a_n4064_39072# 1.46e-20
C5414 a_8128_46384# a_n743_46660# 0.006641f
C5415 a_n881_46662# a_33_46660# 0.002482f
C5416 a_n1613_43370# a_601_46902# 0.178721f
C5417 a_6575_47204# a_6755_46942# 1.56e-19
C5418 a_n1435_47204# a_9863_46634# 2.27e-20
C5419 a_9313_45822# a_10467_46802# 0.009777f
C5420 a_6151_47436# a_7832_46660# 0.016469f
C5421 a_12891_46348# a_n2293_46634# 5.27e-20
C5422 a_5807_45002# a_19321_45002# 0.376188f
C5423 a_10334_44484# a_10405_44172# 0.002711f
C5424 a_n2661_43922# a_n2472_43914# 0.068474f
C5425 a_n2293_43922# a_n2840_43914# 0.001304f
C5426 a_n2661_42834# a_n2065_43946# 0.035267f
C5427 a_8975_43940# a_8333_44056# 7.34e-19
C5428 a_1307_43914# a_n1557_42282# 6.39e-20
C5429 a_11823_42460# a_12379_42858# 0.033971f
C5430 a_10193_42453# a_5534_30871# 0.136243f
C5431 a_18588_44850# a_11967_42832# 8.49e-19
C5432 a_20193_45348# a_14021_43940# 0.118757f
C5433 a_1423_45028# a_4093_43548# 1.31e-20
C5434 a_n2661_44458# a_11341_43940# 0.001405f
C5435 a_n913_45002# a_10341_43396# 0.032712f
C5436 a_3537_45260# a_7274_43762# 4.26e-19
C5437 a_1606_42308# RST_Z 1.44945f
C5438 a_2779_44458# a_2698_46116# 2.15e-19
C5439 a_17970_44736# a_12741_44636# 9.86e-19
C5440 a_18443_44721# a_11415_45002# 7.02e-22
C5441 a_n699_43396# a_167_45260# 6.1e-22
C5442 a_5343_44458# a_1823_45246# 2.1e-19
C5443 a_19478_44306# a_19321_45002# 6.34e-21
C5444 a_20365_43914# a_13661_43548# 0.020045f
C5445 a_3905_42865# a_4646_46812# 1.17e-19
C5446 a_10555_44260# a_768_44030# 0.00973f
C5447 a_15367_44484# a_3090_45724# 5.11e-19
C5448 a_n2293_42834# a_526_44458# 1.7774f
C5449 a_413_45260# a_380_45546# 0.001298f
C5450 a_n37_45144# a_n1099_45572# 1.51e-19
C5451 a_3429_45260# a_n2661_45546# 5.93e-20
C5452 a_1667_45002# a_n863_45724# 0.20954f
C5453 a_2382_45260# a_n2293_45546# 0.078874f
C5454 a_n143_45144# a_310_45028# 1.85e-20
C5455 a_16922_45042# a_18985_46122# 4.99e-21
C5456 a_n2661_44458# a_5497_46414# 6.51e-22
C5457 a_17719_45144# a_18189_46348# 0.002906f
C5458 a_11691_44458# a_11387_46155# 1.27e-22
C5459 a_n97_42460# a_12861_44030# 5.48e-20
C5460 a_648_43396# a_584_46384# 0.050476f
C5461 a_8791_43396# a_n971_45724# 8.26e-19
C5462 a_n1557_42282# a_n443_46116# 0.006023f
C5463 a_17124_42282# a_4958_30871# 0.20224f
C5464 a_14113_42308# a_7174_31319# 4.19e-20
C5465 a_16522_42674# a_17303_42282# 2.42e-20
C5466 a_5934_30871# a_1239_39587# 1.67e-19
C5467 a_5932_42308# a_n3565_39304# 3.95e-21
C5468 a_11459_47204# VDD 0.34771f
C5469 a_5649_42852# CAL_N 0.005399f
C5470 a_13678_32519# a_22521_40599# 2.48e-21
C5471 a_n2661_46634# a_1138_42852# 4.66e-20
C5472 a_n1925_46634# a_n1076_46494# 0.003622f
C5473 a_n1021_46688# a_n901_46420# 0.001157f
C5474 a_n2438_43548# a_n1423_46090# 9.01e-21
C5475 a_11901_46660# a_12251_46660# 0.219633f
C5476 a_11735_46660# a_12816_46660# 0.102325f
C5477 a_5732_46660# a_765_45546# 0.003297f
C5478 a_11813_46116# a_12991_46634# 1.29e-20
C5479 a_6755_46942# a_10861_46660# 2.63e-19
C5480 a_768_44030# a_5937_45572# 0.05116f
C5481 a_n881_46662# a_12005_46116# 1.14e-20
C5482 a_14209_32519# VDAC_N 2.4e-19
C5483 a_4883_46098# a_22959_46124# 1.36e-19
C5484 a_22223_47212# a_6945_45028# 4.85e-19
C5485 a_11453_44696# a_19900_46494# 3.8e-20
C5486 a_12465_44636# a_22223_46124# 7.35e-21
C5487 a_6575_47204# a_8049_45260# 0.002085f
C5488 a_6151_47436# a_10586_45546# 1.83e-20
C5489 a_21811_47423# a_10809_44734# 0.005196f
C5490 a_n1899_43946# a_n1917_43396# 4.39e-19
C5491 a_n809_44244# a_n2129_43609# 3.98e-20
C5492 a_n2065_43946# a_n1352_43396# 0.009873f
C5493 a_18079_43940# a_15493_43940# 0.040279f
C5494 a_18451_43940# a_11341_43940# 0.004129f
C5495 a_19862_44208# a_20365_43914# 0.075162f
C5496 a_n1331_43914# a_n1699_43638# 1.55e-19
C5497 a_n1549_44318# a_n2267_43396# 9.07e-20
C5498 a_n1761_44111# a_n1177_43370# 1.22e-19
C5499 a_n2661_43922# a_10695_43548# 1.39e-20
C5500 a_n1917_44484# a_n1853_43023# 1.77e-20
C5501 a_9313_44734# a_12281_43396# 0.027032f
C5502 a_10193_42453# a_19647_42308# 0.004706f
C5503 a_7499_43078# a_7174_31319# 9.76e-21
C5504 a_11750_44172# a_11816_44260# 0.006978f
C5505 a_10949_43914# a_12603_44260# 0.001915f
C5506 a_14539_43914# a_16855_43396# 9.74e-19
C5507 en_comp a_22400_42852# 0.730145f
C5508 a_22591_44484# VDD 0.223346f
C5509 a_11322_45546# a_11682_45822# 0.034435f
C5510 a_14495_45572# a_15143_45578# 8.73e-19
C5511 a_11652_45724# a_10907_45822# 1.68e-19
C5512 a_2711_45572# a_13297_45572# 8.55e-20
C5513 C7_N_btm C7_P_btm 0.028901f
C5514 C6_N_btm C6_P_btm 0.019861f
C5515 C5_N_btm C5_P_btm 0.03705f
C5516 C4_N_btm C4_P_btm 0.02642f
C5517 C3_N_btm C3_P_btm 2.90911f
C5518 C2_N_btm C2_P_btm 0.026726f
C5519 a_20922_43172# a_16327_47482# 0.001914f
C5520 a_13635_43156# a_12465_44636# 3.45e-20
C5521 a_10405_44172# a_9290_44172# 0.001407f
C5522 a_n2661_43922# a_n357_42282# 0.088336f
C5523 a_1115_44172# a_526_44458# 0.009996f
C5524 a_n2661_42834# a_n755_45592# 0.059506f
C5525 a_3363_44484# a_3503_45724# 8.59e-21
C5526 a_2982_43646# a_3090_45724# 1.98e-20
C5527 a_4361_42308# a_n2293_46634# 5.54e-21
C5528 a_14209_32519# a_21588_30879# 0.056208f
C5529 a_11415_45002# a_17583_46090# 2.43e-20
C5530 a_12741_44636# a_14840_46494# 9.71e-23
C5531 a_3483_46348# a_5164_46348# 0.025074f
C5532 a_22000_46634# a_10809_44734# 0.012475f
C5533 a_20731_47026# a_6945_45028# 0.001536f
C5534 a_4699_43561# a_2813_43396# 1.26e-20
C5535 a_2982_43646# a_6547_43396# 4.43e-21
C5536 a_3626_43646# a_6197_43396# 3.15e-20
C5537 a_n2661_42282# a_5755_42852# 0.006322f
C5538 a_n356_44636# a_961_42354# 0.005209f
C5539 a_n97_42460# a_9803_43646# 1.56e-20
C5540 a_5343_44458# a_5934_30871# 7.67e-19
C5541 a_14021_43940# a_20301_43646# 0.024612f
C5542 a_4093_43548# a_4181_43396# 2.48e-19
C5543 a_16922_45042# a_17303_42282# 1.31e-20
C5544 a_15493_43940# a_14209_32519# 3.85e-21
C5545 a_11341_43940# a_17364_32525# 0.005541f
C5546 a_n971_45724# DATA[3] 0.09508f
C5547 a_n23_47502# DATA[0] 0.022435f
C5548 a_n237_47217# DATA[1] 0.139838f
C5549 a_10193_42453# a_11691_44458# 0.046462f
C5550 a_4099_45572# a_4223_44672# 3.68e-19
C5551 a_2711_45572# a_4743_44484# 4.71e-21
C5552 a_3357_43084# a_5111_44636# 0.318002f
C5553 a_n745_45366# a_n467_45028# 0.110406f
C5554 en_comp a_n967_45348# 0.001993f
C5555 a_2437_43646# a_3232_43370# 2.01e-19
C5556 a_18817_42826# a_17339_46660# 3.49e-19
C5557 a_5934_30871# a_n2956_39768# 6.35e-21
C5558 a_n1352_43396# a_n755_45592# 3.17e-19
C5559 a_n447_43370# a_n357_42282# 0.00435f
C5560 a_5649_42852# a_8199_44636# 9.98e-20
C5561 a_13258_32519# a_13507_46334# 0.049541f
C5562 a_19237_31679# a_22521_39511# 1.89e-20
C5563 a_n863_45724# VDD 1.89058f
C5564 a_16680_45572# a_11599_46634# 0.002914f
C5565 a_15903_45785# a_16327_47482# 0.005367f
C5566 a_16020_45572# a_12861_44030# 9.09e-21
C5567 a_5066_45546# a_n755_45592# 4.16e-20
C5568 a_13483_43940# a_13575_42558# 1.75e-21
C5569 a_n2157_42858# a_n1991_42858# 0.905962f
C5570 a_10341_43396# a_20922_43172# 8.95e-20
C5571 a_743_42282# a_1847_42826# 0.004285f
C5572 a_n97_42460# a_19518_43218# 3.81e-19
C5573 a_17665_42852# VDD 0.006567f
C5574 a_14537_43396# a_14539_43914# 0.135541f
C5575 a_17719_45144# a_18315_45260# 0.017382f
C5576 a_16922_45042# a_19778_44110# 0.026041f
C5577 a_1423_45028# a_10157_44484# 5.42e-19
C5578 a_7499_43078# a_10729_43914# 0.23002f
C5579 a_1307_43914# a_12883_44458# 2.26e-21
C5580 a_n745_45366# a_n2661_43922# 2.34e-20
C5581 a_3537_45260# a_5891_43370# 0.359819f
C5582 a_n913_45002# a_n2293_43922# 0.019153f
C5583 a_5147_45002# a_6109_44484# 7.39e-19
C5584 a_873_42968# a_n863_45724# 0.002982f
C5585 a_n2293_42282# a_n755_45592# 0.208531f
C5586 a_13249_42308# a_11415_45002# 0.071546f
C5587 a_3775_45552# a_3699_46348# 1.45e-19
C5588 a_4880_45572# a_1823_45246# 0.002594f
C5589 a_18341_45572# a_15227_44166# 0.017357f
C5590 a_18175_45572# a_19466_46812# 7.28e-19
C5591 a_18909_45814# a_18834_46812# 9e-22
C5592 a_16115_45572# a_13059_46348# 1.11e-20
C5593 a_2809_45348# a_n2293_46634# 0.001204f
C5594 a_3537_45260# a_4817_46660# 4.15e-22
C5595 a_5147_45002# a_4646_46812# 0.010619f
C5596 a_5111_44636# a_3877_44458# 3.05e-20
C5597 a_3357_43084# a_6086_46660# 3.67e-19
C5598 a_6194_45824# a_5204_45822# 4.22e-20
C5599 a_2711_45572# a_8016_46348# 0.028247f
C5600 a_20193_45348# a_13507_46334# 0.253904f
C5601 a_7_44811# a_n746_45260# 0.001383f
C5602 a_4361_42308# a_13249_42558# 7.13e-20
C5603 a_18525_43370# a_18057_42282# 6.86e-21
C5604 a_22165_42308# a_22400_42852# 0.005425f
C5605 a_743_42282# a_15486_42560# 0.010882f
C5606 a_5649_42852# a_13070_42354# 6.66e-20
C5607 a_4190_30871# a_15803_42450# 1.32e-19
C5608 a_15743_43084# a_17303_42282# 1.95e-20
C5609 a_14209_32519# a_5742_30871# 0.005505f
C5610 a_19987_42826# a_20753_42852# 0.07365f
C5611 a_21671_42860# a_14097_32519# 8.99e-20
C5612 a_5534_30871# a_n784_42308# 9.92256f
C5613 a_17730_32519# VDAC_N 0.008268f
C5614 a_11599_46634# a_13747_46662# 0.25325f
C5615 a_15811_47375# a_5807_45002# 0.004711f
C5616 a_16023_47582# a_16285_47570# 0.001705f
C5617 a_15673_47210# a_16131_47204# 0.034619f
C5618 a_10227_46804# a_16119_47582# 0.004305f
C5619 a_16327_47482# a_16697_47582# 2.95e-19
C5620 a_6151_47436# a_n743_46660# 0.03019f
C5621 a_6491_46660# a_n1925_46634# 0.003135f
C5622 a_n1151_42308# a_288_46660# 8.13e-19
C5623 a_3785_47178# a_2107_46812# 2.1e-20
C5624 a_2124_47436# a_n2661_46098# 1.36e-19
C5625 a_n443_46116# a_33_46660# 1.22e-19
C5626 a_584_46384# a_1799_45572# 0.179456f
C5627 a_n2109_47186# a_4646_46812# 0.021783f
C5628 a_n1917_44484# a_n1899_43946# 0.012479f
C5629 a_n2267_44484# a_n1549_44318# 5.88e-19
C5630 a_n1352_44484# a_n2065_43946# 0.00236f
C5631 a_n1177_44458# a_n1761_44111# 4.25e-20
C5632 a_18443_44721# a_11967_42832# 0.035979f
C5633 a_18287_44626# a_19615_44636# 9.28e-19
C5634 a_n2129_44697# a_n809_44244# 3.14e-20
C5635 a_n2661_44458# a_175_44278# 5.37e-21
C5636 a_n2661_43370# a_10949_43914# 2.82e-20
C5637 a_8696_44636# a_14579_43548# 5.14e-23
C5638 a_10193_42453# a_4190_30871# 0.305842f
C5639 a_3363_44484# a_n2661_43922# 0.005466f
C5640 a_n2017_45002# a_n2012_43396# 0.009581f
C5641 a_3357_43084# a_4235_43370# 0.00216f
C5642 a_n913_45002# a_n97_42460# 0.109647f
C5643 a_n1059_45260# a_104_43370# 1.35e-20
C5644 a_n2293_45010# a_n1190_43762# 4.42e-20
C5645 a_n967_45348# a_n1699_43638# 0.001377f
C5646 a_n2293_45010# VDD 1.885f
C5647 a_18451_43940# a_16327_47482# 0.001635f
C5648 a_15682_43940# a_10227_46804# 0.003864f
C5649 a_21115_43940# a_12861_44030# 0.035299f
C5650 a_6171_45002# a_10809_44734# 0.244599f
C5651 a_5205_44484# a_6945_45028# 0.058545f
C5652 a_7281_43914# a_n1613_43370# 0.030229f
C5653 a_9482_43914# a_2324_44458# 0.009807f
C5654 a_14797_45144# a_13925_46122# 1.91e-20
C5655 a_13556_45296# a_14840_46494# 2.96e-19
C5656 a_6453_43914# a_n881_46662# 2.61e-19
C5657 a_21297_45572# a_8049_45260# 2.09e-19
C5658 a_413_45260# a_526_44458# 0.103799f
C5659 a_17668_45572# a_16375_45002# 2.56e-19
C5660 a_17730_32519# a_21588_30879# 0.05582f
C5661 a_14539_43914# a_3090_45724# 0.040638f
C5662 a_2479_44172# a_768_44030# 0.056833f
C5663 a_5009_45028# a_4185_45028# 0.002751f
C5664 a_5837_45028# a_3483_46348# 0.00532f
C5665 a_17613_45144# a_11415_45002# 0.004987f
C5666 a_n2661_43370# a_376_46348# 1.86e-21
C5667 a_8685_42308# a_10533_42308# 4.55e-21
C5668 a_n1386_35608# VIN_P 0.367112f
C5669 C8_P_btm C2_P_btm 0.138777f
C5670 C7_P_btm C3_P_btm 0.134911f
C5671 C6_P_btm C4_P_btm 0.143514f
C5672 a_22959_47212# a_21076_30879# 0.002641f
C5673 a_6575_47204# a_8953_45546# 4.65e-19
C5674 a_9313_45822# a_8016_46348# 0.02464f
C5675 a_6151_47436# a_11189_46129# 7.98e-21
C5676 a_n1435_47204# a_6165_46155# 1.3e-20
C5677 a_9067_47204# a_5937_45572# 1.6e-19
C5678 a_4915_47217# a_10903_43370# 0.004769f
C5679 SMPL_ON_P a_n2956_39304# 0.039212f
C5680 a_n2497_47436# a_n967_46494# 7.99e-21
C5681 a_n971_45724# a_6945_45028# 0.247957f
C5682 a_2107_46812# a_3090_45724# 0.003997f
C5683 a_5807_45002# a_13059_46348# 0.1145f
C5684 a_12549_44172# a_18285_46348# 0.008787f
C5685 a_16131_47204# a_16388_46812# 2.48e-19
C5686 a_7411_46660# a_7715_46873# 0.162909f
C5687 a_15928_47570# a_765_45546# 0.003038f
C5688 a_3877_44458# a_6086_46660# 0.002133f
C5689 a_4817_46660# a_6969_46634# 5.31e-20
C5690 a_5257_43370# a_7577_46660# 4.41e-20
C5691 a_18911_45144# a_19268_43646# 5.23e-21
C5692 a_1307_43914# a_3935_42891# 0.318189f
C5693 a_17730_32519# a_15493_43940# 0.006052f
C5694 a_n2661_43922# a_n2433_43396# 0.001232f
C5695 a_n2661_42834# a_n2129_43609# 0.009349f
C5696 a_18494_42460# a_18525_43370# 4.73e-19
C5697 a_18184_42460# a_18783_43370# 2.81e-21
C5698 a_7281_43914# a_7584_44260# 0.001377f
C5699 a_n2293_43922# a_n4318_39304# 5.19e-19
C5700 a_n356_44636# a_2982_43646# 0.434193f
C5701 a_n2661_44458# a_10341_43396# 7.76e-20
C5702 a_11691_44458# a_16137_43396# 5.49e-20
C5703 a_19778_44110# a_15743_43084# 0.00304f
C5704 a_n2017_45002# a_n914_42852# 1.25e-19
C5705 en_comp a_22223_42860# 4.89e-22
C5706 a_n2810_45028# a_n2293_42282# 1.93e-20
C5707 a_9313_44734# VDD 0.389068f
C5708 a_n3420_39072# VIN_P 0.031754f
C5709 a_n3420_38528# C5_P_btm 0.001712f
C5710 a_n4064_38528# C7_P_btm 1.64e-19
C5711 a_n3565_39304# VREF 0.098117f
C5712 a_n4209_39304# VCM 0.05604f
C5713 a_6667_45809# a_7227_45028# 4.77e-19
C5714 a_2711_45572# a_4808_45572# 9.57e-19
C5715 a_4093_43548# a_4646_46812# 3.43e-21
C5716 a_9801_43940# a_8270_45546# 0.014887f
C5717 a_14205_43396# a_13661_43548# 2.89e-19
C5718 a_14485_44260# a_15227_44166# 4.39e-21
C5719 a_7274_43762# a_n2293_46634# 1.42e-19
C5720 a_n2661_44458# a_n356_45724# 8.5e-21
C5721 a_17970_44736# a_16375_45002# 0.00591f
C5722 a_18443_44721# a_13259_45724# 0.004991f
C5723 a_n1352_44484# a_n755_45592# 1.52e-20
C5724 a_n699_43396# a_n863_45724# 0.23135f
C5725 a_19006_44850# a_17715_44484# 1.14e-20
C5726 a_4361_42308# a_18597_46090# 0.024928f
C5727 a_4520_42826# a_4791_45118# 1.52e-19
C5728 a_20447_31679# a_22609_37990# 9.79e-21
C5729 a_n3565_38502# a_n4064_38528# 0.228245f
C5730 a_5072_46660# VDD 0.081835f
C5731 a_4958_30871# C2_N_btm 9.53e-20
C5732 COMP_P VDAC_Ni 9.79e-19
C5733 a_765_45546# a_1138_42852# 0.02041f
C5734 a_22365_46825# a_20202_43084# 0.115624f
C5735 a_16388_46812# a_3483_46348# 4.06e-21
C5736 a_n2442_46660# a_n2661_45546# 6.66e-19
C5737 a_768_44030# a_n443_42852# 0.00732f
C5738 a_5257_43370# a_5431_46482# 9.25e-20
C5739 a_n2293_46634# a_n2810_45572# 5.41e-20
C5740 a_n2661_46634# a_n2956_38216# 3.93e-19
C5741 a_15368_46634# a_13759_46122# 1.21e-20
C5742 a_12816_46660# a_2324_44458# 1.64e-21
C5743 a_14976_45028# a_13925_46122# 1.92e-19
C5744 a_n1761_44111# a_n1991_42858# 1.58e-21
C5745 a_n1899_43946# a_n1853_43023# 4.54e-20
C5746 a_18451_43940# a_10341_43396# 1.01e-20
C5747 a_5244_44056# a_743_42282# 1.87e-21
C5748 a_n2267_43396# a_n1177_43370# 0.041762f
C5749 a_n1699_43638# a_n1917_43396# 0.209641f
C5750 a_n2129_43609# a_n1352_43396# 0.041828f
C5751 a_n2433_43396# a_n447_43370# 1.32e-20
C5752 a_11341_43940# a_9145_43396# 0.017582f
C5753 a_15493_43396# a_14955_43396# 0.076347f
C5754 a_n1331_43914# a_n2157_42858# 3.92e-20
C5755 a_1307_43914# a_15890_42674# 3.24e-21
C5756 a_n2810_45028# a_n3565_39590# 0.021277f
C5757 en_comp a_n4209_39590# 7.54e-19
C5758 a_20974_43370# VDD 0.550101f
C5759 a_13527_45546# a_9482_43914# 7.42e-19
C5760 a_13163_45724# a_13556_45296# 0.001027f
C5761 a_11823_42460# a_14180_45002# 6.93e-21
C5762 a_7499_43078# a_1423_45028# 0.020575f
C5763 a_2711_45572# a_8488_45348# 5.77e-19
C5764 a_8192_45572# a_3232_43370# 5.95e-19
C5765 a_8120_45572# a_6171_45002# 6.76e-19
C5766 a_8685_43396# a_8199_44636# 0.03394f
C5767 a_6031_43396# a_2324_44458# 2.16e-20
C5768 a_104_43370# a_n1925_42282# 4.1e-21
C5769 a_20935_43940# a_n357_42282# 2.76e-19
C5770 a_13483_43940# a_n443_42852# 2.18e-20
C5771 a_7871_42858# a_3090_45724# 1.56e-20
C5772 a_14205_43396# a_4185_45028# 4.43e-21
C5773 a_18783_43370# a_12741_44636# 4.28e-21
C5774 a_14955_43396# a_3483_46348# 1.76e-19
C5775 a_10057_43914# CLK 1.02e-19
C5776 a_10053_45546# a_6151_47436# 2.75e-22
C5777 a_8746_45002# a_4915_47217# 9.87e-21
C5778 a_12791_45546# a_n1151_42308# 1.07e-20
C5779 a_17583_46090# a_13259_45724# 0.191869f
C5780 a_14493_46090# a_15002_46116# 2.6e-19
C5781 a_1176_45822# a_n443_42852# 0.071187f
C5782 a_3147_46376# a_3503_45724# 5.03e-19
C5783 a_3483_46348# a_3316_45546# 1.91e-21
C5784 a_7287_43370# a_7227_42852# 0.008095f
C5785 a_16759_43396# a_16823_43084# 0.038761f
C5786 a_2813_43396# a_1847_42826# 2.9e-19
C5787 a_3626_43646# a_10922_42852# 4.54e-20
C5788 a_2982_43646# a_12379_42858# 1.63e-19
C5789 a_n2661_42282# a_1067_42314# 8.97e-20
C5790 a_16137_43396# a_4190_30871# 0.113768f
C5791 a_16977_43638# a_17433_43396# 4.2e-19
C5792 a_10341_43396# a_17364_32525# 5.25e-19
C5793 a_19862_44208# a_22400_42852# 5.55e-21
C5794 a_3080_42308# a_5534_30871# 0.019853f
C5795 a_1123_46634# DATA[1] 0.00365f
C5796 a_18599_43230# VDD 0.197104f
C5797 a_13249_42308# a_11967_42832# 0.023012f
C5798 a_2711_45572# a_1414_42308# 1.75e-21
C5799 a_15595_45028# a_15685_45394# 0.004764f
C5800 a_14537_43396# a_14309_45028# 0.006215f
C5801 a_n745_45366# a_n452_44636# 0.001046f
C5802 a_n143_45144# a_n2661_44458# 4.34e-20
C5803 a_n467_45028# a_n2433_44484# 2.79e-19
C5804 a_n913_45002# a_742_44458# 0.302053f
C5805 a_n1059_45260# a_949_44458# 2.96e-19
C5806 a_n2293_45010# a_n699_43396# 0.005002f
C5807 a_22400_42852# a_4185_45028# 0.105692f
C5808 a_15803_42450# a_15227_44166# 0.006356f
C5809 a_n1641_43230# a_n357_42282# 2.03e-19
C5810 a_13291_42460# a_10903_43370# 0.135558f
C5811 a_14403_45348# a_4915_47217# 1.22e-19
C5812 a_14537_43396# a_11453_44696# 0.029591f
C5813 a_6431_45366# a_n1613_43370# 0.006556f
C5814 a_6171_45002# a_n881_46662# 0.090566f
C5815 a_n2661_45010# a_n2956_39768# 1.22e-20
C5816 a_2437_43646# a_n133_46660# 3.38e-21
C5817 a_2680_45002# a_768_44030# 0.028861f
C5818 a_10193_42453# a_15227_44166# 0.205591f
C5819 a_11823_42460# a_15009_46634# 2.01e-21
C5820 a_743_42282# a_n473_42460# 1.85e-19
C5821 a_22165_42308# a_22223_42860# 0.171681f
C5822 a_3626_43646# a_17531_42308# 0.003944f
C5823 a_2982_43646# a_18727_42674# 1.36e-19
C5824 a_n4318_39304# a_n3420_39616# 0.256393f
C5825 a_8952_43230# a_9114_42852# 0.006453f
C5826 a_4190_30871# a_n784_42308# 0.019472f
C5827 a_8873_43396# a_5934_30871# 4.31e-21
C5828 a_14209_32519# a_22765_42852# 4.61e-20
C5829 a_11133_46155# CLK 0.001561f
C5830 a_14840_46494# RST_Z 2.03e-21
C5831 a_22397_42558# VDD 0.006424f
C5832 a_n815_47178# a_n881_46662# 2.82e-20
C5833 a_n1741_47186# a_5159_47243# 1.44e-19
C5834 a_4915_47217# a_4883_46098# 0.024005f
C5835 a_14955_47212# a_15507_47210# 5.87e-19
C5836 a_14311_47204# a_15811_47375# 6.14e-21
C5837 a_584_46384# a_2747_46873# 2.14e-19
C5838 a_2063_45854# a_2487_47570# 0.003691f
C5839 a_1209_47178# a_3315_47570# 4.55e-20
C5840 a_13717_47436# a_16327_47482# 2.02e-19
C5841 a_12861_44030# a_16241_47178# 3e-20
C5842 a_11031_47542# a_10227_46804# 3.37e-19
C5843 a_n1151_42308# a_n2312_40392# 1.57e-19
C5844 a_17613_45144# a_11967_42832# 8.83e-21
C5845 a_21359_45002# a_17517_44484# 9.2e-20
C5846 a_n2433_44484# a_n2661_43922# 0.075698f
C5847 a_n2129_44697# a_n2661_42834# 0.001254f
C5848 a_8701_44490# a_5891_43370# 0.001099f
C5849 a_742_44458# a_556_44484# 0.044092f
C5850 a_16922_45042# a_20159_44458# 0.012027f
C5851 a_n2661_44458# a_n2293_43922# 1.21e-19
C5852 a_1307_43914# a_6453_43914# 0.006717f
C5853 a_8103_44636# a_8238_44734# 0.008535f
C5854 a_18443_44721# a_18989_43940# 0.0016f
C5855 a_11827_44484# a_17061_44734# 0.0048f
C5856 a_5111_44636# a_9672_43914# 0.001516f
C5857 a_n1059_45260# a_11341_43940# 4.96e-19
C5858 a_5205_44484# a_6756_44260# 1.27e-19
C5859 a_n3420_39072# a_n2956_38680# 0.001161f
C5860 a_n2946_39072# a_n2956_39304# 0.150476f
C5861 a_6123_31319# a_n443_42852# 6.89e-19
C5862 a_15037_45618# VDD 0.08759f
C5863 a_11787_45002# a_11415_45002# 0.072246f
C5864 a_2274_45254# a_1823_45246# 0.255985f
C5865 a_327_44734# a_167_45260# 0.199136f
C5866 a_5891_43370# a_n2293_46634# 0.105307f
C5867 a_9313_44734# a_22612_30879# 1.86e-20
C5868 a_13249_42308# a_13259_45724# 0.358931f
C5869 a_14495_45572# a_14383_46116# 6.09e-19
C5870 a_3775_45552# a_n755_45592# 0.100709f
C5871 a_11136_45572# a_8049_45260# 8.45e-20
C5872 a_11541_44484# a_11309_47204# 3.58e-22
C5873 a_14673_44172# a_n881_46662# 1.47e-19
C5874 a_18909_45814# a_10809_44734# 3.61e-23
C5875 a_3357_43084# a_9290_44172# 5.59e-22
C5876 a_21073_44484# a_18479_47436# 5.66e-19
C5877 a_1606_42308# a_2713_42308# 0.002318f
C5878 a_n2293_42282# a_n2302_40160# 3.05e-20
C5879 a_17538_32519# VDAC_N 0.005064f
C5880 a_12891_46348# a_6755_46942# 0.025465f
C5881 a_5807_45002# a_7577_46660# 0.003957f
C5882 a_n2661_46634# a_5907_46634# 0.006487f
C5883 a_n1925_46634# a_4646_46812# 0.089593f
C5884 a_2107_46812# a_3699_46634# 0.004263f
C5885 a_601_46902# a_1057_46660# 4.2e-19
C5886 a_1110_47026# a_n2661_46098# 3.75e-20
C5887 a_11453_44696# a_3090_45724# 0.232756f
C5888 a_12465_44636# a_16292_46812# 2.02e-20
C5889 a_13507_46334# a_19333_46634# 0.009057f
C5890 a_20990_47178# a_19692_46634# 1.02e-20
C5891 a_14311_47204# a_13059_46348# 7.47e-21
C5892 a_10227_46804# a_12347_46660# 0.004629f
C5893 a_15811_47375# a_14226_46987# 2.43e-21
C5894 a_12861_44030# a_16721_46634# 0.070721f
C5895 a_9863_47436# a_765_45546# 0.001205f
C5896 a_n2109_47186# a_n901_46420# 9.56e-21
C5897 a_n1917_44484# a_n1699_43638# 2.44e-20
C5898 a_n1177_44458# a_n2267_43396# 2.68e-21
C5899 a_15433_44458# a_14955_43940# 0.005438f
C5900 a_n2065_43946# a_n1549_44318# 0.110816f
C5901 a_n1761_44111# a_n1331_43914# 0.043168f
C5902 a_n1699_44726# a_n1917_43396# 8.81e-20
C5903 a_n2661_44458# a_n97_42460# 3.24e-21
C5904 a_10193_42453# a_14635_42282# 0.00461f
C5905 a_18184_42460# a_3626_43646# 0.052679f
C5906 a_11823_42460# a_12800_43218# 0.00522f
C5907 a_9313_44734# a_22959_43948# 5.71e-19
C5908 a_5111_44636# a_743_42282# 0.024053f
C5909 a_n967_45348# a_n2157_42858# 0.02564f
C5910 a_n913_45002# a_n901_43156# 0.075029f
C5911 en_comp a_n1853_43023# 2.91e-19
C5912 a_n1059_45260# a_n1076_43230# 0.001392f
C5913 a_n2017_45002# a_n13_43084# 8.63e-19
C5914 a_413_45260# a_14209_32519# 3.38e-20
C5915 a_n4334_37440# VDD 0.385859f
C5916 a_18114_32519# VDD 0.550312f
C5917 a_22465_38105# a_22821_38993# 0.09356f
C5918 a_4958_30871# C8_P_btm 0.001147f
C5919 a_n1557_42282# a_n1613_43370# 1.85e-19
C5920 a_18374_44850# a_17715_44484# 6.22e-20
C5921 a_12607_44458# a_10809_44734# 0.0024f
C5922 a_8783_44734# a_8199_44636# 0.00224f
C5923 a_18248_44752# a_18819_46122# 2.46e-21
C5924 a_18287_44626# a_17957_46116# 2.68e-21
C5925 a_16501_45348# a_16375_45002# 0.00327f
C5926 a_17613_45144# a_13259_45724# 0.002217f
C5927 a_2779_44458# a_526_44458# 0.090804f
C5928 a_20512_43084# a_17339_46660# 1.02e-19
C5929 a_9165_43940# a_2107_46812# 1.02e-19
C5930 a_17538_32519# a_21588_30879# 0.055813f
C5931 a_n2661_42834# a_3483_46348# 0.0234f
C5932 a_n2661_43922# a_3147_46376# 3.32e-21
C5933 a_10180_45724# CLK 0.095799f
C5934 a_n4315_30879# a_n2946_39866# 4.06e-20
C5935 a_n4064_40160# a_n3690_39616# 2.54e-19
C5936 a_13569_47204# VDD 0.00491f
C5937 a_1606_42308# C8_N_btm 6.73e-20
C5938 a_3090_45724# a_17639_46660# 5.38e-20
C5939 a_15227_44166# a_21363_46634# 1.47e-19
C5940 a_19692_46634# a_20273_46660# 0.02419f
C5941 a_14513_46634# a_16388_46812# 2.55e-21
C5942 a_12891_46348# a_8049_45260# 0.035062f
C5943 a_n2438_43548# a_n2956_39304# 0.014879f
C5944 a_n1925_46634# a_n1545_46494# 6.83e-19
C5945 a_4883_46098# a_20850_46482# 2.25e-19
C5946 a_11813_46116# a_11415_45002# 4.47e-21
C5947 a_15493_43940# a_17538_32519# 0.013565f
C5948 a_11967_42832# a_19700_43370# 1.03e-21
C5949 a_n2661_42834# a_n2840_42826# 0.174935f
C5950 a_3499_42826# a_3540_43646# 0.007239f
C5951 a_3905_42865# a_3457_43396# 5.36e-20
C5952 a_n356_44636# a_7871_42858# 2.26e-20
C5953 a_375_42282# a_n784_42308# 0.004284f
C5954 a_14021_43940# a_13565_43940# 0.001756f
C5955 a_22959_43948# a_20974_43370# 0.005835f
C5956 a_5111_44636# a_5755_42308# 6.35e-19
C5957 a_n913_45002# a_10533_42308# 0.246621f
C5958 a_n1059_45260# a_10723_42308# 5.28e-20
C5959 a_n2017_45002# a_11323_42473# 0.003882f
C5960 a_3537_45260# a_6773_42558# 0.001736f
C5961 a_17737_43940# VDD 0.285511f
C5962 a_15599_45572# a_16223_45938# 9.73e-19
C5963 a_15903_45785# a_16020_45572# 0.157972f
C5964 a_16855_45546# a_16680_45572# 0.233657f
C5965 a_16115_45572# a_8696_44636# 7.81e-20
C5966 a_15765_45572# a_17478_45572# 2.62e-19
C5967 a_10193_42453# a_2437_43646# 2.74e-20
C5968 a_13667_43396# a_13059_46348# 0.00451f
C5969 a_16137_43396# a_15227_44166# 0.002078f
C5970 a_1467_44172# a_n863_45724# 0.021736f
C5971 a_n809_44244# a_n357_42282# 0.001553f
C5972 a_8483_43230# a_n1613_43370# 5.99e-19
C5973 a_19273_43230# a_16327_47482# 9.01e-20
C5974 a_7754_38470# CAL_P 1.73e-19
C5975 a_18114_32519# a_22469_39537# 2.15e-20
C5976 a_2202_46116# VDD 0.20904f
C5977 a_21613_42308# a_22469_40625# 1.4e-21
C5978 a_22775_42308# a_22521_40599# 1.89e-20
C5979 a_n4209_38216# a_n3690_38304# 0.045342f
C5980 a_n3565_39590# a_n2302_37690# 2.81e-19
C5981 a_2112_39137# VDAC_Pi 0.01062f
C5982 a_n3607_38528# a_n3420_37984# 3.77e-20
C5983 C2_N_btm C7_N_btm 0.138288f
C5984 C3_N_btm C6_N_btm 0.133742f
C5985 C4_N_btm C5_N_btm 18.6196f
C5986 C0_dummy_N_btm C10_N_btm 0.749362f
C5987 C0_N_btm C9_N_btm 0.146135f
C5988 C1_N_btm C8_N_btm 0.129306f
C5989 a_3483_46348# a_5066_45546# 0.081087f
C5990 a_10903_43370# a_10809_44734# 0.353301f
C5991 a_17583_46090# a_18189_46348# 7.78e-19
C5992 a_12594_46348# a_6945_45028# 5.55e-20
C5993 a_n1699_43638# a_n1853_43023# 7.66e-20
C5994 a_n2267_43396# a_n1991_42858# 3.69e-20
C5995 a_n1917_43396# a_n2157_42858# 1.43e-19
C5996 a_n2433_43396# a_n1641_43230# 0.001096f
C5997 a_4235_43370# a_743_42282# 1.55e-19
C5998 a_14579_43548# a_14205_43396# 0.066243f
C5999 a_9145_43396# a_10341_43396# 0.085699f
C6000 a_n2129_43609# a_n1423_42826# 1.14e-19
C6001 a_14021_43940# a_5534_30871# 1.65e-19
C6002 a_11341_43940# a_19987_42826# 1.11e-19
C6003 a_21115_43940# a_20922_43172# 6.4e-20
C6004 a_15493_43940# a_19339_43156# 2.37e-20
C6005 a_9313_44734# a_11551_42558# 8.33e-20
C6006 a_n2293_43922# a_8325_42308# 4.97e-20
C6007 a_9803_43646# a_9885_43646# 0.171361f
C6008 a_8685_43396# a_8945_43396# 3.33e-19
C6009 a_3422_30871# COMP_P 0.208163f
C6010 a_3080_42308# a_4190_30871# 0.01835f
C6011 a_13507_46334# CLK 8.83e-20
C6012 a_4883_46098# DATA[5] 2.29e-20
C6013 a_13887_32519# VDD 0.424101f
C6014 a_18341_45572# a_19113_45348# 5.8e-19
C6015 a_19431_45546# a_11827_44484# 1.24e-20
C6016 a_18479_45785# a_11691_44458# 0.025645f
C6017 a_8162_45546# a_8375_44464# 1.5e-21
C6018 a_16147_45260# a_16237_45028# 0.005426f
C6019 a_11963_45334# a_13017_45260# 3.97e-20
C6020 a_4558_45348# a_1423_45028# 1.71e-19
C6021 a_6171_45002# a_1307_43914# 0.037515f
C6022 a_13460_43230# a_10903_43370# 3.23e-19
C6023 a_5342_30871# a_9290_44172# 6.73e-19
C6024 a_6809_43396# a_n443_42852# 5.25e-19
C6025 a_n1076_43230# a_n1925_42282# 1.95e-20
C6026 a_14955_43396# a_n357_42282# 6.56e-20
C6027 a_n13_43084# a_526_44458# 2.42e-19
C6028 a_7174_31319# a_n2312_38680# 3.87e-21
C6029 a_22465_38105# a_21588_30879# 7.99e-19
C6030 a_22223_42860# a_4185_45028# 2.62e-20
C6031 a_8696_44636# a_5807_45002# 0.024228f
C6032 a_7499_43078# a_4646_46812# 0.158236f
C6033 a_2711_45572# a_10428_46928# 4.68e-20
C6034 a_16855_45546# a_13747_46662# 0.02676f
C6035 a_7227_45028# a_5257_43370# 7.21e-21
C6036 a_13485_45572# a_768_44030# 9.77e-20
C6037 a_14033_45572# a_12549_44172# 2.6e-19
C6038 a_18909_45814# a_n881_46662# 1.16e-20
C6039 a_3357_43084# a_20990_47178# 1.67e-19
C6040 a_2437_43646# a_21496_47436# 0.01965f
C6041 a_22223_45572# a_13507_46334# 0.015966f
C6042 a_21513_45002# a_4883_46098# 0.005388f
C6043 a_n1059_45260# a_16327_47482# 0.235708f
C6044 a_413_45260# a_13381_47204# 1.38e-19
C6045 a_8191_45002# a_n1151_42308# 7.92e-19
C6046 a_6431_45366# a_4791_45118# 1.75e-20
C6047 a_n755_45592# a_3218_45724# 0.045755f
C6048 a_380_45546# a_n23_45546# 0.002746f
C6049 a_n1099_45572# a_n356_45724# 0.070228f
C6050 a_n2661_45546# a_1609_45822# 0.02204f
C6051 a_n1079_45724# a_n1013_45572# 0.010598f
C6052 a_n452_45724# a_n310_45899# 0.005572f
C6053 a_4905_42826# a_4921_42308# 0.046918f
C6054 a_8952_43230# a_10518_42984# 0.002305f
C6055 a_9127_43156# a_10835_43094# 4.52e-21
C6056 a_3539_42460# a_2713_42308# 8.99e-20
C6057 a_2982_43646# a_3823_42558# 0.006269f
C6058 a_n97_42460# a_8325_42308# 3e-19
C6059 a_14021_43940# a_19647_42308# 1.51e-21
C6060 a_21076_30879# a_19864_35138# 5.61e-20
C6061 a_18900_46660# START 2.58e-19
C6062 a_21363_46634# EN_OFFSET_CAL 4.24e-21
C6063 a_7754_38470# CAL_N 3.08e-19
C6064 a_8530_39574# a_11206_38545# 0.046219f
C6065 a_8515_42308# VDD 0.194691f
C6066 a_n1741_47186# a_5815_47464# 0.021904f
C6067 a_584_46384# a_2063_45854# 0.406382f
C6068 a_n971_45724# a_4700_47436# 8.66e-19
C6069 a_327_47204# a_n1151_42308# 0.013822f
C6070 a_n237_47217# a_3815_47204# 1.74e-20
C6071 a_1209_47178# a_3160_47472# 1.39e-19
C6072 a_18587_45118# a_18287_44626# 3.25e-20
C6073 a_18911_45144# a_18248_44752# 3.13e-19
C6074 a_n2267_44484# a_n1177_44458# 0.042415f
C6075 a_18315_45260# a_18443_44721# 4.68e-19
C6076 a_n1699_44726# a_n1917_44484# 0.209641f
C6077 a_n2129_44697# a_n1352_44484# 0.048248f
C6078 a_n2433_44484# a_n452_44636# 1.17e-20
C6079 a_n2661_44458# a_742_44458# 0.026794f
C6080 a_11827_44484# a_13076_44458# 0.007928f
C6081 a_1307_43914# a_14673_44172# 0.012594f
C6082 a_14537_43396# a_15146_44484# 0.002264f
C6083 a_11691_44458# a_10057_43914# 1.34e-20
C6084 a_13556_45296# a_16335_44484# 1.13e-19
C6085 a_n2661_43370# a_7640_43914# 1.31e-19
C6086 a_10193_42453# a_11257_43940# 2.15e-19
C6087 a_15861_45028# a_15493_43396# 1.31e-20
C6088 a_n913_45002# a_n984_44318# 0.013973f
C6089 a_n745_45366# a_n809_44244# 1.57e-19
C6090 a_413_45260# a_17730_32519# 0.026007f
C6091 a_n2661_45010# a_453_43940# 0.004674f
C6092 a_3357_43084# a_3905_42865# 0.125186f
C6093 a_n967_45348# a_n1761_44111# 0.015839f
C6094 a_n2293_45010# a_1467_44172# 1.84e-19
C6095 a_19326_42852# a_n357_42282# 1.44e-19
C6096 a_n1736_42282# a_n2810_45572# 2.3e-20
C6097 a_n4318_38216# a_n2956_38216# 0.023519f
C6098 a_2711_45572# VDD 1.22011f
C6099 a_13887_32519# a_22469_39537# 1.15e-20
C6100 a_8746_45002# a_10809_44734# 0.049227f
C6101 a_6709_45028# a_3090_45724# 1.32e-20
C6102 a_2437_43646# a_21363_46634# 2.82e-19
C6103 a_3357_43084# a_20273_46660# 0.02704f
C6104 a_6472_45840# a_5066_45546# 2.68e-19
C6105 a_18114_32519# a_22612_30879# 0.061298f
C6106 a_19721_31679# a_21588_30879# 0.055771f
C6107 a_5518_44484# a_768_44030# 0.00362f
C6108 a_n2661_43370# a_4651_46660# 1.49e-21
C6109 a_18787_45572# a_11415_45002# 7.51e-19
C6110 a_15861_45028# a_3483_46348# 2.64e-19
C6111 a_5342_30871# a_15051_42282# 0.029795f
C6112 a_15567_42826# a_14113_42308# 1.63e-20
C6113 a_5193_42852# a_5267_42460# 3.13e-19
C6114 a_14635_42282# a_n784_42308# 2.26e-20
C6115 a_5193_43172# a_5932_42308# 1.9e-21
C6116 a_768_44030# a_n2661_46634# 5.84e-20
C6117 a_13661_43548# a_13747_46662# 0.095862f
C6118 a_9804_47204# a_n1925_46634# 9.26e-22
C6119 a_n881_46662# a_171_46873# 0.018745f
C6120 a_n1613_43370# a_33_46660# 0.599895f
C6121 a_11031_47542# a_10467_46802# 1.42e-19
C6122 a_7903_47542# a_6755_46942# 9.91e-21
C6123 a_9313_45822# a_10428_46928# 1.12e-19
C6124 a_2063_45854# a_11901_46660# 0.001041f
C6125 a_11691_44458# a_14021_43940# 3.38e-19
C6126 a_17517_44484# a_19279_43940# 0.020718f
C6127 a_n2661_43922# a_n2840_43914# 0.171265f
C6128 a_n2661_42834# a_n2472_43914# 0.012267f
C6129 a_10193_42453# a_14543_43071# 1.03e-21
C6130 a_18479_45785# a_4190_30871# 0.123942f
C6131 a_11827_44484# a_15301_44260# 4.18e-19
C6132 a_7229_43940# a_7287_43370# 8.37e-20
C6133 a_n1059_45260# a_10341_43396# 0.037338f
C6134 a_1606_42308# C2_P_btm 0.021793f
C6135 a_4743_44484# a_1823_45246# 0.001634f
C6136 a_17767_44458# a_12741_44636# 2.58e-19
C6137 a_18287_44626# a_11415_45002# 9.88e-20
C6138 a_15493_43396# a_19321_45002# 1.18e-20
C6139 a_19862_44208# a_13747_46662# 0.15289f
C6140 a_10807_43548# a_n2293_46634# 0.05087f
C6141 a_20269_44172# a_13661_43548# 0.001724f
C6142 a_15146_44484# a_3090_45724# 7.43e-20
C6143 a_9895_44260# a_768_44030# 9.29e-19
C6144 a_n143_45144# a_n1099_45572# 8.04e-20
C6145 a_3065_45002# a_n2661_45546# 0.004264f
C6146 a_327_44734# a_n863_45724# 0.353745f
C6147 a_2274_45254# a_n2293_45546# 0.07158f
C6148 a_n659_45366# a_n755_45592# 4.7e-19
C6149 a_16922_45042# a_18819_46122# 9.18e-21
C6150 a_17719_45144# a_17715_44484# 0.009296f
C6151 a_n2661_44458# a_5204_45822# 5e-21
C6152 a_11827_44484# a_12594_46348# 5.74e-21
C6153 a_8147_43396# a_n971_45724# 0.116186f
C6154 a_548_43396# a_584_46384# 7.2e-19
C6155 a_6123_31319# a_1736_39587# 1.03e-19
C6156 a_n3674_37592# a_n3565_38216# 1.57e-19
C6157 a_n1630_35242# a_n4209_38216# 2.41e-19
C6158 a_16522_42674# a_4958_30871# 0.020415f
C6159 a_9313_45822# VDD 0.5747f
C6160 a_13678_32519# CAL_N 1.36e-19
C6161 a_n2293_46634# a_472_46348# 1.43e-21
C6162 a_171_46873# a_n2157_46122# 3.28e-21
C6163 a_n2661_46634# a_1176_45822# 4.24e-19
C6164 a_n1925_46634# a_n901_46420# 0.004832f
C6165 a_n2438_43548# a_n1991_46122# 0.001576f
C6166 a_33_46660# a_n2293_46098# 1.87e-20
C6167 a_13747_46662# a_4185_45028# 2.24e-20
C6168 a_6755_46942# a_12359_47026# 8.58e-19
C6169 a_11735_46660# a_12991_46634# 0.043475f
C6170 a_11901_46660# a_12469_46902# 0.175891f
C6171 a_5907_46634# a_765_45546# 0.003106f
C6172 a_10554_47026# a_10933_46660# 3.16e-19
C6173 a_11813_46116# a_12251_46660# 3.12e-19
C6174 a_10249_46116# a_10861_46660# 3.67e-19
C6175 a_768_44030# a_8199_44636# 0.026637f
C6176 a_n881_46662# a_10903_43370# 3.24e-19
C6177 a_11453_44696# a_20075_46420# 2.89e-20
C6178 a_12465_44636# a_6945_45028# 0.023497f
C6179 a_n2833_47464# a_n2840_45546# 3.38e-21
C6180 a_4883_46098# a_10809_44734# 0.068164f
C6181 a_7903_47542# a_8049_45260# 2.11e-20
C6182 a_n1899_43946# a_n1699_43638# 2.25e-19
C6183 a_n1761_44111# a_n1917_43396# 2.84e-19
C6184 a_n2065_43946# a_n1177_43370# 2.42e-19
C6185 a_n1549_44318# a_n2129_43609# 1.85e-20
C6186 a_19862_44208# a_20269_44172# 0.049487f
C6187 a_17973_43940# a_15493_43940# 0.028173f
C6188 a_18326_43940# a_11341_43940# 0.003644f
C6189 a_n1331_43914# a_n2267_43396# 0.001024f
C6190 a_n2661_43922# a_9803_43646# 1.71e-20
C6191 a_n2661_42834# a_10695_43548# 2.95e-20
C6192 a_n356_44636# a_17324_43396# 2.85e-21
C6193 a_n2661_44458# a_n901_43156# 5.46e-22
C6194 a_n1917_44484# a_n2157_42858# 1.66e-21
C6195 a_10193_42453# a_19511_42282# 0.133376f
C6196 a_10949_43914# a_12495_44260# 0.002649f
C6197 a_n2293_43922# a_9145_43396# 0.019866f
C6198 a_5343_44458# a_5649_42852# 3.17e-20
C6199 a_14539_43914# a_17486_43762# 1.39e-19
C6200 a_n2017_45002# a_20753_42852# 3.3e-20
C6201 a_19963_31679# COMP_P 2.93e-20
C6202 a_22485_44484# VDD 0.258874f
C6203 a_9049_44484# a_9159_45572# 0.007938f
C6204 a_10490_45724# a_11682_45822# 0.014138f
C6205 a_11525_45546# a_10907_45822# 4.14e-19
C6206 C2_N_btm C3_P_btm 1.33e-19
C6207 C3_N_btm C4_P_btm 1.02e-19
C6208 C1_N_btm C2_P_btm 2.79e-20
C6209 a_19987_42826# a_16327_47482# 0.053812f
C6210 a_9672_43914# a_9290_44172# 0.071844f
C6211 a_n2661_43922# a_310_45028# 2.83e-19
C6212 a_n2661_42834# a_n357_42282# 0.239713f
C6213 a_644_44056# a_526_44458# 3.05e-19
C6214 a_3363_44484# a_3316_45546# 3.64e-20
C6215 a_13887_32519# a_22612_30879# 0.060052f
C6216 a_5934_30871# VDAC_P 0.029185f
C6217 a_12816_46660# a_12839_46116# 1.51e-19
C6218 a_11415_45002# a_15682_46116# 1.66e-19
C6219 a_12741_44636# a_15015_46420# 1.62e-21
C6220 a_3147_46376# a_5164_46348# 1.45e-21
C6221 a_3483_46348# a_5068_46348# 4.35e-20
C6222 a_21188_46660# a_10809_44734# 0.010814f
C6223 a_4185_45028# a_4419_46090# 0.066314f
C6224 a_20935_43940# a_20749_43396# 1.23e-20
C6225 a_3626_43646# a_6293_42852# 6.33e-20
C6226 a_n97_42460# a_9145_43396# 4.77e-19
C6227 a_14021_43940# a_4190_30871# 0.086029f
C6228 a_15493_43940# a_22591_43396# 1.85e-20
C6229 a_n2661_42282# a_5111_42852# 4.21e-20
C6230 a_n356_44636# a_1184_42692# 0.03675f
C6231 a_5343_44458# a_7963_42308# 0.108654f
C6232 a_4093_43548# a_3457_43396# 7.01e-20
C6233 a_5883_43914# a_6481_42558# 9.74e-21
C6234 a_n1741_47186# CLK 0.028114f
C6235 a_n971_45724# DATA[2] 0.099284f
C6236 a_n237_47217# DATA[0] 0.040942f
C6237 a_n746_45260# DATA[1] 5.22e-20
C6238 a_11322_45546# a_11827_44484# 8.07e-20
C6239 a_2711_45572# a_n699_43396# 1.83e-20
C6240 a_n1059_45260# a_n143_45144# 4.32e-20
C6241 a_n2293_45010# a_327_44734# 6.84e-21
C6242 a_3357_43084# a_5147_45002# 0.09352f
C6243 a_n913_45002# a_n467_45028# 1.15e-19
C6244 a_18249_42858# a_17339_46660# 0.008924f
C6245 a_n1352_43396# a_n357_42282# 2.09e-19
C6246 a_n1177_43370# a_n755_45592# 3.74e-19
C6247 a_743_42282# a_9290_44172# 0.117511f
C6248 a_4361_42308# a_8953_45546# 0.012234f
C6249 a_19647_42308# a_13507_46334# 5.23e-19
C6250 a_n1079_45724# VDD 0.172275f
C6251 a_16855_45546# a_11599_46634# 0.002089f
C6252 a_15599_45572# a_16327_47482# 0.331892f
C6253 a_17478_45572# a_12861_44030# 3.55e-19
C6254 a_3357_43084# a_n2109_47186# 0.170493f
C6255 a_7227_45028# a_5807_45002# 6.28e-20
C6256 a_15781_43660# a_15567_42826# 2.55e-19
C6257 a_n2157_42858# a_n1853_43023# 0.290902f
C6258 a_10341_43396# a_19987_42826# 2.55e-19
C6259 a_743_42282# a_791_42968# 5.89e-19
C6260 a_n2472_42826# a_n1991_42858# 9.31e-19
C6261 a_n97_42460# a_19273_43230# 4.33e-20
C6262 a_16877_42852# VDD 0.192454f
C6263 a_14797_45144# a_15004_44636# 2.66e-19
C6264 a_16922_45042# a_18911_45144# 0.042178f
C6265 a_1423_45028# a_9838_44484# 0.254741f
C6266 a_1307_43914# a_12607_44458# 4.31e-20
C6267 a_14537_43396# a_16112_44458# 0.093722f
C6268 a_7499_43078# a_10405_44172# 0.132405f
C6269 a_14180_45002# a_14539_43914# 4.34e-20
C6270 a_n913_45002# a_n2661_43922# 0.024256f
C6271 a_n745_45366# a_n2661_42834# 3.35e-21
C6272 a_3537_45260# a_8375_44464# 0.10437f
C6273 a_n1059_45260# a_n2293_43922# 0.02309f
C6274 a_5111_44636# a_5289_44734# 0.001056f
C6275 a_5147_45002# a_5826_44734# 7.2e-19
C6276 a_n2293_42282# a_n357_42282# 0.01064f
C6277 a_133_42852# a_n863_45724# 1.03e-19
C6278 a_3626_43646# RST_Z 4.03e-19
C6279 a_3775_45552# a_3483_46348# 3.9e-20
C6280 a_18479_45785# a_15227_44166# 0.035756f
C6281 a_2304_45348# a_n2293_46634# 0.00666f
C6282 a_375_42282# a_n2438_43548# 2.84e-20
C6283 a_16147_45260# a_19466_46812# 3.68e-21
C6284 a_16333_45814# a_13059_46348# 3.56e-20
C6285 a_4558_45348# a_4646_46812# 7.53e-22
C6286 a_5147_45002# a_3877_44458# 1.31e-20
C6287 a_3357_43084# a_5841_46660# 1.99e-19
C6288 a_6194_45824# a_5164_46348# 4.82e-20
C6289 a_2711_45572# a_7920_46348# 0.001215f
C6290 a_5263_45724# a_5497_46414# 3.95e-21
C6291 a_11827_44484# a_12465_44636# 0.785011f
C6292 a_11691_44458# a_13507_46334# 3.47e-20
C6293 a_n310_44811# a_n746_45260# 0.002132f
C6294 a_18783_43370# a_17303_42282# 2.56e-21
C6295 a_15743_43084# a_4958_30871# 3.06e-20
C6296 a_19164_43230# a_20753_42852# 9.53e-20
C6297 a_5649_42852# a_12563_42308# 1.31e-19
C6298 a_4361_42308# a_14456_42282# 0.007582f
C6299 a_743_42282# a_15051_42282# 0.011096f
C6300 a_4190_30871# a_15764_42576# 9.01e-20
C6301 a_16137_43396# a_19511_42282# 0.002509f
C6302 a_19987_42826# a_20356_42852# 0.014848f
C6303 a_21195_42852# a_14097_32519# 2.56e-20
C6304 a_21671_42860# a_22400_42852# 8.4e-20
C6305 a_10586_45546# CLK 0.125859f
C6306 a_11599_46634# a_13661_43548# 0.078449f
C6307 a_14955_47212# a_13747_46662# 3.09e-21
C6308 a_15507_47210# a_5807_45002# 0.002062f
C6309 a_18479_47436# a_12549_44172# 0.015281f
C6310 a_10227_46804# a_15928_47570# 0.025137f
C6311 a_16327_47482# a_16285_47570# 0.001903f
C6312 a_16241_47178# a_16697_47582# 4.2e-19
C6313 a_15811_47375# a_16131_47204# 0.002108f
C6314 a_6545_47178# a_n1925_46634# 0.02342f
C6315 a_4883_46098# a_n881_46662# 0.193691f
C6316 a_9067_47204# a_n2661_46634# 1.36e-19
C6317 a_584_46384# a_645_46660# 3.21e-21
C6318 a_1431_47204# a_n2661_46098# 1.15e-19
C6319 a_n1151_42308# a_1983_46706# 4.68e-20
C6320 a_n443_46116# a_171_46873# 0.029327f
C6321 a_n237_47217# a_3524_46660# 1.32e-21
C6322 a_n2109_47186# a_3877_44458# 0.021838f
C6323 a_n1917_44484# a_n1761_44111# 3.33e-19
C6324 a_n2267_44484# a_n1331_43914# 7.69e-19
C6325 a_n1177_44458# a_n2065_43946# 0.001595f
C6326 a_18287_44626# a_11967_42832# 0.789765f
C6327 a_18374_44850# a_18588_44850# 0.097745f
C6328 a_n2661_44458# a_n984_44318# 1.3e-20
C6329 a_n1699_44726# a_n1899_43946# 1.33e-19
C6330 a_n2129_44697# a_n1549_44318# 7.49e-21
C6331 a_n2661_43370# a_10729_43914# 4.79e-19
C6332 a_556_44484# a_n2661_43922# 0.00482f
C6333 a_18443_44721# a_19006_44850# 0.049827f
C6334 a_18248_44752# a_19615_44636# 2.73e-19
C6335 a_3363_44484# a_n2661_42834# 0.003152f
C6336 a_3357_43084# a_4093_43548# 0.031759f
C6337 a_n1059_45260# a_n97_42460# 0.869353f
C6338 a_n2017_45002# a_104_43370# 7.08e-21
C6339 a_n967_45348# a_n2267_43396# 0.001133f
C6340 a_n2472_45002# VDD 0.217954f
C6341 a_18326_43940# a_16327_47482# 2.74e-20
C6342 a_14955_43940# a_10227_46804# 0.004814f
C6343 a_20935_43940# a_12861_44030# 0.02414f
C6344 a_6431_45366# a_6945_45028# 0.00135f
C6345 a_3232_43370# a_10809_44734# 0.158726f
C6346 a_6453_43914# a_n1613_43370# 0.007952f
C6347 a_13556_45296# a_15015_46420# 2.21e-20
C6348 a_13348_45260# a_2324_44458# 0.005924f
C6349 a_14537_43396# a_13925_46122# 6.19e-21
C6350 a_14180_45002# a_14493_46090# 6.1e-20
C6351 a_14797_45144# a_13759_46122# 2.6e-20
C6352 a_9482_43914# a_14840_46494# 6.56e-21
C6353 a_1307_43914# a_10903_43370# 0.065094f
C6354 a_413_45260# a_2981_46116# 0.002451f
C6355 a_20447_31679# a_8049_45260# 0.009404f
C6356 a_15004_44636# a_14976_45028# 0.001535f
C6357 a_2127_44172# a_768_44030# 0.002861f
C6358 a_5093_45028# a_3483_46348# 0.05597f
C6359 a_17023_45118# a_11415_45002# 0.004458f
C6360 a_9223_42460# a_9377_42558# 0.010303f
C6361 COMP_P a_7174_31319# 0.029185f
C6362 a_1606_42308# a_4958_30871# 0.019472f
C6363 a_n1838_35608# VIN_P 0.029423f
C6364 C8_P_btm C3_P_btm 0.134581f
C6365 C9_P_btm C2_P_btm 0.141891f
C6366 C7_P_btm C4_P_btm 0.145303f
C6367 C6_P_btm C5_P_btm 22.305399f
C6368 a_768_44030# a_765_45546# 0.033731f
C6369 a_12549_44172# a_17829_46910# 0.057751f
C6370 a_5257_43370# a_7715_46873# 1.05e-20
C6371 a_5807_45002# a_15227_46910# 1.37e-19
C6372 a_3877_44458# a_5841_46660# 9.39e-19
C6373 a_4817_46660# a_6755_46942# 5.52e-20
C6374 a_4646_46812# a_6999_46987# 4.77e-19
C6375 a_11453_44696# a_21076_30879# 8.96e-19
C6376 a_22959_47212# a_22959_46660# 0.025171f
C6377 a_9067_47204# a_8199_44636# 6.76e-22
C6378 a_6575_47204# a_5937_45572# 1.83e-20
C6379 a_n2497_47436# a_n1379_46482# 5.68e-19
C6380 a_n1151_42308# a_14275_46494# 0.003302f
C6381 a_18911_45144# a_15743_43084# 1.13e-21
C6382 a_22591_44484# a_15493_43940# 2.12e-21
C6383 a_n2661_43922# a_n4318_39304# 8.01e-19
C6384 a_22485_44484# a_22959_43948# 8.19e-19
C6385 a_n2661_42834# a_n2433_43396# 0.02044f
C6386 a_11827_44484# a_16409_43396# 1.18e-21
C6387 a_18184_42460# a_18525_43370# 6.19e-21
C6388 a_1307_43914# a_3681_42891# 0.236785f
C6389 a_18494_42460# a_18429_43548# 2.84e-20
C6390 a_7542_44172# a_n2661_42282# 1.24e-20
C6391 a_5343_44458# a_8685_43396# 2.44e-19
C6392 en_comp a_22165_42308# 4.83e-21
C6393 a_9241_44734# VDD 0.003445f
C6394 a_n3420_38528# C6_P_btm 8.47e-20
C6395 a_n3565_38502# C4_P_btm 0.042623f
C6396 a_n3565_38216# EN_VIN_BSTR_P 0.005343f
C6397 a_n4209_39304# VREF_GND 0.02097f
C6398 a_6667_45809# a_6598_45938# 0.209641f
C6399 a_6511_45714# a_7227_45028# 0.213161f
C6400 a_3175_45822# a_3260_45572# 1.48e-19
C6401 a_2711_45572# a_5024_45822# 3.69e-19
C6402 a_1414_42308# a_1823_45246# 0.002939f
C6403 a_6453_43914# a_n2293_46098# 0.002061f
C6404 a_453_43940# a_1138_42852# 0.018298f
C6405 a_14021_43940# a_15227_44166# 0.052407f
C6406 a_14205_43396# a_5807_45002# 9.38e-20
C6407 a_9420_43940# a_8270_45546# 0.007316f
C6408 a_14358_43442# a_13661_43548# 1.8e-19
C6409 a_5837_43396# a_n2293_46634# 1.35e-19
C6410 a_n2661_44458# a_3503_45724# 4.06e-21
C6411 a_n1177_44458# a_n755_45592# 1.63e-19
C6412 a_17767_44458# a_16375_45002# 0.00258f
C6413 a_18287_44626# a_13259_45724# 0.002131f
C6414 a_5891_43370# a_8049_45260# 0.00367f
C6415 a_n2293_43922# a_n1925_42282# 2.06056f
C6416 a_18588_44850# a_17715_44484# 4.47e-20
C6417 a_4190_30871# a_13507_46334# 0.186424f
C6418 a_13467_32519# a_18597_46090# 0.002694f
C6419 a_5649_42852# a_10227_46804# 2.58e-19
C6420 a_n4334_38528# a_n4064_38528# 0.449049f
C6421 a_n3690_38528# a_n3420_38528# 0.431104f
C6422 a_n3565_38502# a_n2946_38778# 0.406164f
C6423 a_n4209_38502# a_n2302_38778# 0.406492f
C6424 a_6540_46812# VDD 0.084698f
C6425 a_4958_30871# C1_N_btm 9.46e-20
C6426 a_13059_46348# a_3483_46348# 0.319214f
C6427 a_765_45546# a_1176_45822# 0.241847f
C6428 a_20885_46660# a_20202_43084# 2.46e-21
C6429 a_12549_44172# a_n443_42852# 0.069091f
C6430 a_n2442_46660# a_n2810_45572# 0.045104f
C6431 a_n2956_39768# a_n2956_38216# 0.043382f
C6432 a_n2472_46634# a_n2661_45546# 0.001532f
C6433 a_14976_45028# a_13759_46122# 1.44e-20
C6434 a_3090_45724# a_13925_46122# 1.1e-19
C6435 a_n2065_43946# a_n1991_42858# 1.27e-20
C6436 a_n1761_44111# a_n1853_43023# 0.019636f
C6437 a_n1899_43946# a_n2157_42858# 4.17e-19
C6438 a_3905_42865# a_743_42282# 3.39e-19
C6439 a_n2433_43396# a_n1352_43396# 0.102325f
C6440 a_n2267_43396# a_n1917_43396# 0.227165f
C6441 a_n2129_43609# a_n1177_43370# 0.08445f
C6442 a_1307_43914# a_15959_42545# 1.52e-21
C6443 a_15493_43396# a_15095_43370# 1.04e-20
C6444 a_n2956_37592# a_n4209_39590# 0.090416f
C6445 a_14401_32519# VDD 0.562673f
C6446 a_13527_45546# a_13348_45260# 0.002161f
C6447 a_11823_42460# a_13777_45326# 5.57e-20
C6448 a_8746_45002# a_1307_43914# 9.72e-20
C6449 a_13163_45724# a_9482_43914# 8.82e-21
C6450 a_10193_42453# a_16751_45260# 0.048213f
C6451 a_13249_42308# a_13017_45260# 1.91e-19
C6452 a_2711_45572# a_8137_45348# 7.99e-20
C6453 a_n3674_37592# a_n1613_43370# 8.6e-20
C6454 a_n97_42460# a_n1925_42282# 0.021883f
C6455 a_20623_43914# a_n357_42282# 1.2e-20
C6456 a_12429_44172# a_n443_42852# 1.23e-19
C6457 a_7227_42852# a_3090_45724# 3.82e-19
C6458 a_19268_43646# a_11415_45002# 2.56e-21
C6459 a_15095_43370# a_3483_46348# 1.36e-21
C6460 a_10440_44484# CLK 0.013272f
C6461 a_9049_44484# a_6151_47436# 3.15e-20
C6462 a_10193_42453# a_4915_47217# 1.89e-20
C6463 a_11823_42460# a_n1151_42308# 9.67e-20
C6464 a_3483_46348# a_3218_45724# 1.76e-19
C6465 a_3147_46376# a_3316_45546# 0.012262f
C6466 a_1176_45822# a_509_45822# 1.26e-19
C6467 a_15682_46116# a_13259_45724# 0.002706f
C6468 a_13925_46122# a_15002_46116# 1.46e-19
C6469 a_5937_45572# a_n2661_45546# 1.02e-19
C6470 a_20365_43914# a_20256_43172# 4.57e-20
C6471 a_n2433_43396# a_n2293_42282# 7.51e-20
C6472 a_16977_43638# a_16823_43084# 0.022663f
C6473 a_10341_43396# a_22959_43396# 0.001295f
C6474 a_3626_43646# a_10991_42826# 1e-19
C6475 a_2982_43646# a_10341_42308# 4.06e-20
C6476 a_n2661_42282# a_n1630_35242# 0.093522f
C6477 a_11967_42832# a_17124_42282# 0.067231f
C6478 a_17324_43396# a_17486_43762# 0.006453f
C6479 a_16759_43396# a_17021_43396# 0.001705f
C6480 a_16409_43396# a_17433_43396# 2.36e-20
C6481 a_n2293_43922# a_n4315_30879# 2.47e-20
C6482 a_14021_43940# a_14635_42282# 6.42e-20
C6483 a_19862_44208# a_20836_43172# 8.42e-20
C6484 a_n743_46660# CLK 0.028835f
C6485 a_18817_42826# VDD 0.204624f
C6486 a_20447_31679# a_22469_40625# 1.91e-20
C6487 a_1423_45028# a_n2661_43370# 0.027675f
C6488 a_14180_45002# a_14309_45028# 0.062574f
C6489 a_n467_45028# a_n2661_44458# 0.031118f
C6490 a_n1059_45260# a_742_44458# 0.030569f
C6491 a_413_45260# a_19721_31679# 0.116395f
C6492 a_n967_45348# a_n2267_44484# 1.92e-19
C6493 a_15764_42576# a_15227_44166# 0.003122f
C6494 a_n1423_42826# a_n357_42282# 5.7e-19
C6495 a_4156_43218# a_526_44458# 2.93e-19
C6496 a_13003_42852# a_10903_43370# 0.006128f
C6497 a_14401_32519# a_22469_39537# 1.48e-20
C6498 a_3754_38470# w_1575_34946# 6.84e-19
C6499 a_1307_43914# a_4883_46098# 0.026965f
C6500 a_14309_45348# a_4915_47217# 0.002491f
C6501 a_14180_45002# a_11453_44696# 0.005785f
C6502 a_6171_45002# a_n1613_43370# 0.026867f
C6503 a_3232_43370# a_n881_46662# 0.001015f
C6504 a_3357_43084# a_n1925_46634# 0.034378f
C6505 a_2437_43646# a_n2438_43548# 0.045715f
C6506 a_2382_45260# a_768_44030# 0.094536f
C6507 a_13163_45724# a_12816_46660# 1.14e-19
C6508 a_743_42282# a_n961_42308# 1.36e-19
C6509 a_21671_42860# a_22223_42860# 3.81e-19
C6510 a_3626_43646# a_17303_42282# 0.037411f
C6511 a_2982_43646# a_18057_42282# 9.61e-20
C6512 a_10083_42826# a_10553_43218# 0.007399f
C6513 a_11189_46129# CLK 3.69e-19
C6514 a_15015_46420# RST_Z 4.05e-21
C6515 a_n815_47178# a_n1613_43370# 2.12e-19
C6516 a_n971_45724# a_3094_47243# 2.1e-19
C6517 a_14955_47212# a_11599_46634# 0.011007f
C6518 a_14311_47204# a_15507_47210# 8.1e-22
C6519 a_584_46384# a_2487_47570# 0.005904f
C6520 a_1209_47178# a_3094_47570# 7.14e-20
C6521 a_13717_47436# a_16241_47178# 6.54e-20
C6522 a_12861_44030# a_15673_47210# 5.52e-20
C6523 a_n443_46116# a_4883_46098# 0.037308f
C6524 a_17023_45118# a_11967_42832# 5.47e-20
C6525 a_21101_45002# a_17517_44484# 1.93e-19
C6526 a_18287_44626# a_18989_43940# 0.193279f
C6527 a_n2661_44458# a_n2661_43922# 6.64988f
C6528 a_n2433_44484# a_n2661_42834# 0.002352f
C6529 a_8103_44636# a_5891_43370# 0.029956f
C6530 a_1423_45028# a_2998_44172# 0.006884f
C6531 a_8701_44490# a_8375_44464# 0.001158f
C6532 a_18443_44721# a_18374_44850# 0.209641f
C6533 a_1307_43914# a_5663_43940# 0.11718f
C6534 a_5883_43914# a_7640_43914# 0.003384f
C6535 a_5111_44636# a_9028_43914# 3.72e-19
C6536 en_comp a_19862_44208# 4.89e-21
C6537 a_5205_44484# a_n2661_42282# 2.56e-19
C6538 a_n2017_45002# a_11341_43940# 9e-20
C6539 a_17124_42282# a_13259_45724# 0.003167f
C6540 a_n3420_39072# a_n2956_39304# 0.208204f
C6541 a_7227_42308# a_n443_42852# 8.04e-21
C6542 a_5742_30871# a_n863_45724# 2.35e-20
C6543 a_14033_45822# VDD 0.195067f
C6544 a_413_45260# a_167_45260# 0.120357f
C6545 a_1667_45002# a_1823_45246# 0.24808f
C6546 a_6171_45002# a_n2293_46098# 2.23e-21
C6547 a_8375_44464# a_n2293_46634# 1.16e-21
C6548 a_9313_44734# a_21588_30879# 1.69e-20
C6549 en_comp a_4185_45028# 0.001836f
C6550 a_13904_45546# a_13259_45724# 0.007639f
C6551 a_13249_42308# a_14383_46116# 7.26e-20
C6552 a_18341_45572# a_10809_44734# 6.97e-21
C6553 a_2437_43646# a_11133_46155# 3.61e-22
C6554 a_n2661_42282# a_n971_45724# 3.65e-19
C6555 a_n784_42308# a_4921_42308# 4.81e-20
C6556 a_5534_30871# a_n3420_39072# 0.339008f
C6557 COMP_P a_5932_42308# 0.029797f
C6558 a_14635_42282# a_15764_42576# 9.01e-21
C6559 a_5807_45002# a_7715_46873# 0.029268f
C6560 a_n1925_46634# a_3877_44458# 0.070082f
C6561 a_n2661_46634# a_5167_46660# 0.007924f
C6562 a_2107_46812# a_2959_46660# 0.003474f
C6563 a_33_46660# a_1057_46660# 2.36e-20
C6564 a_12891_46348# a_10249_46116# 6.35e-21
C6565 a_11309_47204# a_6755_46942# 0.09972f
C6566 a_n881_46662# a_6682_46660# 3.35e-19
C6567 a_12465_44636# a_15559_46634# 4.15e-21
C6568 a_4883_46098# a_17609_46634# 3.14e-20
C6569 a_13507_46334# a_15227_44166# 0.235687f
C6570 a_20894_47436# a_19692_46634# 4.29e-20
C6571 a_15811_47375# a_14513_46634# 9.55e-20
C6572 a_13717_47436# a_16721_46634# 6.05e-22
C6573 a_12861_44030# a_16388_46812# 0.11634f
C6574 a_9067_47204# a_765_45546# 0.007492f
C6575 a_13487_47204# a_13059_46348# 7.45e-20
C6576 a_n2497_47436# a_n1076_46494# 0.001159f
C6577 a_n815_47178# a_n2293_46098# 5.23e-38
C6578 SMPL_ON_P a_n1853_46287# 8.1e-21
C6579 a_n1741_47186# a_n1991_46122# 1.1e-19
C6580 a_n2267_44484# a_n1917_43396# 2.3e-19
C6581 a_n1917_44484# a_n2267_43396# 5.62e-21
C6582 a_n2433_44484# a_n1352_43396# 3.97e-20
C6583 a_n1761_44111# a_n1899_43946# 0.737653f
C6584 a_n2065_43946# a_n1331_43914# 0.053479f
C6585 a_14815_43914# a_14955_43940# 3.05e-19
C6586 a_n1352_44484# a_n2433_43396# 1.79e-21
C6587 a_18494_42460# a_2982_43646# 8.78e-19
C6588 a_10193_42453# a_13291_42460# 0.050019f
C6589 a_9313_44734# a_15493_43940# 4.02e-19
C6590 a_1307_43914# a_16243_43396# 0.001611f
C6591 a_n1059_45260# a_n901_43156# 0.021049f
C6592 en_comp a_n2157_42858# 0.005749f
C6593 a_n2017_45002# a_n1076_43230# 0.006096f
C6594 a_3065_45002# a_4361_42308# 8.6e-19
C6595 a_n913_45002# a_n1641_43230# 3.71e-20
C6596 a_n4209_37414# VDD 0.817347f
C6597 a_20205_45028# VDD 0.005516f
C6598 a_4958_30871# C9_P_btm 0.209166f
C6599 a_22465_38105# a_22545_38993# 0.253407f
C6600 a_9396_43370# a_4883_46098# 0.172323f
C6601 a_8685_43396# a_10227_46804# 0.227547f
C6602 a_14955_43396# a_12861_44030# 0.024664f
C6603 a_13467_32519# w_11334_34010# 3.26e-19
C6604 a_18443_44721# a_17715_44484# 3.58e-20
C6605 a_8333_44734# a_8199_44636# 0.002302f
C6606 a_18287_44626# a_18189_46348# 1.01e-19
C6607 a_5891_43370# a_8953_45546# 0.321625f
C6608 a_8975_43940# a_10809_44734# 0.169586f
C6609 a_18248_44752# a_17957_46116# 6.35e-20
C6610 a_16405_45348# a_16375_45002# 0.012425f
C6611 a_742_44458# a_n1925_42282# 1.15e-20
C6612 a_n2293_42834# a_n863_45724# 0.107229f
C6613 a_949_44458# a_526_44458# 0.03455f
C6614 a_2779_44458# a_2981_46116# 2e-21
C6615 a_17023_45118# a_13259_45724# 1.58e-19
C6616 a_2304_45348# a_2277_45546# 7.72e-19
C6617 a_11691_44458# a_10586_45546# 1e-20
C6618 a_14401_32519# a_22612_30879# 0.062739f
C6619 a_10053_45546# CLK 0.001305f
C6620 a_10193_42453# DATA[5] 4.15e-19
C6621 a_n4315_30879# a_n3420_39616# 0.03477f
C6622 a_n4064_40160# a_n3565_39590# 0.031111f
C6623 a_7174_31319# a_n4209_39304# 4.73e-21
C6624 a_1606_42308# C7_N_btm 0.00238f
C6625 a_7577_46660# a_3483_46348# 7.22e-22
C6626 a_11735_46660# a_11415_45002# 9.22e-21
C6627 a_15227_44166# a_20623_46660# 0.008959f
C6628 a_14513_46634# a_13059_46348# 0.006934f
C6629 a_14180_46812# a_16388_46812# 1.67e-20
C6630 a_19692_46634# a_20411_46873# 0.215749f
C6631 a_19466_46812# a_20273_46660# 7.76e-20
C6632 a_14976_45028# a_16434_46660# 5.98e-20
C6633 a_n1925_46634# a_n1736_46482# 0.002936f
C6634 a_11309_47204# a_8049_45260# 5.06e-19
C6635 a_9804_47204# a_10044_46482# 9.19e-19
C6636 a_13507_46334# a_21071_46482# 7.31e-19
C6637 a_4883_46098# a_19443_46116# 0.002033f
C6638 a_5257_43370# a_4419_46090# 8.58e-19
C6639 a_11967_42832# a_19268_43646# 4.72e-19
C6640 a_19615_44636# a_15743_43084# 9.04e-21
C6641 a_7542_44172# a_7112_43396# 0.001277f
C6642 a_7845_44172# a_7287_43370# 0.011834f
C6643 a_15493_43940# a_20974_43370# 0.069596f
C6644 a_22959_43948# a_14401_32519# 0.006409f
C6645 a_18326_43940# a_n97_42460# 7.83e-21
C6646 a_3499_42826# a_2982_43646# 0.018486f
C6647 a_375_42282# a_196_42282# 0.165785f
C6648 a_18479_45785# a_19511_42282# 5.07e-20
C6649 a_22223_43948# a_17538_32519# 0.001143f
C6650 a_18681_44484# a_16137_43396# 5.5e-22
C6651 a_11341_43940# a_21845_43940# 4.76e-19
C6652 a_2382_45260# a_6123_31319# 9e-21
C6653 a_5147_45002# a_5755_42308# 1.29e-20
C6654 a_n1059_45260# a_10533_42308# 6.69e-21
C6655 a_n2017_45002# a_10723_42308# 0.003736f
C6656 en_comp a_9803_42558# 4.34e-21
C6657 a_5111_44636# a_5421_42558# 0.003313f
C6658 a_n913_45002# a_10545_42558# 0.001151f
C6659 a_15682_43940# VDD 1.22657f
C6660 a_16333_45814# a_8696_44636# 5.96e-20
C6661 a_15599_45572# a_16020_45572# 0.086708f
C6662 a_15765_45572# a_15861_45028# 9.85e-20
C6663 a_16115_45572# a_16680_45572# 7.99e-20
C6664 a_3175_45822# a_413_45260# 0.011644f
C6665 a_175_44278# a_380_45546# 5.93e-21
C6666 a_1115_44172# a_n863_45724# 0.008873f
C6667 a_2479_44172# a_n2661_45546# 6.41e-21
C6668 a_10867_43940# a_10903_43370# 0.004161f
C6669 a_8292_43218# a_n1613_43370# 0.011565f
C6670 a_18861_43218# a_16327_47482# 0.004178f
C6671 a_961_42354# a_n1151_42308# 2.65e-22
C6672 a_1823_45246# VDD 1.7584f
C6673 a_21613_42308# a_22521_40599# 2.02e-20
C6674 a_1343_38525# VDAC_Ni 0.006713f
C6675 a_n3565_39590# a_n4064_37440# 0.031724f
C6676 a_n4064_39616# a_n3565_37414# 0.029074f
C6677 a_n3420_39616# a_n3420_37440# 0.053603f
C6678 C1_N_btm C7_N_btm 0.128479f
C6679 C2_N_btm C6_N_btm 0.137206f
C6680 C0_dummy_N_btm C9_N_btm 0.111645f
C6681 C0_N_btm C8_N_btm 0.146541f
C6682 C3_N_btm C5_N_btm 0.135528f
C6683 C0_dummy_P_btm C10_N_btm 7.53e-19
C6684 a_3147_46376# a_5066_45546# 5.42e-21
C6685 a_13059_46348# a_n357_42282# 1.98e-19
C6686 a_17583_46090# a_17715_44484# 0.22771f
C6687 a_20935_43940# a_20922_43172# 4.63e-19
C6688 a_n1699_43638# a_n2157_42858# 0.008327f
C6689 a_n2267_43396# a_n1853_43023# 0.003945f
C6690 a_n2433_43396# a_n1423_42826# 1.44e-19
C6691 a_14579_43548# a_14358_43442# 0.142377f
C6692 a_13667_43396# a_14205_43396# 0.076384f
C6693 a_4093_43548# a_743_42282# 4.56e-21
C6694 a_n2129_43609# a_n1991_42858# 2.81e-19
C6695 a_14021_43940# a_14543_43071# 4.97e-20
C6696 a_15493_43940# a_18599_43230# 1.61e-20
C6697 a_11341_43940# a_19164_43230# 1.25e-20
C6698 a_9313_44734# a_5742_30871# 9.25e-19
C6699 a_8685_43396# a_8873_43396# 0.001422f
C6700 a_9145_43396# a_9885_43646# 0.052876f
C6701 a_n4318_40392# a_n3420_39616# 4.98e-21
C6702 a_11453_44696# SINGLE_ENDED 0.001844f
C6703 a_13507_46334# EN_OFFSET_CAL 0.00115f
C6704 a_4883_46098# DATA[4] 2.04e-21
C6705 a_22223_43396# VDD 0.279195f
C6706 a_5907_45546# a_n2661_43922# 2.29e-20
C6707 a_18175_45572# a_11691_44458# 7.13e-20
C6708 a_18479_45785# a_19113_45348# 0.013845f
C6709 a_11787_45002# a_13017_45260# 4.5e-20
C6710 a_4574_45260# a_1423_45028# 1.58e-19
C6711 a_3232_43370# a_1307_43914# 0.14252f
C6712 a_8953_45002# a_9482_43914# 0.010057f
C6713 a_6171_45002# a_16019_45002# 0.01229f
C6714 a_2680_45002# a_2903_45348# 0.011458f
C6715 a_n2293_45010# a_n2293_42834# 0.001084f
C6716 a_n2302_38778# a_n2312_39304# 5.35e-19
C6717 a_6643_43396# a_n443_42852# 9.4e-19
C6718 a_n901_43156# a_n1925_42282# 4.57e-20
C6719 a_15095_43370# a_n357_42282# 0.034944f
C6720 a_22165_42308# a_4185_45028# 6.61e-20
C6721 a_16680_45572# a_5807_45002# 0.006746f
C6722 a_8568_45546# a_4646_46812# 1.23e-19
C6723 a_6598_45938# a_5257_43370# 2.41e-19
C6724 a_2711_45572# a_10150_46912# 1.65e-20
C6725 a_6511_45714# a_7715_46873# 9.45e-19
C6726 a_16115_45572# a_13747_46662# 0.029803f
C6727 a_13485_45572# a_12549_44172# 0.004173f
C6728 a_18341_45572# a_n881_46662# 1.2e-19
C6729 a_3357_43084# a_20894_47436# 0.002793f
C6730 a_2437_43646# a_13507_46334# 0.117533f
C6731 a_n2017_45002# a_16327_47482# 0.209709f
C6732 a_413_45260# a_11459_47204# 4.35e-19
C6733 a_11787_45002# a_2063_45854# 2.33e-20
C6734 a_1423_45028# a_n2497_47436# 1.36987f
C6735 a_3232_43370# a_n443_46116# 0.059286f
C6736 a_6171_45002# a_4791_45118# 0.031317f
C6737 a_7705_45326# a_n1151_42308# 0.042252f
C6738 a_n755_45592# a_2957_45546# 0.044162f
C6739 a_n2661_45546# a_n443_42852# 0.141363f
C6740 a_380_45546# a_n356_45724# 0.088749f
C6741 a_n2956_38216# a_n906_45572# 1.15e-19
C6742 a_8952_43230# a_10083_42826# 6.11e-20
C6743 a_9127_43156# a_10518_42984# 6.11e-20
C6744 a_3626_43646# a_2713_42308# 2.32e-20
C6745 a_2982_43646# a_3318_42354# 9.73e-19
C6746 a_3080_42308# a_4921_42308# 1e-19
C6747 a_15037_43940# a_15051_42282# 2.46e-20
C6748 a_14021_43940# a_19511_42282# 1.9e-21
C6749 a_4905_42826# a_4933_42558# 4.27e-19
C6750 a_1512_43396# a_1606_42308# 9.64e-21
C6751 a_18280_46660# START 1.24e-19
C6752 a_8530_39574# VDAC_P 0.064895f
C6753 a_7754_38470# a_11206_38545# 7.39e-19
C6754 a_5934_30871# VDD 0.431204f
C6755 a_18114_32519# VDAC_N 0.003502f
C6756 a_n1741_47186# a_5129_47502# 0.012935f
C6757 a_n2109_47186# a_6151_47436# 9.88e-20
C6758 a_n971_45724# a_4007_47204# 0.01992f
C6759 a_n785_47204# a_n1151_42308# 0.07743f
C6760 a_2124_47436# a_2063_45854# 0.074695f
C6761 a_n237_47217# a_3785_47178# 1.77e-21
C6762 a_1209_47178# a_2905_45572# 1.33e-19
C6763 a_16019_45002# a_14673_44172# 5.98e-19
C6764 a_8696_44636# a_15493_43396# 4.65e-20
C6765 a_18315_45260# a_18287_44626# 0.005579f
C6766 a_18587_45118# a_18248_44752# 6.46e-20
C6767 a_n2433_44484# a_n1352_44484# 0.102355f
C6768 a_n2267_44484# a_n1917_44484# 0.212549f
C6769 a_n2129_44697# a_n1177_44458# 0.027646f
C6770 a_n2661_44458# a_n452_44636# 0.006933f
C6771 a_11827_44484# a_12883_44458# 0.003401f
C6772 a_n2661_43370# a_6109_44484# 1.34e-19
C6773 a_11691_44458# a_10440_44484# 2.28e-20
C6774 a_13556_45296# a_16241_44484# 1.49e-19
C6775 a_10193_42453# a_11173_43940# 2.8e-20
C6776 a_n1059_45260# a_n984_44318# 0.001489f
C6777 a_413_45260# a_22591_44484# 0.024147f
C6778 a_n967_45348# a_n2065_43946# 0.02253f
C6779 a_n913_45002# a_n809_44244# 0.002076f
C6780 a_n2661_45010# a_1414_42308# 0.059385f
C6781 en_comp a_n1761_44111# 2.29e-21
C6782 a_n2293_45010# a_1115_44172# 0.09282f
C6783 a_n2472_42282# a_n2956_38216# 2.12e-20
C6784 a_n3674_38216# a_n2810_45572# 0.023322f
C6785 a_17364_32525# a_22459_39145# 1.15e-20
C6786 a_14209_32519# a_22521_39511# 8.25e-21
C6787 a_n2661_42834# a_12861_44030# 1.42e-20
C6788 a_6229_45572# a_2324_44458# 3.26e-19
C6789 a_11682_45822# a_10903_43370# 0.071222f
C6790 a_10193_42453# a_10809_44734# 0.02204f
C6791 a_3357_43084# a_20411_46873# 0.157199f
C6792 a_7229_43940# a_3090_45724# 0.054969f
C6793 a_2437_43646# a_20623_46660# 4.3e-20
C6794 a_6194_45824# a_5066_45546# 5.14e-20
C6795 a_18114_32519# a_21588_30879# 0.055884f
C6796 a_5343_44458# a_768_44030# 0.066821f
C6797 a_11691_44458# a_n743_46660# 5.94e-20
C6798 a_n2661_43370# a_4646_46812# 0.028718f
C6799 a_8696_44636# a_3483_46348# 0.06521f
C6800 a_15279_43071# a_15051_42282# 0.006313f
C6801 a_5342_30871# a_14113_42308# 0.203397f
C6802 a_13291_42460# a_n784_42308# 1.58e-20
C6803 a_4190_30871# a_n3420_39072# 0.10848f
C6804 a_5807_45002# a_13747_46662# 0.103485f
C6805 a_12549_44172# a_n2661_46634# 0.024531f
C6806 a_8128_46384# a_n1925_46634# 0.21095f
C6807 a_n881_46662# a_n133_46660# 0.005885f
C6808 a_n1613_43370# a_171_46873# 0.11335f
C6809 a_2266_47243# a_2107_46812# 2.19e-19
C6810 a_9313_45822# a_10150_46912# 3.39e-20
C6811 a_n1435_47204# a_8667_46634# 3.08e-20
C6812 a_6851_47204# a_6969_46634# 1.59e-19
C6813 a_7227_47204# a_6755_46942# 1.17e-19
C6814 a_11031_47542# a_10428_46928# 8.15e-19
C6815 a_6545_47178# a_6999_46987# 3.51e-19
C6816 a_n237_47217# a_3090_45724# 3.45e-19
C6817 a_2063_45854# a_11813_46116# 0.093948f
C6818 a_17517_44484# a_20766_44850# 0.018462f
C6819 a_n2661_42834# a_n2840_43914# 0.014735f
C6820 a_1307_43914# a_4905_42826# 7.98e-19
C6821 a_5883_43914# a_10729_43914# 5.61e-21
C6822 a_18114_32519# a_15493_43940# 0.001192f
C6823 a_11827_44484# a_15037_44260# 4.08e-19
C6824 a_3232_43370# a_9396_43370# 5.79e-19
C6825 a_n1059_45260# a_9885_43646# 7.13e-20
C6826 a_n913_45002# a_14955_43396# 6.71e-21
C6827 a_n2017_45002# a_10341_43396# 2.51e-19
C6828 a_1606_42308# C3_P_btm 5.68e-19
C6829 a_n699_43396# a_1823_45246# 0.08003f
C6830 a_16979_44734# a_12741_44636# 0.008336f
C6831 a_18248_44752# a_11415_45002# 3.19e-20
C6832 a_19328_44172# a_19321_45002# 1.77e-19
C6833 a_3600_43914# a_3877_44458# 0.001072f
C6834 a_10949_43914# a_n2293_46634# 0.001108f
C6835 a_12429_44172# a_n2661_46634# 1.5e-21
C6836 a_19862_44208# a_13661_43548# 2.53e-20
C6837 a_9801_44260# a_768_44030# 8.82e-19
C6838 a_14180_45002# a_14180_46482# 2.55e-21
C6839 a_2680_45002# a_n2661_45546# 0.004432f
C6840 a_n967_45348# a_n755_45592# 2.3e-19
C6841 a_413_45260# a_n863_45724# 0.140312f
C6842 a_1667_45002# a_n2293_45546# 0.07132f
C6843 a_n467_45028# a_n1099_45572# 0.007609f
C6844 a_16922_45042# a_17957_46116# 2.12e-21
C6845 a_17613_45144# a_17715_44484# 0.012898f
C6846 a_11691_44458# a_11189_46129# 1.61e-19
C6847 a_n2661_44458# a_5164_46348# 0.001579f
C6848 a_6123_31319# a_1239_39587# 1.95e-19
C6849 a_n3674_37592# a_n4334_38304# 7.84e-20
C6850 a_16104_42674# a_4958_30871# 0.029272f
C6851 a_16522_42674# a_16269_42308# 4.61e-19
C6852 a_1606_42308# a_n4064_38528# 1.87e-20
C6853 a_5932_42308# a_n4209_39304# 4.36e-21
C6854 a_11031_47542# VDD 0.214104f
C6855 a_5649_42852# VDAC_P 3.45e-20
C6856 a_13467_32519# a_22469_40625# 1.21e-20
C6857 a_13887_32519# VDAC_N 2.99e-19
C6858 a_n2293_46634# a_376_46348# 2.26e-21
C6859 a_n1925_46634# a_n1641_46494# 0.005997f
C6860 a_n2661_46634# a_1208_46090# 8.96e-21
C6861 a_n2438_43548# a_n1853_46287# 0.001451f
C6862 a_171_46873# a_n2293_46098# 0.001626f
C6863 a_13661_43548# a_4185_45028# 2.36e-21
C6864 a_6755_46942# a_12156_46660# 0.013732f
C6865 a_11735_46660# a_12251_46660# 0.105995f
C6866 a_5167_46660# a_765_45546# 0.003506f
C6867 a_8270_45546# a_3090_45724# 0.046518f
C6868 a_10623_46897# a_10933_46660# 0.013793f
C6869 a_10554_47026# a_10861_46660# 3.69e-19
C6870 a_10249_46116# a_12359_47026# 1.42e-19
C6871 a_11813_46116# a_12469_46902# 2.33e-20
C6872 a_9804_47204# a_9823_46155# 0.063581f
C6873 a_13507_46334# a_22959_46124# 5.09e-19
C6874 a_n1151_42308# a_14371_46494# 2.26e-19
C6875 a_21811_47423# a_6945_45028# 4.87e-19
C6876 a_4883_46098# a_22223_46124# 0.001059f
C6877 a_21496_47436# a_10809_44734# 0.0112f
C6878 a_11453_44696# a_19335_46494# 6.23e-20
C6879 a_12465_44636# a_21137_46414# 5.25e-22
C6880 a_20640_44752# a_2982_43646# 1.2e-20
C6881 a_n1899_43946# a_n2267_43396# 1.93e-19
C6882 a_n2065_43946# a_n1917_43396# 0.003538f
C6883 a_n1761_44111# a_n1699_43638# 0.003713f
C6884 a_10807_43548# a_11173_44260# 0.05223f
C6885 a_14815_43914# a_8685_43396# 3.62e-20
C6886 a_17737_43940# a_15493_43940# 0.037029f
C6887 a_18079_43940# a_11341_43940# 0.00423f
C6888 a_n1331_43914# a_n2129_43609# 3.76e-21
C6889 a_n1549_44318# a_n2433_43396# 3.69e-20
C6890 a_n2661_42834# a_9803_43646# 5.53e-20
C6891 a_n356_44636# a_17499_43370# 2.72e-19
C6892 a_n2267_44484# a_n1853_43023# 7.38e-22
C6893 a_n2661_44458# a_n1641_43230# 2.46e-22
C6894 a_5891_43370# a_10149_43396# 3.71e-19
C6895 a_n2661_43922# a_9145_43396# 3.97e-20
C6896 a_10193_42453# a_18548_42308# 5.7e-19
C6897 a_n2017_45002# a_20356_42852# 5.14e-20
C6898 a_20512_43084# VDD 0.317257f
C6899 a_13249_42308# a_14495_45572# 0.027073f
C6900 a_11322_45546# a_10907_45822# 0.012408f
C6901 a_2711_45572# a_12649_45572# 4.51e-19
C6902 C1_N_btm C3_P_btm 5.17e-19
C6903 C3_N_btm C5_P_btm 1.02e-19
C6904 C2_N_btm C4_P_btm 3.54e-20
C6905 C0_N_btm C2_P_btm 2.79e-20
C6906 a_19164_43230# a_16327_47482# 0.292734f
C6907 a_10807_43548# a_8953_45546# 5.44e-21
C6908 a_9028_43914# a_9290_44172# 0.169653f
C6909 a_22315_44484# a_8049_45260# 2.42e-21
C6910 a_n2661_43922# a_n1099_45572# 2.98e-21
C6911 a_20749_43396# a_19321_45002# 2.22e-19
C6912 a_13887_32519# a_21588_30879# 0.056445f
C6913 a_19862_44208# a_4185_45028# 1.38e-20
C6914 a_12991_46634# a_12839_46116# 2.15e-19
C6915 a_11415_45002# a_2324_44458# 0.097878f
C6916 a_12741_44636# a_14275_46494# 1.03e-20
C6917 a_3483_46348# a_4704_46090# 2.61e-19
C6918 a_22000_46634# a_6945_45028# 2.76e-19
C6919 a_21363_46634# a_10809_44734# 0.012784f
C6920 a_9313_44734# a_22765_42852# 2.97e-19
C6921 a_3626_43646# a_6031_43396# 3.24e-20
C6922 a_2982_43646# a_6197_43396# 7.06e-21
C6923 a_14021_43940# a_21259_43561# 0.021338f
C6924 a_n2661_42282# a_4520_42826# 1.86e-20
C6925 a_n356_44636# a_1576_42282# 0.003861f
C6926 a_5343_44458# a_6123_31319# 0.003724f
C6927 w_11334_34010# VCM 0.001153f
C6928 a_n746_45260# DATA[0] 0.03466f
C6929 a_n971_45724# DATA[1] 0.050116f
C6930 a_2711_45572# a_4223_44672# 1.51e-20
C6931 a_n2293_45010# a_413_45260# 9.42e-22
C6932 a_n1059_45260# a_n467_45028# 0.229142f
C6933 a_n745_45366# a_n659_45366# 0.006584f
C6934 a_3357_43084# a_4558_45348# 2.13e-21
C6935 a_n2956_37592# en_comp 0.013325f
C6936 a_n913_45002# a_n955_45028# 6.28e-19
C6937 a_6123_31319# a_n2956_39768# 5.77e-21
C6938 a_10341_43396# a_526_44458# 0.005028f
C6939 a_n1917_43396# a_n755_45592# 9.06e-20
C6940 a_n1177_43370# a_n357_42282# 7.33e-19
C6941 a_19511_42282# a_13507_46334# 0.004827f
C6942 a_21335_42336# a_18597_46090# 6.48e-21
C6943 a_19237_31679# a_22459_39145# 1.6e-20
C6944 a_17730_32519# a_22521_39511# 1.16e-20
C6945 a_n2293_45546# VDD 2.06545f
C6946 a_16115_45572# a_11599_46634# 8.83e-19
C6947 a_15903_45785# a_15673_47210# 4.56e-21
C6948 a_15861_45028# a_12861_44030# 0.015193f
C6949 a_2437_43646# a_n1741_47186# 4.86702f
C6950 a_10193_42453# a_n881_46662# 6.12e-20
C6951 a_6598_45938# a_5807_45002# 0.002355f
C6952 a_15681_43442# a_15567_42826# 3.35e-19
C6953 a_n2472_42826# a_n1853_43023# 0.00154f
C6954 a_743_42282# a_685_42968# 0.001652f
C6955 a_10341_43396# a_19164_43230# 1.41e-20
C6956 a_n2840_42826# a_n1991_42858# 1.88e-19
C6957 a_n97_42460# a_18861_43218# 0.001021f
C6958 a_16245_42852# VDD 0.205729f
C6959 a_19431_45546# a_19279_43940# 1.77e-21
C6960 a_17613_45144# a_17719_45144# 0.080654f
C6961 a_16922_45042# a_18587_45118# 0.021516f
C6962 a_14537_43396# a_15004_44636# 0.047224f
C6963 a_1423_45028# a_5883_43914# 0.067915f
C6964 a_1307_43914# a_8975_43940# 0.00588f
C6965 a_9049_44484# a_9028_43914# 7.44e-19
C6966 a_2711_45572# a_15493_43940# 0.128282f
C6967 a_n1059_45260# a_n2661_43922# 0.034597f
C6968 a_n913_45002# a_n2661_42834# 0.027216f
C6969 a_3537_45260# a_7640_43914# 0.006345f
C6970 a_n2017_45002# a_n2293_43922# 0.654835f
C6971 a_5111_44636# a_5205_44734# 1.91e-19
C6972 a_413_45260# a_9313_44734# 4.55e-20
C6973 a_22959_42860# a_n357_42282# 2.46e-20
C6974 a_9803_42558# a_4185_45028# 8.71e-20
C6975 a_13527_45546# a_11415_45002# 3.65e-20
C6976 a_11823_42460# a_12741_44636# 0.031865f
C6977 a_7227_45028# a_3483_46348# 0.00331f
C6978 a_5024_45822# a_1823_45246# 6.21e-21
C6979 a_15765_45572# a_13059_46348# 1.96e-19
C6980 a_18175_45572# a_15227_44166# 0.018929f
C6981 a_18596_45572# a_3090_45724# 1.73e-19
C6982 a_17786_45822# a_19466_46812# 9.25e-23
C6983 a_375_42282# a_n743_46660# 8.64e-21
C6984 a_2232_45348# a_n2293_46634# 8.56e-19
C6985 a_3537_45260# a_4651_46660# 4.86e-21
C6986 a_4574_45260# a_4646_46812# 1.08e-20
C6987 a_4558_45348# a_3877_44458# 0.028316f
C6988 a_5907_45546# a_5164_46348# 5.55e-20
C6989 a_2711_45572# a_6419_46155# 0.002668f
C6990 a_5263_45724# a_5204_45822# 0.109078f
C6991 a_18494_42460# a_11453_44696# 5.41e-22
C6992 a_n23_44458# a_n746_45260# 0.046452f
C6993 a_5111_42852# a_5379_42460# 1.62e-19
C6994 a_4190_30871# a_15486_42560# 2.48e-19
C6995 a_4361_42308# a_13575_42558# 0.006929f
C6996 a_16867_43762# a_17124_42282# 8.78e-22
C6997 a_743_42282# a_14113_42308# 0.015227f
C6998 a_13887_32519# a_5742_30871# 0.004679f
C6999 a_19987_42826# a_20256_42852# 0.015204f
C7000 a_21356_42826# a_14097_32519# 2.8e-20
C7001 a_21195_42852# a_22400_42852# 4.89e-20
C7002 a_11387_46482# DATA[5] 5.29e-20
C7003 a_14311_47204# a_13747_46662# 2.25e-21
C7004 a_11599_46634# a_5807_45002# 0.303048f
C7005 a_15507_47210# a_16131_47204# 9.73e-19
C7006 a_18143_47464# a_12549_44172# 0.0015f
C7007 a_10227_46804# a_768_44030# 0.050994f
C7008 a_16241_47178# a_16285_47570# 3.69e-19
C7009 a_15673_47210# a_16697_47582# 2.36e-20
C7010 a_584_46384# a_479_46660# 1.75e-20
C7011 a_n971_45724# a_2864_46660# 1.42e-20
C7012 a_n1151_42308# a_2107_46812# 0.073605f
C7013 a_1431_47204# a_1799_45572# 3.57e-19
C7014 a_1239_47204# a_n2661_46098# 0.004048f
C7015 a_n443_46116# a_n133_46660# 1e-19
C7016 a_n237_47217# a_3699_46634# 1.03e-19
C7017 a_4883_46098# a_n1613_43370# 0.025959f
C7018 a_12861_44030# a_19321_45002# 0.10527f
C7019 a_6575_47204# a_n2661_46634# 6.01e-19
C7020 a_6151_47436# a_n1925_46634# 0.052327f
C7021 a_13717_47436# a_19594_46812# 3.95e-20
C7022 a_n1699_44726# a_n1761_44111# 0.008854f
C7023 a_n2267_44484# a_n1899_43946# 5.37e-19
C7024 a_n1917_44484# a_n2065_43946# 6.49e-19
C7025 a_n2433_44484# a_n1549_44318# 1.09e-19
C7026 a_18248_44752# a_11967_42832# 0.500539f
C7027 a_18287_44626# a_19006_44850# 0.086658f
C7028 a_n2129_44697# a_n1331_43914# 1.13e-20
C7029 a_n2661_44458# a_n809_44244# 8.95e-20
C7030 a_n2661_43370# a_10405_44172# 2.85e-21
C7031 a_7499_43078# a_743_42282# 0.087933f
C7032 a_8696_44636# a_10695_43548# 6.31e-21
C7033 a_18443_44721# a_18588_44850# 0.057222f
C7034 a_484_44484# a_n2661_43922# 6.52e-19
C7035 a_556_44484# a_n2661_42834# 2.49e-19
C7036 a_n913_45002# a_n1352_43396# 0.002153f
C7037 a_n1059_45260# a_n447_43370# 0.018401f
C7038 a_n2017_45002# a_n97_42460# 0.169401f
C7039 a_n967_45348# a_n2129_43609# 0.021282f
C7040 en_comp a_n2267_43396# 0.028399f
C7041 a_n2661_45010# VDD 0.842431f
C7042 a_18079_43940# a_16327_47482# 0.001128f
C7043 a_13483_43940# a_10227_46804# 8.62e-19
C7044 a_14021_43940# a_4915_47217# 4.68e-20
C7045 a_20623_43914# a_12861_44030# 0.033132f
C7046 a_6171_45002# a_6945_45028# 0.032875f
C7047 a_13159_45002# a_2324_44458# 0.00216f
C7048 a_14180_45002# a_13925_46122# 2.26e-20
C7049 a_9482_43914# a_15015_46420# 1.28e-20
C7050 a_14537_43396# a_13759_46122# 1.79e-20
C7051 a_13556_45296# a_14275_46494# 3.84e-21
C7052 a_2437_43646# a_10586_45546# 2.49e-20
C7053 a_22959_45572# a_8049_45260# 0.176374f
C7054 a_8696_44636# a_n357_42282# 4.53e-21
C7055 a_18545_45144# a_17339_46660# 2.2e-19
C7056 a_453_43940# a_768_44030# 0.110708f
C7057 a_15004_44636# a_3090_45724# 0.010872f
C7058 a_5009_45028# a_3483_46348# 0.029292f
C7059 a_16922_45042# a_11415_45002# 0.012903f
C7060 a_n2661_43370# a_n901_46420# 2.09e-20
C7061 a_8515_42308# a_5742_30871# 1.16e-20
C7062 a_9223_42460# a_9293_42558# 0.011552f
C7063 C8_P_btm C4_P_btm 0.145646f
C7064 C9_P_btm C3_P_btm 0.137552f
C7065 C7_P_btm C5_P_btm 0.151416f
C7066 C10_P_btm C2_P_btm 0.327137f
C7067 a_5257_43370# a_7411_46660# 1.2e-20
C7068 a_4651_46660# a_6969_46634# 2.71e-21
C7069 a_12549_44172# a_765_45546# 0.118284f
C7070 a_n743_46660# a_15227_44166# 3.07e-19
C7071 a_4646_46812# a_6682_46987# 8.46e-19
C7072 a_13747_46662# a_14226_46987# 4.64e-19
C7073 a_5807_45002# a_13693_46688# 5.45e-19
C7074 a_22959_47212# a_12741_44636# 3.06e-19
C7075 a_11453_44696# a_22959_46660# 4.6e-19
C7076 SMPL_ON_N a_21076_30879# 0.030428f
C7077 a_4883_46098# a_n2293_46098# 0.009323f
C7078 a_n1435_47204# a_5204_45822# 1.65e-20
C7079 a_6575_47204# a_8199_44636# 1.83e-20
C7080 a_9863_47436# a_8016_46348# 8.34e-20
C7081 a_n2497_47436# a_n1545_46494# 0.001346f
C7082 a_n2661_43922# a_n2840_43370# 3.06e-19
C7083 a_626_44172# a_685_42968# 9.72e-19
C7084 a_22485_44484# a_15493_43940# 0.087012f
C7085 a_8975_43940# a_9396_43370# 1.2e-20
C7086 a_1307_43914# a_2905_42968# 0.003188f
C7087 a_6453_43914# a_6756_44260# 0.001377f
C7088 a_n2661_42834# a_n4318_39304# 0.041301f
C7089 a_7281_43914# a_n2661_42282# 8.78e-20
C7090 a_11827_44484# a_16547_43609# 5.55e-20
C7091 en_comp a_21671_42860# 4.89e-21
C7092 a_n913_45002# a_n2293_42282# 0.028018f
C7093 a_8855_44734# VDD 4.01e-19
C7094 a_n4209_39304# VREF 0.195875f
C7095 a_n3565_39304# VIN_P 0.039159f
C7096 a_n3565_38502# C5_P_btm 0.00105f
C7097 a_n3420_38528# C7_P_btm 7.66e-20
C7098 a_6472_45840# a_7227_45028# 0.208286f
C7099 a_6511_45714# a_6598_45938# 0.06628f
C7100 a_2711_45572# a_3260_45572# 3.63e-19
C7101 a_5663_43940# a_n2293_46098# 0.142661f
C7102 a_1414_42308# a_1138_42852# 4.35e-19
C7103 a_9165_43940# a_8270_45546# 0.063297f
C7104 a_14358_43442# a_5807_45002# 4.13e-19
C7105 a_14579_43548# a_13661_43548# 8.17e-20
C7106 a_5565_43396# a_n2293_46634# 2.79e-20
C7107 a_n2661_44458# a_3316_45546# 0.003189f
C7108 a_18248_44752# a_13259_45724# 0.003522f
C7109 a_16979_44734# a_16375_45002# 4.01e-20
C7110 a_8375_44464# a_8049_45260# 8.15e-22
C7111 a_2779_44458# a_n863_45724# 4.69e-21
C7112 a_n699_43396# a_n2293_45546# 4.61e-21
C7113 a_n2293_43922# a_526_44458# 1.43e-19
C7114 a_n2661_43922# a_n1925_42282# 0.028186f
C7115 a_17517_44484# a_19900_46494# 2.41e-21
C7116 a_11967_42832# a_2324_44458# 0.005512f
C7117 a_17325_44484# a_17715_44484# 1.25e-19
C7118 a_21259_43561# a_13507_46334# 1.05e-20
C7119 a_2905_42968# a_n443_46116# 2.28e-19
C7120 a_19963_31679# a_22609_37990# 8.31e-21
C7121 a_20447_31679# a_22609_38406# 4.44e-21
C7122 a_1736_39043# a_2684_37794# 0.193802f
C7123 comp_n a_1177_38525# 0.003093f
C7124 a_n4209_38502# a_n4064_38528# 0.265711f
C7125 a_n3565_38502# a_n3420_38528# 0.278952f
C7126 a_n4064_39072# a_n3565_38216# 0.030681f
C7127 a_5732_46660# VDD 0.277366f
C7128 a_4958_30871# C0_N_btm 9.29e-20
C7129 a_765_45546# a_1208_46090# 0.134766f
C7130 a_20719_46660# a_20202_43084# 4.3e-21
C7131 a_12891_46348# a_n443_42852# 7.66e-20
C7132 a_n2661_46634# a_n2661_45546# 5.96e-19
C7133 a_n2840_46634# a_n2956_38216# 0.001369f
C7134 a_3090_45724# a_13759_46122# 5.3e-22
C7135 a_15009_46634# a_13925_46122# 1.53e-19
C7136 a_15368_46634# a_12594_46348# 1.41e-21
C7137 a_1606_42308# a_7754_40130# 0.001975f
C7138 a_n2065_43946# a_n1853_43023# 2.64e-21
C7139 a_n1761_44111# a_n2157_42858# 2.98e-19
C7140 a_18079_43940# a_10341_43396# 3.24e-20
C7141 a_n2267_43396# a_n1699_43638# 0.179796f
C7142 a_n2129_43609# a_n1917_43396# 0.036131f
C7143 a_n2433_43396# a_n1177_43370# 0.043475f
C7144 a_n4318_39304# a_n1352_43396# 4.15e-20
C7145 a_15493_43396# a_14205_43396# 5.22e-20
C7146 a_1307_43914# a_15803_42450# 7.31e-22
C7147 a_3537_45260# a_7174_31319# 4.88e-21
C7148 a_n2810_45028# a_n4209_39590# 0.021994f
C7149 a_n2956_37592# a_n2216_40160# 1.2e-19
C7150 a_21381_43940# VDD 0.344882f
C7151 a_10193_42453# a_1307_43914# 0.054328f
C7152 a_8162_45546# a_1423_45028# 5.61e-21
C7153 a_13904_45546# a_13017_45260# 1.12e-19
C7154 a_11823_42460# a_13556_45296# 0.001625f
C7155 a_5907_45546# a_5837_45028# 9.32e-20
C7156 a_13163_45724# a_13348_45260# 8.77e-21
C7157 a_2711_45572# a_n2293_42834# 0.002511f
C7158 a_18175_45572# a_2437_43646# 1.98e-21
C7159 a_11682_45822# a_3232_43370# 1.34e-19
C7160 a_19256_45572# a_19365_45572# 0.007416f
C7161 a_19431_45546# a_19610_45572# 0.007399f
C7162 a_8685_43396# a_8016_46348# 7.84e-20
C7163 a_n97_42460# a_526_44458# 0.277959f
C7164 a_16795_42852# a_6755_46942# 1.85e-20
C7165 a_5755_42852# a_3090_45724# 8.56e-21
C7166 a_14579_43548# a_4185_45028# 3.54e-21
C7167 a_10334_44484# CLK 0.012484f
C7168 a_n914_46116# VDD 7.75e-19
C7169 a_7499_43078# a_6151_47436# 1.49e-19
C7170 a_7230_45938# a_6851_47204# 4.87e-21
C7171 a_10180_45724# a_4915_47217# 1.08e-20
C7172 a_8746_45002# a_4791_45118# 0.001033f
C7173 a_167_45260# a_n23_45546# 0.001656f
C7174 a_3147_46376# a_3218_45724# 0.0111f
C7175 a_805_46414# a_n443_42852# 0.003153f
C7176 a_2324_44458# a_13259_45724# 0.068761f
C7177 a_4419_46090# a_n755_45592# 0.0037f
C7178 a_20269_44172# a_20256_43172# 5.7e-20
C7179 a_5013_44260# a_4921_42308# 7.51e-21
C7180 a_15781_43660# a_743_42282# 1.91e-20
C7181 a_16409_43396# a_16823_43084# 0.020816f
C7182 a_10341_43396# a_14209_32519# 0.006519f
C7183 a_n97_42460# a_19164_43230# 0.005382f
C7184 a_3626_43646# a_10796_42968# 8.42e-20
C7185 a_2982_43646# a_10922_42852# 4.62e-20
C7186 a_n2661_42282# a_564_42282# 2.77e-19
C7187 a_12281_43396# a_5649_42852# 1.3e-19
C7188 a_16759_43396# a_16855_43396# 0.013793f
C7189 a_16977_43638# a_17021_43396# 3.69e-19
C7190 a_11967_42832# a_16522_42674# 5.62e-19
C7191 a_14021_43940# a_13291_42460# 3.77e-20
C7192 a_383_46660# DATA[0] 2.11e-19
C7193 a_18249_42858# VDD 0.250132f
C7194 a_20447_31679# a_22521_40599# 2.27e-20
C7195 a_n2956_37592# a_n2216_37690# 0.001674f
C7196 a_10193_42453# a_18579_44172# 0.12582f
C7197 a_n913_45002# a_n1352_44484# 0.003041f
C7198 a_n1059_45260# a_n452_44636# 0.010366f
C7199 a_n745_45366# a_n1177_44458# 1.89e-21
C7200 a_6171_45002# a_11827_44484# 0.09294f
C7201 a_413_45260# a_18114_32519# 0.053981f
C7202 a_n2661_45010# a_n699_43396# 3.08e-20
C7203 a_n2017_45002# a_742_44458# 2.47e-19
C7204 en_comp a_n2267_44484# 0.029536f
C7205 a_n967_45348# a_n2129_44697# 0.017689f
C7206 a_n955_45028# a_n2661_44458# 2.09e-19
C7207 a_15486_42560# a_15227_44166# 7.01e-19
C7208 a_n1991_42858# a_n357_42282# 8.06e-19
C7209 a_n13_43084# a_n863_45724# 0.041588f
C7210 a_4361_42308# a_n443_42852# 0.016253f
C7211 a_n1853_43023# a_n755_45592# 0.002072f
C7212 a_3935_43218# a_526_44458# 6.08e-19
C7213 a_17538_32519# a_22521_39511# 1.06e-20
C7214 a_13777_45326# a_11453_44696# 0.004241f
C7215 a_n2661_43370# a_6545_47178# 3.03e-20
C7216 a_14309_45028# a_n1151_42308# 2.59e-21
C7217 a_3232_43370# a_n1613_43370# 0.091534f
C7218 a_5691_45260# a_n881_46662# 1.46e-19
C7219 a_2437_43646# a_n743_46660# 0.031693f
C7220 a_2274_45254# a_768_44030# 0.001893f
C7221 a_2711_45572# a_14226_46660# 3.51e-22
C7222 a_8697_45822# a_8270_45546# 0.001837f
C7223 a_13163_45724# a_12991_46634# 3.39e-20
C7224 a_12791_45546# a_12816_46660# 3.25e-20
C7225 a_9290_44172# CLK 0.151406f
C7226 a_11133_46155# DATA[5] 2.67e-20
C7227 a_21671_42860# a_22165_42308# 0.009789f
C7228 a_21195_42852# a_22223_42860# 1.88e-19
C7229 a_3626_43646# a_4958_30871# 0.087921f
C7230 a_2982_43646# a_17531_42308# 1.21e-19
C7231 a_13887_32519# a_22765_42852# 8.08e-19
C7232 a_21125_42558# VDD 0.004371f
C7233 a_n2109_47186# a_5159_47243# 0.00107f
C7234 a_n1741_47186# a_7989_47542# 4.61e-19
C7235 a_4915_47217# a_13507_46334# 0.032373f
C7236 a_14311_47204# a_11599_46634# 4.05e-22
C7237 a_584_46384# a_2266_47570# 9.67e-19
C7238 a_13717_47436# a_15673_47210# 1.97e-19
C7239 a_12861_44030# a_15811_47375# 0.144648f
C7240 a_n1151_42308# a_11453_44696# 2.35e-21
C7241 a_4791_45118# a_4883_46098# 0.135093f
C7242 a_8746_45002# a_8791_43396# 6.27e-21
C7243 a_16922_45042# a_11967_42832# 0.019919f
C7244 a_21005_45260# a_17517_44484# 5.11e-20
C7245 a_18287_44626# a_18374_44850# 0.053385f
C7246 a_18248_44752# a_18989_43940# 0.207562f
C7247 a_8103_44636# a_8375_44464# 0.13675f
C7248 a_6298_44484# a_5891_43370# 1.52e-21
C7249 a_11827_44484# a_14673_44172# 0.150125f
C7250 a_1307_43914# a_5495_43940# 0.024105f
C7251 a_5883_43914# a_6109_44484# 0.078113f
C7252 a_8701_44490# a_7640_43914# 2.97e-19
C7253 a_n2661_44458# a_n2661_42834# 0.008313f
C7254 a_1423_45028# a_2889_44172# 4.49e-19
C7255 a_n4318_40392# a_n2661_43922# 3.97e-19
C7256 a_5111_44636# a_8333_44056# 0.280148f
C7257 a_16522_42674# a_13259_45724# 9.98e-20
C7258 a_n3565_39304# a_n2956_38680# 0.068534f
C7259 a_n3690_39392# a_n2956_39304# 0.016795f
C7260 a_6761_42308# a_n443_42852# 0.00173f
C7261 a_n37_45144# a_167_45260# 0.277898f
C7262 a_3232_43370# a_n2293_46098# 0.054403f
C7263 a_15433_44458# a_12549_44172# 4.8e-20
C7264 a_7640_43914# a_n2293_46634# 7.73e-20
C7265 a_5883_43914# a_4646_46812# 0.019308f
C7266 a_700_44734# a_n2438_43548# 9.12e-20
C7267 a_327_44734# a_1823_45246# 6.91e-21
C7268 a_13527_45546# a_13259_45724# 0.00477f
C7269 a_18909_45814# a_6945_45028# 2.55e-22
C7270 a_18479_45785# a_10809_44734# 1.4e-21
C7271 a_3357_43084# a_9823_46155# 3.52e-21
C7272 a_3422_30871# a_18597_46090# 0.030159f
C7273 a_14635_42282# a_15486_42560# 0.002155f
C7274 a_2123_42473# a_2351_42308# 0.084895f
C7275 a_5807_45002# a_7411_46660# 0.006898f
C7276 a_n2661_46634# a_5385_46902# 0.007092f
C7277 a_2107_46812# a_3177_46902# 0.001642f
C7278 a_491_47026# a_n2661_46098# 6.63e-19
C7279 a_n1925_46634# a_3221_46660# 6.56e-19
C7280 a_11309_47204# a_10249_46116# 0.033926f
C7281 a_n881_46662# a_8035_47026# 0.003736f
C7282 a_n1613_43370# a_6682_46660# 7.54e-19
C7283 a_12465_44636# a_15368_46634# 7.1e-20
C7284 a_14401_32519# VDAC_N 2.6e-19
C7285 a_13507_46334# a_18834_46812# 0.004721f
C7286 a_4883_46098# a_16292_46812# 1.69e-20
C7287 a_21177_47436# a_15227_44166# 9.06e-22
C7288 a_15811_47375# a_14180_46812# 2.14e-19
C7289 a_19787_47423# a_19692_46634# 5.22e-20
C7290 a_10227_46804# a_10933_46660# 0.00489f
C7291 a_n1741_47186# a_n1853_46287# 1.65e-19
C7292 a_12861_44030# a_13059_46348# 0.504219f
C7293 a_6575_47204# a_765_45546# 0.061901f
C7294 a_13717_47436# a_16388_46812# 4.02e-20
C7295 a_n2267_44484# a_n1699_43638# 6.29e-20
C7296 a_n2065_43946# a_n1899_43946# 0.614122f
C7297 a_5891_43370# a_10555_44260# 0.015358f
C7298 a_18184_42460# a_2982_43646# 0.020575f
C7299 a_1307_43914# a_16137_43396# 4.75e-21
C7300 a_n2293_45010# a_n13_43084# 3.54e-20
C7301 en_comp a_n2472_42826# 0.019667f
C7302 a_n2017_45002# a_n901_43156# 0.005917f
C7303 a_n913_45002# a_n1423_42826# 2.51e-19
C7304 a_n1059_45260# a_n1641_43230# 1.74e-19
C7305 a_2437_43646# a_1847_42826# 1.57e-20
C7306 a_8530_39574# VDD 0.346613f
C7307 a_19929_45028# VDD 0.005632f
C7308 a_4958_30871# C10_P_btm 6.95e-19
C7309 a_22465_38105# a_22521_39511# 0.902378f
C7310 a_8791_43396# a_4883_46098# 0.001239f
C7311 a_15095_43370# a_12861_44030# 6.6e-19
C7312 a_8238_44734# a_8199_44636# 0.003158f
C7313 a_18287_44626# a_17715_44484# 6.13e-20
C7314 a_18248_44752# a_18189_46348# 0.002127f
C7315 a_10057_43914# a_10809_44734# 0.060542f
C7316 a_5891_43370# a_5937_45572# 5.83e-19
C7317 a_2304_45348# a_1609_45822# 0.002594f
C7318 a_16321_45348# a_16375_45002# 0.009082f
C7319 a_742_44458# a_526_44458# 0.54618f
C7320 a_16922_45042# a_13259_45724# 0.401687f
C7321 a_n2661_44458# a_5066_45546# 8.22e-20
C7322 a_14401_32519# a_21588_30879# 0.058775f
C7323 a_7845_44172# a_3090_45724# 0.001391f
C7324 a_15367_44484# a_12741_44636# 5.35e-20
C7325 a_9049_44484# CLK 7.29e-22
C7326 a_11823_42460# RST_Z 1.21e-19
C7327 a_n2302_40160# a_n4209_39590# 9.15e-19
C7328 a_n4064_40160# a_n4334_39616# 0.014656f
C7329 a_7174_31319# a_1343_38525# 2.49e-19
C7330 a_15928_47570# VDD 0.08228f
C7331 a_1606_42308# C6_N_btm 2.33e-19
C7332 a_17701_42308# CAL_N 8.77e-20
C7333 a_5257_43370# a_4185_45028# 9.55e-20
C7334 a_7715_46873# a_3483_46348# 2.08e-20
C7335 a_19692_46634# a_20107_46660# 0.126737f
C7336 a_19466_46812# a_20411_46873# 0.001378f
C7337 a_15227_44166# a_20841_46902# 1.43e-19
C7338 a_14180_46812# a_13059_46348# 0.074456f
C7339 a_19333_46634# a_20273_46660# 1.31e-19
C7340 a_768_44030# a_8034_45724# 4.91e-21
C7341 a_n2312_38680# a_n1736_46482# 1.05e-19
C7342 a_9804_47204# a_9823_46482# 0.006171f
C7343 a_5275_47026# a_5497_46414# 7.81e-20
C7344 a_6540_46812# a_6419_46155# 7.76e-19
C7345 a_13507_46334# a_20850_46482# 9.11e-19
C7346 a_4883_46098# a_20254_46482# 1.42e-19
C7347 a_11967_42832# a_15743_43084# 0.180938f
C7348 a_7281_43914# a_7112_43396# 0.001258f
C7349 a_7542_44172# a_7287_43370# 0.003428f
C7350 a_18079_43940# a_n97_42460# 3.05e-20
C7351 a_15493_43940# a_14401_32519# 0.052433f
C7352 a_22223_43948# a_20974_43370# 7.69e-19
C7353 a_1307_43914# a_n784_42308# 2.99e-19
C7354 a_n356_44636# a_5755_42852# 5.65e-21
C7355 a_13076_44458# a_12545_42858# 1.33e-20
C7356 a_n2661_42282# a_n1557_42282# 4.93e-19
C7357 a_375_42282# a_n473_42460# 8.64e-19
C7358 a_11341_43940# a_17538_32519# 4.23e-19
C7359 a_18579_44172# a_16137_43396# 9.57e-20
C7360 a_3537_45260# a_5932_42308# 0.008724f
C7361 a_n2017_45002# a_10533_42308# 0.003333f
C7362 en_comp a_9223_42460# 4.34e-21
C7363 a_n913_45002# a_9885_42558# 0.001674f
C7364 a_14955_43940# VDD 0.253201f
C7365 a_15903_45785# a_15861_45028# 0.232345f
C7366 a_15765_45572# a_8696_44636# 6.07e-19
C7367 a_15599_45572# a_17478_45572# 1.88e-20
C7368 a_16333_45814# a_16680_45572# 0.051162f
C7369 a_10053_45546# a_2437_43646# 8.54e-21
C7370 a_2711_45572# a_413_45260# 0.022324f
C7371 a_4905_42826# a_n2293_46098# 0.004f
C7372 a_16759_43396# a_3090_45724# 7.41e-22
C7373 a_n809_44244# a_n1099_45572# 2.33e-20
C7374 a_644_44056# a_n863_45724# 6.33e-20
C7375 a_n1899_43946# a_n755_45592# 3.13e-19
C7376 a_13565_43940# a_9290_44172# 1.77e-20
C7377 a_15597_42852# a_10227_46804# 6.37e-19
C7378 a_n784_42308# a_n443_46116# 2.29e-21
C7379 a_19721_31679# a_22521_39511# 2.63e-20
C7380 a_1138_42852# VDD 0.397518f
C7381 C0_N_btm C7_N_btm 0.140846f
C7382 C0_dummy_N_btm C8_N_btm 0.234177f
C7383 C1_N_btm C6_N_btm 0.127656f
C7384 C3_N_btm C4_N_btm 9.61674f
C7385 C2_N_btm C5_N_btm 0.13795f
C7386 C0_dummy_P_btm C9_N_btm 4.11e-19
C7387 C0_P_btm C10_N_btm 8.52e-19
C7388 a_21613_42308# CAL_N 1.44e-19
C7389 a_765_45546# a_n2661_45546# 0.006374f
C7390 a_5164_46348# a_n1925_42282# 3.73e-20
C7391 a_5204_45822# a_526_44458# 0.001107f
C7392 a_10903_43370# a_6945_45028# 1.05e-19
C7393 a_15682_46116# a_17715_44484# 0.003258f
C7394 a_1736_39587# a_3754_38470# 0.002438f
C7395 a_n4209_39590# a_n2302_37690# 2.4e-19
C7396 a_n3565_39590# a_n2946_37690# 1.92e-19
C7397 a_n4064_39616# a_n4334_37440# 8.04e-19
C7398 a_n4064_40160# a_n3607_37440# 5.58e-20
C7399 a_n2433_43396# a_n1991_42858# 6.51e-19
C7400 a_n2267_43396# a_n2157_42858# 6.7e-20
C7401 a_13667_43396# a_14358_43442# 0.001448f
C7402 a_9145_43396# a_14955_43396# 0.06858f
C7403 a_n2129_43609# a_n1853_43023# 1.06e-19
C7404 a_11341_43940# a_19339_43156# 1.47e-20
C7405 a_9313_44734# a_11323_42473# 5.36e-20
C7406 a_14539_43914# a_17531_42308# 5.33e-20
C7407 a_8685_43396# a_12281_43396# 0.038443f
C7408 a_11453_44696# START 8.37e-19
C7409 a_22959_47212# RST_Z 0.001482f
C7410 a_4883_46098# DATA[3] 2.04e-21
C7411 a_5649_42852# VDD 0.438443f
C7412 a_20273_45572# a_16922_45042# 4.48e-20
C7413 a_5907_45546# a_n2661_42834# 1.65e-20
C7414 a_18175_45572# a_19113_45348# 3.29e-19
C7415 a_11787_45002# a_11963_45334# 0.185422f
C7416 a_16147_45260# a_11691_44458# 7.44e-20
C7417 a_11682_45822# a_8975_43940# 1.53e-20
C7418 a_3537_45260# a_1423_45028# 0.046355f
C7419 a_5691_45260# a_1307_43914# 1.36e-19
C7420 a_6171_45002# a_15595_45028# 0.012742f
C7421 a_2680_45002# a_2809_45348# 0.010132f
C7422 a_3357_43084# a_n2661_43370# 0.030835f
C7423 a_5534_30871# a_9290_44172# 0.472376f
C7424 a_12895_43230# a_10903_43370# 0.011631f
C7425 a_n4064_38528# a_n2312_39304# 1.13e-20
C7426 a_15743_43084# a_13259_45724# 0.021493f
C7427 a_n1641_43230# a_n1925_42282# 1.11e-20
C7428 a_14205_43396# a_n357_42282# 6.12e-20
C7429 a_21671_42860# a_4185_45028# 2.44e-20
C7430 a_16333_45814# a_13747_46662# 0.018523f
C7431 a_16855_45546# a_5807_45002# 7.38e-19
C7432 a_8162_45546# a_4646_46812# 8.55e-19
C7433 a_6667_45809# a_5257_43370# 5.18e-20
C7434 a_2711_45572# a_9863_46634# 4.34e-20
C7435 a_16115_45572# a_13661_43548# 3.92e-20
C7436 a_13385_45572# a_12549_44172# 0.001759f
C7437 a_13485_45572# a_12891_46348# 4.18e-19
C7438 a_18479_45785# a_n881_46662# 9.48e-20
C7439 a_2437_43646# a_21177_47436# 0.014824f
C7440 a_21513_45002# a_13507_46334# 5.14e-19
C7441 a_3357_43084# a_19787_47423# 0.001723f
C7442 a_413_45260# a_9313_45822# 2.11e-19
C7443 a_10951_45334# a_2063_45854# 0.016425f
C7444 a_3232_43370# a_4791_45118# 0.268929f
C7445 a_6709_45028# a_n1151_42308# 0.286957f
C7446 a_n755_45592# a_1848_45724# 0.030306f
C7447 a_n863_45724# a_n23_45546# 4.47e-19
C7448 a_n452_45724# a_n356_45724# 0.318161f
C7449 a_n2661_45546# a_509_45822# 4.99e-19
C7450 a_n2956_38216# a_n1013_45572# 2.26e-19
C7451 a_9127_43156# a_10083_42826# 0.011187f
C7452 a_2982_43646# a_2903_42308# 4.44e-21
C7453 a_14401_32519# a_5742_30871# 0.005978f
C7454 a_4905_42826# a_3905_42558# 3.25e-20
C7455 a_20820_30879# a_21589_35634# 5.09e-20
C7456 a_7754_38470# VDAC_P 0.063714f
C7457 a_8530_39574# a_8912_37509# 0.426772f
C7458 a_n4064_37440# a_n3607_37440# 7.1e-19
C7459 a_7963_42308# VDD 0.266057f
C7460 a_n1741_47186# a_4915_47217# 0.128899f
C7461 a_n2109_47186# a_5815_47464# 0.00257f
C7462 a_n971_45724# a_3815_47204# 0.04068f
C7463 a_n23_47502# a_n1151_42308# 0.005195f
C7464 a_2124_47436# a_584_46384# 0.220021f
C7465 a_1209_47178# a_2952_47436# 4.55e-19
C7466 a_1431_47204# a_2063_45854# 1.97e-19
C7467 a_15595_45028# a_14673_44172# 2.84e-20
C7468 a_18315_45260# a_18248_44752# 3.25e-19
C7469 a_n2661_44458# a_n1352_44484# 0.00782f
C7470 a_16922_45042# a_18989_43940# 3.37e-19
C7471 a_n2267_44484# a_n1699_44726# 0.172319f
C7472 a_n2129_44697# a_n1917_44484# 0.030172f
C7473 a_n2433_44484# a_n1177_44458# 0.043567f
C7474 a_11691_44458# a_10334_44484# 2.3e-20
C7475 a_11827_44484# a_12607_44458# 0.023193f
C7476 a_13556_45296# a_15367_44484# 0.003919f
C7477 a_14537_43396# a_17517_44484# 6.26e-21
C7478 a_413_45260# a_22485_44484# 6.37e-21
C7479 a_n1059_45260# a_n809_44244# 0.021842f
C7480 a_n2661_45010# a_1467_44172# 0.001683f
C7481 en_comp a_n2065_43946# 2.47e-19
C7482 a_n2017_45002# a_n984_44318# 3.14e-21
C7483 a_n2293_45010# a_644_44056# 0.014621f
C7484 a_3357_43084# a_2998_44172# 0.119142f
C7485 a_n2104_42282# a_n2810_45572# 2.3e-20
C7486 a_1606_42308# a_13259_45724# 3.55e-20
C7487 a_n3674_38680# a_n2956_38216# 0.022975f
C7488 a_22400_42852# a_n357_42282# 1.12e-19
C7489 COMP_P a_20692_30879# 6.17e-20
C7490 a_3422_30871# w_11334_34010# 1.91172f
C7491 a_15143_45578# a_2324_44458# 0.002313f
C7492 a_11682_45822# a_11387_46155# 2.23e-19
C7493 a_11136_45572# a_8199_44636# 0.001393f
C7494 a_10180_45724# a_10809_44734# 0.007361f
C7495 a_11280_45822# a_10903_43370# 6.44e-19
C7496 a_8975_43940# a_n1613_43370# 4.75e-21
C7497 a_7276_45260# a_3090_45724# 8.07e-21
C7498 a_n913_45002# a_13059_46348# 2.23e-19
C7499 a_3357_43084# a_20107_46660# 0.025828f
C7500 a_2437_43646# a_20841_46902# 1.33e-20
C7501 a_6171_45002# a_15559_46634# 3.5e-22
C7502 a_2711_45572# a_5527_46155# 1.62e-19
C7503 a_3733_45822# a_526_44458# 3.36e-19
C7504 a_5907_45546# a_5066_45546# 9e-19
C7505 a_4743_44484# a_768_44030# 0.002819f
C7506 a_11963_45334# a_11813_46116# 2.51e-19
C7507 a_n2661_43370# a_3877_44458# 0.038641f
C7508 a_17668_45572# a_11415_45002# 0.002419f
C7509 a_16789_45572# a_12741_44636# 1.15e-19
C7510 a_5534_30871# a_15051_42282# 2e-19
C7511 a_12891_46348# a_n2661_46634# 1.07e-19
C7512 a_5807_45002# a_13661_43548# 0.062335f
C7513 a_n881_46662# a_n2438_43548# 0.080298f
C7514 a_n1613_43370# a_n133_46660# 0.347805f
C7515 a_n2312_39304# a_n2661_46098# 0.006111f
C7516 a_n1435_47204# a_7927_46660# 2.14e-20
C7517 a_9313_45822# a_9863_46634# 1.77e-19
C7518 a_6851_47204# a_6755_46942# 8.96e-19
C7519 a_6151_47436# a_6999_46987# 0.001316f
C7520 a_2063_45854# a_11735_46660# 8.71e-19
C7521 a_9838_44484# a_9672_43914# 7.43e-19
C7522 a_17517_44484# a_20835_44721# 0.029603f
C7523 a_18114_32519# a_22223_43948# 0.003272f
C7524 a_1307_43914# a_3080_42308# 0.01819f
C7525 a_10193_42453# a_13635_43156# 0.001112f
C7526 a_5883_43914# a_10405_44172# 6.88e-21
C7527 a_n1655_44484# a_n4318_39768# 1.21e-19
C7528 a_11827_44484# a_14761_44260# 1.07e-19
C7529 a_3232_43370# a_8791_43396# 1.36e-20
C7530 a_n1059_45260# a_14955_43396# 4.49e-20
C7531 a_n913_45002# a_15095_43370# 0.00588f
C7532 COMP_P VIN_N 0.001768f
C7533 a_1606_42308# C4_P_btm 3.05e-19
C7534 a_4223_44672# a_1823_45246# 0.008169f
C7535 a_949_44458# a_167_45260# 0.021626f
C7536 a_14539_43914# a_12741_44636# 0.09527f
C7537 a_n699_43396# a_1138_42852# 0.024181f
C7538 a_17517_44484# a_3090_45724# 0.020082f
C7539 a_2998_44172# a_3877_44458# 3.23e-20
C7540 a_15493_43396# a_13747_46662# 8.51e-22
C7541 a_10729_43914# a_n2293_46634# 0.004608f
C7542 a_19478_44306# a_13661_43548# 5.27e-20
C7543 a_9248_44260# a_768_44030# 2.63e-19
C7544 a_13159_45002# a_12839_46116# 4.85e-20
C7545 a_n37_45144# a_n863_45724# 0.056531f
C7546 a_2382_45260# a_n2661_45546# 8.68e-19
C7547 a_n143_45144# a_n452_45724# 3.05e-21
C7548 a_327_44734# a_n2293_45546# 0.027309f
C7549 a_n967_45348# a_n357_42282# 0.003964f
C7550 en_comp a_n755_45592# 1.09e-20
C7551 a_11827_44484# a_10903_43370# 0.021644f
C7552 a_17613_45144# a_17583_46090# 4.26e-20
C7553 a_11691_44458# a_9290_44172# 3.23e-20
C7554 a_16922_45042# a_18189_46348# 0.015824f
C7555 a_3080_42308# a_n443_46116# 3.12e-21
C7556 a_4905_42826# a_4791_45118# 0.516502f
C7557 a_5932_42308# a_1343_38525# 2.86e-19
C7558 a_n3674_37592# a_n4209_38216# 1.31e-19
C7559 a_9863_47436# VDD 0.207794f
C7560 a_4361_42308# CAL_N 0.003501f
C7561 a_13467_32519# a_22521_40599# 1.43e-20
C7562 a_13747_46662# a_3483_46348# 3.96e-19
C7563 a_n2293_46634# a_n1076_46494# 2.06e-20
C7564 a_n1021_46688# a_n1991_46122# 1.13e-19
C7565 a_n2438_43548# a_n2157_46122# 0.270054f
C7566 a_n133_46660# a_n2293_46098# 8.67e-21
C7567 a_n743_46660# a_n1853_46287# 6.94e-19
C7568 a_5807_45002# a_4185_45028# 5.59e-20
C7569 a_n1925_46634# a_n1423_46090# 0.005255f
C7570 a_n2312_38680# a_n1641_46494# 2.29e-20
C7571 a_10249_46116# a_12156_46660# 1.26e-19
C7572 a_11813_46116# a_11901_46660# 0.211542f
C7573 a_11735_46660# a_12469_46902# 0.053479f
C7574 a_5385_46902# a_765_45546# 0.001698f
C7575 a_10623_46897# a_10861_46660# 0.001705f
C7576 a_6755_46942# a_10425_46660# 2.19e-19
C7577 a_768_44030# a_8016_46348# 0.034453f
C7578 a_9804_47204# a_9569_46155# 0.040648f
C7579 a_n881_46662# a_11133_46155# 4.96e-21
C7580 a_13507_46334# a_10809_44734# 0.603934f
C7581 a_4883_46098# a_6945_45028# 0.083863f
C7582 a_4915_47217# a_10586_45546# 2.07e-20
C7583 a_12465_44636# a_20708_46348# 4.4e-21
C7584 a_18989_43940# a_15743_43084# 3.46e-19
C7585 a_n2065_43946# a_n1699_43638# 1.48e-19
C7586 a_n1761_44111# a_n2267_43396# 1.9e-19
C7587 a_n1899_43946# a_n2129_43609# 4.63e-20
C7588 a_n1331_43914# a_n2433_43396# 0.003897f
C7589 a_15682_43940# a_15493_43940# 0.067033f
C7590 a_17973_43940# a_11341_43940# 0.005348f
C7591 a_10807_43548# a_10555_44260# 9.97e-20
C7592 a_n356_44636# a_16759_43396# 3.62e-21
C7593 a_n2129_44697# a_n1853_43023# 6.76e-22
C7594 a_10193_42453# a_18310_42308# 0.004586f
C7595 a_10949_43914# a_11173_44260# 6.19e-19
C7596 a_10729_43914# a_11816_44260# 0.003322f
C7597 a_19478_44306# a_19862_44208# 0.001187f
C7598 a_5891_43370# a_9885_43396# 7.85e-20
C7599 a_n2661_42834# a_9145_43396# 1.09e-19
C7600 a_n1549_44318# a_n4318_39304# 1.68e-19
C7601 a_n2017_45002# a_20256_42852# 4.86e-19
C7602 a_10193_42453# a_11682_45822# 0.032292f
C7603 a_10490_45724# a_10907_45822# 0.229517f
C7604 a_7499_43078# a_8791_45572# 0.004777f
C7605 a_8568_45546# a_9159_45572# 0.011449f
C7606 a_13904_45546# a_14495_45572# 0.092344f
C7607 a_2711_45572# a_12561_45572# 4.68e-19
C7608 C0_N_btm C3_P_btm 3.06e-19
C7609 C3_N_btm C6_P_btm 2.03e-19
C7610 C2_N_btm C5_P_btm 3.54e-20
C7611 C1_N_btm C4_P_btm 8.82e-20
C7612 C0_dummy_N_btm C2_P_btm 2.79e-20
C7613 a_12545_42858# a_12465_44636# 1.55e-20
C7614 a_19339_43156# a_16327_47482# 0.346029f
C7615 a_3422_30871# a_8049_45260# 2.49e-20
C7616 a_5891_43370# a_n443_42852# 0.175668f
C7617 a_n2661_42834# a_n1099_45572# 2.37e-21
C7618 a_n2661_43922# a_380_45546# 1e-20
C7619 a_12978_47026# VDD 7.19e-19
C7620 a_3699_46348# a_4185_45028# 0.001724f
C7621 a_20623_46660# a_10809_44734# 0.008272f
C7622 a_21188_46660# a_6945_45028# 0.004363f
C7623 a_5934_30871# VDAC_N 0.007175f
C7624 a_3483_46348# a_4419_46090# 0.218073f
C7625 a_6123_31319# VDAC_P 0.009598f
C7626 a_22223_43948# a_13887_32519# 4.31e-19
C7627 a_2982_43646# a_6293_42852# 5.06e-20
C7628 a_15493_43940# a_22223_43396# 2.09e-20
C7629 a_n2661_42282# a_3935_42891# 2.51e-22
C7630 a_n356_44636# a_1067_42314# 0.019369f
C7631 a_5883_43914# a_6171_42473# 6.43e-23
C7632 a_4223_44672# a_5934_30871# 1.39e-21
C7633 a_9313_44734# a_20753_42852# 4.13e-19
C7634 a_5343_44458# a_7227_42308# 2.39e-19
C7635 a_14021_43940# a_19177_43646# 8.27e-19
C7636 a_n1741_47186# DATA[5] 0.069294f
C7637 w_1575_34946# VCM 0.001153f
C7638 a_n971_45724# DATA[0] 0.213213f
C7639 a_8685_43396# VDD 0.261626f
C7640 a_3775_45552# a_n2661_44458# 6.23e-21
C7641 a_2711_45572# a_2779_44458# 2.23e-20
C7642 a_8746_45002# a_11827_44484# 1.23e-19
C7643 a_n1059_45260# a_n955_45028# 4.12e-19
C7644 a_n2810_45028# en_comp 4.45e-19
C7645 a_n745_45366# a_n967_45348# 0.010748f
C7646 a_3357_43084# a_4574_45260# 2.55e-21
C7647 a_n2661_45010# a_327_44734# 0.04375f
C7648 a_n2293_45010# a_n37_45144# 7.8e-21
C7649 a_n2017_45002# a_n467_45028# 8.92e-22
C7650 a_18083_42858# a_17339_46660# 0.001069f
C7651 a_5932_42308# a_n2293_46634# 3.78e-20
C7652 a_12563_42308# a_12549_44172# 1.25e-20
C7653 a_104_43370# a_n863_45724# 0.046664f
C7654 a_9885_43646# a_526_44458# 0.008704f
C7655 a_n1699_43638# a_n755_45592# 1.23e-19
C7656 a_n1917_43396# a_n357_42282# 6.93e-20
C7657 a_4361_42308# a_8199_44636# 0.024061f
C7658 a_n3565_38216# SMPL_ON_P 6.6e-19
C7659 a_n2956_38216# VDD 0.484692f
C7660 a_16333_45814# a_11599_46634# 3.08e-19
C7661 a_15903_45785# a_15811_47375# 3.35e-20
C7662 a_8696_44636# a_12861_44030# 0.046746f
C7663 a_6667_45809# a_5807_45002# 2.91e-19
C7664 a_526_44458# a_3503_45724# 0.06484f
C7665 a_1337_46116# a_997_45618# 0.001151f
C7666 a_8049_45260# a_21167_46155# 3.64e-19
C7667 a_20974_43370# a_20753_42852# 2.74e-20
C7668 a_n2472_42826# a_n2157_42858# 0.080495f
C7669 a_n2840_42826# a_n1853_43023# 3.22e-19
C7670 a_10341_43396# a_19339_43156# 9.56e-19
C7671 a_6293_42852# a_5837_42852# 0.001685f
C7672 a_15953_42852# VDD 0.005646f
C7673 a_18479_45785# a_18579_44172# 0.045071f
C7674 a_16922_45042# a_18315_45260# 0.065907f
C7675 a_1423_45028# a_8701_44490# 0.063232f
C7676 a_1307_43914# a_10057_43914# 0.03199f
C7677 a_9482_43914# a_16979_44734# 5.28e-20
C7678 a_13556_45296# a_14539_43914# 0.025347f
C7679 a_7499_43078# a_9028_43914# 5.08e-20
C7680 a_5093_45028# a_n2661_44458# 0.002375f
C7681 a_n2017_45002# a_n2661_43922# 0.034672f
C7682 a_3537_45260# a_6109_44484# 1.75e-19
C7683 a_n1059_45260# a_n2661_42834# 0.029616f
C7684 a_n467_45028# a_n89_44484# 0.003687f
C7685 a_n2109_45247# a_n2293_43922# 7.56e-20
C7686 a_22223_42860# a_n357_42282# 4.11e-19
C7687 a_9223_42460# a_4185_45028# 8.35e-20
C7688 a_5742_30871# a_1823_45246# 4.25e-20
C7689 a_2982_43646# RST_Z 0.015013f
C7690 a_6598_45938# a_3483_46348# 3.25e-21
C7691 a_15903_45785# a_13059_46348# 9.2e-19
C7692 a_18479_45785# a_17609_46634# 4.93e-20
C7693 a_16751_45260# a_n743_46660# 0.028358f
C7694 a_16147_45260# a_15227_44166# 0.282941f
C7695 a_1423_45028# a_n2293_46634# 0.025918f
C7696 a_1307_43914# a_n2438_43548# 0.006717f
C7697 a_19256_45572# a_3090_45724# 7.35e-19
C7698 a_3537_45260# a_4646_46812# 0.361823f
C7699 a_413_45260# a_6540_46812# 1.57e-21
C7700 a_4574_45260# a_3877_44458# 0.010367f
C7701 a_n2661_43370# a_8128_46384# 3.48e-20
C7702 a_5263_45724# a_5164_46348# 0.005959f
C7703 a_2711_45572# a_6165_46155# 9.84e-19
C7704 a_19721_31679# a_16327_47482# 1.56e-20
C7705 a_n356_44636# a_n746_45260# 0.418585f
C7706 a_n23_44458# a_n971_45724# 1.18e-20
C7707 a_8975_43940# a_4791_45118# 2.73e-20
C7708 a_17499_43370# a_18057_42282# 4.45e-19
C7709 a_5111_42852# a_5267_42460# 6.12e-19
C7710 a_13635_43156# a_n784_42308# 1.68e-20
C7711 a_5649_42852# a_11551_42558# 6.94e-20
C7712 a_4361_42308# a_13070_42354# 0.007985f
C7713 a_4190_30871# a_15051_42282# 5.46e-20
C7714 a_17324_43396# a_17531_42308# 2.3e-21
C7715 a_743_42282# a_13657_42558# 0.007754f
C7716 a_21356_42826# a_22400_42852# 3.91e-20
C7717 a_5342_30871# COMP_P 0.027184f
C7718 a_3160_47472# a_2107_46812# 0.041673f
C7719 a_1209_47178# a_n2661_46098# 2.85e-19
C7720 a_n1151_42308# a_948_46660# 0.002412f
C7721 a_n443_46116# a_n2438_43548# 0.070894f
C7722 a_n971_45724# a_3524_46660# 0.016598f
C7723 a_n237_47217# a_2959_46660# 8.83e-21
C7724 a_n2497_47436# a_3877_44458# 0.024435f
C7725 a_13717_47436# a_19321_45002# 1.59e-19
C7726 a_13487_47204# a_13747_46662# 2.35e-19
C7727 a_4915_47217# a_n743_46660# 0.026159f
C7728 a_7903_47542# a_n2661_46634# 1.47e-20
C7729 a_5815_47464# a_n1925_46634# 5.57e-20
C7730 a_13507_46334# a_n881_46662# 0.019152f
C7731 a_14955_47212# a_5807_45002# 2.52e-20
C7732 a_10227_46804# a_12549_44172# 0.360691f
C7733 a_n1699_44726# a_n2065_43946# 7.01e-20
C7734 a_n2267_44484# a_n1761_44111# 1.89e-19
C7735 a_n2433_44484# a_n1331_43914# 0.001693f
C7736 a_17970_44736# a_11967_42832# 0.00733f
C7737 a_18287_44626# a_18588_44850# 9.73e-19
C7738 a_18248_44752# a_19006_44850# 0.056391f
C7739 a_n2129_44697# a_n1899_43946# 2.08e-20
C7740 a_n2661_44458# a_n1549_44318# 1.29e-20
C7741 a_n2661_43370# a_9672_43914# 1.19e-37
C7742 a_8696_44636# a_9803_43646# 5.08e-21
C7743 a_1307_43914# a_14021_43940# 0.017312f
C7744 a_n89_44484# a_n2661_43922# 3.35e-19
C7745 a_484_44484# a_n2661_42834# 4.92e-19
C7746 a_n967_45348# a_n2433_43396# 0.00115f
C7747 en_comp a_n2129_43609# 0.008951f
C7748 a_n913_45002# a_n1177_43370# 0.014185f
C7749 a_n2293_45010# a_104_43370# 2.23e-19
C7750 a_n1059_45260# a_n1352_43396# 3.37e-20
C7751 a_n2661_45010# a_n1809_43762# 9.47e-20
C7752 a_413_45260# a_14401_32519# 5.55e-20
C7753 a_n2840_45002# VDD 0.289706f
C7754 a_17973_43940# a_16327_47482# 0.001972f
C7755 a_15493_43396# a_11599_46634# 2.13e-21
C7756 a_20365_43914# a_12861_44030# 0.044371f
C7757 a_9482_43914# a_14275_46494# 8.66e-21
C7758 a_14180_45002# a_13759_46122# 1.47e-20
C7759 a_13017_45260# a_2324_44458# 0.021259f
C7760 a_5495_43940# a_n1613_43370# 8.26e-21
C7761 a_3232_43370# a_6945_45028# 2.77e-19
C7762 a_n467_45028# a_526_44458# 1.12e-20
C7763 a_19963_31679# a_8049_45260# 0.2062f
C7764 a_17668_45572# a_13259_45724# 0.050071f
C7765 a_20193_45348# a_20411_46873# 0.002202f
C7766 a_18450_45144# a_17339_46660# 3.54e-19
C7767 a_13720_44458# a_3090_45724# 2.05e-21
C7768 a_5708_44484# a_5257_43370# 0.056224f
C7769 a_1414_42308# a_768_44030# 0.072003f
C7770 a_16501_45348# a_11415_45002# 9.97e-19
C7771 a_16922_45042# a_20202_43084# 1.58e-19
C7772 a_n2293_42834# a_1823_45246# 0.031316f
C7773 a_n2661_43370# a_n1641_46494# 2.3e-20
C7774 a_8325_42308# a_9885_42558# 1.55e-21
C7775 a_5934_30871# a_5742_30871# 16.7261f
C7776 a_8685_42308# a_9377_42558# 0.003285f
C7777 a_9223_42460# a_9803_42558# 0.001368f
C7778 C9_P_btm C4_P_btm 0.154834f
C7779 C8_P_btm C5_P_btm 0.145019f
C7780 C7_P_btm C6_P_btm 26.0771f
C7781 C10_P_btm C3_P_btm 0.321945f
C7782 a_12891_46348# a_765_45546# 0.041192f
C7783 a_12549_44172# a_17339_46660# 0.081298f
C7784 a_13747_46662# a_14513_46634# 6.82e-19
C7785 a_4646_46812# a_6969_46634# 0.072545f
C7786 a_4651_46660# a_6755_46942# 5.05e-21
C7787 a_22959_47212# a_20820_30879# 0.004677f
C7788 a_11453_44696# a_12741_44636# 1.02327f
C7789 a_22731_47423# a_21076_30879# 0.001083f
C7790 a_11599_46634# a_3483_46348# 3.49e-19
C7791 a_4915_47217# a_11189_46129# 3.08e-22
C7792 a_6151_47436# a_9823_46155# 0.001307f
C7793 a_n1435_47204# a_5164_46348# 1.08e-20
C7794 a_n2497_47436# a_n1736_46482# 0.005472f
C7795 a_2063_45854# a_2324_44458# 0.028153f
C7796 a_n1151_42308# a_13925_46122# 4.64e-19
C7797 a_n1741_47186# a_10809_44734# 0.332771f
C7798 a_22485_44484# a_22223_43948# 0.016889f
C7799 a_6453_43914# a_n2661_42282# 0.122766f
C7800 a_18579_44172# a_14021_43940# 0.033047f
C7801 a_1307_43914# a_2075_43172# 0.077359f
C7802 a_n2661_42834# a_n2840_43370# 0.026572f
C7803 a_8975_43940# a_8791_43396# 4e-20
C7804 a_11827_44484# a_16243_43396# 1.51e-20
C7805 a_20512_43084# a_15493_43940# 0.021257f
C7806 a_10057_43914# a_9396_43370# 1.26e-19
C7807 a_n1059_45260# a_n2293_42282# 0.033257f
C7808 en_comp a_21195_42852# 4.83e-21
C7809 a_8783_44734# VDD 4.43e-19
C7810 a_n3565_38502# C6_P_btm 1.26e-20
C7811 a_n3565_38216# a_n1532_35090# 1e-19
C7812 a_n4209_38216# EN_VIN_BSTR_P 0.004167f
C7813 a_6472_45840# a_6598_45938# 0.178024f
C7814 a_6511_45714# a_6667_45809# 0.113977f
C7815 a_175_44278# a_167_45260# 5.9e-20
C7816 a_5495_43940# a_n2293_46098# 0.096987f
C7817 a_1467_44172# a_1138_42852# 0.034446f
C7818 a_13667_43396# a_13661_43548# 0.168674f
C7819 a_8487_44056# a_8270_45546# 1.88e-19
C7820 a_4181_43396# a_n2293_46634# 3.92e-20
C7821 a_n2661_43922# a_526_44458# 0.154533f
C7822 a_n2661_44458# a_3218_45724# 3.08e-20
C7823 a_949_44458# a_n863_45724# 0.034335f
C7824 a_7640_43914# a_8049_45260# 0.003041f
C7825 a_14539_43914# a_16375_45002# 3.75e-20
C7826 a_17970_44736# a_13259_45724# 0.011308f
C7827 a_5343_44458# a_n2661_45546# 1.16e-20
C7828 a_n2661_42834# a_n1925_42282# 0.029302f
C7829 a_17517_44484# a_20075_46420# 6e-21
C7830 a_2075_43172# a_n443_46116# 0.002146f
C7831 a_n3565_38502# a_n3690_38528# 0.246863f
C7832 a_1736_39043# a_1177_38525# 1.72e-19
C7833 a_n4334_38528# a_n3420_38528# 0.015595f
C7834 a_n4209_38502# a_n2946_38778# 0.022704f
C7835 a_n4064_39072# a_n4334_38304# 3.17e-19
C7836 a_5907_46634# VDD 0.341121f
C7837 a_4958_30871# C0_dummy_N_btm 1.65e-20
C7838 a_765_45546# a_805_46414# 8.01e-20
C7839 a_n2956_39768# a_n2661_45546# 6.28e-20
C7840 a_14084_46812# a_13925_46122# 9.14e-19
C7841 a_n2065_43946# a_n2157_42858# 6.86e-21
C7842 a_17973_43940# a_10341_43396# 1.83e-20
C7843 a_n2433_43396# a_n1917_43396# 0.108815f
C7844 a_n2129_43609# a_n1699_43638# 0.022218f
C7845 a_2998_44172# a_743_42282# 1.28e-20
C7846 a_1307_43914# a_15764_42576# 8.77e-22
C7847 en_comp a_n2302_40160# 2.07e-19
C7848 a_19741_43940# VDD 0.153579f
C7849 a_13527_45546# a_13017_45260# 9.04e-20
C7850 a_11823_42460# a_9482_43914# 0.033152f
C7851 a_13163_45724# a_13159_45002# 0.010135f
C7852 a_10193_42453# a_16019_45002# 6.67e-19
C7853 a_2711_45572# a_7639_45394# 2.87e-19
C7854 a_10907_45822# a_6171_45002# 0.024408f
C7855 a_8696_44636# a_n913_45002# 2.6e-20
C7856 a_7174_31319# w_11334_34010# 7.7e-19
C7857 a_n784_42308# a_n1613_43370# 0.002725f
C7858 a_20269_44172# a_n357_42282# 1.22e-20
C7859 a_10807_43548# a_n443_42852# 0.173997f
C7860 a_5111_42852# a_3090_45724# 5.57e-21
C7861 a_20256_43172# a_13661_43548# 5.04e-19
C7862 a_15743_43084# a_20202_43084# 0.021267f
C7863 a_14358_43442# a_3483_46348# 1.32e-20
C7864 a_10157_44484# CLK 0.002339f
C7865 a_2711_45572# a_16023_47582# 8.57e-20
C7866 a_10053_45546# a_4915_47217# 3.01e-22
C7867 a_8568_45546# a_6151_47436# 6.1e-21
C7868 a_11962_45724# a_n1151_42308# 8.76e-37
C7869 a_4185_45028# a_n755_45592# 0.024134f
C7870 a_167_45260# a_n356_45724# 9.47e-19
C7871 a_3147_46376# a_2957_45546# 8.73e-20
C7872 a_472_46348# a_n443_42852# 4.66e-19
C7873 a_n1925_42282# a_5066_45546# 3.2e-20
C7874 a_10809_44734# a_10586_45546# 5.07e-19
C7875 a_14840_46494# a_13259_45724# 0.002156f
C7876 a_2324_44458# a_14383_46116# 1.41e-19
C7877 a_5244_44056# a_4921_42308# 1.76e-21
C7878 a_6197_43396# a_7227_42852# 3.42e-20
C7879 a_11967_42832# a_16104_42674# 4.18e-19
C7880 a_10341_43396# a_22591_43396# 0.172197f
C7881 a_n97_42460# a_19339_43156# 0.012502f
C7882 a_2982_43646# a_10991_42826# 1.03e-19
C7883 a_3626_43646# a_10835_43094# 2.04e-20
C7884 a_16547_43609# a_16823_43084# 0.08061f
C7885 a_n2661_42282# a_n3674_37592# 0.12829f
C7886 a_15743_43084# a_16867_43762# 8.49e-19
C7887 a_16977_43638# a_16855_43396# 3.16e-19
C7888 a_16243_43396# a_17433_43396# 2.56e-19
C7889 a_601_46902# DATA[0] 2.35e-19
C7890 a_n743_46660# DATA[5] 5.08e-21
C7891 a_17333_42852# VDD 0.525529f
C7892 a_19963_31679# a_22469_40625# 1.59e-20
C7893 a_n2810_45028# a_n2216_37690# 0.003507f
C7894 a_n2956_37592# a_n2860_37690# 0.001388f
C7895 a_626_44172# a_n2661_43370# 0.008858f
C7896 a_14797_45144# a_15060_45348# 0.010598f
C7897 a_10193_42453# a_18245_44484# 1.51e-19
C7898 a_n1059_45260# a_n1352_44484# 2.66e-19
C7899 a_n913_45002# a_n1177_44458# 0.017911f
C7900 a_n967_45348# a_n2433_44484# 3.53e-20
C7901 en_comp a_n2129_44697# 0.00879f
C7902 a_n2293_45010# a_949_44458# 0.001253f
C7903 a_3232_43370# a_11827_44484# 0.094278f
C7904 a_3357_43084# a_5883_43914# 0.046158f
C7905 a_15051_42282# a_15227_44166# 2.31e-20
C7906 a_n2157_42858# a_n755_45592# 1.64e-22
C7907 a_n1076_43230# a_n863_45724# 1.91e-20
C7908 a_n2293_42282# a_n1925_42282# 0.234055f
C7909 a_n1853_43023# a_n357_42282# 0.04297f
C7910 a_n4318_38680# a_n2956_38216# 0.023204f
C7911 a_3445_43172# a_526_44458# 2.76e-19
C7912 a_14635_42282# a_9290_44172# 3.64e-19
C7913 VDAC_Ni w_1575_34946# 7.89e-19
C7914 a_13556_45296# a_11453_44696# 0.027553f
C7915 a_14797_45144# a_12465_44636# 0.002814f
C7916 a_1307_43914# a_13507_46334# 3.03e-20
C7917 a_n2661_43370# a_6151_47436# 0.003024f
C7918 a_4927_45028# a_n881_46662# 0.001762f
C7919 a_5691_45260# a_n1613_43370# 5.61e-21
C7920 a_8336_45822# a_8270_45546# 0.009698f
C7921 a_11823_42460# a_12816_46660# 1.3e-20
C7922 a_12791_45546# a_12991_46634# 5.89e-20
C7923 a_21195_42852# a_22165_42308# 0.007883f
C7924 a_2982_43646# a_17303_42282# 0.139588f
C7925 a_n4318_39304# a_n4334_39616# 7.95e-19
C7926 a_17364_32525# a_14097_32519# 0.059348f
C7927 a_8605_42826# a_9114_42852# 2.6e-19
C7928 a_3626_43646# a_16269_42308# 0.001405f
C7929 a_10355_46116# CLK 0.002305f
C7930 a_11189_46129# DATA[5] 1.65e-20
C7931 a_n1741_47186# a_n881_46662# 0.179671f
C7932 a_n2109_47186# a_4842_47243# 0.002652f
C7933 SMPL_ON_P a_n1613_43370# 5.27e-21
C7934 a_14311_47204# a_14955_47212# 3.11e-20
C7935 a_2124_47436# a_2266_47570# 0.007833f
C7936 a_13717_47436# a_15811_47375# 1.75e-19
C7937 a_13487_47204# a_11599_46634# 9.96e-21
C7938 a_12861_44030# a_15507_47210# 2.51e-20
C7939 a_4700_47436# a_4883_46098# 1.43e-19
C7940 a_20567_45036# a_17517_44484# 7.16e-20
C7941 a_18287_44626# a_18443_44721# 0.10279f
C7942 a_8103_44636# a_7640_43914# 0.101633f
C7943 a_6298_44484# a_8375_44464# 8.94e-21
C7944 a_18248_44752# a_18374_44850# 0.170059f
C7945 a_1423_45028# a_2675_43914# 4.85e-20
C7946 a_n2840_44458# a_n2661_43922# 0.001534f
C7947 a_1307_43914# a_5013_44260# 0.358053f
C7948 a_5518_44484# a_5891_43370# 2.14e-20
C7949 a_n2661_44458# a_11649_44734# 8.36e-19
C7950 a_17970_44736# a_18989_43940# 1.91e-21
C7951 a_5343_44458# a_8238_44734# 1.98e-21
C7952 a_11827_44484# a_14581_44484# 1.34e-19
C7953 a_5111_44636# a_8018_44260# 4.54e-19
C7954 a_3232_43370# a_6756_44260# 6.17e-21
C7955 a_n3565_39304# a_n2956_39304# 0.307358f
C7956 a_413_45260# a_1823_45246# 0.043122f
C7957 a_n143_45144# a_167_45260# 0.03701f
C7958 a_5708_44484# a_5807_45002# 3.53e-20
C7959 a_6109_44484# a_n2293_46634# 2.18e-19
C7960 a_14815_43914# a_12549_44172# 0.026324f
C7961 a_15060_45348# a_14976_45028# 0.005133f
C7962 a_14112_44734# a_768_44030# 0.004013f
C7963 a_327_44734# a_1138_42852# 1.41e-19
C7964 a_15685_45394# a_3090_45724# 4.27e-20
C7965 a_13163_45724# a_13259_45724# 0.166368f
C7966 a_4099_45572# a_3503_45724# 1.81e-19
C7967 a_4880_45572# a_n2661_45546# 0.003682f
C7968 a_18175_45572# a_10809_44734# 1.39e-20
C7969 a_3357_43084# a_9569_46155# 1.93e-20
C7970 a_18579_44172# a_13507_46334# 2e-20
C7971 a_21398_44850# a_18597_46090# 0.002638f
C7972 a_5013_44260# a_n443_46116# 7.51e-21
C7973 a_5495_43940# a_4791_45118# 8.22e-20
C7974 a_1755_42282# a_2351_42308# 3.31e-19
C7975 a_14635_42282# a_15051_42282# 0.007421f
C7976 a_n2293_42282# a_n4315_30879# 3.44e-21
C7977 a_5807_45002# a_5257_43370# 0.683815f
C7978 a_n2661_46634# a_4817_46660# 0.047477f
C7979 a_1983_46706# a_2443_46660# 2.86e-19
C7980 a_2107_46812# a_2609_46660# 0.003525f
C7981 a_n2293_46634# a_4646_46812# 0.135642f
C7982 a_n133_46660# a_1057_46660# 2.56e-19
C7983 a_288_46660# a_n2661_46098# 2.31e-20
C7984 a_n2438_43548# a_1302_46660# 5.38e-19
C7985 a_n1925_46634# a_3055_46660# 0.001224f
C7986 a_n743_46660# a_2162_46660# 3.68e-19
C7987 a_n881_46662# a_7832_46660# 7.95e-20
C7988 a_12465_44636# a_14976_45028# 4.97e-20
C7989 a_3080_42308# a_3754_39134# 1.67e-20
C7990 a_13507_46334# a_17609_46634# 0.01055f
C7991 a_4883_46098# a_15559_46634# 7.47e-20
C7992 a_20990_47178# a_15227_44166# 4.31e-19
C7993 a_n1741_47186# a_n2157_46122# 2.78e-19
C7994 SMPL_ON_P a_n2293_46098# 7.56e-20
C7995 a_n2497_47436# a_n1641_46494# 0.020605f
C7996 a_n1920_47178# a_n1853_46287# 0.001135f
C7997 a_n2109_47186# a_n1991_46122# 8.21e-21
C7998 a_12861_44030# a_15227_46910# 0.050112f
C7999 a_13717_47436# a_13059_46348# 5.91e-19
C8000 a_7903_47542# a_765_45546# 0.001413f
C8001 a_19787_47423# a_19466_46812# 1.48e-19
C8002 a_10227_46804# a_10861_46660# 0.003218f
C8003 a_19386_47436# a_19692_46634# 2.42e-20
C8004 a_11599_46634# a_14513_46634# 1.15e-20
C8005 a_n2433_44484# a_n1917_43396# 2.93e-20
C8006 a_n2267_44484# a_n2267_43396# 0.001024f
C8007 a_n2065_43946# a_n1761_44111# 0.617556f
C8008 a_n1917_44484# a_n2433_43396# 2.16e-20
C8009 a_9313_44734# a_11341_43940# 1.41e-19
C8010 a_n2293_45010# a_n1076_43230# 3.21e-21
C8011 a_n2017_45002# a_n1641_43230# 0.011397f
C8012 a_n913_45002# a_n1991_42858# 0.024791f
C8013 a_2382_45260# a_4361_42308# 3.26e-20
C8014 a_n1059_45260# a_n1423_42826# 2.7e-19
C8015 en_comp a_n2840_42826# 0.002468f
C8016 a_7754_38470# VDD 0.302129f
C8017 a_18545_45144# VDD 3.69e-20
C8018 a_8147_43396# a_4883_46098# 6.45e-20
C8019 a_14205_43396# a_12861_44030# 6.35e-20
C8020 a_743_42282# a_n2497_47436# 2.68e-22
C8021 a_5891_43370# a_8199_44636# 0.399007f
C8022 a_8375_44464# a_5937_45572# 1.42e-20
C8023 a_10440_44484# a_10809_44734# 0.002452f
C8024 a_18248_44752# a_17715_44484# 5.78e-20
C8025 a_7640_43914# a_8953_45546# 1.62e-20
C8026 a_17970_44736# a_18189_46348# 5.88e-19
C8027 a_n452_44636# a_526_44458# 3.8e-20
C8028 a_1423_45028# a_2277_45546# 9.3e-22
C8029 a_7542_44172# a_3090_45724# 0.137368f
C8030 a_7499_43078# CLK 9.27e-21
C8031 a_n4334_40480# a_n4334_39616# 0.050585f
C8032 a_n4064_40160# a_n4209_39590# 0.059936f
C8033 a_n2302_40160# a_n2216_40160# 0.011479f
C8034 a_n4315_30879# a_n3565_39590# 0.027163f
C8035 a_768_44030# VDD 1.53454f
C8036 a_1606_42308# C5_N_btm 1.89e-19
C8037 a_7411_46660# a_3483_46348# 2.45e-19
C8038 a_14035_46660# a_13059_46348# 0.072321f
C8039 a_15227_44166# a_20273_46660# 2.91e-19
C8040 a_19466_46812# a_20107_46660# 1.31e-20
C8041 a_19692_46634# a_19551_46910# 0.0536f
C8042 a_19333_46634# a_20411_46873# 2.17e-20
C8043 a_14180_46812# a_15227_46910# 3.46e-19
C8044 a_12359_47026# a_765_45546# 3.39e-21
C8045 a_n2312_38680# a_n2956_38680# 6.25577f
C8046 a_n2293_46634# a_n1545_46494# 1.01e-19
C8047 a_n1925_46634# a_n2956_39304# 2.57e-19
C8048 a_9804_47204# a_9241_46436# 4.41e-20
C8049 a_n881_46662# a_10586_45546# 1.46e-20
C8050 a_5275_47026# a_5204_45822# 4.42e-20
C8051 a_n743_46660# a_10809_44734# 0.032324f
C8052 a_11453_44696# a_16375_45002# 0.104273f
C8053 a_4883_46098# a_20009_46494# 1.23e-19
C8054 a_n443_46116# a_603_45572# 0.004683f
C8055 a_7281_43914# a_7287_43370# 0.003639f
C8056 a_11341_43940# a_20974_43370# 0.013722f
C8057 a_22223_43948# a_14401_32519# 0.157135f
C8058 a_17973_43940# a_n97_42460# 1.1e-21
C8059 a_11967_42832# a_18783_43370# 0.001091f
C8060 a_22591_44484# a_10341_43396# 3.21e-19
C8061 a_n356_44636# a_5111_42852# 1.83e-20
C8062 a_15493_43940# a_21381_43940# 0.02116f
C8063 a_375_42282# a_n961_42308# 3.02e-20
C8064 a_2998_44172# a_2813_43396# 2e-19
C8065 a_5111_44636# a_4921_42308# 0.004461f
C8066 a_3537_45260# a_6171_42473# 3.79e-20
C8067 a_3232_43370# a_3581_42558# 7.4e-20
C8068 a_n913_45002# a_9377_42558# 2.17e-19
C8069 a_n2017_45002# a_10545_42558# 9.16e-19
C8070 a_13483_43940# VDD 0.219591f
C8071 a_15599_45572# a_15861_45028# 1.72e-20
C8072 a_15903_45785# a_8696_44636# 1.89e-19
C8073 a_15765_45572# a_16680_45572# 0.118759f
C8074 a_3080_42308# a_n2293_46098# 5.04e-19
C8075 a_9145_43396# a_13059_46348# 0.028786f
C8076 a_21356_42826# a_13747_46662# 1.41e-19
C8077 a_19987_42826# a_19321_45002# 5.73e-20
C8078 a_175_44278# a_n863_45724# 0.113317f
C8079 a_n1549_44318# a_n1099_45572# 2.98e-21
C8080 a_n1761_44111# a_n755_45592# 0.015303f
C8081 a_11257_43940# a_9290_44172# 6.04e-19
C8082 a_7309_43172# a_n1613_43370# 7.87e-19
C8083 a_1755_42282# a_584_46384# 8.38e-21
C8084 a_n784_42308# a_4791_45118# 4.27e-20
C8085 a_5932_42308# w_11334_34010# 9.2e-19
C8086 a_18114_32519# a_22521_39511# 1.28e-20
C8087 a_1176_45822# VDD 0.781481f
C8088 C0_dummy_N_btm C7_N_btm 0.119061f
C8089 C0_N_btm C6_N_btm 0.139059f
C8090 C1_N_btm C5_N_btm 0.127408f
C8091 C2_N_btm C4_N_btm 7.72909f
C8092 C0_dummy_P_btm C8_N_btm 3.42e-19
C8093 C1_P_btm C10_N_btm 9.71e-19
C8094 C0_P_btm C9_N_btm 4.64e-19
C8095 a_21887_42336# CAL_N 8.2e-19
C8096 a_3483_46348# a_4365_46436# 3.61e-19
C8097 a_1823_45246# a_5527_46155# 3.02e-21
C8098 a_17639_46660# a_16375_45002# 8.23e-20
C8099 a_5164_46348# a_526_44458# 2.61e-20
C8100 a_11189_46129# a_10809_44734# 3.89e-20
C8101 a_15682_46116# a_17583_46090# 0.013015f
C8102 a_n2302_38778# a_n2302_37984# 0.052227f
C8103 a_n3565_39590# a_n3420_37440# 0.035128f
C8104 a_n4209_39590# a_n4064_37440# 0.033425f
C8105 a_n4064_39616# a_n4209_37414# 0.028043f
C8106 a_n3420_39616# a_n3565_37414# 0.028804f
C8107 a_n4064_40160# a_n4251_37440# 0.001069f
C8108 a_20623_43914# a_19987_42826# 1.37e-19
C8109 a_n2129_43609# a_n2157_42858# 0.007212f
C8110 a_n2433_43396# a_n1853_43023# 4.61e-19
C8111 a_1568_43370# a_743_42282# 2.22e-19
C8112 a_9145_43396# a_15095_43370# 0.213415f
C8113 a_14021_43940# a_13635_43156# 0.001414f
C8114 a_15493_43940# a_18249_42858# 2.89e-20
C8115 a_11341_43940# a_18599_43230# 3.88e-20
C8116 a_9313_44734# a_10723_42308# 1.32e-20
C8117 a_19237_31679# a_14097_32519# 0.052198f
C8118 a_19862_44208# a_21195_42852# 0.002065f
C8119 a_13667_43396# a_14579_43548# 5.78e-19
C8120 a_11453_44696# RST_Z 0.004685f
C8121 a_13678_32519# VDD 0.454512f
C8122 a_4099_45572# a_n2661_43922# 2.36e-20
C8123 a_18341_45572# a_11827_44484# 6.05e-21
C8124 a_20107_45572# a_16922_45042# 1.06e-19
C8125 a_8696_44636# a_n2661_44458# 1.37553f
C8126 a_6171_45002# a_15415_45028# 0.008633f
C8127 a_4927_45028# a_1307_43914# 8.94e-21
C8128 a_2680_45002# a_2304_45348# 1.96e-19
C8129 a_2274_45254# a_2903_45348# 6.01e-19
C8130 a_n2661_45010# a_n2293_42834# 2.08e-20
C8131 a_14543_43071# a_9290_44172# 0.005728f
C8132 a_13113_42826# a_10903_43370# 0.011891f
C8133 a_5837_43396# a_n443_42852# 2.02e-19
C8134 a_n1423_42826# a_n1925_42282# 1.97e-20
C8135 a_17324_43396# a_16375_45002# 1.24e-20
C8136 a_14358_43442# a_n357_42282# 3e-20
C8137 a_7174_31319# a_n2442_46660# 5.91e-21
C8138 a_21195_42852# a_4185_45028# 2.22e-20
C8139 a_16333_45814# a_13661_43548# 8.09e-19
C8140 a_15765_45572# a_13747_46662# 0.5661f
C8141 a_6511_45714# a_5257_43370# 9.68e-20
C8142 a_2711_45572# a_8492_46660# 8.18e-21
C8143 a_7230_45938# a_4646_46812# 0.005389f
C8144 a_13297_45572# a_12549_44172# 5.89e-19
C8145 a_13385_45572# a_12891_46348# 0.001139f
C8146 a_18175_45572# a_n881_46662# 1.17e-19
C8147 a_2437_43646# a_20990_47178# 0.008979f
C8148 a_3357_43084# a_19386_47436# 4.09e-19
C8149 a_413_45260# a_11031_47542# 1.03e-19
C8150 a_10775_45002# a_2063_45854# 0.012226f
C8151 a_626_44172# a_n2497_47436# 0.249352f
C8152 a_4927_45028# a_n443_46116# 5.42e-19
C8153 a_5691_45260# a_4791_45118# 0.001279f
C8154 a_7229_43940# a_n1151_42308# 0.036511f
C8155 a_n863_45724# a_n356_45724# 0.003189f
C8156 a_n755_45592# a_997_45618# 0.133124f
C8157 a_n2661_45546# a_n906_45572# 6.4e-19
C8158 a_9127_43156# a_8952_43230# 0.234322f
C8159 a_17364_32525# a_22959_42860# 5e-19
C8160 a_2982_43646# a_2713_42308# 1.35e-21
C8161 a_2896_43646# a_2903_42308# 7.11e-21
C8162 a_3080_42308# a_3905_42558# 0.008414f
C8163 a_4905_42826# a_3581_42558# 8.56e-21
C8164 a_20820_30879# a_19864_35138# 1.44e-20
C8165 a_20273_46660# EN_OFFSET_CAL 3.18e-20
C8166 a_3754_38470# a_11206_38545# 0.078412f
C8167 a_8530_39574# VDAC_N 0.06498f
C8168 a_7754_38470# a_8912_37509# 0.575911f
C8169 a_n2302_37690# a_n2216_37690# 0.011479f
C8170 a_n4064_37440# a_n4251_37440# 0.00105f
C8171 a_6123_31319# VDD 0.532709f
C8172 a_n2109_47186# a_5129_47502# 0.021297f
C8173 a_n971_45724# a_3785_47178# 0.032234f
C8174 a_n237_47217# a_n1151_42308# 0.63407f
C8175 a_1431_47204# a_584_46384# 0.005844f
C8176 a_n1741_47186# a_n443_46116# 0.053258f
C8177 a_1209_47178# a_2553_47502# 8.64e-19
C8178 a_1239_47204# a_2063_45854# 3.11e-20
C8179 a_15037_45618# a_11341_43940# 2.21e-21
C8180 a_15415_45028# a_14673_44172# 9.28e-20
C8181 a_18315_45260# a_17970_44736# 6.02e-19
C8182 a_n2433_44484# a_n1917_44484# 0.113784f
C8183 a_16922_45042# a_18374_44850# 9.15e-20
C8184 a_n2129_44697# a_n1699_44726# 0.018607f
C8185 a_n2661_44458# a_n1177_44458# 0.006328f
C8186 a_11827_44484# a_8975_43940# 0.076327f
C8187 a_11691_44458# a_10157_44484# 1.48e-20
C8188 a_13556_45296# a_15146_44484# 4.94e-20
C8189 a_n2661_43370# a_5289_44734# 3.39e-19
C8190 a_n913_45002# a_n1331_43914# 3.47e-19
C8191 a_n2293_45010# a_175_44278# 0.030523f
C8192 a_n2017_45002# a_n809_44244# 1.63e-21
C8193 en_comp a_n2472_43914# 0.014244f
C8194 a_n2661_45010# a_1115_44172# 0.003124f
C8195 a_n1059_45260# a_n1549_44318# 3.77e-19
C8196 a_n2840_42282# a_n2956_38216# 2.12e-20
C8197 a_n4318_38216# a_n2810_45572# 0.023144f
C8198 a_20836_43172# a_n357_42282# 9.04e-20
C8199 COMP_P a_20205_31679# 3.65e-20
C8200 a_9313_44734# a_16327_47482# 0.169217f
C8201 a_3422_30871# w_1575_34946# 1.88476f
C8202 a_14495_45572# a_2324_44458# 0.00152f
C8203 a_10907_45822# a_10903_43370# 0.199567f
C8204 a_10193_42453# a_6945_45028# 9.46e-20
C8205 a_15143_45578# a_14840_46494# 1.28e-19
C8206 a_11064_45572# a_8199_44636# 7.43e-21
C8207 a_3357_43084# a_19551_46910# 5.32e-20
C8208 a_n1059_45260# a_13059_46348# 2.69e-20
C8209 a_5205_44484# a_3090_45724# 0.005908f
C8210 a_6171_45002# a_15368_46634# 1.38e-19
C8211 a_2437_43646# a_20273_46660# 4.41e-20
C8212 a_3638_45822# a_526_44458# 3.45e-19
C8213 a_5263_45724# a_5066_45546# 0.022243f
C8214 a_3775_45552# a_n1925_42282# 2.95e-21
C8215 a_n699_43396# a_768_44030# 1.37533f
C8216 a_11787_45002# a_11813_46116# 1.43e-19
C8217 a_11963_45334# a_11735_46660# 1.91e-21
C8218 a_17568_45572# a_11415_45002# 9.66e-19
C8219 a_20256_43172# a_20573_43172# 0.001295f
C8220 a_10341_42308# a_10149_42308# 1.97e-19
C8221 a_5534_30871# a_14113_42308# 5.72e-21
C8222 a_11309_47204# a_n2661_46634# 0.042272f
C8223 a_n881_46662# a_n743_46660# 0.527182f
C8224 a_n1613_43370# a_n2438_43548# 1.04064f
C8225 a_n2312_40392# a_n2661_46098# 1.45e-20
C8226 a_9313_45822# a_8492_46660# 8.95e-19
C8227 a_6545_47178# a_6969_46634# 0.002934f
C8228 a_9863_47436# a_10150_46912# 4.65e-21
C8229 a_n1435_47204# a_8145_46902# 4.03e-21
C8230 a_6491_46660# a_6755_46942# 0.007927f
C8231 a_6151_47436# a_6682_46987# 0.003543f
C8232 a_2063_45854# a_11186_47026# 0.012485f
C8233 a_n971_45724# a_3090_45724# 0.071442f
C8234 a_n1151_42308# a_8270_45546# 0.01803f
C8235 a_17517_44484# a_20679_44626# 0.031895f
C8236 a_1307_43914# a_4699_43561# 1.54e-19
C8237 a_10193_42453# a_12895_43230# 1.15e-20
C8238 a_11823_42460# a_10796_42968# 5.88e-19
C8239 a_5883_43914# a_9672_43914# 4.69e-19
C8240 a_626_44172# a_1568_43370# 1.82e-21
C8241 a_n1821_44484# a_n4318_39768# 3.01e-19
C8242 a_3537_45260# a_3457_43396# 3.07e-20
C8243 a_5205_44484# a_6547_43396# 1.82e-19
C8244 a_7229_43940# a_6197_43396# 0.001981f
C8245 a_n913_45002# a_14205_43396# 3.11e-19
C8246 a_n1059_45260# a_15095_43370# 0.108103f
C8247 a_5111_44636# a_6452_43396# 0.024938f
C8248 a_3232_43370# a_8147_43396# 1.83e-19
C8249 a_1606_42308# C5_P_btm 1.89e-19
C8250 a_2779_44458# a_1823_45246# 0.00892f
C8251 a_742_44458# a_167_45260# 9.2e-20
C8252 a_949_44458# a_2202_46116# 7.07e-21
C8253 a_17767_44458# a_11415_45002# 4.21e-20
C8254 a_16112_44458# a_12741_44636# 0.019518f
C8255 a_19478_44306# a_5807_45002# 0.001092f
C8256 a_10405_44172# a_n2293_46634# 0.002468f
C8257 a_15493_43396# a_13661_43548# 0.491785f
C8258 a_13017_45260# a_12839_46116# 5.04e-21
C8259 a_1423_45028# a_8049_45260# 1.12e-19
C8260 a_n2661_43370# a_n2956_38680# 2.4e-20
C8261 a_1307_43914# a_10586_45546# 1.48e-20
C8262 a_n467_45028# a_n452_45724# 0.001128f
C8263 a_n143_45144# a_n863_45724# 0.033306f
C8264 a_2274_45254# a_n2661_45546# 0.002096f
C8265 a_413_45260# a_n2293_45546# 0.066602f
C8266 en_comp a_n357_42282# 2.96e-20
C8267 a_16922_45042# a_17715_44484# 0.039816f
C8268 a_20974_43370# a_16327_47482# 0.004018f
C8269 a_3080_42308# a_4791_45118# 1.96e-19
C8270 a_4699_43561# a_n443_46116# 9.16e-21
C8271 a_14456_42282# a_7174_31319# 9.76e-21
C8272 a_1606_42308# a_n3420_38528# 2.3e-20
C8273 a_9067_47204# VDD 0.47483f
C8274 a_13467_32519# CAL_N 2.02e-19
C8275 a_13661_43548# a_3483_46348# 0.381471f
C8276 a_n2293_46634# a_n901_46420# 3.18e-20
C8277 a_n2661_46634# a_472_46348# 1.17e-20
C8278 a_n1021_46688# a_n1853_46287# 2.81e-20
C8279 a_n2438_43548# a_n2293_46098# 0.409291f
C8280 a_n1925_46634# a_n1991_46122# 0.008581f
C8281 a_11735_46660# a_11901_46660# 0.579036f
C8282 a_4817_46660# a_765_45546# 0.010165f
C8283 a_10428_46928# a_10933_46660# 2.28e-19
C8284 a_10249_46116# a_10425_46660# 3.17e-19
C8285 a_6755_46942# a_10185_46660# 3.5e-19
C8286 a_9804_47204# a_9625_46129# 0.037672f
C8287 a_n881_46662# a_11189_46129# 2.91e-19
C8288 a_8128_46384# a_9569_46155# 3.31e-20
C8289 a_5649_42852# VDAC_N 3.45e-20
C8290 a_21177_47436# a_10809_44734# 0.009997f
C8291 a_21496_47436# a_6945_45028# 0.001335f
C8292 a_13507_46334# a_22223_46124# 0.024274f
C8293 a_4883_46098# a_21137_46414# 0.010468f
C8294 a_6575_47204# a_8034_45724# 2.35e-20
C8295 a_11453_44696# a_18985_46122# 9.23e-20
C8296 a_n2065_43946# a_n2267_43396# 0.009359f
C8297 a_n1761_44111# a_n2129_43609# 0.029483f
C8298 a_n1899_43946# a_n2433_43396# 6.91e-19
C8299 a_10729_43914# a_11173_44260# 0.057346f
C8300 a_10949_43914# a_10555_44260# 0.034175f
C8301 a_14955_43940# a_15493_43940# 0.110232f
C8302 a_17737_43940# a_11341_43940# 0.004705f
C8303 a_n356_44636# a_16977_43638# 1.19e-21
C8304 a_9313_44734# a_10341_43396# 0.175125f
C8305 a_n2433_44484# a_n1853_43023# 2.06e-21
C8306 a_11967_42832# a_3626_43646# 0.001552f
C8307 a_10193_42453# a_18220_42308# 0.004148f
C8308 a_5343_44458# a_4361_42308# 0.004068f
C8309 a_15493_43396# a_19862_44208# 8.78e-19
C8310 a_5891_43370# a_8945_43396# 2.41e-19
C8311 a_11823_42460# a_4958_30871# 4.65e-19
C8312 a_5883_43914# a_743_42282# 3.05e-20
C8313 a_18989_43940# a_18783_43370# 4.79e-19
C8314 a_19479_31679# COMP_P 2e-20
C8315 a_n913_45002# a_22400_42852# 0.002067f
C8316 a_n2017_45002# a_19326_42852# 3.73e-19
C8317 a_13904_45546# a_13249_42308# 0.13587f
C8318 a_10490_45724# a_10210_45822# 0.014252f
C8319 a_8568_45546# a_8791_45572# 0.011458f
C8320 a_7499_43078# a_8697_45572# 0.004673f
C8321 a_8746_45002# a_10907_45822# 1.47e-19
C8322 C0_dummy_P_btm C2_P_btm 7.14548f
C8323 C0_dummy_N_btm C3_P_btm 2.08e-19
C8324 C3_N_btm C7_P_btm 3.05e-19
C8325 C2_N_btm C6_P_btm 7.09e-20
C8326 C1_N_btm C5_P_btm 8.82e-20
C8327 C0_N_btm C4_P_btm 7.74e-20
C8328 a_18599_43230# a_16327_47482# 0.182696f
C8329 a_10807_43548# a_8199_44636# 6.84e-21
C8330 a_n2293_43922# a_n863_45724# 7.65e-20
C8331 a_8375_44464# a_n443_42852# 6.71e-19
C8332 a_n2661_42834# a_380_45546# 3.2e-21
C8333 a_13678_32519# a_22612_30879# 0.060546f
C8334 a_5934_30871# a_6886_37412# 3.68e-19
C8335 a_3483_46348# a_4185_45028# 0.430982f
C8336 a_5257_43370# a_n755_45592# 2.64e-20
C8337 a_11415_45002# a_15015_46420# 4.21e-20
C8338 a_12741_44636# a_13925_46122# 7.71e-21
C8339 a_1823_45246# a_6165_46155# 3.85e-21
C8340 a_21188_46660# a_21137_46414# 4.35e-19
C8341 a_21363_46634# a_6945_45028# 1.28e-19
C8342 a_20841_46902# a_10809_44734# 0.006187f
C8343 a_22223_43948# a_22223_43396# 0.025171f
C8344 a_2982_43646# a_6031_43396# 8.49e-21
C8345 a_20974_43370# a_10341_43396# 0.08579f
C8346 a_15493_43940# a_5649_42852# 3.25e-20
C8347 a_n2661_42282# a_3681_42891# 1.24e-20
C8348 a_5883_43914# a_5755_42308# 4.69e-21
C8349 a_5343_44458# a_6761_42308# 1.34e-19
C8350 a_4223_44672# a_7963_42308# 2.12e-21
C8351 a_1568_43370# a_2813_43396# 4.85e-19
C8352 a_n356_44636# a_n1630_35242# 5.72e-21
C8353 a_n1741_47186# DATA[4] 0.020035f
C8354 a_n452_47436# DATA[0] 0.039965f
C8355 a_16147_45260# a_16751_45260# 0.054632f
C8356 a_10193_42453# a_11827_44484# 0.121679f
C8357 a_7499_43078# a_11691_44458# 0.007969f
C8358 a_n1059_45260# a_n659_45366# 0.001645f
C8359 a_n2810_45028# a_n2956_37592# 6.13705f
C8360 a_n2661_45010# a_413_45260# 0.003446f
C8361 a_3357_43084# a_3537_45260# 0.026461f
C8362 a_n2293_45010# a_n143_45144# 7.12e-21
C8363 a_n913_45002# a_n967_45348# 1.00127f
C8364 a_6171_42473# a_n2293_46634# 2.55e-21
C8365 a_5932_42308# a_n2442_46660# 5.39e-21
C8366 a_n97_42460# a_n863_45724# 0.581863f
C8367 a_3626_43646# a_13259_45724# 0.037016f
C8368 a_n2267_43396# a_n755_45592# 2.31e-20
C8369 a_n1699_43638# a_n357_42282# 4.63e-20
C8370 a_15743_43084# a_17715_44484# 1.72e-19
C8371 a_20712_42282# a_18597_46090# 8.69e-19
C8372 a_17730_32519# a_22459_39145# 1.35e-20
C8373 a_n2472_45546# VDD 0.290266f
C8374 a_10907_45822# a_4883_46098# 1.59e-21
C8375 a_15765_45572# a_11599_46634# 0.001673f
C8376 a_2437_43646# a_n2109_47186# 0.027184f
C8377 a_10053_45546# a_n881_46662# 4.53e-21
C8378 a_8162_45546# a_8128_46384# 2.64e-19
C8379 a_6511_45714# a_5807_45002# 0.012932f
C8380 a_526_44458# a_3316_45546# 0.128261f
C8381 a_1337_46116# a_n755_45592# 8.94e-20
C8382 a_8049_45260# a_20850_46155# 3.79e-19
C8383 a_6031_43396# a_5837_42852# 5.29e-20
C8384 a_n2840_42826# a_n2157_42858# 7.58e-21
C8385 a_10341_43396# a_18599_43230# 1.21e-19
C8386 a_15597_42852# VDD 0.239357f
C8387 a_18175_45572# a_18579_44172# 5.04e-22
C8388 a_14180_45002# a_13720_44458# 4.96e-19
C8389 a_2711_45572# a_11341_43940# 1.54309f
C8390 a_16922_45042# a_17719_45144# 0.22253f
C8391 a_1423_45028# a_8103_44636# 0.064947f
C8392 a_1307_43914# a_10440_44484# 5.64e-20
C8393 a_9482_43914# a_14539_43914# 2.22e-19
C8394 a_7499_43078# a_8333_44056# 0.005667f
C8395 a_17023_45118# a_17613_45144# 0.001643f
C8396 a_13556_45296# a_16112_44458# 0.001671f
C8397 a_5009_45028# a_n2661_44458# 0.002424f
C8398 a_n2293_45010# a_n2293_43922# 0.00103f
C8399 a_n2017_45002# a_n2661_42834# 0.037965f
C8400 a_n467_45028# a_n310_44484# 2.23e-19
C8401 a_22165_42308# a_n357_42282# 1.25e-19
C8402 a_n1329_42308# a_n2956_39304# 6.85e-20
C8403 COMP_P a_n2956_38680# 0.001147f
C8404 a_8791_42308# a_4185_45028# 1.64e-19
C8405 a_6667_45809# a_3483_46348# 3.14e-22
C8406 a_15599_45572# a_13059_46348# 5.07e-19
C8407 a_8696_44636# a_14035_46660# 6.34e-21
C8408 a_19431_45546# a_3090_45724# 4.09e-21
C8409 a_1307_43914# a_n743_46660# 0.002676f
C8410 a_9482_43914# a_2107_46812# 0.109711f
C8411 a_1145_45348# a_n2293_46634# 1.48e-19
C8412 a_3537_45260# a_3877_44458# 0.12249f
C8413 a_3357_43084# a_6969_46634# 3.01e-20
C8414 a_413_45260# a_5732_46660# 8.11e-21
C8415 a_5263_45724# a_5068_46348# 2.95e-19
C8416 a_2711_45572# a_5497_46414# 0.001047f
C8417 a_19778_44110# a_11453_44696# 8.76e-20
C8418 a_21359_45002# a_4883_46098# 5.09e-22
C8419 a_22223_45036# a_13507_46334# 0.005873f
C8420 a_18114_32519# a_16327_47482# 5.2e-20
C8421 a_5883_43914# a_6151_47436# 8.07e-21
C8422 a_n356_44636# a_n971_45724# 1.4e-19
C8423 a_6194_45824# a_4419_46090# 7.7e-20
C8424 a_17324_43396# a_17303_42282# 2.04e-20
C8425 a_17499_43370# a_17531_42308# 9.86e-20
C8426 a_5649_42852# a_5742_30871# 0.059614f
C8427 a_4361_42308# a_12563_42308# 0.009982f
C8428 a_4190_30871# a_14113_42308# 6.14e-20
C8429 a_19164_43230# a_19326_42852# 0.006453f
C8430 a_20922_43172# a_22400_42852# 1.28e-20
C8431 a_743_42282# a_13333_42558# 0.001019f
C8432 a_20692_30879# a_22609_37990# 1.07e-20
C8433 a_2905_45572# a_2107_46812# 0.031826f
C8434 a_327_47204# a_n2661_46098# 2.08e-20
C8435 a_n1151_42308# a_1123_46634# 0.002563f
C8436 a_1209_47178# a_1799_45572# 1.57e-19
C8437 a_n971_45724# a_3699_46634# 0.024384f
C8438 a_n443_46116# a_n743_46660# 0.532861f
C8439 a_12861_44030# a_13747_46662# 0.139424f
C8440 a_7227_47204# a_n2661_46634# 1.7e-19
C8441 a_15507_47210# a_16697_47582# 2.56e-19
C8442 a_16023_47582# a_16119_47582# 0.013793f
C8443 a_17591_47464# a_12549_44172# 0.001606f
C8444 a_14311_47204# a_5807_45002# 3.38e-19
C8445 a_10227_46804# a_12891_46348# 0.058451f
C8446 a_n2433_44484# a_n1899_43946# 2.69e-19
C8447 a_n2267_44484# a_n2065_43946# 1.98e-19
C8448 a_17767_44458# a_11967_42832# 0.003339f
C8449 a_n2661_44458# a_n1331_43914# 8.46e-21
C8450 a_n2129_44697# a_n1761_44111# 5.53e-19
C8451 a_n2661_43370# a_9028_43914# 5.67e-21
C8452 a_8696_44636# a_9145_43396# 2.59e-20
C8453 a_5608_44484# a_5708_44484# 0.005294f
C8454 a_18248_44752# a_18588_44850# 0.027606f
C8455 a_9313_44734# a_n2293_43922# 0.026681f
C8456 a_14537_43396# a_15301_44260# 2.79e-19
C8457 a_n310_44484# a_n2661_43922# 1.2e-19
C8458 a_n89_44484# a_n2661_42834# 2.61e-19
C8459 a_n2017_45002# a_n1352_43396# 8.78e-19
C8460 a_n2293_45010# a_n97_42460# 4.81e-19
C8461 en_comp a_n2433_43396# 0.036527f
C8462 a_n2302_39866# a_n2956_38216# 3.61e-19
C8463 a_17737_43940# a_16327_47482# 3e-21
C8464 a_20269_44172# a_12861_44030# 0.047709f
C8465 a_3737_43940# a_584_46384# 8.18e-19
C8466 a_22591_45572# a_8049_45260# 0.036446f
C8467 a_5244_44056# a_n881_46662# 1.42e-21
C8468 a_13556_45296# a_13925_46122# 2.8e-21
C8469 a_13777_45326# a_13759_46122# 9.69e-19
C8470 a_11963_45334# a_2324_44458# 0.001724f
C8471 a_1423_45028# a_8953_45546# 0.021907f
C8472 a_5365_45348# a_5164_46348# 5.46e-19
C8473 a_17568_45572# a_13259_45724# 0.005159f
C8474 a_1467_44172# a_768_44030# 0.022755f
C8475 a_21359_45002# a_21188_46660# 4.5e-21
C8476 a_20567_45036# a_20731_47026# 2.2e-21
C8477 a_16405_45348# a_11415_45002# 9.91e-19
C8478 a_n2293_42834# a_1138_42852# 0.015752f
C8479 a_7963_42308# a_5742_30871# 1.16e-20
C8480 COMP_P a_13258_32519# 0.010297f
C8481 a_8685_42308# a_9293_42558# 0.003228f
C8482 C8_P_btm C6_P_btm 0.163943f
C8483 C9_P_btm C5_P_btm 0.150576f
C8484 C10_P_btm C4_P_btm 0.703336f
C8485 a_13747_46662# a_14180_46812# 0.021289f
C8486 a_4646_46812# a_6755_46942# 0.362783f
C8487 a_3877_44458# a_6969_46634# 0.101189f
C8488 a_n2661_46634# a_12156_46660# 0.009815f
C8489 a_5429_46660# a_5257_43370# 2.57e-20
C8490 a_12549_44172# a_15312_46660# 5.76e-20
C8491 a_11309_47204# a_765_45546# 0.03506f
C8492 a_11453_44696# a_20820_30879# 0.002153f
C8493 SMPL_ON_N a_12741_44636# 8.39e-20
C8494 a_22223_47212# a_21076_30879# 7.91e-19
C8495 a_6151_47436# a_9569_46155# 2.49e-19
C8496 a_6575_47204# a_8016_46348# 5.51e-20
C8497 a_n1435_47204# a_5068_46348# 3.74e-21
C8498 a_4915_47217# a_9290_44172# 0.002979f
C8499 a_n2497_47436# a_n2956_38680# 2.47e-20
C8500 a_n1151_42308# a_13759_46122# 2.36e-19
C8501 a_584_46384# a_2324_44458# 2.7e-19
C8502 a_18587_45118# a_18525_43370# 1.2e-22
C8503 a_5663_43940# a_n2661_42282# 0.00715f
C8504 a_22485_44484# a_11341_43940# 0.006131f
C8505 a_1307_43914# a_1847_42826# 0.428505f
C8506 a_20512_43084# a_22223_43948# 0.001071f
C8507 a_18184_42460# a_17499_43370# 2.47e-20
C8508 a_375_42282# a_685_42968# 2.44e-19
C8509 a_9313_44734# a_n97_42460# 1.76217f
C8510 a_n2293_42834# a_5649_42852# 0.002922f
C8511 a_10057_43914# a_8791_43396# 2.04e-20
C8512 a_n356_44636# a_1427_43646# 0.00321f
C8513 a_11827_44484# a_16137_43396# 8.22e-20
C8514 a_18114_32519# a_10341_43396# 4.67e-19
C8515 a_n913_45002# a_22223_42860# 0.011179f
C8516 en_comp a_21356_42826# 4.89e-21
C8517 a_n2017_45002# a_n2293_42282# 0.095773f
C8518 a_3357_43084# a_4649_43172# 1.01e-20
C8519 a_n4209_39304# VIN_P 0.049722f
C8520 a_n4209_38502# C5_P_btm 0.040445f
C8521 a_n3565_38502# C7_P_btm 1.43e-20
C8522 a_n3565_38216# a_n1386_35608# 1.22e-21
C8523 a_6472_45840# a_6667_45809# 0.215953f
C8524 a_6194_45824# a_6598_45938# 0.051162f
C8525 a_1115_44172# a_1138_42852# 0.012127f
C8526 a_5013_44260# a_n2293_46098# 0.040459f
C8527 a_3457_43396# a_n2293_46634# 8.01e-19
C8528 a_8415_44056# a_8270_45546# 1.57e-19
C8529 a_15301_44260# a_3090_45724# 9.33e-19
C8530 a_12281_43396# a_12549_44172# 0.004094f
C8531 a_n2661_42834# a_526_44458# 0.06021f
C8532 a_n2661_44458# a_2957_45546# 5.79e-21
C8533 a_n452_44636# a_n452_45724# 6.69e-19
C8534 a_16112_44458# a_16375_45002# 4.06e-20
C8535 a_n1177_44458# a_n1099_45572# 2.8e-19
C8536 a_17767_44458# a_13259_45724# 0.026768f
C8537 a_742_44458# a_n863_45724# 0.629795f
C8538 a_4743_44484# a_n2661_45546# 0.004404f
C8539 a_17517_44484# a_19335_46494# 2.71e-21
C8540 a_4361_42308# a_10227_46804# 0.073929f
C8541 a_20556_43646# a_18597_46090# 1.94e-19
C8542 a_1847_42826# a_n443_46116# 0.00118f
C8543 a_19963_31679# a_22609_38406# 3.67e-21
C8544 a_1239_39043# a_1177_38525# 0.031327f
C8545 a_n4209_38502# a_n3420_38528# 0.230544f
C8546 a_n4064_39072# a_n4209_38216# 0.03057f
C8547 a_n3420_39072# a_n3565_38216# 0.030682f
C8548 a_n4334_38528# a_n3690_38528# 8.67e-19
C8549 a_5167_46660# VDD 0.203378f
C8550 a_4958_30871# C0_dummy_P_btm 1.65e-20
C8551 a_765_45546# a_472_46348# 6.08e-19
C8552 a_4646_46812# a_8049_45260# 0.001749f
C8553 a_13661_43548# a_n357_42282# 2.24e-19
C8554 a_n2956_39768# a_n2810_45572# 0.043168f
C8555 a_n2840_46634# a_n2661_45546# 6.53e-19
C8556 a_14084_46812# a_13759_46122# 0.001243f
C8557 a_11901_46660# a_2324_44458# 9.43e-21
C8558 a_15368_46634# a_10903_43370# 4.05e-21
C8559 a_12429_44172# a_12281_43396# 1.87e-20
C8560 a_17737_43940# a_10341_43396# 4.05e-20
C8561 a_n2433_43396# a_n1699_43638# 0.062578f
C8562 a_n2129_43609# a_n2267_43396# 0.230013f
C8563 a_15493_43940# a_8685_43396# 6.24e-19
C8564 a_n2293_42834# a_7963_42308# 7.42e-19
C8565 a_1307_43914# a_15486_42560# 9.69e-21
C8566 a_n4318_39304# a_n1917_43396# 1.69e-19
C8567 a_n2956_37592# a_n2302_40160# 0.006106f
C8568 en_comp a_n4064_40160# 1.93e-20
C8569 a_3065_45002# a_7174_31319# 4.88e-21
C8570 a_13163_45724# a_13017_45260# 2.76e-20
C8571 a_5263_45724# a_5093_45028# 4.44e-20
C8572 a_11823_42460# a_13348_45260# 4.52e-20
C8573 a_2711_45572# a_7418_45394# 9.37e-20
C8574 a_19256_45572# a_20528_45572# 1.03e-20
C8575 a_10907_45822# a_3232_43370# 4.17e-19
C8576 a_8696_44636# a_n1059_45260# 2.7e-21
C8577 a_7174_31319# w_1575_34946# 0.001988f
C8578 a_n1177_43370# a_n1925_42282# 1.62e-22
C8579 a_19862_44208# a_n357_42282# 0.138067f
C8580 a_10949_43914# a_n443_42852# 3.54e-20
C8581 a_4361_42308# a_17339_46660# 3.78e-20
C8582 a_4520_42826# a_3090_45724# 2.44e-19
C8583 a_18707_42852# a_13661_43548# 1.38e-19
C8584 a_15567_42826# a_6755_46942# 7.16e-21
C8585 a_518_46482# VDD 3.14e-19
C8586 a_2711_45572# a_16327_47482# 0.101699f
C8587 a_6812_45938# a_6491_46660# 1.44e-21
C8588 a_8162_45546# a_6151_47436# 6.52e-20
C8589 a_9049_44484# a_4915_47217# 1.19e-20
C8590 a_11652_45724# a_n1151_42308# 4.93e-20
C8591 a_8697_45822# a_n971_45724# 0.002809f
C8592 a_167_45260# a_3503_45724# 1.15e-19
C8593 a_3699_46348# a_n755_45592# 0.003336f
C8594 a_2804_46116# a_2957_45546# 0.009196f
C8595 a_472_46348# a_509_45822# 2.66e-19
C8596 a_376_46348# a_n443_42852# 7.22e-19
C8597 a_4185_45028# a_n357_42282# 0.023019f
C8598 a_526_44458# a_5066_45546# 0.009401f
C8599 a_15015_46420# a_13259_45724# 0.001291f
C8600 a_n743_46660# DATA[4] 1.69e-21
C8601 a_19268_43646# a_19700_43370# 0.017165f
C8602 a_16243_43396# a_16823_43084# 0.05964f
C8603 a_10341_43396# a_13887_32519# 0.030175f
C8604 a_6197_43396# a_5755_42852# 4.26e-20
C8605 a_n97_42460# a_18599_43230# 0.006824f
C8606 a_3905_42865# a_4921_42308# 1.92e-19
C8607 a_3626_43646# a_10518_42984# 2.25e-20
C8608 a_2982_43646# a_10796_42968# 8.58e-20
C8609 a_15743_43084# a_16664_43396# 0.01372f
C8610 a_16977_43638# a_17486_43762# 2.6e-19
C8611 a_16409_43396# a_16855_43396# 2.28e-19
C8612 a_33_46660# DATA[0] 1.05e-20
C8613 a_18083_42858# VDD 0.408512f
C8614 a_19963_31679# a_22521_40599# 1.85e-20
C8615 a_n2810_45028# a_n2860_37690# 6.28e-19
C8616 a_n2956_37592# a_n2302_37690# 0.04217f
C8617 a_9482_43914# a_14309_45028# 3.6e-19
C8618 a_14797_45144# a_14976_45348# 0.007688f
C8619 a_14537_43396# a_15060_45348# 0.001339f
C8620 a_13556_45296# a_13807_45067# 2.63e-19
C8621 a_n967_45348# a_n2661_44458# 0.0255f
C8622 a_n2661_45010# a_2779_44458# 4.72e-20
C8623 a_n2293_45010# a_742_44458# 3.27e-20
C8624 en_comp a_n2433_44484# 0.029809f
C8625 a_n1059_45260# a_n1177_44458# 9.59e-19
C8626 a_n1630_35242# a_21076_30879# 0.034943f
C8627 a_14113_42308# a_15227_44166# 4.65e-20
C8628 a_n2157_42858# a_n357_42282# 1.01e-19
C8629 a_n2293_42282# a_526_44458# 0.010969f
C8630 a_n3674_39304# a_n2956_38216# 0.023342f
C8631 a_n901_43156# a_n863_45724# 1.75e-19
C8632 a_13291_42460# a_9290_44172# 0.078684f
C8633 a_17538_32519# a_22459_39145# 1.25e-20
C8634 a_14401_32519# a_22521_39511# 8.94e-21
C8635 a_14537_43396# a_12465_44636# 0.031033f
C8636 a_9482_43914# a_11453_44696# 0.042575f
C8637 a_15415_45028# a_4883_46098# 1.77e-20
C8638 a_5111_44636# a_n881_46662# 0.00608f
C8639 a_3537_45260# a_8128_46384# 0.001708f
C8640 a_4927_45028# a_n1613_43370# 6.4e-22
C8641 a_2437_43646# a_n1925_46634# 0.02753f
C8642 a_3357_43084# a_n2293_46634# 0.963711f
C8643 a_327_44734# a_768_44030# 0.00311f
C8644 a_11136_45572# a_10467_46802# 1.63e-20
C8645 a_22959_43396# a_14097_32519# 0.00104f
C8646 a_21195_42852# a_21671_42860# 0.177876f
C8647 a_2982_43646# a_4958_30871# 0.136637f
C8648 a_8037_42858# a_9114_42852# 1.46e-19
C8649 a_21356_42826# a_22165_42308# 5.1e-21
C8650 a_8685_43396# a_5742_30871# 4.78e-19
C8651 a_17364_32525# a_22400_42852# 1.05e-20
C8652 a_3626_43646# a_16197_42308# 7.17e-19
C8653 a_13925_46122# RST_Z 4.05e-21
C8654 a_22775_42308# VDD 0.426018f
C8655 a_n1741_47186# a_n1613_43370# 0.018791f
C8656 a_n971_45724# a_2583_47243# 0.006608f
C8657 a_n785_47204# a_7_47243# 7.85e-19
C8658 a_1209_47178# a_2747_46873# 2.14e-19
C8659 a_13717_47436# a_15507_47210# 2.86e-19
C8660 a_12861_44030# a_11599_46634# 0.169929f
C8661 a_18494_42460# a_17517_44484# 0.022635f
C8662 a_6298_44484# a_7640_43914# 0.031665f
C8663 a_5343_44458# a_5891_43370# 1.06553f
C8664 a_18248_44752# a_18443_44721# 0.206455f
C8665 a_1307_43914# a_5244_44056# 0.025291f
C8666 a_2711_45572# a_10341_43396# 0.03441f
C8667 a_n452_44636# a_n310_44484# 0.007833f
C8668 a_n2661_44458# a_9159_44484# 1.56e-19
C8669 a_17970_44736# a_18374_44850# 0.051162f
C8670 a_17767_44458# a_18989_43940# 3.82e-21
C8671 a_n2840_44458# a_n2661_42834# 8.29e-19
C8672 a_11827_44484# a_13940_44484# 4.46e-19
C8673 a_3232_43370# a_n2661_42282# 0.005579f
C8674 a_n4334_39392# a_n2956_39304# 6.77e-20
C8675 a_9223_42460# a_n755_45592# 1.28e-19
C8676 a_6481_42558# a_n443_42852# 0.001736f
C8677 a_n4209_39304# a_n2956_38680# 0.021073f
C8678 a_13921_42308# a_13259_45724# 9.76e-19
C8679 a_9803_42558# a_n357_42282# 4.98e-21
C8680 a_8103_44636# a_4646_46812# 0.002138f
C8681 a_13857_44734# a_768_44030# 0.011246f
C8682 a_4927_45028# a_n2293_46098# 0.015237f
C8683 a_14976_45348# a_14976_45028# 0.002418f
C8684 a_n467_45028# a_167_45260# 1.04e-19
C8685 a_413_45260# a_1138_42852# 0.026098f
C8686 a_12791_45546# a_13259_45724# 0.001427f
C8687 a_11682_45822# a_10586_45546# 0.014019f
C8688 a_4808_45572# a_n2661_45546# 0.001338f
C8689 a_13249_42308# a_14537_46482# 1.3e-20
C8690 a_17668_45572# a_17715_44484# 0.006757f
C8691 a_19256_45572# a_19335_46494# 5.26e-20
C8692 a_18479_45785# a_6945_45028# 4.52e-21
C8693 a_3357_43084# a_9625_46129# 1.12e-20
C8694 a_19279_43940# a_4883_46098# 3.51e-21
C8695 a_3422_30871# a_18479_47436# 1.58e-20
C8696 a_20980_44850# a_18597_46090# 0.005953f
C8697 a_5013_44260# a_4791_45118# 0.02062f
C8698 a_1184_42692# a_2713_42308# 4.61e-20
C8699 a_1755_42282# a_2123_42473# 0.014573f
C8700 a_1606_42308# a_2351_42308# 0.191324f
C8701 a_14635_42282# a_14113_42308# 0.052122f
C8702 a_n2661_46634# a_4955_46873# 0.03751f
C8703 a_2107_46812# a_2443_46660# 0.013591f
C8704 a_1983_46706# a_n2661_46098# 0.147223f
C8705 a_948_46660# a_2609_46660# 2.98e-20
C8706 a_n2293_46634# a_3877_44458# 1.3e-21
C8707 a_n743_46660# a_1302_46660# 0.002121f
C8708 a_288_46660# a_1799_45572# 7.3e-22
C8709 a_5807_45002# a_5429_46660# 1.03e-19
C8710 a_9804_47204# a_6755_46942# 0.028571f
C8711 a_11453_44696# a_12816_46660# 8.81e-22
C8712 a_12465_44636# a_3090_45724# 1.51e-19
C8713 a_n1741_47186# a_n2293_46098# 2.17e-20
C8714 SMPL_ON_P a_n2472_46090# 2.92e-19
C8715 a_n1920_47178# a_n2157_46122# 7.93e-21
C8716 a_n2109_47186# a_n1853_46287# 3.06e-20
C8717 a_n2497_47436# a_n1423_46090# 0.008067f
C8718 a_12861_44030# a_13693_46688# 5.48e-19
C8719 a_n1435_47204# a_13059_46348# 2.88e-21
C8720 a_7227_47204# a_765_45546# 0.005844f
C8721 a_15811_47375# a_13885_46660# 0.0013f
C8722 a_19386_47436# a_19466_46812# 2.89e-19
C8723 a_10227_46804# a_12359_47026# 0.012196f
C8724 a_11599_46634# a_14180_46812# 2.26e-20
C8725 a_18597_46090# a_19692_46634# 0.019861f
C8726 a_20894_47436# a_15227_44166# 9.3e-22
C8727 a_4883_46098# a_15368_46634# 0.023335f
C8728 a_13507_46334# a_16292_46812# 3.92e-19
C8729 a_n2129_44697# a_n2267_43396# 1.8e-20
C8730 a_n2472_43914# a_n1761_44111# 1.8e-19
C8731 a_13857_44734# a_13483_43940# 3.4e-20
C8732 a_9313_44734# a_21115_43940# 9.92e-21
C8733 a_10057_43914# a_10651_43940# 0.003719f
C8734 a_n2293_42834# a_8685_43396# 1.23e-19
C8735 a_n1059_45260# a_n1991_42858# 8.68e-20
C8736 a_n913_45002# a_n1853_43023# 0.094845f
C8737 a_3537_45260# a_743_42282# 0.033447f
C8738 a_n2017_45002# a_n1423_42826# 0.008318f
C8739 a_n2661_45010# a_n13_43084# 4.49e-21
C8740 a_n2293_45010# a_n901_43156# 2.97e-20
C8741 a_18450_45144# VDD 2.13e-19
C8742 a_22465_38105# a_22459_39145# 0.98555f
C8743 a_14358_43442# a_12861_44030# 1.87e-20
C8744 a_8375_44464# a_8199_44636# 0.043989f
C8745 a_17767_44458# a_18189_46348# 3.29e-19
C8746 a_5891_43370# a_8349_46414# 7.96e-21
C8747 a_10334_44484# a_10809_44734# 0.002242f
C8748 a_17970_44736# a_17715_44484# 0.001614f
C8749 a_7640_43914# a_5937_45572# 2.38e-19
C8750 a_1423_45028# a_1609_45822# 2.44e-19
C8751 a_7281_43914# a_3090_45724# 0.170855f
C8752 a_5708_44484# a_3483_46348# 0.005523f
C8753 a_n2661_43922# a_167_45260# 2.12e-19
C8754 a_n4315_30879# a_n4334_39616# 6.38e-20
C8755 a_n4334_40480# a_n4209_39590# 6.38e-20
C8756 a_n4064_40160# a_n2216_40160# 0.005638f
C8757 a_12549_44172# VDD 3.08339f
C8758 a_1606_42308# C4_N_btm 3.05e-19
C8759 a_5257_43370# a_3483_46348# 0.028522f
C8760 a_19333_46634# a_20107_46660# 1.09e-20
C8761 a_15227_44166# a_20411_46873# 0.041968f
C8762 a_13885_46660# a_13059_46348# 9.73e-19
C8763 a_19466_46812# a_19551_46910# 0.008633f
C8764 a_18834_46812# a_20273_46660# 4.32e-20
C8765 a_19692_46634# a_19123_46287# 0.00443f
C8766 a_12156_46660# a_765_45546# 0.001818f
C8767 a_n2312_38680# a_n2956_39304# 5.96956f
C8768 a_n2293_46634# a_n1736_46482# 0.004173f
C8769 a_9804_47204# a_8049_45260# 8.45e-19
C8770 a_8128_46384# a_9241_46436# 1.58e-20
C8771 a_4646_46812# a_8953_45546# 2.27e-20
C8772 a_5732_46660# a_6165_46155# 0.001142f
C8773 a_11453_44696# a_18243_46436# 1.02e-19
C8774 a_13507_46334# a_20254_46482# 3.81e-19
C8775 a_4883_46098# a_19597_46482# 1.2e-19
C8776 a_18479_47436# a_21167_46155# 5.49e-19
C8777 a_n443_46116# a_509_45572# 0.003835f
C8778 a_2889_44172# a_2813_43396# 4.01e-20
C8779 a_21115_43940# a_20974_43370# 2.85e-19
C8780 a_11341_43940# a_14401_32519# 0.008534f
C8781 a_17737_43940# a_n97_42460# 1.26e-20
C8782 a_n2661_42282# a_4905_42826# 5.42e-20
C8783 a_11967_42832# a_18525_43370# 0.010117f
C8784 a_22485_44484# a_10341_43396# 4.73e-20
C8785 a_13076_44458# a_12379_42858# 1.36e-20
C8786 a_n356_44636# a_4520_42826# 2.14e-20
C8787 a_12607_44458# a_12545_42858# 5.22e-21
C8788 a_15493_43940# a_19741_43940# 0.027038f
C8789 a_3537_45260# a_5755_42308# 0.002651f
C8790 a_5147_45002# a_4921_42308# 2e-19
C8791 a_3065_45002# a_5932_42308# 4.34e-21
C8792 en_comp a_8685_42308# 4.34e-21
C8793 a_n2017_45002# a_9885_42558# 0.006803f
C8794 a_3232_43370# a_3497_42558# 7.4e-20
C8795 a_n913_45002# a_9293_42558# 2.08e-19
C8796 a_12429_44172# VDD 0.169047f
C8797 a_15903_45785# a_16680_45572# 5.47e-21
C8798 a_15765_45572# a_16855_45546# 0.042415f
C8799 a_16333_45814# a_16115_45572# 0.209641f
C8800 a_15599_45572# a_8696_44636# 5.37e-19
C8801 a_4699_43561# a_n2293_46098# 0.001614f
C8802 a_15781_43660# a_15227_44166# 0.016739f
C8803 a_16409_43396# a_3090_45724# 4.65e-21
C8804 a_5342_30871# a_n2293_46634# 3.03e-20
C8805 a_n984_44318# a_n863_45724# 0.002194f
C8806 a_n809_44244# a_n452_45724# 4.69e-20
C8807 a_n2065_43946# a_n755_45592# 3.71e-20
C8808 a_1414_42308# a_n2661_45546# 3.34e-20
C8809 a_n1761_44111# a_n357_42282# 0.004602f
C8810 a_11173_43940# a_9290_44172# 0.001076f
C8811 a_16877_42852# a_16327_47482# 7.73e-21
C8812 a_5932_42308# w_1575_34946# 0.0018f
C8813 a_1606_42308# a_584_46384# 2.19e-19
C8814 a_19721_31679# a_22459_39145# 1.93e-20
C8815 a_n2661_43370# CLK 0.011991f
C8816 a_1208_46090# VDD 0.178097f
C8817 a_21335_42336# CAL_N 9.12e-19
C8818 a_n3420_38528# a_n3607_38304# 6.01e-19
C8819 a_n3420_39616# a_n4334_37440# 4.91e-19
C8820 a_n4209_39590# a_n2946_37690# 1.64e-19
C8821 a_n3565_39590# a_n3690_37440# 1.95e-19
C8822 a_1736_39043# VDAC_Pi 0.001304f
C8823 a_1736_39587# VDAC_Ni 5.68e-19
C8824 C0_dummy_N_btm C6_N_btm 0.1194f
C8825 C2_N_btm C3_N_btm 5.99608f
C8826 C0_N_btm C5_N_btm 0.138093f
C8827 C1_N_btm C4_N_btm 0.128167f
C8828 C0_dummy_P_btm C7_N_btm 2.05e-19
C8829 C1_P_btm C9_N_btm 5.29e-19
C8830 C0_P_btm C8_N_btm 3.87e-19
C8831 a_1823_45246# a_5210_46155# 1.93e-20
C8832 a_20411_46873# a_21071_46482# 2.24e-19
C8833 a_4704_46090# a_n1925_42282# 2.45e-19
C8834 a_9290_44172# a_10809_44734# 0.239594f
C8835 a_19237_31679# a_22400_42852# 2.13e-20
C8836 a_14539_43914# a_4958_30871# 0.00214f
C8837 a_n2293_43922# a_8515_42308# 3.54e-20
C8838 a_9313_44734# a_10533_42308# 8.54e-19
C8839 a_19862_44208# a_21356_42826# 0.001265f
C8840 a_15493_43940# a_17333_42852# 1.29e-20
C8841 a_9145_43396# a_14205_43396# 0.13322f
C8842 a_n2433_43396# a_n2157_42858# 2.73e-19
C8843 a_20365_43914# a_19987_42826# 4.65e-20
C8844 a_22223_47212# SINGLE_ENDED 6.55e-19
C8845 SMPL_ON_N RST_Z 2.43362f
C8846 a_21855_43396# VDD 0.289066f
C8847 a_4099_45572# a_n2661_42834# 4.28e-22
C8848 a_18479_45785# a_11827_44484# 0.03055f
C8849 a_10907_45822# a_8975_43940# 1.46e-19
C8850 a_2382_45260# a_2304_45348# 0.045704f
C8851 a_3065_45002# a_1423_45028# 0.017813f
C8852 a_5111_44636# a_1307_43914# 0.114933f
C8853 a_6171_45002# a_14797_45144# 0.00824f
C8854 a_2274_45254# a_2809_45348# 9.76e-19
C8855 a_13460_43230# a_9290_44172# 0.005304f
C8856 a_12545_42858# a_10903_43370# 0.026404f
C8857 a_5565_43396# a_n443_42852# 1.34e-19
C8858 a_n1991_42858# a_n1925_42282# 1.72e-19
C8859 a_18525_43370# a_13259_45724# 5.74e-20
C8860 a_17499_43370# a_16375_45002# 1.41e-19
C8861 a_14579_43548# a_n357_42282# 0.049501f
C8862 a_22775_42308# a_22612_30879# 8.11e-21
C8863 a_21356_42826# a_4185_45028# 1.61e-20
C8864 a_15903_45785# a_13747_46662# 0.022255f
C8865 a_6472_45840# a_5257_43370# 0.012073f
C8866 a_2711_45572# a_8667_46634# 3.36e-20
C8867 a_12749_45572# a_12549_44172# 0.004689f
C8868 a_8192_45572# a_n1925_46634# 0.03394f
C8869 a_13297_45572# a_12891_46348# 3.27e-19
C8870 a_16333_45814# a_5807_45002# 3.87e-19
C8871 a_15765_45572# a_13661_43548# 1.83e-20
C8872 a_16147_45260# a_n881_46662# 3.57e-19
C8873 a_2437_43646# a_20894_47436# 0.007723f
C8874 a_3357_43084# a_18597_46090# 0.160577f
C8875 a_413_45260# a_9863_47436# 1.03e-19
C8876 a_7276_45260# a_n1151_42308# 0.062423f
C8877 a_8953_45002# a_2063_45854# 2.32e-19
C8878 a_4927_45028# a_4791_45118# 0.03353f
C8879 a_n1079_45724# a_n356_45724# 9.52e-19
C8880 a_n357_42282# a_997_45618# 0.023595f
C8881 a_n2661_45546# a_n1013_45572# 0.001202f
C8882 a_22959_43396# a_22959_42860# 0.026152f
C8883 a_n97_42460# a_8515_42308# 2.07e-19
C8884 a_22959_43948# a_22775_42308# 3.38e-21
C8885 a_8387_43230# a_8952_43230# 7.99e-20
C8886 a_8037_42858# a_10518_42984# 2e-20
C8887 a_3080_42308# a_3581_42558# 3.31e-19
C8888 a_20731_47026# SINGLE_ENDED 1.3e-20
C8889 a_3754_38470# VDAC_P 0.323951f
C8890 a_n4064_37440# a_n2216_37690# 0.005567f
C8891 a_8530_39574# a_6886_37412# 0.616015f
C8892 a_n3420_37440# a_n3607_37440# 0.001516f
C8893 a_7754_38470# VDAC_N 0.110573f
C8894 a_7227_42308# VDD 0.296912f
C8895 a_n2109_47186# a_4915_47217# 0.352259f
C8896 a_1209_47178# a_2063_45854# 0.00786f
C8897 a_1431_47204# a_2124_47436# 0.010942f
C8898 a_n971_45724# a_3381_47502# 0.008848f
C8899 a_n746_45260# a_n1151_42308# 0.116939f
C8900 a_1239_47204# a_584_46384# 1.75e-19
C8901 a_n1741_47186# a_4791_45118# 0.024211f
C8902 a_n237_47217# a_3160_47472# 0.037234f
C8903 a_n2293_45010# a_n984_44318# 0.048428f
C8904 a_n2017_45002# a_n1549_44318# 9.31e-19
C8905 a_n2956_37592# a_n2472_43914# 9.42e-21
C8906 a_n2661_45010# a_644_44056# 8.47e-20
C8907 a_n745_45366# a_n1761_44111# 5.25e-20
C8908 a_n913_45002# a_n1899_43946# 0.017336f
C8909 a_n1059_45260# a_n1331_43914# 4.5e-20
C8910 a_11827_44484# a_10057_43914# 2.12e-19
C8911 a_n2661_43370# a_5205_44734# 1.1e-19
C8912 a_7499_43078# a_11257_43940# 6.52e-20
C8913 a_2711_45572# a_n97_42460# 0.137121f
C8914 a_8560_45348# a_5891_43370# 7.06e-20
C8915 a_16922_45042# a_18443_44721# 6.14e-20
C8916 a_n2129_44697# a_n2267_44484# 0.698671f
C8917 a_n2433_44484# a_n1699_44726# 0.058433f
C8918 a_n2661_44458# a_n1917_44484# 0.008101f
C8919 a_17719_45144# a_17970_44736# 4.66e-19
C8920 a_14797_45144# a_14673_44172# 9.74e-20
C8921 a_n2472_42282# a_n2810_45572# 2.3e-20
C8922 a_9885_42558# a_526_44458# 9.36e-19
C8923 a_5891_43370# a_10227_46804# 0.2393f
C8924 a_3775_45552# a_526_44458# 0.015665f
C8925 a_4099_45572# a_5066_45546# 4.69e-20
C8926 a_3357_43084# a_19123_46287# 1.6e-20
C8927 a_n2017_45002# a_13059_46348# 3.52e-20
C8928 a_6171_45002# a_14976_45028# 0.024858f
C8929 a_2437_43646# a_20411_46873# 7.51e-20
C8930 a_13249_42308# a_2324_44458# 0.072143f
C8931 a_15143_45578# a_15015_46420# 0.011172f
C8932 a_11682_45822# a_11189_46129# 0.00283f
C8933 a_10210_45822# a_10903_43370# 0.001155f
C8934 a_10544_45572# a_8199_44636# 1.89e-19
C8935 a_9049_44484# a_10809_44734# 9.15e-21
C8936 a_10180_45724# a_6945_45028# 2.08e-20
C8937 a_7735_45067# a_4646_46812# 2.05e-19
C8938 a_4223_44672# a_768_44030# 0.136643f
C8939 a_11787_45002# a_11735_46660# 1.9e-19
C8940 a_17034_45572# a_11415_45002# 2.62e-19
C8941 a_5534_30871# a_13657_42558# 1.73e-19
C8942 a_16131_47204# a_5807_45002# 6.5e-19
C8943 a_n881_46662# a_n1021_46688# 0.15991f
C8944 a_n1613_43370# a_n743_46660# 0.521102f
C8945 a_n1435_47204# a_7577_46660# 5.91e-21
C8946 a_6151_47436# a_6969_46634# 0.030417f
C8947 a_6545_47178# a_6755_46942# 0.022995f
C8948 a_9863_47436# a_9863_46634# 0.003636f
C8949 a_9313_45822# a_8667_46634# 0.004188f
C8950 a_2063_45854# a_10768_47026# 0.005084f
C8951 a_5883_43914# a_9028_43914# 0.05428f
C8952 a_17517_44484# a_20640_44752# 0.54753f
C8953 a_1307_43914# a_4235_43370# 0.016608f
C8954 a_11823_42460# a_10835_43094# 0.006753f
C8955 a_10193_42453# a_13113_42826# 4.41e-21
C8956 a_626_44172# a_1049_43396# 2.99e-19
C8957 a_11827_44484# a_14021_43940# 3.51e-19
C8958 a_5205_44484# a_6765_43638# 8.52e-19
C8959 a_5111_44636# a_9396_43370# 0.203348f
C8960 a_n913_45002# a_14358_43442# 3.05e-20
C8961 a_n1059_45260# a_14205_43396# 4.2e-20
C8962 a_n2017_45002# a_15095_43370# 0.002423f
C8963 a_5147_45002# a_6452_43396# 2.05e-19
C8964 a_1606_42308# C6_P_btm 2.33e-19
C8965 a_949_44458# a_1823_45246# 0.005758f
C8966 a_16979_44734# a_11415_45002# 3.74e-20
C8967 a_15004_44636# a_12741_44636# 0.008679f
C8968 a_15493_43396# a_5807_45002# 0.002975f
C8969 a_9672_43914# a_n2293_46634# 4.81e-20
C8970 a_19328_44172# a_13661_43548# 2.29e-19
C8971 a_22959_43948# a_12549_44172# 2.47e-20
C8972 a_14673_44172# a_14976_45028# 8.68e-20
C8973 a_n2661_43370# a_n2956_39304# 1.05e-20
C8974 a_1667_45002# a_n2661_45546# 0.003128f
C8975 a_n37_45144# a_n2293_45546# 0.042299f
C8976 a_n467_45028# a_n863_45724# 0.037721f
C8977 a_n967_45348# a_n1099_45572# 3.54e-20
C8978 a_17023_45118# a_15682_46116# 5.09e-19
C8979 a_9801_43940# a_4883_46098# 0.001598f
C8980 a_14401_32519# a_16327_47482# 2.02e-20
C8981 a_4699_43561# a_4791_45118# 1.93e-20
C8982 a_3539_42460# a_584_46384# 9.82e-19
C8983 a_n2661_44458# a_4419_46090# 6.4e-20
C8984 a_13575_42558# a_7174_31319# 4.88e-21
C8985 a_6575_47204# VDD 1.32036f
C8986 a_5807_45002# a_3483_46348# 0.018693f
C8987 a_n743_46660# a_n2293_46098# 0.213418f
C8988 a_n2293_46634# a_n1641_46494# 0.002502f
C8989 a_n2438_43548# a_n2472_46090# 0.020059f
C8990 a_n1021_46688# a_n2157_46122# 0.00108f
C8991 a_n1925_46634# a_n1853_46287# 0.012373f
C8992 a_n2312_38680# a_n1991_46122# 2.37e-19
C8993 a_11735_46660# a_11813_46116# 0.162547f
C8994 a_4955_46873# a_765_45546# 0.008652f
C8995 a_10554_47026# a_10425_46660# 4.2e-19
C8996 a_10249_46116# a_10185_46660# 7.29e-19
C8997 a_9804_47204# a_8953_45546# 3.84e-19
C8998 a_8128_46384# a_9625_46129# 3.11e-20
C8999 a_20990_47178# a_10809_44734# 0.00204f
C9000 a_13507_46334# a_6945_45028# 0.187229f
C9001 a_4883_46098# a_20708_46348# 0.014516f
C9002 a_7903_47542# a_8034_45724# 8.49e-21
C9003 a_11453_44696# a_18819_46122# 7.1e-20
C9004 a_12465_44636# a_20075_46420# 5.91e-21
C9005 a_13678_32519# VDAC_N 3.33e-19
C9006 a_n1899_43946# a_n4318_39304# 2.93e-19
C9007 a_7542_44172# a_8487_44056# 2.54e-20
C9008 a_19328_44172# a_19862_44208# 0.002604f
C9009 a_7845_44172# a_8415_44056# 9.13e-21
C9010 a_5891_43370# a_8873_43396# 0.001547f
C9011 a_10193_42453# a_18214_42558# 0.028997f
C9012 a_n2433_44484# a_n2157_42858# 1.17e-21
C9013 a_n2661_44458# a_n1853_43023# 1.84e-21
C9014 a_n356_44636# a_16409_43396# 3.54e-20
C9015 a_15682_43940# a_11341_43940# 0.021147f
C9016 a_10729_43914# a_10555_44260# 0.038445f
C9017 a_15493_43396# a_19478_44306# 0.154347f
C9018 a_n1761_44111# a_n2433_43396# 5.56e-19
C9019 a_n2065_43946# a_n2129_43609# 7.7e-19
C9020 a_18287_44626# a_19268_43646# 6.61e-20
C9021 a_18443_44721# a_15743_43084# 1.36e-21
C9022 a_8746_45002# a_10210_45822# 0.013725f
C9023 a_10193_42453# a_10907_45822# 6.45e-20
C9024 a_8568_45546# a_8697_45572# 0.010132f
C9025 a_8162_45546# a_8791_45572# 6.1e-19
C9026 a_2711_45572# a_16020_45572# 0.006155f
C9027 a_7499_43078# a_8192_45572# 9.59e-19
C9028 C0_dummy_P_btm C3_P_btm 0.087354f
C9029 C3_N_btm C8_P_btm 5.08e-19
C9030 C2_N_btm C7_P_btm 1.06e-19
C9031 C1_N_btm C6_P_btm 1.76e-19
C9032 C0_N_btm C5_P_btm 7.74e-20
C9033 C0_dummy_N_btm C4_P_btm 6.85e-20
C9034 C10_N_btm EN_VIN_BSTR_N 0.320569f
C9035 C0_P_btm C2_P_btm 0.827449f
C9036 a_12379_42858# a_12465_44636# 4.6e-19
C9037 a_18817_42826# a_16327_47482# 0.215236f
C9038 a_n2661_43922# a_n863_45724# 0.115404f
C9039 a_7640_43914# a_n443_42852# 4e-21
C9040 a_10949_43914# a_8199_44636# 4.16e-20
C9041 a_743_42282# a_n2293_46634# 4.23e-20
C9042 a_18533_43940# a_17339_46660# 0.006189f
C9043 a_13678_32519# a_21588_30879# 0.056847f
C9044 a_4958_30871# a_n4064_37984# 0.030919f
C9045 a_6123_31319# VDAC_N 0.006993f
C9046 a_3483_46348# a_3699_46348# 0.06281f
C9047 a_19692_46634# a_8049_45260# 0.045516f
C9048 a_11901_46660# a_12839_46116# 3.72e-20
C9049 a_5257_43370# a_n357_42282# 3.28e-19
C9050 a_11415_45002# a_14275_46494# 1.84e-19
C9051 a_12741_44636# a_13759_46122# 1e-20
C9052 a_1823_45246# a_5497_46414# 1.22e-20
C9053 a_20528_46660# a_20075_46420# 4.61e-19
C9054 a_18280_46660# a_17957_46116# 1.49e-19
C9055 a_21363_46634# a_21137_46414# 0.001902f
C9056 a_20623_46660# a_6945_45028# 0.004994f
C9057 a_20273_46660# a_10809_44734# 0.027345f
C9058 a_11341_43940# a_22223_43396# 0.00507f
C9059 a_14401_32519# a_10341_43396# 0.133035f
C9060 a_22223_43948# a_5649_42852# 3.06e-19
C9061 a_19862_44208# a_20749_43396# 0.008749f
C9062 a_n2661_42282# a_2905_42968# 1.83e-20
C9063 a_n356_44636# a_564_42282# 9.95e-19
C9064 a_4223_44672# a_6123_31319# 4.56e-21
C9065 a_1568_43370# a_2437_43396# 7.56e-20
C9066 a_5343_44458# a_6773_42558# 4.65e-20
C9067 a_15493_43940# a_13678_32519# 7.99e-22
C9068 a_n1741_47186# DATA[3] 0.033504f
C9069 w_11334_34010# VIN_N 2.57e-20
C9070 a_n815_47178# DATA[0] 0.068508f
C9071 a_n913_45002# en_comp 7.44e-20
C9072 a_n2293_45010# a_n467_45028# 5.33e-20
C9073 a_n2661_45010# a_n37_45144# 6.21e-20
C9074 a_n1059_45260# a_n967_45348# 0.081574f
C9075 a_16147_45260# a_1307_43914# 0.150161f
C9076 a_6598_45938# a_n2661_44458# 5.14e-21
C9077 a_n13_43084# a_1138_42852# 3.75e-20
C9078 a_5755_42308# a_n2293_46634# 2.62e-20
C9079 a_16877_43172# a_6755_46942# 2.09e-19
C9080 a_n2129_43609# a_n755_45592# 0.001714f
C9081 a_n447_43370# a_n863_45724# 7e-19
C9082 a_n2267_43396# a_n357_42282# 8.73e-20
C9083 a_n4209_38216# SMPL_ON_P 8.15e-19
C9084 a_3422_30871# CAL_P 0.083836f
C9085 a_n2661_45546# VDD 0.733118f
C9086 a_10210_45822# a_4883_46098# 6.13e-19
C9087 a_15903_45785# a_11599_46634# 0.00101f
C9088 a_11064_45572# a_10227_46804# 6.09e-20
C9089 a_16855_45546# a_12861_44030# 4.91e-19
C9090 a_9049_44484# a_n881_46662# 4.56e-21
C9091 a_6472_45840# a_5807_45002# 0.016039f
C9092 a_526_44458# a_3218_45724# 0.032949f
C9093 a_8049_45260# a_20692_30879# 5.54e-20
C9094 a_10807_43548# a_12563_42308# 4.73e-21
C9095 a_21381_43940# a_20753_42852# 2.35e-19
C9096 a_n97_42460# a_16877_42852# 0.011527f
C9097 a_n2840_42826# a_n2472_42826# 7.52e-19
C9098 a_11750_44172# a_11633_42558# 6.73e-22
C9099 a_14853_42852# VDD 0.004079f
C9100 a_18341_45572# a_19279_43940# 1.85e-20
C9101 a_13777_45326# a_13720_44458# 1.97e-19
C9102 a_16922_45042# a_17613_45144# 0.10967f
C9103 a_1423_45028# a_6298_44484# 0.103777f
C9104 a_1307_43914# a_10334_44484# 3.55e-20
C9105 a_9482_43914# a_16112_44458# 3.24e-19
C9106 a_13556_45296# a_15004_44636# 0.127354f
C9107 a_7499_43078# a_8018_44260# 9.13e-21
C9108 a_2711_45572# a_21115_43940# 7.44e-20
C9109 a_n2293_45010# a_n2661_43922# 0.030818f
C9110 a_n2472_45002# a_n2293_43922# 7.11e-20
C9111 COMP_P a_n2956_39304# 8.08e-19
C9112 a_n4318_37592# a_n2956_38680# 0.02321f
C9113 a_21671_42860# a_n357_42282# 0.001708f
C9114 a_8685_42308# a_4185_45028# 6.95e-20
C9115 a_11823_42460# a_11415_45002# 0.349238f
C9116 a_6511_45714# a_3483_46348# 8.76e-21
C9117 a_1990_45572# a_1823_45246# 0.001177f
C9118 a_16147_45260# a_17609_46634# 2.56e-21
C9119 a_18691_45572# a_3090_45724# 3.57e-19
C9120 a_16019_45002# a_n743_46660# 0.002622f
C9121 a_n2293_42834# a_768_44030# 0.036156f
C9122 a_15297_45822# a_13059_46348# 0.002837f
C9123 a_626_44172# a_n2293_46634# 0.005771f
C9124 a_3357_43084# a_6755_46942# 6.8e-20
C9125 a_413_45260# a_5907_46634# 1.96e-20
C9126 a_3429_45260# a_3877_44458# 0.02987f
C9127 a_2711_45572# a_5204_45822# 0.021829f
C9128 a_18911_45144# a_11453_44696# 4.04e-19
C9129 a_11827_44484# a_13507_46334# 0.384415f
C9130 a_10440_44484# a_4791_45118# 1.07e-20
C9131 a_4361_42308# a_11633_42558# 4.09e-20
C9132 a_17499_43370# a_17303_42282# 4.37e-20
C9133 a_16823_43084# a_15803_42450# 0.008769f
C9134 a_5649_42852# a_11323_42473# 5.44e-20
C9135 a_16137_43396# a_18214_42558# 0.0459f
C9136 a_13678_32519# a_5742_30871# 0.004679f
C9137 a_20922_43172# a_20836_43172# 0.001377f
C9138 a_1847_42826# a_3905_42558# 1.42e-20
C9139 a_5534_30871# COMP_P 0.027557f
C9140 a_743_42282# a_13249_42558# 0.001357f
C9141 a_20205_31679# a_22609_37990# 9e-21
C9142 a_3422_30871# CAL_N 0.236929f
C9143 a_n785_47204# a_n2661_46098# 3.17e-20
C9144 a_4791_45118# a_n743_46660# 0.080217f
C9145 a_n1151_42308# a_383_46660# 0.002404f
C9146 a_n237_47217# a_2609_46660# 4.06e-20
C9147 a_n971_45724# a_2959_46660# 2.33e-19
C9148 a_584_46384# a_491_47026# 5.54e-20
C9149 a_4883_46098# a_5063_47570# 2.16e-22
C9150 a_13487_47204# a_5807_45002# 5.04e-20
C9151 a_13717_47436# a_13747_46662# 0.003701f
C9152 a_6851_47204# a_n2661_46634# 9.8e-20
C9153 a_4915_47217# a_n1925_46634# 1.12e-19
C9154 a_12861_44030# a_13661_43548# 0.8566f
C9155 a_10227_46804# a_11309_47204# 0.026748f
C9156 a_16327_47482# a_16119_47582# 1.79e-19
C9157 a_16023_47582# a_15928_47570# 0.049827f
C9158 a_16588_47582# a_12549_44172# 2.25e-20
C9159 en_comp a_n4318_39304# 1.82e-19
C9160 a_7229_43940# a_7499_43940# 6.92e-19
C9161 a_n2017_45002# a_n1177_43370# 4.91e-19
C9162 a_2437_43646# a_1756_43548# 8.79e-19
C9163 a_n2661_45010# a_104_43370# 1.69e-20
C9164 a_n2293_45010# a_n447_43370# 1.3e-19
C9165 a_n310_44484# a_n2661_42834# 9.37e-20
C9166 a_14537_43396# a_15037_44260# 0.001968f
C9167 a_9313_44734# a_n2661_43922# 0.028486f
C9168 a_10193_42453# a_16823_43084# 0.03411f
C9169 a_n2661_43370# a_8333_44056# 5.2e-21
C9170 a_n2661_44458# a_n1899_43946# 3.15e-20
C9171 a_16979_44734# a_11967_42832# 3.65e-19
C9172 a_n2433_44484# a_n1761_44111# 7.96e-20
C9173 a_n2129_44697# a_n2065_43946# 7.26e-19
C9174 a_7174_31319# a_n443_42852# 4.88e-21
C9175 a_15682_43940# a_16327_47482# 0.002941f
C9176 a_10807_43548# a_10227_46804# 0.025916f
C9177 a_19862_44208# a_12861_44030# 0.721035f
C9178 a_8487_44056# a_n971_45724# 2.58e-21
C9179 a_17034_45572# a_13259_45724# 0.002067f
C9180 a_3357_43084# a_8049_45260# 0.08902f
C9181 a_n967_45348# a_n1925_42282# 0.004046f
C9182 a_13556_45296# a_13759_46122# 1.81e-20
C9183 a_9482_43914# a_13925_46122# 1.87e-19
C9184 a_11787_45002# a_2324_44458# 0.002598f
C9185 a_1423_45028# a_5937_45572# 0.083936f
C9186 a_1307_43914# a_9290_44172# 0.122831f
C9187 a_5105_45348# a_5164_46348# 6.6e-20
C9188 a_1115_44172# a_768_44030# 0.003218f
C9189 a_16321_45348# a_11415_45002# 0.001041f
C9190 a_n2661_43370# a_n1991_46122# 8.66e-21
C9191 a_2809_45028# a_2804_46116# 6.45e-21
C9192 a_8325_42308# a_9293_42558# 7.62e-20
C9193 a_6123_31319# a_5742_30871# 0.106954f
C9194 a_8791_42308# a_9223_42460# 0.014257f
C9195 C8_P_btm C7_P_btm 31.072699f
C9196 C9_P_btm C6_P_btm 0.165353f
C9197 C10_P_btm C5_P_btm 0.51798f
C9198 a_n743_46660# a_16292_46812# 0.064277f
C9199 a_5807_45002# a_14513_46634# 0.006821f
C9200 a_13747_46662# a_14035_46660# 0.040628f
C9201 a_3877_44458# a_6755_46942# 0.388535f
C9202 a_5263_46660# a_5257_43370# 2.87e-20
C9203 a_13759_47204# a_13059_46348# 1.99e-19
C9204 a_12549_44172# a_14447_46660# 9.1e-20
C9205 a_11453_44696# a_22591_46660# 7.09e-19
C9206 SMPL_ON_N a_20820_30879# 0.029764f
C9207 a_12465_44636# a_21076_30879# 2.7e-19
C9208 a_4883_46098# a_21542_46660# 5.31e-19
C9209 a_12861_44030# a_4185_45028# 2.17e-20
C9210 a_6151_47436# a_9625_46129# 2.77e-19
C9211 a_7903_47542# a_8016_46348# 1.87e-20
C9212 a_6575_47204# a_7920_46348# 3.65e-19
C9213 a_n2833_47464# a_n2956_38680# 1.71e-20
C9214 a_n2497_47436# a_n2956_39304# 2.52e-20
C9215 a_n1151_42308# a_13351_46090# 5.07e-20
C9216 a_n1741_47186# a_6945_45028# 2.51584f
C9217 a_17613_45144# a_15743_43084# 1.82e-22
C9218 a_18587_45118# a_18429_43548# 1.57e-21
C9219 a_20512_43084# a_11341_43940# 0.02996f
C9220 a_5663_43940# a_6101_44260# 0.013015f
C9221 a_n356_44636# a_n1557_42282# 0.017569f
C9222 a_5495_43940# a_n2661_42282# 0.003301f
C9223 a_375_42282# a_421_43172# 0.00164f
C9224 a_13249_42308# a_1606_42308# 1.12e-20
C9225 a_n913_45002# a_22165_42308# 0.074472f
C9226 en_comp a_20922_43172# 3.26e-22
C9227 a_n4209_38502# C6_P_btm 0.001141f
C9228 a_n3565_38502# C8_P_btm 1.65e-20
C9229 a_n3565_38216# a_n1838_35608# 1.01e-19
C9230 a_n4209_38216# a_n1532_35090# 1.2e-19
C9231 a_22469_40625# a_20692_30879# 2.12e-20
C9232 a_6194_45824# a_6667_45809# 7.99e-20
C9233 a_6472_45840# a_6511_45714# 0.781352f
C9234 a_4099_45572# a_3775_45552# 0.003943f
C9235 a_5244_44056# a_n2293_46098# 6.1e-19
C9236 a_2813_43396# a_n2293_46634# 8.36e-19
C9237 a_7499_43940# a_8270_45546# 5.55e-20
C9238 a_18533_44260# a_6755_46942# 9.89e-21
C9239 a_n2661_44458# a_1848_45724# 3.76e-22
C9240 a_n2129_44697# a_n755_45592# 9.75e-19
C9241 a_n452_44636# a_n863_45724# 0.01836f
C9242 a_949_44458# a_n2293_45546# 0.004678f
C9243 a_n699_43396# a_n2661_45546# 0.022358f
C9244 a_16979_44734# a_13259_45724# 3.78e-21
C9245 a_743_42282# a_18597_46090# 3.54e-19
C9246 a_5342_30871# w_11334_34010# 0.00275f
C9247 a_n4209_38502# a_n3690_38528# 0.045251f
C9248 a_n3420_39072# a_n4334_38304# 2.34e-19
C9249 a_n4334_38528# a_n3565_38502# 2e-19
C9250 a_5385_46902# VDD 0.203316f
C9251 a_4958_30871# C0_P_btm 9.29e-20
C9252 a_765_45546# a_376_46348# 1.21e-19
C9253 a_5807_45002# a_n357_42282# 6.44e-20
C9254 a_n2956_39768# a_n2840_45546# 7e-20
C9255 a_13607_46688# a_13759_46122# 0.004856f
C9256 a_11813_46116# a_2324_44458# 1.71e-20
C9257 a_n2810_45028# a_n2302_40160# 0.001344f
C9258 a_n2956_37592# a_n4064_40160# 0.012264f
C9259 a_n4318_39304# a_n1699_43638# 8.9e-20
C9260 a_1307_43914# a_15051_42282# 1.26e-20
C9261 a_n2293_42834# a_6123_31319# 4.85e-19
C9262 a_n2433_43396# a_n2267_43396# 0.756435f
C9263 a_15682_43940# a_10341_43396# 3.89e-19
C9264 a_n2472_43914# a_n2472_42826# 0.001034f
C9265 a_11823_42460# a_13159_45002# 7.87e-19
C9266 a_12791_45546# a_13017_45260# 3.34e-19
C9267 a_2711_45572# a_6945_45348# 9.26e-20
C9268 a_18909_45814# a_19365_45572# 4.2e-19
C9269 a_10729_43914# a_n443_42852# 1.44e-20
C9270 a_19478_44306# a_n357_42282# 2.51e-20
C9271 a_n1917_43396# a_n1925_42282# 2.35e-19
C9272 a_10651_43940# a_10586_45546# 6.43e-22
C9273 a_3626_43646# a_17715_44484# 3.08e-21
C9274 a_9396_43370# a_9290_44172# 5.85e-20
C9275 a_3935_42891# a_3090_45724# 5.91e-20
C9276 a_16759_43396# a_12741_44636# 1.39e-19
C9277 a_13667_43396# a_3483_46348# 1.35e-19
C9278 a_22469_40625# VIN_N 2.79e-20
C9279 a_n1533_46116# VDD 0.143145f
C9280 a_7230_45938# a_6151_47436# 1.1e-20
C9281 a_6812_45938# a_6545_47178# 1.37e-19
C9282 a_11525_45546# a_n1151_42308# 2.76e-20
C9283 a_3483_46348# a_n755_45592# 5.99e-19
C9284 a_n1853_46287# a_n310_45572# 2.88e-19
C9285 a_14275_46494# a_13259_45724# 2.55e-19
C9286 a_6945_45028# a_10586_45546# 3.78e-20
C9287 a_6031_43396# a_7227_42852# 1.51e-19
C9288 a_15743_43084# a_19700_43370# 0.004331f
C9289 a_10341_43396# a_22223_43396# 0.038582f
C9290 a_6293_42852# a_5755_42852# 0.114235f
C9291 a_n97_42460# a_18817_42826# 0.003814f
C9292 a_3626_43646# a_10083_42826# 9.29e-20
C9293 a_2982_43646# a_10835_43094# 2.09e-20
C9294 a_16137_43396# a_16823_43084# 0.038492f
C9295 a_n2661_42282# a_n784_42308# 0.062364f
C9296 a_12281_43396# a_4361_42308# 0.021275f
C9297 a_16409_43396# a_17486_43762# 1.46e-19
C9298 a_n743_46660# DATA[3] 1.69e-21
C9299 a_171_46873# DATA[0] 9.78e-20
C9300 a_17701_42308# VDD 0.243354f
C9301 a_n2956_37592# a_n4064_37440# 0.070596f
C9302 a_n2810_45028# a_n2302_37690# 0.162246f
C9303 a_n2661_45010# a_949_44458# 0.071688f
C9304 a_n2293_45010# a_n452_44636# 3.23e-20
C9305 en_comp a_n2661_44458# 0.030481f
C9306 a_10193_42453# a_19279_43940# 4.41e-19
C9307 a_14537_43396# a_14976_45348# 9.13e-19
C9308 a_375_42282# a_n2661_43370# 0.012518f
C9309 a_9482_43914# a_13807_45067# 0.00608f
C9310 a_11823_42460# a_11967_42832# 0.573139f
C9311 a_n1641_43230# a_n863_45724# 2.33e-21
C9312 a_13003_42852# a_9290_44172# 7.01e-20
C9313 a_13157_43218# a_10903_43370# 6.01e-19
C9314 a_5111_44636# a_n1613_43370# 0.601769f
C9315 a_13348_45260# a_11453_44696# 0.005514f
C9316 a_14180_45002# a_12465_44636# 0.015526f
C9317 a_15595_45028# a_13507_46334# 1.41e-20
C9318 a_413_45260# a_768_44030# 0.182253f
C9319 a_n913_45002# a_13661_43548# 6.88e-20
C9320 a_5147_45002# a_n881_46662# 3.9e-19
C9321 a_10490_45724# a_3090_45724# 1.78e-21
C9322 a_11823_42460# a_12251_46660# 2.92e-20
C9323 a_3626_43646# a_15761_42308# 1.94e-19
C9324 a_4190_30871# COMP_P 0.027242f
C9325 a_8387_43230# a_8495_42852# 0.057222f
C9326 a_9127_43156# a_9306_43218# 0.007399f
C9327 a_8952_43230# a_9061_43230# 0.007416f
C9328 a_14209_32519# a_14097_32519# 10.7606f
C9329 a_21356_42826# a_21671_42860# 0.084365f
C9330 a_13759_46122# RST_Z 8.63e-20
C9331 a_21613_42308# VDD 0.273985f
C9332 a_n2109_47186# a_n881_46662# 0.023562f
C9333 a_n971_45724# a_2266_47243# 0.00941f
C9334 a_n785_47204# a_n310_47243# 0.001173f
C9335 a_1209_47178# a_2487_47570# 2.94e-19
C9336 a_13717_47436# a_11599_46634# 3.05e-19
C9337 a_12861_44030# a_14955_47212# 6.92e-20
C9338 a_13487_47204# a_14311_47204# 0.00114f
C9339 a_18184_42460# a_17517_44484# 0.020871f
C9340 a_18248_44752# a_18287_44626# 0.633819f
C9341 a_6298_44484# a_6109_44484# 0.068396f
C9342 a_5343_44458# a_8375_44464# 0.007376f
C9343 a_1307_43914# a_3905_42865# 0.224019f
C9344 a_n2661_44458# a_10617_44484# 0.003557f
C9345 a_17970_44736# a_18443_44721# 7.99e-20
C9346 a_7499_43078# a_6452_43396# 1.51e-20
C9347 a_1423_45028# a_2479_44172# 3.74e-20
C9348 a_11827_44484# a_13296_44484# 6.45e-19
C9349 a_3537_45260# a_9028_43914# 1.3e-19
C9350 a_n913_45002# a_19862_44208# 3.9e-20
C9351 a_3232_43370# a_6101_44260# 0.001648f
C9352 a_5932_42308# a_n443_42852# 4.07e-19
C9353 a_9223_42460# a_n357_42282# 3.69e-20
C9354 a_n4209_39304# a_n2956_39304# 0.328727f
C9355 a_8791_42308# a_n755_45592# 7.02e-19
C9356 a_13657_42308# a_13259_45724# 6.47e-20
C9357 a_11136_45572# VDD 0.004463f
C9358 a_6298_44484# a_4646_46812# 1.65052f
C9359 a_413_45260# a_1176_45822# 3.98e-20
C9360 a_5111_44636# a_n2293_46098# 0.086926f
C9361 a_n913_45002# a_4185_45028# 0.855072f
C9362 a_13468_44734# a_768_44030# 0.001477f
C9363 a_11823_42460# a_13259_45724# 0.626941f
C9364 a_3175_45822# a_3316_45546# 0.05019f
C9365 a_2711_45572# a_3503_45724# 0.058013f
C9366 a_8696_44636# a_526_44458# 5.2e-21
C9367 a_9159_45572# a_8049_45260# 1.83e-19
C9368 a_11280_45822# a_10586_45546# 1.28e-20
C9369 a_19256_45572# a_19553_46090# 1.97e-19
C9370 a_17668_45572# a_17583_46090# 5.29e-21
C9371 a_19431_45546# a_19335_46494# 0.002697f
C9372 a_18799_45938# a_18819_46122# 2.22e-19
C9373 a_18175_45572# a_6945_45028# 3.9e-21
C9374 a_17568_45572# a_17715_44484# 0.001302f
C9375 a_2437_43646# a_9823_46155# 1.23e-20
C9376 a_3357_43084# a_8953_45546# 2.47e-20
C9377 a_20512_43084# a_16327_47482# 0.118893f
C9378 a_7542_44172# a_n1151_42308# 2.32e-19
C9379 a_n2661_42282# SMPL_ON_P 0.003852f
C9380 a_5244_44056# a_4791_45118# 0.003487f
C9381 a_1606_42308# a_2123_42473# 0.011716f
C9382 a_1576_42282# a_2713_42308# 1.15e-20
C9383 a_14635_42282# a_13657_42558# 4.38e-21
C9384 a_13291_42460# a_14113_42308# 0.025652f
C9385 a_1184_42692# a_2725_42558# 1.23e-20
C9386 a_n2661_46634# a_4651_46660# 0.020633f
C9387 a_2107_46812# a_n2661_46098# 0.037509f
C9388 a_1983_46706# a_1799_45572# 0.089984f
C9389 a_948_46660# a_2443_46660# 4.94e-20
C9390 a_n743_46660# a_1057_46660# 9.22e-19
C9391 a_1123_46634# a_2609_46660# 3.37e-20
C9392 a_n2293_46634# a_3221_46660# 2.47e-21
C9393 a_n1925_46634# a_2162_46660# 4.85e-19
C9394 a_5807_45002# a_5263_46660# 1.75e-19
C9395 a_11309_47204# a_10467_46802# 0.023291f
C9396 a_9804_47204# a_10249_46116# 0.034717f
C9397 a_8128_46384# a_6755_46942# 0.01823f
C9398 a_n1613_43370# a_6086_46660# 0.001965f
C9399 SMPL_ON_P a_n2840_46090# 7.81e-19
C9400 a_n2109_47186# a_n2157_46122# 1.26e-21
C9401 a_n2497_47436# a_n1991_46122# 0.037858f
C9402 a_12861_44030# a_14543_46987# 6.49e-19
C9403 a_13381_47204# a_13059_46348# 3.39e-21
C9404 a_6851_47204# a_765_45546# 0.006814f
C9405 a_10227_46804# a_12156_46660# 0.025653f
C9406 a_19386_47436# a_19333_46634# 0.001224f
C9407 a_18597_46090# a_19466_46812# 0.074092f
C9408 a_11599_46634# a_14035_46660# 0.021792f
C9409 a_13507_46334# a_15559_46634# 0.216791f
C9410 a_4883_46098# a_14976_45028# 0.019383f
C9411 a_12465_44636# a_15009_46634# 2.01e-20
C9412 en_comp a_17364_32525# 8.05e-20
C9413 a_n2293_45010# a_n1641_43230# 2.03e-19
C9414 a_n1059_45260# a_n1853_43023# 0.03561f
C9415 a_n913_45002# a_n2157_42858# 0.00135f
C9416 a_n2017_45002# a_n1991_42858# 0.053113f
C9417 a_14537_43396# a_16547_43609# 2.37e-20
C9418 a_10057_43914# a_10555_43940# 0.001842f
C9419 a_n2840_43914# a_n1761_44111# 1.61e-20
C9420 a_n2472_43914# a_n2065_43946# 0.039807f
C9421 a_n2267_44484# a_n2433_43396# 0.00138f
C9422 a_n2433_44484# a_n2267_43396# 2.4e-19
C9423 a_n2129_44697# a_n2129_43609# 9.9e-19
C9424 a_3754_38470# VDD 2.52245f
C9425 a_22465_38105# a_22521_40055# 0.214039f
C9426 a_14579_43548# a_12861_44030# 1.6e-20
C9427 a_1423_45028# a_n443_42852# 1.15e-19
C9428 a_5891_43370# a_8016_46348# 0.183035f
C9429 a_17767_44458# a_17715_44484# 0.07408f
C9430 a_7640_43914# a_8199_44636# 0.003096f
C9431 a_6109_44484# a_5937_45572# 0.163331f
C9432 a_10157_44484# a_10809_44734# 3.6e-19
C9433 a_15037_43940# a_n2293_46634# 0.001262f
C9434 a_6453_43914# a_3090_45724# 0.00316f
C9435 a_17517_44484# a_12741_44636# 0.01998f
C9436 a_5608_44484# a_3483_46348# 0.001851f
C9437 a_n2293_43922# a_1823_45246# 1.33e-19
C9438 a_3363_44484# a_3699_46348# 1.94e-21
C9439 a_9049_44484# DATA[4] 1.59e-19
C9440 a_12891_46348# VDD 1.01428f
C9441 a_n4064_40160# a_n4251_40480# 0.00119f
C9442 a_7174_31319# a_1736_39587# 1.22e-19
C9443 a_n4315_30879# a_n4209_39590# 4.31257f
C9444 a_1606_42308# C3_N_btm 5.68e-19
C9445 a_15227_44166# a_20107_46660# 4.52e-19
C9446 a_18834_46812# a_20411_46873# 4.86e-22
C9447 a_14180_46812# a_14543_46987# 0.005265f
C9448 a_19333_46634# a_19551_46910# 0.08213f
C9449 a_19466_46812# a_19123_46287# 0.007907f
C9450 a_13885_46660# a_15227_46910# 1.69e-19
C9451 a_17609_46634# a_20273_46660# 3.59e-21
C9452 a_19692_46634# a_18285_46348# 5.98e-20
C9453 a_n2293_46634# a_n2956_38680# 1.99e-19
C9454 a_n2104_46634# a_n2956_39304# 6.41e-19
C9455 a_9804_47204# a_8781_46436# 1.48e-20
C9456 a_8128_46384# a_8049_45260# 0.00208f
C9457 a_n881_46662# a_8062_46155# 1.93e-19
C9458 a_4646_46812# a_5937_45572# 0.105447f
C9459 a_n743_46660# a_6945_45028# 0.029165f
C9460 a_5907_46634# a_6165_46155# 0.003895f
C9461 a_4883_46098# a_18051_46116# 0.003099f
C9462 a_13507_46334# a_20009_46494# 1.94e-19
C9463 a_18479_47436# a_20850_46155# 0.003424f
C9464 a_n443_46116# a_n89_45572# 0.006092f
C9465 a_15682_43940# a_n97_42460# 0.002081f
C9466 a_20935_43940# a_20974_43370# 0.005283f
C9467 a_11341_43940# a_21381_43940# 0.034147f
C9468 a_11967_42832# a_18429_43548# 0.019775f
C9469 a_18588_44850# a_18783_43370# 7.03e-21
C9470 a_n2661_42282# a_3080_42308# 0.161683f
C9471 a_20512_43084# a_10341_43396# 0.758407f
C9472 a_n356_44636# a_3935_42891# 2.82e-22
C9473 a_3737_43940# a_3992_43940# 0.005172f
C9474 a_n913_45002# a_9803_42558# 0.001906f
C9475 a_n2017_45002# a_9377_42558# 0.001128f
C9476 a_11750_44172# VDD 0.131662f
C9477 a_15903_45785# a_16855_45546# 9.79e-21
C9478 a_15599_45572# a_16680_45572# 0.102355f
C9479 a_15765_45572# a_16115_45572# 0.20669f
C9480 a_n97_42460# a_1823_45246# 0.006778f
C9481 a_15681_43442# a_15227_44166# 0.015868f
C9482 a_16547_43609# a_3090_45724# 3.84e-21
C9483 a_n809_44244# a_n863_45724# 0.016179f
C9484 a_10867_43940# a_9290_44172# 2.47e-19
C9485 a_12800_43218# a_12465_44636# 4.53e-20
C9486 a_n1630_35242# a_n1151_42308# 0.056434f
C9487 a_n4064_37984# C3_P_btm 0.030933f
C9488 a_18114_32519# a_22459_39145# 1.47e-20
C9489 a_19721_31679# a_22521_40055# 7.56e-21
C9490 a_11361_45348# CLK 3.72e-20
C9491 a_805_46414# VDD 0.154663f
C9492 a_7174_31319# CAL_N 0.018266f
C9493 a_n3420_38528# a_n4251_38304# 8.88e-19
C9494 a_n3420_39616# a_n4209_37414# 0.027966f
C9495 a_n4209_39590# a_n3420_37440# 0.038354f
C9496 a_n3565_39590# a_n3565_37414# 0.032079f
C9497 a_n4064_38528# a_n4064_37984# 0.057015f
C9498 a_4419_46090# a_n1925_42282# 0.056546f
C9499 C1_N_btm C3_N_btm 8.06688f
C9500 C0_dummy_N_btm C5_N_btm 0.11375f
C9501 C0_N_btm C4_N_btm 0.138331f
C9502 C0_dummy_P_btm C6_N_btm 1.37e-19
C9503 C1_P_btm C8_N_btm 4.41e-19
C9504 C0_P_btm C7_N_btm 2.32e-19
C9505 a_20411_46873# a_20850_46482# 9.61e-19
C9506 a_4704_46090# a_526_44458# 2.04e-19
C9507 a_11189_46129# a_6945_45028# 9.57e-21
C9508 a_2324_44458# a_15682_46116# 0.343876f
C9509 a_9313_44734# a_10545_42558# 6.42e-19
C9510 a_17730_32519# a_14097_32519# 0.053763f
C9511 a_n356_44636# a_15890_42674# 2.92e-19
C9512 a_n2293_43922# a_5934_30871# 0.079987f
C9513 a_19862_44208# a_20922_43172# 0.164553f
C9514 a_11341_43940# a_18249_42858# 4.65e-20
C9515 a_15493_43940# a_18083_42858# 1.12e-20
C9516 a_9145_43396# a_14358_43442# 0.053427f
C9517 a_1209_43370# a_743_42282# 3.61e-21
C9518 a_n2433_43396# a_n2472_42826# 9.53e-19
C9519 a_20269_44172# a_19987_42826# 8.09e-21
C9520 a_12465_44636# SINGLE_ENDED 0.067716f
C9521 a_22731_47423# RST_Z 4.82e-19
C9522 a_4361_42308# VDD 0.42717f
C9523 a_18175_45572# a_11827_44484# 1.29e-20
C9524 a_17668_45572# a_17613_45144# 5.67e-19
C9525 a_18799_45938# a_18911_45144# 4.07e-20
C9526 a_2711_45572# a_n2661_43922# 4.93e-20
C9527 a_2274_45254# a_2304_45348# 0.062682f
C9528 a_2680_45002# a_1423_45028# 0.003069f
C9529 a_6171_45002# a_14537_43396# 0.054973f
C9530 a_5147_45002# a_1307_43914# 0.032106f
C9531 a_2437_43646# a_n2661_43370# 0.033415f
C9532 a_22775_42308# a_21588_30879# 7.29e-21
C9533 a_n1853_43023# a_n1925_42282# 0.003483f
C9534 a_4181_43396# a_n443_42852# 1.39e-19
C9535 a_13635_43156# a_9290_44172# 0.394766f
C9536 a_12089_42308# a_10903_43370# 3.79e-19
C9537 a_20922_43172# a_4185_45028# 9.67e-21
C9538 a_15903_45785# a_13661_43548# 0.001692f
C9539 a_15599_45572# a_13747_46662# 0.041358f
C9540 a_15765_45572# a_5807_45002# 0.003059f
C9541 a_6194_45824# a_5257_43370# 0.029055f
C9542 a_6812_45938# a_3877_44458# 4.82e-21
C9543 a_4880_45572# a_4955_46873# 1.35e-20
C9544 a_8120_45572# a_n1925_46634# 0.004093f
C9545 a_12649_45572# a_12549_44172# 0.004247f
C9546 a_17786_45822# a_n881_46662# 4.61e-20
C9547 a_21350_45938# a_13507_46334# 2.55e-20
C9548 a_3357_43084# a_18780_47178# 2.77e-19
C9549 a_2437_43646# a_19787_47423# 0.006262f
C9550 a_19479_31679# a_18597_46090# 3e-20
C9551 a_413_45260# a_9067_47204# 4.35e-19
C9552 a_5205_44484# a_n1151_42308# 1.12e-20
C9553 a_5111_44636# a_4791_45118# 1.11355f
C9554 a_375_42282# a_n2497_47436# 0.018989f
C9555 a_n357_42282# a_n755_45592# 0.664842f
C9556 a_n2293_45546# a_n356_45724# 6.95e-20
C9557 a_310_45028# a_997_45618# 3.77e-20
C9558 a_n863_45724# a_3316_45546# 8.84e-21
C9559 a_4905_42826# a_5379_42460# 0.077171f
C9560 a_14209_32519# a_22959_42860# 0.007868f
C9561 a_n97_42460# a_5934_30871# 0.221607f
C9562 a_15493_43940# a_22775_42308# 6.96e-21
C9563 a_8605_42826# a_8952_43230# 0.051162f
C9564 a_8037_42858# a_10083_42826# 1.62e-19
C9565 a_3080_42308# a_3497_42558# 4.3e-19
C9566 a_20820_30879# a_18194_35068# 1.52e-19
C9567 a_n3420_37440# a_n4251_37440# 0.001432f
C9568 a_n4064_37440# a_n2860_37690# 0.003766f
C9569 a_3754_38470# a_8912_37509# 1.88278f
C9570 a_n3690_37440# a_n3607_37440# 0.007692f
C9571 a_7754_38470# a_6886_37412# 0.180842f
C9572 a_8530_39574# a_5700_37509# 0.947638f
C9573 a_6761_42308# VDD 0.259312f
C9574 a_n971_45724# a_n1151_42308# 0.682801f
C9575 a_1209_47178# a_584_46384# 0.104123f
C9576 a_n237_47217# a_2905_45572# 0.025329f
C9577 a_n1741_47186# a_4700_47436# 0.008526f
C9578 a_n2109_47186# a_n443_46116# 0.080373f
C9579 en_comp a_19237_31679# 1.18e-19
C9580 a_2437_43646# a_2998_44172# 1.59e-20
C9581 a_n2293_45010# a_n809_44244# 0.041966f
C9582 a_n2661_45010# a_175_44278# 6.99e-20
C9583 a_n1059_45260# a_n1899_43946# 5.95e-19
C9584 a_n913_45002# a_n1761_44111# 0.036392f
C9585 a_11827_44484# a_10440_44484# 1.55e-19
C9586 a_n2661_43370# a_4181_44734# 4.39e-19
C9587 a_7499_43078# a_11173_43940# 5.28e-20
C9588 a_n4318_40392# a_n1917_44484# 3.81e-20
C9589 a_17478_45572# a_17737_43940# 7.33e-21
C9590 a_14537_43396# a_14673_44172# 0.044194f
C9591 a_16922_45042# a_18287_44626# 1.76e-19
C9592 a_n2433_44484# a_n2267_44484# 0.730194f
C9593 a_n2661_44458# a_n1699_44726# 0.009008f
C9594 a_17719_45144# a_17767_44458# 0.001046f
C9595 a_20256_43172# a_n357_42282# 3.27e-19
C9596 a_n3674_38680# a_n2810_45572# 0.023027f
C9597 a_7174_31319# a_8199_44636# 4.88e-21
C9598 a_13904_45546# a_2324_44458# 0.004897f
C9599 a_10053_45546# a_6945_45028# 5.1e-22
C9600 a_10907_45822# a_11133_46155# 8.41e-19
C9601 a_9159_45572# a_8953_45546# 0.004909f
C9602 a_7499_43078# a_10809_44734# 0.053075f
C9603 a_11280_45822# a_11189_46129# 0.001906f
C9604 a_10306_45572# a_8199_44636# 5.75e-19
C9605 a_11682_45822# a_9290_44172# 0.00219f
C9606 a_n2661_43922# a_9313_45822# 3.03e-20
C9607 a_11827_44484# a_n743_46660# 2.74e-20
C9608 a_2779_44458# a_768_44030# 0.014949f
C9609 a_9482_43914# a_8270_45546# 0.004867f
C9610 a_7418_45067# a_4646_46812# 0.001853f
C9611 a_6171_45002# a_3090_45724# 0.030689f
C9612 a_2437_43646# a_20107_46660# 5.01e-21
C9613 a_3357_43084# a_18285_46348# 1.63e-20
C9614 a_8103_44636# a_8128_46384# 8.65e-21
C9615 a_16789_45572# a_11415_45002# 1.55e-19
C9616 a_5534_30871# a_13333_42558# 0.002157f
C9617 a_5342_30871# a_14456_42282# 0.160195f
C9618 a_n881_46662# a_n1925_46634# 0.467945f
C9619 a_n1613_43370# a_n1021_46688# 0.006304f
C9620 a_2747_46873# a_1983_46706# 3.11e-19
C9621 a_n1435_47204# a_7715_46873# 8.51e-20
C9622 a_6151_47436# a_6755_46942# 0.361724f
C9623 a_9313_45822# a_7927_46660# 9.18e-20
C9624 a_21359_45002# a_14021_43940# 5.71e-21
C9625 a_8701_44490# a_9028_43914# 0.008509f
C9626 a_17517_44484# a_20362_44736# 0.047565f
C9627 a_1307_43914# a_4093_43548# 0.002897f
C9628 a_5883_43914# a_8333_44056# 0.152643f
C9629 a_10193_42453# a_12545_42858# 8.12e-20
C9630 a_375_42282# a_1568_43370# 3.7e-21
C9631 a_5205_44484# a_6197_43396# 1.83e-19
C9632 a_7229_43940# a_6031_43396# 1.49e-19
C9633 a_5111_44636# a_8791_43396# 0.05316f
C9634 a_n913_45002# a_14579_43548# 0.239851f
C9635 a_n1059_45260# a_14358_43442# 1.98e-20
C9636 a_n2017_45002# a_14205_43396# 6.74e-21
C9637 a_3065_45002# a_3457_43396# 0.005043f
C9638 a_1606_42308# C7_P_btm 0.00238f
C9639 a_n2661_44458# a_4185_45028# 0.030414f
C9640 a_742_44458# a_1823_45246# 4.02e-19
C9641 a_949_44458# a_1138_42852# 0.013552f
C9642 a_14539_43914# a_11415_45002# 0.010769f
C9643 a_13720_44458# a_12741_44636# 0.00841f
C9644 a_18451_43940# a_13661_43548# 0.129334f
C9645 a_19328_44172# a_5807_45002# 7.07e-21
C9646 a_15493_43940# a_12549_44172# 0.932577f
C9647 a_14673_44172# a_3090_45724# 0.018197f
C9648 a_n2661_42282# a_n2438_43548# 4.44e-20
C9649 a_5105_45348# a_5066_45546# 1.87e-19
C9650 a_n2661_45010# a_n356_45724# 6.56e-21
C9651 a_n745_45366# a_n755_45592# 0.014023f
C9652 a_n143_45144# a_n2293_45546# 0.012062f
C9653 a_327_44734# a_n2661_45546# 7.19e-19
C9654 a_2437_43646# a_2307_45899# 4.14e-19
C9655 a_16922_45042# a_15682_46116# 6.61e-19
C9656 a_9420_43940# a_4883_46098# 0.001234f
C9657 a_21381_43940# a_16327_47482# 0.001197f
C9658 a_3626_43646# a_584_46384# 0.195961f
C9659 a_13070_42354# a_7174_31319# 4.88e-21
C9660 a_5932_42308# a_1736_39587# 1.46e-19
C9661 a_7903_47542# VDD 0.202868f
C9662 a_n2438_43548# a_n2840_46090# 0.002055f
C9663 a_n2661_46634# a_n1076_46494# 1.61e-20
C9664 a_n1021_46688# a_n2293_46098# 6.25e-19
C9665 a_n1925_46634# a_n2157_46122# 0.00977f
C9666 a_n2104_46634# a_n1991_46122# 2.68e-19
C9667 a_n2312_38680# a_n1853_46287# 3.4e-19
C9668 a_11186_47026# a_11813_46116# 2.23e-20
C9669 a_10467_46802# a_12156_46660# 3.88e-21
C9670 a_4651_46660# a_765_45546# 0.004164f
C9671 a_9804_47204# a_5937_45572# 5.55e-20
C9672 a_8128_46384# a_8953_45546# 5.55e-20
C9673 a_n1151_42308# a_12005_46436# 1.31e-20
C9674 a_2063_45854# a_11315_46155# 2.18e-19
C9675 a_20894_47436# a_10809_44734# 0.003478f
C9676 a_21177_47436# a_6945_45028# 0.008435f
C9677 a_13507_46334# a_21137_46414# 0.007257f
C9678 a_4883_46098# a_19900_46494# 0.008904f
C9679 a_6151_47436# a_8049_45260# 1.58e-19
C9680 a_11453_44696# a_17957_46116# 0.0084f
C9681 a_12465_44636# a_19335_46494# 6.74e-21
C9682 a_n1613_43370# a_9290_44172# 0.003987f
C9683 a_20512_43084# a_n97_42460# 2.54e-19
C9684 a_n1761_44111# a_n4318_39304# 3.05e-19
C9685 a_14539_43914# a_15037_43396# 8.32e-22
C9686 a_7542_44172# a_8415_44056# 2.49e-20
C9687 a_10405_44172# a_10555_44260# 0.085098f
C9688 a_10193_42453# a_19332_42282# 0.004163f
C9689 a_11967_42832# a_2982_43646# 5.64e-19
C9690 a_n356_44636# a_16547_43609# 3.88e-21
C9691 a_18443_44721# a_18783_43370# 1.12e-19
C9692 a_9313_44734# a_14955_43396# 0.001014f
C9693 a_19328_44172# a_19478_44306# 0.188181f
C9694 a_14955_43940# a_11341_43940# 0.005859f
C9695 a_n2065_43946# a_n2433_43396# 6.16e-19
C9696 a_18374_44850# a_18525_43370# 8.44e-21
C9697 a_18287_44626# a_15743_43084# 3.79e-20
C9698 a_11823_42460# a_15143_45578# 0.120787f
C9699 a_10193_42453# a_10210_45822# 0.026406f
C9700 a_8568_45546# a_8192_45572# 1.96e-19
C9701 a_8162_45546# a_8697_45572# 0.001108f
C9702 a_13527_45546# a_13904_45546# 3.21e-19
C9703 a_7499_43078# a_8120_45572# 1.34e-20
C9704 a_10180_45724# a_10907_45822# 6.72e-20
C9705 C0_dummy_P_btm C4_P_btm 0.113156f
C9706 C3_N_btm C9_P_btm 6.09e-19
C9707 C2_N_btm C8_P_btm 1.77e-19
C9708 C1_N_btm C7_P_btm 2.65e-19
C9709 C0_N_btm C6_P_btm 1.55e-19
C9710 C0_dummy_N_btm C5_P_btm 6.85e-20
C9711 C9_N_btm EN_VIN_BSTR_N 0.226529f
C9712 C1_P_btm C2_P_btm 5.24136f
C9713 C0_P_btm C3_P_btm 0.409238f
C9714 a_9672_43914# a_8953_45546# 1.03e-19
C9715 a_10729_43914# a_8199_44636# 3.27e-20
C9716 a_10807_43548# a_8016_46348# 1.5e-19
C9717 a_18249_42858# a_16327_47482# 0.315855f
C9718 a_21671_42860# a_12861_44030# 5.22e-22
C9719 a_19319_43548# a_17339_46660# 2.03e-19
C9720 a_3363_44484# a_n755_45592# 8.3e-21
C9721 a_n2661_42834# a_n863_45724# 0.094705f
C9722 a_n2661_43922# a_n1079_45724# 9.64e-21
C9723 a_17517_44484# a_16375_45002# 4.98e-19
C9724 a_n1899_43946# a_n1925_42282# 1.14e-19
C9725 a_6109_44484# a_n443_42852# 0.002868f
C9726 a_15493_43396# a_3483_46348# 1.59e-19
C9727 a_12359_47026# VDD 0.142103f
C9728 a_6123_31319# a_6886_37412# 4.22e-19
C9729 a_3147_46376# a_3699_46348# 0.001175f
C9730 a_19466_46812# a_8049_45260# 0.061209f
C9731 a_4646_46812# a_n443_42852# 0.038263f
C9732 a_11415_45002# a_14493_46090# 2.96e-20
C9733 a_12741_44636# a_13351_46090# 5.89e-22
C9734 a_1823_45246# a_5204_45822# 1.73e-19
C9735 a_20623_46660# a_21137_46414# 0.001102f
C9736 a_20841_46902# a_6945_45028# 0.013693f
C9737 a_20411_46873# a_10809_44734# 0.010692f
C9738 a_11341_43940# a_5649_42852# 0.01232f
C9739 a_15493_43940# a_21855_43396# 2.4e-19
C9740 a_14021_43940# a_16823_43084# 0.005626f
C9741 a_21381_43940# a_10341_43396# 0.03047f
C9742 a_4223_44672# a_7227_42308# 3.26e-37
C9743 a_n356_44636# a_n3674_37592# 4.6e-21
C9744 a_n97_42460# a_7221_43396# 1.23e-19
C9745 a_n1741_47186# DATA[2] 0.017604f
C9746 a_n1605_47204# DATA[0] 4.69e-19
C9747 a_7274_43762# VDD 4.6e-19
C9748 a_n2293_45010# a_n955_45028# 8.22e-21
C9749 a_n1059_45260# en_comp 8.56e-20
C9750 a_3357_43084# a_3065_45002# 0.316449f
C9751 a_n2661_45010# a_n143_45144# 5.24e-21
C9752 a_n2017_45002# a_n967_45348# 0.095287f
C9753 a_16147_45260# a_16019_45002# 0.186254f
C9754 a_6667_45809# a_n2661_44458# 6.66e-21
C9755 a_17364_32525# a_4185_45028# 0.046035f
C9756 a_n97_42460# a_n2293_45546# 2.89e-21
C9757 a_n1352_43396# a_n863_45724# 9.43e-21
C9758 a_n2433_43396# a_n755_45592# 5.17e-20
C9759 a_2982_43646# a_13259_45724# 0.06616f
C9760 a_n2129_43609# a_n357_42282# 0.001046f
C9761 a_743_42282# a_8953_45546# 0.032209f
C9762 a_18214_42558# a_13507_46334# 1.84e-19
C9763 a_20712_42282# a_18479_47436# 1.22e-20
C9764 a_13258_32519# a_18597_46090# 0.023292f
C9765 a_21125_42558# a_16327_47482# 5.5e-19
C9766 a_17517_44484# RST_Z 0.004664f
C9767 a_n2810_45572# VDD 0.557886f
C9768 a_15599_45572# a_11599_46634# 0.26676f
C9769 a_10544_45572# a_10227_46804# 0.00205f
C9770 a_2437_43646# a_n2497_47436# 0.027407f
C9771 a_6194_45824# a_5807_45002# 0.02442f
C9772 a_8049_45260# a_20205_31679# 0.301209f
C9773 a_526_44458# a_2957_45546# 1.97e-19
C9774 a_10807_43548# a_11633_42558# 8.38e-19
C9775 a_17538_32519# a_14097_32519# 0.050981f
C9776 a_n97_42460# a_16245_42852# 0.088473f
C9777 a_10341_43396# a_18249_42858# 9.84e-20
C9778 a_11750_44172# a_11551_42558# 8.92e-22
C9779 a_13622_42852# VDD 4.6e-19
C9780 a_13556_45296# a_13720_44458# 0.212774f
C9781 a_16922_45042# a_17023_45118# 0.099834f
C9782 a_1423_45028# a_5518_44484# 0.047243f
C9783 a_1307_43914# a_10157_44484# 6.43e-20
C9784 a_9482_43914# a_15004_44636# 0.34299f
C9785 a_7499_43078# a_7911_44260# 7.28e-19
C9786 a_18479_45785# a_19279_43940# 0.019159f
C9787 a_14537_43396# a_12607_44458# 1.38e-21
C9788 a_2711_45572# a_20935_43940# 1.09e-19
C9789 a_n2472_45002# a_n2661_43922# 6.45e-19
C9790 a_n2661_45010# a_n2293_43922# 2.75e-20
C9791 a_n2293_45010# a_n2661_42834# 0.083461f
C9792 a_3537_45260# a_5205_44734# 6.62e-22
C9793 a_6171_42473# a_5937_45572# 8.33e-22
C9794 a_n2293_42282# a_n863_45724# 0.028166f
C9795 a_15567_42826# a_n443_42852# 3.58e-19
C9796 a_n1736_42282# a_n2956_38680# 2.5e-20
C9797 a_21195_42852# a_n357_42282# 0.09377f
C9798 a_n4318_37592# a_n2956_39304# 0.023347f
C9799 a_8325_42308# a_4185_45028# 9.41e-20
C9800 a_12427_45724# a_11415_45002# 1.12e-20
C9801 a_6472_45840# a_3483_46348# 1.46e-20
C9802 a_3775_45552# a_167_45260# 1.19e-20
C9803 a_3733_45822# a_1823_45246# 0.003114f
C9804 a_18909_45814# a_3090_45724# 7.08e-19
C9805 a_15595_45028# a_n743_46660# 2.81e-20
C9806 a_15225_45822# a_13059_46348# 0.002175f
C9807 a_6517_45366# a_5807_45002# 5.73e-19
C9808 a_501_45348# a_n2293_46634# 1.32e-19
C9809 a_3065_45002# a_3877_44458# 0.287919f
C9810 a_3357_43084# a_10249_46116# 5.65e-20
C9811 a_413_45260# a_5167_46660# 1.29e-20
C9812 a_n913_45002# a_5257_43370# 9.26e-20
C9813 a_2711_45572# a_5164_46348# 0.031464f
C9814 a_21359_45002# a_13507_46334# 6.77e-19
C9815 a_20193_45348# a_18597_46090# 0.021804f
C9816 a_6298_44484# a_6545_47178# 2.86e-20
C9817 a_4181_44734# a_n2497_47436# 0.01129f
C9818 a_10334_44484# a_4791_45118# 1.31e-20
C9819 a_17499_43370# a_4958_30871# 0.001145f
C9820 a_3935_42891# a_3823_42558# 0.012124f
C9821 a_16823_43084# a_15764_42576# 0.0016f
C9822 a_12545_42858# a_n784_42308# 5.9e-21
C9823 a_5649_42852# a_10723_42308# 1.31e-19
C9824 a_4361_42308# a_11551_42558# 0.011423f
C9825 a_743_42282# a_14456_42282# 0.006738f
C9826 a_15743_43084# a_17124_42282# 1.95e-21
C9827 a_19987_42826# a_20836_43172# 1.48e-20
C9828 a_1847_42826# a_3581_42558# 2.17e-20
C9829 a_16137_43396# a_19332_42282# 2.66e-19
C9830 a_20692_30879# a_22609_38406# 4.83e-21
C9831 a_3422_30871# a_11206_38545# 1.36e-20
C9832 a_n971_45724# a_3177_46902# 0.001193f
C9833 a_584_46384# a_288_46660# 1.99e-21
C9834 a_n443_46116# a_n1925_46634# 0.080855f
C9835 a_2553_47502# a_2107_46812# 1.02e-21
C9836 a_n1151_42308# a_601_46902# 0.001897f
C9837 a_2063_45854# a_1983_46706# 0.001595f
C9838 a_n237_47217# a_2443_46660# 6.7e-20
C9839 a_10227_46804# a_11117_47542# 5.57e-20
C9840 a_12861_44030# a_5807_45002# 0.214011f
C9841 a_6491_46660# a_n2661_46634# 0.013828f
C9842 a_13717_47436# a_13661_43548# 2.13e-20
C9843 a_16327_47482# a_15928_47570# 0.001167f
C9844 a_16241_47178# a_16119_47582# 3.16e-19
C9845 a_16763_47508# a_12549_44172# 2.49e-19
C9846 a_n2956_37592# a_n4318_39304# 0.023222f
C9847 a_2437_43646# a_1568_43370# 0.058471f
C9848 a_n2017_45002# a_n1917_43396# 0.01343f
C9849 a_n2661_45010# a_n97_42460# 8.74e-21
C9850 a_n2293_45010# a_n1352_43396# 0.002774f
C9851 en_comp a_n2840_43370# 7.28e-20
C9852 a_n745_45366# a_n2129_43609# 6.64e-20
C9853 a_9241_44734# a_n2661_43922# 1.54e-35
C9854 a_9313_44734# a_n2661_42834# 0.02321f
C9855 a_n2661_44458# a_n1761_44111# 1.08e-19
C9856 a_14539_43914# a_11967_42832# 0.512158f
C9857 a_n2433_44484# a_n2065_43946# 0.008496f
C9858 a_15415_45028# a_14021_43940# 6.12e-21
C9859 a_n2946_39866# a_n2956_38216# 4.86e-20
C9860 a_20447_31679# VDD 0.665681f
C9861 a_1423_45028# a_8199_44636# 0.088277f
C9862 a_9482_43914# a_13759_46122# 1e-20
C9863 a_10951_45334# a_2324_44458# 0.002224f
C9864 a_13777_45326# a_12594_46348# 0.00118f
C9865 a_4640_45348# a_5164_46348# 1.3e-19
C9866 a_10949_43914# a_10227_46804# 2.49e-20
C9867 a_19478_44306# a_12861_44030# 2.84e-20
C9868 a_18315_45260# a_18280_46660# 4.34e-22
C9869 a_644_44056# a_768_44030# 0.177755f
C9870 a_16789_45572# a_13259_45724# 9.06e-19
C9871 a_19479_31679# a_8049_45260# 0.022565f
C9872 en_comp a_n1925_42282# 4.02e-19
C9873 a_413_45260# a_518_46482# 1.79e-21
C9874 a_14309_45028# a_11415_45002# 0.040538f
C9875 a_2809_45028# a_2698_46116# 2.22e-20
C9876 a_14097_32519# a_22465_38105# 0.002065f
C9877 a_5934_30871# a_10533_42308# 7.8e-20
C9878 a_7227_42308# a_5742_30871# 2.87e-20
C9879 a_8685_42308# a_9223_42460# 0.166964f
C9880 a_8325_42308# a_9803_42558# 5.62e-20
C9881 C9_P_btm C7_P_btm 0.22201f
C9882 C10_P_btm C6_P_btm 0.895671f
C9883 a_n743_46660# a_15559_46634# 2.71e-19
C9884 a_5807_45002# a_14180_46812# 0.007999f
C9885 a_13747_46662# a_13885_46660# 0.028801f
C9886 a_13675_47204# a_13059_46348# 8.27e-20
C9887 a_11453_44696# a_11415_45002# 0.123733f
C9888 SMPL_ON_N a_22591_46660# 0.011048f
C9889 a_22731_47423# a_20820_30879# 0.001051f
C9890 a_22223_47212# a_12741_44636# 7.08e-20
C9891 a_4883_46098# a_21297_46660# 1.2e-19
C9892 a_21811_47423# a_21076_30879# 1.63e-19
C9893 a_13487_47204# a_3483_46348# 4.28e-19
C9894 a_4915_47217# a_9823_46155# 1.19e-20
C9895 a_6151_47436# a_8953_45546# 8.27e-19
C9896 a_7903_47542# a_7920_46348# 2.96e-21
C9897 a_6545_47178# a_5937_45572# 1.49e-20
C9898 a_n1151_42308# a_12594_46348# 4.07e-19
C9899 a_n1435_47204# a_4419_46090# 1.69e-20
C9900 a_19279_43940# a_14021_43940# 2.21e-19
C9901 a_20512_43084# a_21115_43940# 1.49e-21
C9902 a_16922_45042# a_19268_43646# 1.77e-21
C9903 a_5663_43940# a_5841_44260# 0.007617f
C9904 a_5013_44260# a_n2661_42282# 1.85e-20
C9905 a_n356_44636# a_766_43646# 9.89e-19
C9906 a_375_42282# a_133_43172# 7.97e-20
C9907 a_n913_45002# a_21671_42860# 8.31e-20
C9908 en_comp a_19987_42826# 9.77e-21
C9909 a_5891_43370# VDD 2.12137f
C9910 a_n4209_38502# C7_P_btm 7.54e-20
C9911 a_n3565_38502# C9_P_btm 1.91e-20
C9912 a_n4209_38216# a_n1386_35608# 1.32e-19
C9913 a_22469_40625# a_20205_31679# 1.74e-20
C9914 a_22521_40599# a_20692_30879# 2.53e-20
C9915 a_6194_45824# a_6511_45714# 0.102325f
C9916 a_19237_31679# a_4185_45028# 0.004066f
C9917 a_3905_42865# a_n2293_46098# 0.237656f
C9918 a_9145_43396# a_13661_43548# 0.135139f
C9919 a_14539_43914# a_13259_45724# 0.002022f
C9920 a_742_44458# a_n2293_45546# 1.34e-19
C9921 a_4223_44672# a_n2661_45546# 0.041115f
C9922 a_n1352_44484# a_n863_45724# 1.83e-21
C9923 a_n2433_44484# a_n755_45592# 4.6e-21
C9924 a_17517_44484# a_18985_46122# 2.43e-21
C9925 a_12189_44484# a_10809_44734# 1.06e-19
C9926 a_20556_43646# a_18479_47436# 9.29e-19
C9927 a_5649_42852# a_16327_47482# 9.95e-20
C9928 a_5342_30871# w_1575_34946# 0.002142f
C9929 a_20447_31679# a_22469_39537# 5.38e-20
C9930 a_n4209_38502# a_n3565_38502# 6.84323f
C9931 a_n3565_39304# a_n3565_38216# 0.02823f
C9932 a_n3420_39072# a_n4209_38216# 0.030577f
C9933 a_4817_46660# VDD 0.370615f
C9934 a_4958_30871# C1_P_btm 9.46e-20
C9935 a_21188_46660# a_21297_46660# 0.007416f
C9936 a_21363_46634# a_21542_46660# 0.007399f
C9937 a_20731_47026# a_12741_44636# 8.49e-19
C9938 a_5072_46660# a_5066_45546# 3.51e-21
C9939 a_11735_46660# a_2324_44458# 1.17e-20
C9940 a_3090_45724# a_10903_43370# 0.031245f
C9941 a_n1630_35242# VDAC_Pi 1.06e-19
C9942 en_comp a_n4315_30879# 0.001378f
C9943 a_n2810_45028# a_n4064_40160# 0.001122f
C9944 a_n2956_37592# a_n4334_40480# 0.0011f
C9945 a_2382_45260# a_7174_31319# 4.88e-21
C9946 a_895_43940# a_743_42282# 2.08e-20
C9947 a_n4318_39304# a_n2267_43396# 4.55e-19
C9948 a_19721_31679# a_14097_32519# 0.051111f
C9949 a_10807_43548# a_12281_43396# 7.83e-20
C9950 a_n2293_42834# a_7227_42308# 7.22e-20
C9951 a_11341_43940# a_8685_43396# 2.48e-19
C9952 a_n2433_43396# a_n2129_43609# 0.283605f
C9953 a_14955_43940# a_10341_43396# 6.65e-21
C9954 a_18533_43940# VDD 0.182147f
C9955 a_11823_42460# a_13017_45260# 0.030503f
C9956 a_7499_43078# a_1307_43914# 0.109806f
C9957 a_11322_45546# a_13777_45326# 2.22e-21
C9958 a_18341_45572# a_19365_45572# 2.36e-20
C9959 a_18479_45785# a_19610_45572# 8.18e-19
C9960 a_n961_42308# a_n1613_43370# 0.0058f
C9961 a_13258_32519# w_11334_34010# 2.64e-19
C9962 a_19095_43396# a_17339_46660# 0.049229f
C9963 a_10405_44172# a_n443_42852# 7.35e-20
C9964 a_15493_43396# a_n357_42282# 9.67e-20
C9965 VDAC_P VCM 11.743501f
C9966 a_n722_46482# VDD 1.22e-19
C9967 a_2711_45572# a_15673_47210# 2.77e-20
C9968 a_6812_45938# a_6151_47436# 0.018338f
C9969 a_6977_45572# a_n971_45724# 4.78e-20
C9970 a_9049_44484# a_4791_45118# 0.009879f
C9971 a_11322_45546# a_n1151_42308# 0.001795f
C9972 a_11823_42460# a_2063_45854# 8.26e-19
C9973 a_1823_45246# a_3503_45724# 0.295715f
C9974 a_167_45260# a_3218_45724# 1.73e-19
C9975 a_1138_42852# a_n356_45724# 1.67e-20
C9976 a_3147_46376# a_n755_45592# 1.44e-19
C9977 a_3483_46348# a_n357_42282# 5.91e-21
C9978 a_n1925_42282# a_4365_46436# 0.009374f
C9979 a_14493_46090# a_13259_45724# 7.12e-20
C9980 a_14840_46494# a_14949_46494# 0.007416f
C9981 a_15015_46420# a_15194_46482# 0.007399f
C9982 a_14275_46494# a_14383_46116# 0.057222f
C9983 a_2324_44458# a_14537_46482# 2.56e-21
C9984 a_6031_43396# a_5755_42852# 4.17e-19
C9985 a_15743_43084# a_19268_43646# 0.010228f
C9986 a_10341_43396# a_5649_42852# 0.049047f
C9987 a_n97_42460# a_18249_42858# 0.003512f
C9988 a_3905_42865# a_3905_42558# 2.95e-19
C9989 a_3626_43646# a_8952_43230# 9.54e-21
C9990 a_2982_43646# a_10518_42984# 2.29e-20
C9991 a_n2661_42282# a_196_42282# 2.77e-19
C9992 a_16243_43396# a_16855_43396# 3.82e-19
C9993 a_n743_46660# DATA[2] 1.69e-21
C9994 a_n133_46660# DATA[0] 1.6e-19
C9995 a_n2438_43548# DATA[1] 5.69e-20
C9996 a_n2293_46634# CLK 1.2e-20
C9997 a_17595_43084# VDD 0.168112f
C9998 a_19479_31679# a_22469_40625# 1.34e-20
C9999 a_n2956_37592# a_n2946_37690# 0.148852f
C10000 a_n2810_45028# a_n4064_37440# 0.22413f
C10001 a_3357_43084# a_6298_44484# 3.5e-19
C10002 a_n913_45002# a_n2267_44484# 1.1e-19
C10003 en_comp a_n4318_40392# 3.37e-20
C10004 a_n2017_45002# a_n1917_44484# 0.012037f
C10005 a_n2661_45010# a_742_44458# 0.694478f
C10006 a_n2293_45010# a_n1352_44484# 0.020183f
C10007 a_n2956_37592# a_n2661_44458# 0.003435f
C10008 a_n745_45366# a_n2129_44697# 0.00194f
C10009 a_14537_43396# a_14403_45348# 2.86e-19
C10010 a_13348_45260# a_13807_45067# 6.64e-19
C10011 a_9482_43914# a_13490_45067# 0.007606f
C10012 a_n4318_38680# a_n2810_45572# 0.023234f
C10013 a_n1423_42826# a_n863_45724# 4.06e-21
C10014 a_12991_43230# a_10903_43370# 0.001102f
C10015 a_4558_45348# a_n881_46662# 3.03e-21
C10016 a_5147_45002# a_n1613_43370# 1.57e-20
C10017 a_13159_45002# a_11453_44696# 0.006266f
C10018 a_13777_45326# a_12465_44636# 4.66e-20
C10019 a_15415_45028# a_13507_46334# 1.22e-20
C10020 a_11823_42460# a_12469_46902# 2.61e-20
C10021 a_12791_45546# a_11901_46660# 8.23e-19
C10022 a_12427_45724# a_12251_46660# 1.4e-20
C10023 a_8746_45002# a_3090_45724# 1.22e-19
C10024 a_10193_42453# a_14976_45028# 1.31e-20
C10025 a_413_45260# a_12549_44172# 2.22e-19
C10026 a_n913_45002# a_5807_45002# 2.94e-20
C10027 a_n1059_45260# a_13661_43548# 0.004019f
C10028 a_20447_31679# a_22612_30879# 0.107874f
C10029 a_3626_43646# a_15521_42308# 3.81e-19
C10030 a_14209_32519# a_22400_42852# 8.65e-21
C10031 a_21356_42826# a_21195_42852# 0.03853f
C10032 a_8605_42826# a_8495_42852# 0.097745f
C10033 a_9625_46129# CLK 2.09e-20
C10034 a_21887_42336# VDD 0.210392f
C10035 a_n2109_47186# a_n1613_43370# 0.054203f
C10036 a_1209_47178# a_2266_47570# 9.52e-19
C10037 a_n971_45724# a_3315_47570# 3.15e-19
C10038 a_n1435_47204# a_11599_46634# 3.32e-20
C10039 a_13717_47436# a_14955_47212# 1.64e-19
C10040 a_12861_44030# a_14311_47204# 0.037394f
C10041 a_n1151_42308# a_12465_44636# 0.02014f
C10042 a_19778_44110# a_17517_44484# 0.018823f
C10043 a_5518_44484# a_6109_44484# 0.050093f
C10044 a_11691_44458# a_11541_44484# 0.037586f
C10045 a_17970_44736# a_18287_44626# 0.102355f
C10046 a_1307_43914# a_3600_43914# 0.153686f
C10047 a_5343_44458# a_7640_43914# 0.152634f
C10048 a_9049_44484# a_8791_43396# 1.63e-20
C10049 a_7499_43078# a_9396_43370# 2.11e-19
C10050 a_626_44172# a_895_43940# 0.038336f
C10051 a_13249_42308# a_3626_43646# 0.007551f
C10052 a_9482_43914# a_7845_44172# 5.64e-21
C10053 a_11827_44484# a_12829_44484# 2.53e-19
C10054 a_3537_45260# a_8333_44056# 0.012371f
C10055 a_3232_43370# a_5841_44260# 5.8e-19
C10056 a_6171_42473# a_n443_42852# 6.33e-20
C10057 a_8791_42308# a_n357_42282# 6.28e-20
C10058 a_8685_42308# a_n755_45592# 0.001582f
C10059 a_n2661_44458# a_5257_43370# 0.027109f
C10060 a_1423_45028# a_765_45546# 3.01e-22
C10061 a_5147_45002# a_n2293_46098# 0.211057f
C10062 a_5518_44484# a_4646_46812# 2.19e-19
C10063 a_13213_44734# a_768_44030# 0.00651f
C10064 a_n1059_45260# a_4185_45028# 0.027781f
C10065 a_13857_44734# a_12891_46348# 7.81e-20
C10066 a_327_44734# a_805_46414# 2.28e-19
C10067 a_9313_44734# a_19321_45002# 7.03e-21
C10068 a_10907_45822# a_10586_45546# 0.05477f
C10069 a_2711_45572# a_3316_45546# 0.065336f
C10070 a_3175_45822# a_3218_45724# 0.132424f
C10071 a_12427_45724# a_13259_45724# 6.07e-19
C10072 a_3260_45572# a_n2661_45546# 6.42e-20
C10073 a_19431_45546# a_19553_46090# 8.55e-19
C10074 a_19256_45572# a_18985_46122# 5.12e-19
C10075 a_2437_43646# a_9569_46155# 2.04e-20
C10076 a_3357_43084# a_5937_45572# 0.257963f
C10077 a_11967_42832# a_11453_44696# 6.13e-20
C10078 a_19279_43940# a_13507_46334# 1.3e-20
C10079 a_20980_44850# a_18479_47436# 0.002954f
C10080 a_3422_30871# a_10227_46804# 2.07e-19
C10081 a_21145_44484# a_16327_47482# 1.79e-19
C10082 a_3905_42865# a_4791_45118# 0.208831f
C10083 a_22959_42860# a_22465_38105# 9e-19
C10084 a_1606_42308# a_1755_42282# 0.278431f
C10085 a_n784_42308# a_5379_42460# 1.36e-19
C10086 a_13291_42460# a_13657_42558# 0.026223f
C10087 a_n2661_46634# a_4646_46812# 0.087334f
C10088 a_1123_46634# a_2443_46660# 2.91e-21
C10089 a_2107_46812# a_1799_45572# 0.079386f
C10090 a_948_46660# a_n2661_46098# 0.018472f
C10091 a_288_46660# a_479_46660# 4.61e-19
C10092 a_n2438_43548# a_2864_46660# 3.97e-20
C10093 a_n1925_46634# a_1302_46660# 1.88e-19
C10094 a_11309_47204# a_10428_46928# 0.025525f
C10095 a_n1613_43370# a_5841_46660# 2.95e-19
C10096 a_n2109_47186# a_n2293_46098# 1.23e-19
C10097 a_n2288_47178# a_n2157_46122# 1.61e-20
C10098 a_n2497_47436# a_n1853_46287# 0.029452f
C10099 a_12861_44030# a_14226_46987# 2.1e-19
C10100 a_n1435_47204# a_13693_46688# 1.97e-20
C10101 a_6491_46660# a_765_45546# 0.042766f
C10102 a_10227_46804# a_10425_46660# 6.24e-19
C10103 a_14311_47204# a_14180_46812# 5.09e-19
C10104 a_19386_47436# a_15227_44166# 2.72e-20
C10105 a_18597_46090# a_19333_46634# 1.8e-19
C10106 a_18479_47436# a_19692_46634# 0.078022f
C10107 a_11599_46634# a_13885_46660# 1.52e-20
C10108 a_4883_46098# a_3090_45724# 0.052016f
C10109 a_13507_46334# a_15368_46634# 0.023781f
C10110 a_12465_44636# a_14084_46812# 2.03e-19
C10111 a_n2293_45010# a_n1423_42826# 4.06e-19
C10112 a_n913_45002# a_n2472_42826# 7.39e-21
C10113 a_3065_45002# a_743_42282# 0.040577f
C10114 a_n1059_45260# a_n2157_42858# 1.41e-19
C10115 a_n2661_45010# a_n901_43156# 1.36e-21
C10116 a_n2017_45002# a_n1853_43023# 0.03086f
C10117 a_2711_45572# a_19326_42852# 1.2e-19
C10118 a_10057_43914# a_9801_43940# 0.006215f
C10119 a_8975_43940# a_9420_43940# 2.6e-19
C10120 a_1307_43914# a_15781_43660# 2.51e-20
C10121 a_n2433_44484# a_n2129_43609# 4.74e-21
C10122 a_9313_44734# a_20623_43914# 4.63e-20
C10123 a_n2840_43914# a_n2065_43946# 6.33e-21
C10124 a_8375_44464# a_8016_46348# 1.63e-20
C10125 a_16979_44734# a_17715_44484# 0.005407f
C10126 a_6109_44484# a_8199_44636# 1.61e-22
C10127 a_17767_44458# a_17583_46090# 1.63e-20
C10128 a_n356_44636# a_10903_43370# 2.05e-19
C10129 a_9838_44484# a_10809_44734# 1.37e-19
C10130 a_13667_43396# a_12861_44030# 5.08e-21
C10131 a_5663_43940# a_3090_45724# 0.001711f
C10132 a_14309_45028# a_13259_45724# 0.063402f
C10133 a_117_45144# a_310_45028# 2.88e-35
C10134 a_20193_45348# a_8049_45260# 6.42e-20
C10135 a_1145_45348# a_n443_42852# 2.98e-20
C10136 a_n2293_43922# a_1138_42852# 9.77e-21
C10137 a_17061_44734# a_12741_44636# 0.003447f
C10138 a_n2661_43922# a_1823_45246# 0.441151f
C10139 a_11309_47204# VDD 0.358104f
C10140 a_n4315_30879# a_n2216_40160# 0.001403f
C10141 a_n4334_40480# a_n4251_40480# 0.007692f
C10142 a_7174_31319# a_1239_39587# 2.3e-19
C10143 a_n4064_40160# a_n2302_40160# 0.249627f
C10144 a_1606_42308# C2_N_btm 0.021793f
C10145 a_18834_46812# a_20107_46660# 2.51e-21
C10146 a_19333_46634# a_19123_46287# 0.113955f
C10147 a_14180_46812# a_14226_46987# 0.006879f
C10148 a_13885_46660# a_13693_46688# 5.76e-19
C10149 a_15227_44166# a_19551_46910# 0.018691f
C10150 a_19466_46812# a_18285_46348# 7.08e-22
C10151 a_n2442_46660# a_n2956_38680# 0.047296f
C10152 a_n2293_46634# a_n2956_39304# 3.78e-19
C10153 a_8128_46384# a_8781_46436# 4.93e-20
C10154 a_4646_46812# a_8199_44636# 9.29e-19
C10155 a_5072_46660# a_5068_46348# 5.86e-19
C10156 a_3877_44458# a_5937_45572# 2.07e-20
C10157 a_11453_44696# a_13259_45724# 0.251534f
C10158 a_13507_46334# a_19597_46482# 7.17e-19
C10159 a_14955_43940# a_n97_42460# 6.16e-22
C10160 a_21115_43940# a_21381_43940# 0.073198f
C10161 a_7281_43914# a_6197_43396# 3.25e-19
C10162 a_n2661_42282# a_4699_43561# 1.76e-21
C10163 a_11967_42832# a_17324_43396# 8.32e-19
C10164 a_12607_44458# a_12379_42858# 3.9e-21
C10165 a_n356_44636# a_3681_42891# 1.42e-20
C10166 a_18479_45785# a_19332_42282# 2.44e-19
C10167 a_11341_43940# a_19741_43940# 0.003328f
C10168 a_15493_43940# a_19478_44056# 6.87e-19
C10169 a_n2293_43922# a_5649_42852# 1.78418f
C10170 a_n913_45002# a_9223_42460# 8.58e-19
C10171 a_n1059_45260# a_9803_42558# 8.94e-21
C10172 a_2382_45260# a_5932_42308# 4.34e-21
C10173 a_n2017_45002# a_9293_42558# 0.001147f
C10174 a_10807_43548# VDD 0.68049f
C10175 a_15903_45785# a_16115_45572# 3.12e-19
C10176 a_15599_45572# a_16855_45546# 0.043567f
C10177 a_15765_45572# a_16333_45814# 0.17072f
C10178 a_n3420_37984# C2_P_btm 0.03058f
C10179 a_n4064_37984# C4_P_btm 0.001746f
C10180 a_2982_43646# a_20202_43084# 0.034798f
C10181 a_n97_42460# a_1138_42852# 0.015603f
C10182 a_19987_42826# a_13661_43548# 1.73e-19
C10183 a_5534_30871# a_n2293_46634# 9.88e-20
C10184 a_16243_43396# a_3090_45724# 1.04e-20
C10185 a_n809_44244# a_n1079_45724# 8.53e-21
C10186 a_n984_44318# a_n2293_45546# 1.81e-20
C10187 a_10651_43940# a_9290_44172# 3.97e-19
C10188 a_564_42282# a_n1151_42308# 3.17e-20
C10189 a_472_46348# VDD 0.706547f
C10190 C0_dummy_N_btm C4_N_btm 0.113156f
C10191 C1_N_btm C2_N_btm 5.24136f
C10192 C0_N_btm C3_N_btm 0.409238f
C10193 C0_dummy_P_btm C5_N_btm 6.85e-20
C10194 C1_P_btm C7_N_btm 2.65e-19
C10195 C0_P_btm C6_N_btm 1.55e-19
C10196 a_20712_42282# CAL_N 0.001755f
C10197 a_13258_32519# a_22469_40625# 6.65e-19
C10198 a_n4209_39590# a_n3690_37440# 1.67e-19
C10199 a_n3565_39590# a_n4334_37440# 3.56e-19
C10200 a_4419_46090# a_526_44458# 0.099848f
C10201 a_4185_45028# a_n1925_42282# 0.638728f
C10202 a_3699_46348# a_3873_46454# 0.006584f
C10203 a_17639_46660# a_13259_45724# 5.11e-19
C10204 a_14840_46494# a_15682_46116# 3.86e-19
C10205 a_17730_32519# a_22400_42852# 1.31e-20
C10206 a_n2661_42282# a_6101_43172# 7.12e-20
C10207 a_n356_44636# a_15959_42545# 0.001149f
C10208 a_n2293_43922# a_7963_42308# 3.54e-20
C10209 a_n97_42460# a_5649_42852# 0.008438f
C10210 a_19862_44208# a_19987_42826# 2.09e-19
C10211 a_11341_43940# a_17333_42852# 1.63e-20
C10212 a_15493_43940# a_17701_42308# 2.87e-20
C10213 a_3626_43646# a_19700_43370# 7.81e-19
C10214 a_8685_43396# a_10341_43396# 2.41562f
C10215 a_9145_43396# a_14579_43548# 0.024497f
C10216 a_458_43396# a_743_42282# 3.19e-21
C10217 a_21811_47423# SINGLE_ENDED 0.215228f
C10218 a_12465_44636# START 0.065727f
C10219 a_22223_47212# RST_Z 2.25e-19
C10220 a_13467_32519# VDD 0.353373f
C10221 a_10775_45002# a_10951_45334# 0.185422f
C10222 a_16147_45260# a_11827_44484# 7.51e-20
C10223 a_2711_45572# a_n2661_42834# 2.44e-21
C10224 a_2382_45260# a_1423_45028# 0.036767f
C10225 a_4558_45348# a_1307_43914# 1.16e-20
C10226 a_6171_45002# a_14180_45002# 0.012672f
C10227 a_2274_45254# a_2232_45348# 0.002765f
C10228 a_413_45260# a_2903_45348# 4.7e-19
C10229 a_12379_42858# a_10903_43370# 0.02509f
C10230 a_12895_43230# a_9290_44172# 3.44e-20
C10231 a_19987_42826# a_4185_45028# 3.48e-20
C10232 a_18504_43218# a_17339_46660# 6.4e-19
C10233 a_7174_31319# a_n2956_39768# 5.27e-21
C10234 a_17324_43396# a_13259_45724# 2.64e-19
C10235 a_n2157_42858# a_n1925_42282# 1.51e-19
C10236 a_3457_43396# a_n443_42852# 0.009582f
C10237 a_15599_45572# a_13661_43548# 0.01321f
C10238 a_15903_45785# a_5807_45002# 5.55e-20
C10239 a_5907_45546# a_5257_43370# 0.064039f
C10240 a_4880_45572# a_4651_46660# 1.53e-20
C10241 a_15297_45822# a_13747_46662# 0.001012f
C10242 a_12561_45572# a_12549_44172# 0.001714f
C10243 a_3357_43084# a_18479_47436# 0.292061f
C10244 a_2437_43646# a_19386_47436# 0.00484f
C10245 a_413_45260# a_6575_47204# 2.11e-19
C10246 a_5147_45002# a_4791_45118# 0.10845f
C10247 a_7705_45326# a_2063_45854# 5.97e-19
C10248 a_4558_45348# a_n443_46116# 1.56e-19
C10249 a_310_45028# a_n755_45592# 0.02846f
C10250 a_n1099_45572# a_997_45618# 5.02e-19
C10251 a_4905_42826# a_5267_42460# 0.146764f
C10252 a_4093_43548# a_3905_42558# 4.12e-21
C10253 a_8037_42858# a_8952_43230# 0.118759f
C10254 a_3539_42460# a_1755_42282# 3.25e-19
C10255 a_n97_42460# a_7963_42308# 0.002153f
C10256 a_3080_42308# a_5379_42460# 1.73e-20
C10257 a_14621_43646# a_14635_42282# 1.99e-20
C10258 VDAC_Ni VDAC_P 1.02e-19
C10259 a_n3565_37414# a_n3607_37440# 0.001003f
C10260 a_n2946_37690# a_n2860_37690# 0.011479f
C10261 a_7754_38470# a_5700_37509# 0.971846f
C10262 a_3754_38470# VDAC_N 0.169096f
C10263 a_n4064_37440# a_n2302_37690# 0.239588f
C10264 a_8530_39574# a_5088_37509# 0.166912f
C10265 a_6773_42558# VDD 0.006434f
C10266 a_1239_47204# a_1431_47204# 0.219138f
C10267 a_n971_45724# a_3160_47472# 0.011577f
C10268 a_n452_47436# a_n1151_42308# 0.0065f
C10269 a_327_47204# a_584_46384# 6.38e-19
C10270 a_1209_47178# a_2124_47436# 0.095065f
C10271 a_n1741_47186# a_4007_47204# 0.012359f
C10272 a_n2109_47186# a_4791_45118# 0.34446f
C10273 a_n1059_45260# a_n1761_44111# 0.535535f
C10274 a_3357_43084# a_2479_44172# 0.0305f
C10275 a_n2017_45002# a_n1899_43946# 0.017371f
C10276 a_n2661_45010# a_n984_44318# 2.17e-20
C10277 a_n2293_45010# a_n1549_44318# 0.014826f
C10278 a_n913_45002# a_n2065_43946# 0.018244f
C10279 a_8137_45348# a_5891_43370# 4.09e-20
C10280 a_n2293_42834# a_8238_44734# 2.49e-21
C10281 a_n4318_40392# a_n1699_44726# 2.56e-21
C10282 a_7499_43078# a_10867_43940# 0.004845f
C10283 a_11827_44484# a_10334_44484# 1.87e-19
C10284 a_16922_45042# a_18248_44752# 7.57e-20
C10285 a_n2433_44484# a_n2129_44697# 0.130072f
C10286 a_n2661_44458# a_n2267_44484# 0.046548f
C10287 a_17613_45144# a_17767_44458# 0.003f
C10288 a_n2840_42282# a_n2810_45572# 2.3e-20
C10289 a_18707_42852# a_n357_42282# 0.003328f
C10290 a_13527_45546# a_2324_44458# 0.001831f
C10291 a_9159_45572# a_5937_45572# 0.048183f
C10292 a_14495_45572# a_14275_46494# 0.003638f
C10293 a_10907_45822# a_11189_46129# 0.021145f
C10294 a_10216_45572# a_8199_44636# 4.45e-19
C10295 a_9049_44484# a_6945_45028# 2.27e-20
C10296 a_11280_45822# a_9290_44172# 2.36e-19
C10297 a_19431_45546# a_12741_44636# 3.15e-20
C10298 a_n2661_44458# a_5807_45002# 1.89e-19
C10299 a_949_44458# a_768_44030# 0.002011f
C10300 a_18114_32519# a_19321_45002# 1.08e-21
C10301 a_2711_45572# a_5066_45546# 0.090644f
C10302 a_3232_43370# a_3090_45724# 0.024183f
C10303 a_5534_30871# a_13249_42558# 0.002316f
C10304 a_5342_30871# a_13575_42558# 4.35e-19
C10305 a_13460_43230# a_13657_42558# 2.98e-19
C10306 a_13635_43156# a_14113_42308# 0.002123f
C10307 a_16697_47582# a_5807_45002# 1.37e-19
C10308 a_9804_47204# a_n2661_46634# 0.02862f
C10309 a_n881_46662# a_n2312_38680# 4.41e-20
C10310 a_n1613_43370# a_n1925_46634# 0.33524f
C10311 a_2747_46873# a_2107_46812# 0.0019f
C10312 a_6151_47436# a_10249_46116# 0.056387f
C10313 a_n1435_47204# a_7411_46660# 3.15e-20
C10314 a_9313_45822# a_8145_46902# 3.14e-19
C10315 a_17517_44484# a_20159_44458# 0.026718f
C10316 a_626_44172# a_458_43396# 0.065365f
C10317 a_1307_43914# a_1756_43548# 0.267667f
C10318 a_10193_42453# a_12089_42308# 0.005996f
C10319 a_5883_43914# a_8018_44260# 2.21e-19
C10320 a_n2012_44484# a_n4318_39768# 4.36e-19
C10321 a_11827_44484# a_13565_44260# 4.08e-19
C10322 a_3065_45002# a_2813_43396# 3.35e-21
C10323 a_5111_44636# a_8147_43396# 0.08322f
C10324 a_6431_45366# a_6197_43396# 9.15e-21
C10325 a_n1059_45260# a_14579_43548# 0.250544f
C10326 a_n2017_45002# a_14358_43442# 2.42e-20
C10327 a_3537_45260# a_6655_43762# 0.031868f
C10328 a_2304_45348# VDD 0.004463f
C10329 a_n1630_35242# RST_Z 0.001585f
C10330 a_1606_42308# C8_P_btm 6.73e-20
C10331 a_n2661_44458# a_3699_46348# 3.05e-21
C10332 a_949_44458# a_1176_45822# 4.19e-19
C10333 a_16112_44458# a_11415_45002# 2.93e-20
C10334 a_13076_44458# a_12741_44636# 0.010522f
C10335 a_742_44458# a_1138_42852# 0.040731f
C10336 a_11341_43940# a_768_44030# 0.005879f
C10337 a_8333_44056# a_n2293_46634# 2.16e-20
C10338 a_9313_44734# a_13059_46348# 3.57e-19
C10339 a_18326_43940# a_13661_43548# 0.024789f
C10340 a_22223_43948# a_12549_44172# 6.97e-19
C10341 a_2809_45028# a_526_44458# 0.033247f
C10342 a_413_45260# a_n2661_45546# 0.022797f
C10343 a_n913_45002# a_n755_45592# 0.347782f
C10344 a_n467_45028# a_n2293_45546# 0.067105f
C10345 a_3357_43084# a_n443_42852# 0.042246f
C10346 a_16922_45042# a_2324_44458# 6.23e-21
C10347 a_11827_44484# a_9290_44172# 1.72e-19
C10348 a_n2661_43370# a_10809_44734# 0.077978f
C10349 a_9165_43940# a_4883_46098# 0.00241f
C10350 a_n1557_42282# a_n1151_42308# 0.214486f
C10351 a_3540_43646# a_584_46384# 0.045907f
C10352 a_1756_43548# a_n443_46116# 0.046156f
C10353 a_7227_47204# VDD 0.430714f
C10354 a_12563_42308# a_7174_31319# 9.76e-21
C10355 a_5932_42308# a_1239_39587# 2.77e-19
C10356 a_14113_42308# a_18310_42308# 4.09e-21
C10357 a_n2293_46634# a_n1991_46122# 0.0181f
C10358 a_n2104_46634# a_n1853_46287# 1.31e-20
C10359 a_n2661_46634# a_n901_46420# 9.25e-21
C10360 a_n2312_38680# a_n2157_46122# 0.001134f
C10361 a_n1925_46634# a_n2293_46098# 0.077794f
C10362 a_11186_47026# a_11735_46660# 3.88e-21
C10363 a_4646_46812# a_765_45546# 0.001856f
C10364 a_10467_46802# a_10425_46660# 2.56e-19
C10365 a_9804_47204# a_8199_44636# 8.66e-19
C10366 a_19787_47423# a_10809_44734# 0.002525f
C10367 a_20990_47178# a_6945_45028# 0.026188f
C10368 a_21177_47436# a_21137_46414# 1.13e-19
C10369 a_13507_46334# a_20708_46348# 0.007683f
C10370 a_4883_46098# a_20075_46420# 0.014562f
C10371 a_9313_45822# a_5066_45546# 0.019449f
C10372 a_11453_44696# a_18189_46348# 0.534507f
C10373 a_12465_44636# a_19553_46090# 6.8e-21
C10374 a_n881_46662# a_9823_46155# 1.37e-20
C10375 a_8128_46384# a_5937_45572# 1.99e-19
C10376 a_n2065_43946# a_n4318_39304# 3.62e-19
C10377 a_n2293_43922# a_8685_43396# 0.026511f
C10378 a_4223_44672# a_4361_42308# 7.99e-22
C10379 a_14539_43914# a_16867_43762# 0.004505f
C10380 a_10193_42453# a_18907_42674# 0.002509f
C10381 a_n356_44636# a_16243_43396# 4.44e-20
C10382 a_18374_44850# a_18429_43548# 2e-20
C10383 a_9313_44734# a_15095_43370# 0.039448f
C10384 a_18451_43940# a_19478_44306# 1.92e-19
C10385 a_19328_44172# a_15493_43396# 0.019584f
C10386 a_13483_43940# a_11341_43940# 0.005417f
C10387 a_7542_44172# a_7499_43940# 0.157633f
C10388 a_n2472_43914# a_n2433_43396# 7.88e-19
C10389 a_18287_44626# a_18783_43370# 4.14e-20
C10390 a_18443_44721# a_18525_43370# 0.001063f
C10391 a_18248_44752# a_15743_43084# 8.41e-20
C10392 a_22315_44484# VDD 0.213791f
C10393 a_11823_42460# a_14495_45572# 0.023559f
C10394 a_10180_45724# a_10210_45822# 0.006836f
C10395 a_8162_45546# a_8192_45572# 0.134163f
C10396 a_8746_45002# a_8697_45822# 3e-20
C10397 a_2711_45572# a_15861_45028# 0.02395f
C10398 a_10053_45546# a_10907_45822# 0.003363f
C10399 C3_N_btm C10_P_btm 0.001117f
C10400 C0_dummy_P_btm C5_P_btm 0.11375f
C10401 C2_N_btm C9_P_btm 2.13e-19
C10402 C1_N_btm C8_P_btm 4.41e-19
C10403 C0_N_btm C7_P_btm 2.32e-19
C10404 C0_dummy_N_btm C6_P_btm 1.37e-19
C10405 C8_N_btm EN_VIN_BSTR_N 0.090252f
C10406 C1_P_btm C3_P_btm 8.06688f
C10407 C0_P_btm C4_P_btm 0.138331f
C10408 a_9028_43914# a_8953_45546# 0.01093f
C10409 a_10949_43914# a_8016_46348# 3.79e-20
C10410 a_10405_44172# a_8199_44636# 1.31e-19
C10411 a_685_42968# a_n1613_43370# 2.27e-20
C10412 a_16414_43172# a_10227_46804# 4.57e-21
C10413 a_17333_42852# a_16327_47482# 0.006539f
C10414 a_21195_42852# a_12861_44030# 1.78e-21
C10415 a_5457_43172# a_4791_45118# 2.47e-19
C10416 a_4905_42826# a_3090_45724# 4.85e-19
C10417 a_13467_32519# a_22612_30879# 0.061222f
C10418 a_n1761_44111# a_n1925_42282# 5.08e-20
C10419 a_n2661_43922# a_n2293_45546# 2.12e-19
C10420 a_n2293_43922# a_n2956_38216# 2.59e-20
C10421 a_12156_46660# VDD 0.082428f
C10422 a_n4064_38528# C1_P_btm 4.13e-20
C10423 a_2698_46116# a_4185_45028# 5.29e-21
C10424 a_3147_46376# a_3483_46348# 0.207919f
C10425 a_12991_46634# a_12638_46436# 2.6e-19
C10426 a_11735_46660# a_12839_46116# 3.01e-20
C10427 a_3877_44458# a_n443_42852# 2.84e-23
C10428 a_11415_45002# a_13925_46122# 3.85e-20
C10429 a_1823_45246# a_5164_46348# 3.04e-19
C10430 a_20841_46902# a_21137_46414# 2.33e-19
C10431 a_20623_46660# a_20708_46348# 6.62e-19
C10432 a_20273_46660# a_6945_45028# 0.02808f
C10433 a_20107_46660# a_10809_44734# 0.026612f
C10434 a_5742_30871# a_3754_38470# 1.66e-19
C10435 a_4958_30871# a_n3420_37984# 0.031033f
C10436 a_n97_42460# a_8685_43396# 1.81e-19
C10437 a_15493_43940# a_4361_42308# 7.71e-20
C10438 a_n2661_42282# a_1847_42826# 2.73e-20
C10439 a_3499_42826# a_3935_42891# 7.16e-19
C10440 a_9313_44734# a_14097_32519# 0.053061f
C10441 a_11341_43940# a_13678_32519# 0.001425f
C10442 a_n1605_47204# CLK_DATA 1.66e-20
C10443 SMPL_ON_P DATA[0] 2.42e-19
C10444 a_n1741_47186# DATA[1] 0.021536f
C10445 w_1575_34946# VIN_P 2.57e-20
C10446 a_n2109_45247# a_n967_45348# 1e-19
C10447 a_2437_43646# a_3537_45260# 2.74e-21
C10448 a_n1059_45260# a_n2956_37592# 2.56e-20
C10449 a_n2017_45002# en_comp 0.004677f
C10450 a_n2661_45010# a_n467_45028# 0.227953f
C10451 a_16147_45260# a_15595_45028# 0.00203f
C10452 a_6511_45714# a_n2661_44458# 1.46e-20
C10453 a_22959_43396# a_4185_45028# 0.01521f
C10454 a_5932_42308# a_n2956_39768# 4.83e-21
C10455 a_n2433_43396# a_n357_42282# 2.74e-19
C10456 a_n1177_43370# a_n863_45724# 5.65e-20
C10457 a_15743_43084# a_2324_44458# 9.18e-19
C10458 a_19332_42282# a_13507_46334# 0.001224f
C10459 a_7174_31319# a_10227_46804# 2.63e-20
C10460 a_n2840_45546# VDD 0.302566f
C10461 a_7499_43078# a_n1613_43370# 0.324998f
C10462 a_5907_45546# a_5807_45002# 0.013402f
C10463 a_2711_45572# a_19321_45002# 1.76e-19
C10464 a_2981_46116# a_2957_45546# 6.65e-19
C10465 a_8049_45260# a_20062_46116# 1.01e-19
C10466 a_17538_32519# a_22400_42852# 1.17e-20
C10467 a_n97_42460# a_15953_42852# 0.001782f
C10468 a_10807_43548# a_11551_42558# 0.001883f
C10469 a_10341_43396# a_17333_42852# 3.64e-20
C10470 a_6755_46942# CLK 0.031541f
C10471 a_18175_45572# a_19279_43940# 9.28e-21
C10472 a_13556_45296# a_13076_44458# 8.16e-20
C10473 a_9482_43914# a_13720_44458# 0.188323f
C10474 a_1423_45028# a_5343_44458# 0.128331f
C10475 a_1307_43914# a_9838_44484# 5.82e-22
C10476 a_2711_45572# a_20623_43914# 2.17e-19
C10477 a_20623_45572# a_17517_44484# 1.02e-20
C10478 a_3232_43370# a_n356_44636# 1.34e-20
C10479 a_n2661_45010# a_n2661_43922# 0.111071f
C10480 a_5342_30871# a_n443_42852# 2.41e-19
C10481 a_21356_42826# a_n357_42282# 0.156735f
C10482 a_n1736_42282# a_n2956_39304# 2.99e-20
C10483 a_n3674_38216# a_n2956_38680# 0.02335f
C10484 a_3638_45822# a_1823_45246# 0.003923f
C10485 a_15037_45618# a_13059_46348# 0.064109f
C10486 a_18341_45572# a_3090_45724# 0.016963f
C10487 a_15415_45028# a_n743_46660# 3.05e-20
C10488 a_375_42282# a_n2293_46634# 0.004296f
C10489 a_6125_45348# a_5807_45002# 0.00337f
C10490 a_2437_43646# a_6969_46634# 5.02e-20
C10491 a_3357_43084# a_10554_47026# 2.24e-20
C10492 a_413_45260# a_5385_46902# 1.97e-20
C10493 a_n1059_45260# a_5257_43370# 2.6e-19
C10494 a_2680_45002# a_3877_44458# 2.18e-20
C10495 a_n2661_43370# a_n881_46662# 0.020731f
C10496 a_2711_45572# a_5068_46348# 9.3e-19
C10497 a_18315_45260# a_11453_44696# 0.010513f
C10498 a_20567_45036# a_4883_46098# 1.52e-20
C10499 a_11691_44458# a_18597_46090# 2.38e-20
C10500 a_6298_44484# a_6151_47436# 1.58e-19
C10501 a_4099_45572# a_4419_46090# 0.002575f
C10502 VCM VDD 1.50561f
C10503 a_700_44734# a_n2497_47436# 3.92e-21
C10504 a_10157_44484# a_4791_45118# 5.67e-20
C10505 a_16759_43396# a_4958_30871# 1.9e-19
C10506 a_3681_42891# a_3823_42558# 0.001239f
C10507 a_4361_42308# a_5742_30871# 0.071684f
C10508 a_5649_42852# a_10533_42308# 7.52e-20
C10509 a_743_42282# a_13575_42558# 0.009742f
C10510 a_19987_42826# a_20573_43172# 0.006947f
C10511 a_18817_42826# a_19326_42852# 2.6e-19
C10512 a_1847_42826# a_3497_42558# 2.53e-20
C10513 a_16137_43396# a_18907_42674# 0.001947f
C10514 a_8049_45260# CLK 0.033207f
C10515 a_20205_31679# a_22609_38406# 4.1e-21
C10516 a_3422_30871# VDAC_P 0.476125f
C10517 a_584_46384# a_1983_46706# 0.062968f
C10518 a_n1151_42308# a_33_46660# 0.005251f
C10519 a_n237_47217# a_n2661_46098# 0.01906f
C10520 a_2063_45854# a_2107_46812# 0.214026f
C10521 a_n971_45724# a_2609_46660# 0.004485f
C10522 a_4007_47204# a_n743_46660# 4.48e-20
C10523 a_4791_45118# a_n1925_46634# 0.026798f
C10524 a_13717_47436# a_5807_45002# 2.74e-19
C10525 a_6545_47178# a_n2661_46634# 0.022455f
C10526 a_15673_47210# a_16119_47582# 2.28e-19
C10527 a_16023_47582# a_12549_44172# 7.14e-20
C10528 a_n913_45002# a_n2129_43609# 0.023791f
C10529 a_n2810_45028# a_n4318_39304# 0.023142f
C10530 a_n2661_45010# a_n447_43370# 3.19e-22
C10531 a_n2017_45002# a_n1699_43638# 0.004053f
C10532 a_n2293_45010# a_n1177_43370# 0.001252f
C10533 a_1307_43914# a_12603_44260# 2.49e-19
C10534 a_8855_44734# a_n2661_43922# 1.87e-20
C10535 a_n2661_44458# a_n2065_43946# 8.48e-20
C10536 a_16112_44458# a_11967_42832# 2.42e-19
C10537 a_n2433_44484# a_n2472_43914# 9.53e-19
C10538 a_n2302_39866# a_n2810_45572# 2.61e-19
C10539 a_n3420_39616# a_n2956_38216# 1.85e-19
C10540 a_22959_45572# VDD 0.304443f
C10541 a_22223_45572# a_8049_45260# 0.013885f
C10542 a_n2956_37592# a_n1925_42282# 2.26e-20
C10543 a_14180_45002# a_10903_43370# 0.008124f
C10544 a_9482_43914# a_13351_46090# 2.3e-19
C10545 a_10775_45002# a_2324_44458# 0.003159f
C10546 a_13556_45296# a_12594_46348# 1.95e-21
C10547 a_4185_45348# a_5164_46348# 4.37e-22
C10548 a_18079_43940# a_11599_46634# 3.46e-21
C10549 a_10729_43914# a_10227_46804# 3.09e-19
C10550 a_15493_43396# a_12861_44030# 0.254093f
C10551 a_13807_45067# a_11415_45002# 0.001105f
C10552 a_8975_43940# a_3090_45724# 0.003577f
C10553 a_175_44278# a_768_44030# 6.16e-19
C10554 a_18691_45572# a_19240_46482# 2.45e-19
C10555 a_22400_42852# a_22465_38105# 0.199207f
C10556 a_8685_42308# a_8791_42308# 0.147376f
C10557 a_8325_42308# a_9223_42460# 8.85e-19
C10558 a_6761_42308# a_5742_30871# 1.69e-20
C10559 a_11530_34132# RST_Z 0.01695f
C10560 CAL_P VIN_N 0.001176f
C10561 C10_P_btm C7_P_btm 1.39624f
C10562 C9_P_btm C8_P_btm 39.4538f
C10563 a_5807_45002# a_14035_46660# 0.025174f
C10564 a_n743_46660# a_15368_46634# 0.026392f
C10565 a_n2293_46634# a_15227_44166# 3.53e-19
C10566 a_12549_44172# a_16751_46987# 3.29e-19
C10567 a_9804_47204# a_765_45546# 0.028432f
C10568 a_22731_47423# a_22591_46660# 0.011433f
C10569 a_12465_44636# a_12741_44636# 0.914049f
C10570 a_11453_44696# a_20202_43084# 0.002113f
C10571 SMPL_ON_N a_11415_45002# 4.16e-20
C10572 a_13507_46334# a_21542_46660# 0.001196f
C10573 a_4883_46098# a_21076_30879# 2.94e-20
C10574 a_12861_44030# a_3483_46348# 0.06952f
C10575 a_4915_47217# a_9569_46155# 1.77e-20
C10576 a_6151_47436# a_5937_45572# 0.008183f
C10577 a_n1151_42308# a_12005_46116# 3.22e-19
C10578 a_16922_45042# a_15743_43084# 0.00548f
C10579 a_20512_43084# a_20935_43940# 1.43e-20
C10580 a_n356_44636# a_4905_42826# 6.1e-20
C10581 a_5244_44056# a_n2661_42282# 1.4e-20
C10582 a_n2293_42834# a_4361_42308# 2.59e-19
C10583 a_5883_43914# a_6452_43396# 0.001768f
C10584 a_n913_45002# a_21195_42852# 0.002742f
C10585 en_comp a_19164_43230# 1.47e-21
C10586 a_8375_44464# VDD 0.086619f
C10587 a_n3565_38502# C10_P_btm 2.25e-20
C10588 a_n4209_38502# C8_P_btm 5.41e-20
C10589 a_n4209_38216# a_n1838_35608# 1.13e-19
C10590 a_2711_45572# a_3775_45552# 0.044123f
C10591 a_5907_45546# a_6511_45714# 0.043475f
C10592 a_6194_45824# a_6472_45840# 0.118423f
C10593 a_22521_40599# a_20205_31679# 2.04e-20
C10594 a_22959_44484# a_4185_45028# 0.011365f
C10595 a_10341_43396# a_768_44030# 1.28e-19
C10596 a_9145_43396# a_5807_45002# 1.15e-19
C10597 a_6655_43762# a_n2293_46634# 0.003277f
C10598 a_14021_43940# a_14976_45028# 2.27e-20
C10599 a_7640_43914# a_8034_45724# 1.7e-20
C10600 a_n2661_44458# a_n755_45592# 0.023853f
C10601 a_n1177_44458# a_n863_45724# 1.65e-20
C10602 a_n1352_44484# a_n1079_45724# 1.48e-20
C10603 a_n452_44636# a_n2293_45546# 1.06e-19
C10604 a_2779_44458# a_n2661_45546# 4.85e-20
C10605 a_16112_44458# a_13259_45724# 1.59e-20
C10606 a_17517_44484# a_18819_46122# 5.47e-21
C10607 a_4190_30871# a_18597_46090# 0.022042f
C10608 a_5534_30871# w_11334_34010# 0.002185f
C10609 a_20447_31679# a_22821_38993# 7.74e-20
C10610 a_n4209_38502# a_n4334_38528# 0.25243f
C10611 a_n3420_39072# a_n3607_38528# 2.09e-19
C10612 a_4955_46873# VDD 0.467566f
C10613 a_21188_46660# a_21076_30879# 9.43e-21
C10614 a_20528_46660# a_12741_44636# 0.018376f
C10615 a_5257_43370# a_n1925_42282# 1.27e-20
C10616 a_n2810_45028# a_n4334_40480# 8.59e-19
C10617 a_n2956_37592# a_n4315_30879# 0.107228f
C10618 a_19721_31679# a_22400_42852# 3.49e-20
C10619 a_10949_43914# a_12281_43396# 5.57e-19
C10620 a_n2840_43370# a_n2267_43396# 6.1e-19
C10621 a_18114_32519# a_14097_32519# 0.054468f
C10622 a_n2293_42834# a_6761_42308# 3.63e-21
C10623 a_9313_44734# a_22959_42860# 0.174475f
C10624 a_15433_44458# a_15567_42826# 4.21e-21
C10625 a_2479_44172# a_743_42282# 2.08e-20
C10626 a_n4318_39304# a_n2129_43609# 5.32e-19
C10627 a_13483_43940# a_10341_43396# 3.72e-20
C10628 a_19319_43548# VDD 0.561461f
C10629 a_11823_42460# a_11963_45334# 0.110904f
C10630 a_11962_45724# a_13159_45002# 2.65e-19
C10631 a_10193_42453# a_14537_43396# 1.09e-19
C10632 a_11322_45546# a_13556_45296# 1.25e-20
C10633 a_8192_45572# a_3537_45260# 2.88e-19
C10634 a_18479_45785# a_19365_45572# 0.001158f
C10635 a_n1329_42308# a_n1613_43370# 0.001867f
C10636 VDAC_P VREF_GND 0.203715f
C10637 a_9803_43646# a_3483_46348# 5.4e-19
C10638 a_16409_43396# a_12741_44636# 2.16e-19
C10639 a_20753_42852# a_12549_44172# 8.1e-20
C10640 a_14635_42282# a_n2293_46634# 2.07e-20
C10641 a_9672_43914# a_n443_42852# 8.44e-20
C10642 a_n2267_43396# a_n1925_42282# 6.35e-19
C10643 a_n967_46494# VDD 2.82e-20
C10644 a_2711_45572# a_15811_47375# 1.5e-20
C10645 a_7499_43078# a_4791_45118# 0.024468f
C10646 a_10490_45724# a_n1151_42308# 2.28e-20
C10647 a_1823_45246# a_3316_45546# 0.099099f
C10648 a_167_45260# a_2957_45546# 7.72e-19
C10649 a_1176_45822# a_n356_45724# 1.67e-19
C10650 a_2804_46116# a_n755_45592# 2.12e-20
C10651 a_14493_46090# a_14383_46116# 0.097745f
C10652 a_13925_46122# a_13259_45724# 0.003795f
C10653 a_10341_43396# a_13678_32519# 0.011962f
C10654 a_n97_42460# a_17333_42852# 0.003266f
C10655 a_3626_43646# a_9127_43156# 2.22e-19
C10656 a_2982_43646# a_10083_42826# 9.5e-20
C10657 a_n2661_42282# a_n473_42460# 1.46e-19
C10658 a_18783_43370# a_19268_43646# 0.001296f
C10659 a_15493_43396# a_19518_43218# 8.64e-20
C10660 a_22612_30879# VCM 0.473529f
C10661 a_n1925_46634# DATA[3] 4.06e-21
C10662 a_n2438_43548# DATA[0] 5.04e-19
C10663 a_n743_46660# DATA[1] 1.69e-21
C10664 a_16795_42852# VDD 0.179044f
C10665 a_19479_31679# a_22521_40599# 1.54e-20
C10666 a_n2810_45028# a_n2946_37690# 0.024678f
C10667 a_n2956_37592# a_n3420_37440# 0.233174f
C10668 a_n2017_45002# a_n1699_44726# 0.002575f
C10669 a_n2956_37592# a_n4318_40392# 2.71462f
C10670 a_n2661_45010# a_n452_44636# 0.020671f
C10671 a_3357_43084# a_5518_44484# 0.009558f
C10672 a_n2293_45010# a_n1177_44458# 0.00518f
C10673 a_n913_45002# a_n2129_44697# 0.017685f
C10674 a_18799_45938# a_18989_43940# 1.13e-19
C10675 a_14537_43396# a_14309_45348# 2.07e-19
C10676 a_8696_44636# a_9313_44734# 0.003528f
C10677 a_14180_45002# a_14403_45348# 0.011458f
C10678 a_13348_45260# a_13490_45067# 0.005572f
C10679 a_1307_43914# a_n2661_43370# 1.06e-19
C10680 a_10193_42453# a_20835_44721# 2.06e-19
C10681 a_n1630_35242# a_20820_30879# 2.91e-19
C10682 a_743_42282# a_n443_42852# 0.03363f
C10683 a_20749_43396# a_n357_42282# 0.001735f
C10684 a_n3674_39304# a_n2810_45572# 0.023379f
C10685 a_n1991_42858# a_n863_45724# 3.37e-21
C10686 a_4574_45260# a_n881_46662# 1.99e-20
C10687 a_13017_45260# a_11453_44696# 0.004658f
C10688 a_13556_45296# a_12465_44636# 0.248126f
C10689 a_14180_45002# a_4883_46098# 7.48e-22
C10690 a_n2661_43370# a_n443_46116# 0.030763f
C10691 a_10193_42453# a_3090_45724# 0.027088f
C10692 a_2711_45572# a_13059_46348# 0.075233f
C10693 a_11823_42460# a_11901_46660# 2.29e-20
C10694 a_11962_45724# a_12251_46660# 1.12e-21
C10695 a_413_45260# a_12891_46348# 5.52e-20
C10696 a_n1059_45260# a_5807_45002# 5.37e-20
C10697 a_n2017_45002# a_13661_43548# 9.71e-20
C10698 a_2437_43646# a_n2293_46634# 0.030387f
C10699 a_20447_31679# a_21588_30879# 0.055937f
C10700 a_3357_43084# a_n2661_46634# 0.032385f
C10701 a_22591_43396# a_22400_42852# 5.76e-19
C10702 a_8037_42858# a_8495_42852# 0.027317f
C10703 a_13887_32519# a_14097_32519# 10.5943f
C10704 a_3626_43646# a_17124_42282# 0.004372f
C10705 a_8685_43396# a_10533_42308# 6.52e-23
C10706 a_9145_43396# a_9223_42460# 1.05e-20
C10707 a_20922_43172# a_21195_42852# 0.119168f
C10708 a_21335_42336# VDD 0.199586f
C10709 a_n2497_47436# a_n881_46662# 2.87e-19
C10710 a_n2109_47186# a_3411_47243# 0.001394f
C10711 a_n1741_47186# a_5063_47570# 2.13e-19
C10712 a_n746_45260# a_7_47243# 1.85e-19
C10713 a_n971_45724# a_3094_47570# 5.15e-19
C10714 a_13717_47436# a_14311_47204# 0.00371f
C10715 a_13381_47204# a_11599_46634# 2.3e-21
C10716 a_12861_44030# a_13487_47204# 0.127147f
C10717 a_2063_45854# a_11453_44696# 6.07e-19
C10718 a_18911_45144# a_17517_44484# 2.31e-19
C10719 a_17767_44458# a_18287_44626# 0.043567f
C10720 a_17970_44736# a_18248_44752# 0.117156f
C10721 a_1307_43914# a_2998_44172# 0.233292f
C10722 a_5343_44458# a_6109_44484# 0.285594f
C10723 a_4223_44672# a_5891_43370# 0.020744f
C10724 a_7499_43078# a_8791_43396# 0.04623f
C10725 a_5518_44484# a_5826_44734# 0.017351f
C10726 a_14539_43914# a_18374_44850# 9.06e-21
C10727 a_626_44172# a_2479_44172# 1.03e-20
C10728 a_11827_44484# a_12553_44484# 2.82e-19
C10729 a_n2017_45002# a_19862_44208# 1e-20
C10730 a_20447_31679# a_15493_43940# 1.09e-20
C10731 a_5111_44636# a_n2661_42282# 0.025961f
C10732 a_3232_43370# a_3820_44260# 0.003566f
C10733 a_5755_42308# a_n443_42852# 4.68e-21
C10734 a_8325_42308# a_n755_45592# 0.040306f
C10735 a_8685_42308# a_n357_42282# 1.11e-20
C10736 a_5742_30871# a_n2810_45572# 4.02e-21
C10737 a_5342_30871# CAL_P 0.007017f
C10738 a_327_44734# a_472_46348# 1.53e-19
C10739 a_4558_45348# a_n2293_46098# 0.030863f
C10740 a_11691_44458# a_6755_46942# 0.192426f
C10741 a_5343_44458# a_4646_46812# 0.24395f
C10742 a_n913_45002# a_3483_46348# 1.56e-20
C10743 a_13468_44734# a_12891_46348# 0.001942f
C10744 a_n2293_43922# a_768_44030# 0.027199f
C10745 a_n2017_45002# a_4185_45028# 0.029634f
C10746 a_11962_45724# a_13259_45724# 0.026896f
C10747 a_10210_45822# a_10586_45546# 0.042978f
C10748 a_2711_45572# a_3218_45724# 0.1731f
C10749 a_3175_45822# a_2957_45546# 0.08213f
C10750 a_2211_45572# a_n2661_45546# 3.69e-19
C10751 a_19431_45546# a_18985_46122# 0.00184f
C10752 a_19256_45572# a_18819_46122# 9.17e-19
C10753 a_2437_43646# a_9625_46129# 5.97e-20
C10754 a_3357_43084# a_8199_44636# 9.87e-21
C10755 a_20679_44626# a_4883_46098# 8.04e-21
C10756 a_21073_44484# a_16327_47482# 0.001903f
C10757 a_2998_44172# a_n443_46116# 0.001009f
C10758 a_n784_42308# a_5267_42460# 1.96e-20
C10759 a_13291_42460# a_13333_42558# 0.001565f
C10760 a_22165_42308# a_21973_42336# 5.76e-19
C10761 a_n2661_46634# a_3877_44458# 0.010452f
C10762 a_948_46660# a_1799_45572# 5.85e-19
C10763 a_1123_46634# a_n2661_46098# 0.041919f
C10764 a_n2438_43548# a_3524_46660# 7.85e-21
C10765 a_n1925_46634# a_1057_46660# 1.6e-19
C10766 a_n881_46662# a_6682_46987# 1.68e-19
C10767 a_n2497_47436# a_n2157_46122# 0.034181f
C10768 a_n2288_47178# a_n2293_46098# 1.13e-19
C10769 a_13487_47204# a_14180_46812# 0.001914f
C10770 a_6545_47178# a_765_45546# 0.035873f
C10771 a_12861_44030# a_14513_46634# 0.036912f
C10772 a_10227_46804# a_10185_46660# 0.002879f
C10773 a_18597_46090# a_15227_44166# 0.150202f
C10774 a_18479_47436# a_19466_46812# 0.007963f
C10775 a_13507_46334# a_14976_45028# 0.020647f
C10776 a_3080_42308# a_3754_39466# 2.89e-20
C10777 en_comp a_14209_32519# 6.81e-20
C10778 a_n2293_45010# a_n1991_42858# 7.5e-20
C10779 a_n2661_45010# a_n1641_43230# 4.2e-20
C10780 a_n2017_45002# a_n2157_42858# 0.040763f
C10781 a_14537_43396# a_16137_43396# 2.96e-20
C10782 a_8975_43940# a_9165_43940# 0.004776f
C10783 a_1307_43914# a_15681_43442# 2.36e-20
C10784 a_9313_44734# a_20365_43914# 1.7e-20
C10785 a_n2840_43914# a_n2472_43914# 7.52e-19
C10786 a_n2433_44484# a_n2433_43396# 0.001566f
C10787 VDAC_Ni VDD 0.288547f
C10788 a_17801_45144# VDD 2.88e-19
C10789 a_4958_30871# EN_VIN_BSTR_N 0.021638f
C10790 a_15720_42674# RST_Z 6.53e-21
C10791 a_7640_43914# a_8016_46348# 2.21e-22
C10792 a_14539_43914# a_17715_44484# 6.56e-19
C10793 a_4190_30871# w_11334_34010# 0.006418f
C10794 a_n2661_42834# a_1823_45246# 0.174801f
C10795 a_3363_44484# a_3147_46376# 4e-21
C10796 a_16241_44734# a_12741_44636# 0.006663f
C10797 a_n2661_43922# a_1138_42852# 0.027736f
C10798 a_n97_42460# a_768_44030# 0.034422f
C10799 a_5495_43940# a_3090_45724# 0.004468f
C10800 a_17538_32519# a_13747_46662# 1.11e-19
C10801 a_11257_43940# a_n2293_46634# 1.65e-19
C10802 a_626_44172# a_n443_42852# 0.028669f
C10803 a_11691_44458# a_8049_45260# 7.14e-20
C10804 a_13807_45067# a_13259_45724# 1.17e-19
C10805 a_n4315_30879# a_n4251_40480# 0.00226f
C10806 a_1606_42308# C1_N_btm 0.096405f
C10807 a_5342_30871# CAL_N 0.004302f
C10808 a_15227_44166# a_19123_46287# 0.069758f
C10809 a_14180_46812# a_14513_46634# 0.253235f
C10810 a_13885_46660# a_14543_46987# 7.87e-19
C10811 a_14035_46660# a_14226_46987# 3.26e-19
C10812 a_n2472_46634# a_n2956_38680# 4.88e-19
C10813 a_n2442_46660# a_n2956_39304# 0.046604f
C10814 a_5167_46660# a_5497_46414# 0.003426f
C10815 a_n1925_46634# a_6945_45028# 0.028603f
C10816 a_12465_44636# a_16375_45002# 4.56e-21
C10817 a_4883_46098# a_19431_46494# 2.01e-19
C10818 a_18479_47436# a_20205_31679# 0.001643f
C10819 a_10227_46804# a_20850_46155# 2.21e-19
C10820 a_12861_44030# a_n357_42282# 2.04e-19
C10821 a_n443_46116# a_2307_45899# 0.001194f
C10822 a_6453_43914# a_6197_43396# 0.001638f
C10823 a_2479_44172# a_2813_43396# 0.115852f
C10824 a_n2661_42282# a_4235_43370# 3.96e-21
C10825 a_11967_42832# a_17499_43370# 0.006642f
C10826 a_n356_44636# a_2905_42968# 2.11e-20
C10827 a_13483_43940# a_n97_42460# 1.05e-21
C10828 a_15493_43940# a_18533_43940# 0.052096f
C10829 a_19862_44208# a_21845_43940# 7.54e-21
C10830 a_20935_43940# a_21381_43940# 1.53e-19
C10831 a_11341_43940# a_21205_44306# 3.95e-19
C10832 a_3537_45260# a_4921_42308# 0.01091f
C10833 a_n913_45002# a_8791_42308# 0.005212f
C10834 a_n1059_45260# a_9223_42460# 1.29e-20
C10835 a_n2017_45002# a_9803_42558# 0.003827f
C10836 a_10949_43914# VDD 0.797824f
C10837 a_15903_45785# a_16333_45814# 2.33e-20
C10838 a_15599_45572# a_16115_45572# 0.105995f
C10839 a_15037_45618# a_8696_44636# 3.1e-21
C10840 a_n4064_37984# C5_P_btm 1.01e-19
C10841 a_n3420_37984# C3_P_btm 0.001771f
C10842 a_19164_43230# a_13661_43548# 3.49e-19
C10843 a_14543_43071# a_n2293_46634# 9.13e-20
C10844 a_16137_43396# a_3090_45724# 1.3e-20
C10845 a_n1549_44318# a_n1079_45724# 1.64e-19
C10846 a_n809_44244# a_n2293_45546# 5.56e-20
C10847 a_n1331_43914# a_n863_45724# 1.23e-20
C10848 a_10555_43940# a_9290_44172# 4.56e-19
C10849 a_n3674_37592# a_n1151_42308# 0.007818f
C10850 a_961_42354# a_584_46384# 9.03e-21
C10851 a_376_46348# VDD 0.116284f
C10852 C0_dummy_N_btm C3_N_btm 0.087354f
C10853 C0_N_btm C2_N_btm 0.827449f
C10854 C0_dummy_P_btm C4_N_btm 6.85e-20
C10855 C1_P_btm C6_N_btm 1.76e-19
C10856 C0_P_btm C5_N_btm 7.74e-20
C10857 a_20107_42308# CAL_N 0.001744f
C10858 a_7174_31319# VDAC_P 0.009133f
C10859 a_13258_32519# a_22521_40599# 4.4e-19
C10860 a_4185_45028# a_526_44458# 0.162857f
C10861 a_3699_46348# a_n1925_42282# 0.011511f
C10862 a_3483_46348# a_3873_46454# 6.61e-19
C10863 a_1823_45246# a_5066_45546# 5.66e-19
C10864 a_n3420_38528# a_n4064_37984# 7.35343f
C10865 a_n4064_38528# a_n3420_37984# 0.044626f
C10866 a_n4064_40160# a_n4064_37440# 0.056406f
C10867 a_n3565_39590# a_n4209_37414# 0.031279f
C10868 a_n4209_39590# a_n3565_37414# 0.032656f
C10869 a_n2946_38778# a_n2946_37984# 0.052227f
C10870 a_14840_46494# a_2324_44458# 0.002377f
C10871 a_n2661_42282# a_5837_43172# 7.96e-20
C10872 a_n4318_40392# a_n4251_40480# 0.001483f
C10873 a_n356_44636# a_15803_42450# 0.078793f
C10874 a_5891_43370# a_5742_30871# 1.08e-19
C10875 a_n2293_43922# a_6123_31319# 0.080985f
C10876 a_n2661_42834# a_5934_30871# 1.84e-21
C10877 a_19862_44208# a_19164_43230# 1.82e-21
C10878 a_11341_43940# a_18083_42858# 7.11e-21
C10879 a_15493_43940# a_17595_43084# 1.73e-20
C10880 a_n4318_39304# a_n2840_42826# 4.88e-19
C10881 a_3626_43646# a_19268_43646# 7.05e-22
C10882 a_9145_43396# a_13667_43396# 0.074541f
C10883 a_9803_43646# a_10695_43548# 0.007519f
C10884 a_4883_46098# SINGLE_ENDED 0.1664f
C10885 a_12465_44636# RST_Z 0.002855f
C10886 a_19095_43396# VDD 0.003529f
C10887 a_14495_45572# a_14539_43914# 9.15e-22
C10888 a_19431_45546# a_19778_44110# 0.010264f
C10889 a_17668_45572# a_16922_45042# 4.77e-19
C10890 a_18596_45572# a_18587_45118# 4.99e-19
C10891 a_19256_45572# a_18911_45144# 3.16e-19
C10892 a_10193_42453# a_n356_44636# 2.49128f
C10893 a_2274_45254# a_1423_45028# 8.25e-20
C10894 a_6171_45002# a_13777_45326# 0.010994f
C10895 a_4574_45260# a_1307_43914# 1.78e-21
C10896 a_13113_42826# a_9290_44172# 0.003778f
C10897 a_19164_43230# a_4185_45028# 6.39e-21
C10898 a_n2293_42282# a_1823_45246# 0.03994f
C10899 a_17499_43370# a_13259_45724# 0.018042f
C10900 a_2813_43396# a_n443_42852# 0.017355f
C10901 a_15599_45572# a_5807_45002# 0.002399f
C10902 a_5263_45724# a_5257_43370# 0.088982f
C10903 a_2711_45572# a_7577_46660# 4.24e-20
C10904 a_15225_45822# a_13747_46662# 6.29e-19
C10905 a_3357_43084# a_18143_47464# 5.7e-19
C10906 a_2437_43646# a_18597_46090# 0.006962f
C10907 a_21542_45572# a_16327_47482# 0.002879f
C10908 a_19479_31679# a_18479_47436# 2.29e-20
C10909 a_413_45260# a_7903_47542# 1.03e-19
C10910 a_4558_45348# a_4791_45118# 0.077256f
C10911 a_6709_45028# a_2063_45854# 4.65e-20
C10912 a_4574_45260# a_n443_46116# 5.16e-20
C10913 a_6171_45002# a_n1151_42308# 0.02292f
C10914 a_9482_43914# a_n971_45724# 8.96e-21
C10915 a_1307_43914# a_n2497_47436# 0.069365f
C10916 a_n2661_45546# a_n23_45546# 0.006975f
C10917 a_n1099_45572# a_n755_45592# 0.193775f
C10918 a_310_45028# a_n357_42282# 0.113929f
C10919 a_380_45546# a_997_45618# 0.070624f
C10920 a_n2293_45546# a_3316_45546# 1.26e-20
C10921 a_n97_42460# a_6123_31319# 0.182488f
C10922 a_8605_42826# a_8387_43230# 0.209641f
C10923 a_7871_42858# a_10083_42826# 4.52e-21
C10924 a_8037_42858# a_9127_43156# 0.042737f
C10925 a_13887_32519# a_22959_42860# 0.012735f
C10926 a_3539_42460# a_1606_42308# 2.57e-20
C10927 a_15493_43940# a_21887_42336# 6.82e-21
C10928 a_7765_42852# a_8952_43230# 3.38e-20
C10929 a_4905_42826# a_3823_42558# 3.67e-20
C10930 a_3626_43646# a_1755_42282# 0.119352f
C10931 a_21188_46660# SINGLE_ENDED 4.66e-21
C10932 a_7754_38636# VDAC_P 3.34e-19
C10933 VDAC_Ni a_8912_37509# 4.77e-20
C10934 a_8530_39574# a_4338_37500# 0.093669f
C10935 a_n3420_37440# a_n2860_37690# 0.002301f
C10936 a_n2946_37690# a_n2302_37690# 6.68e-19
C10937 a_7754_38470# a_5088_37509# 0.394117f
C10938 a_3754_38470# a_6886_37412# 7.59e-20
C10939 a_n2497_47436# a_n443_46116# 0.026321f
C10940 a_n971_45724# a_2905_45572# 0.118495f
C10941 a_n815_47178# a_n1151_42308# 0.011772f
C10942 a_1209_47178# a_1431_47204# 0.095209f
C10943 a_n237_47217# a_2553_47502# 4.45e-21
C10944 a_n1741_47186# a_3815_47204# 0.023296f
C10945 a_n2109_47186# a_4700_47436# 0.038955f
C10946 a_n785_47204# a_584_46384# 0.002399f
C10947 a_6481_42558# VDD 0.006426f
C10948 en_comp a_17730_32519# 9.67e-20
C10949 a_2437_43646# a_2675_43914# 3.12e-21
C10950 a_n2293_45010# a_n1331_43914# 0.02919f
C10951 a_n2017_45002# a_n1761_44111# 0.02974f
C10952 a_n2661_45010# a_n809_44244# 2.22e-19
C10953 a_n1059_45260# a_n2065_43946# 7.97e-21
C10954 a_11827_44484# a_10157_44484# 6.15e-20
C10955 a_n4318_40392# a_n2267_44484# 0.004061f
C10956 a_9482_43914# a_17061_44734# 2.21e-21
C10957 a_n2293_42834# a_5891_43370# 0.669411f
C10958 a_16922_45042# a_17970_44736# 2.81e-20
C10959 a_n2661_44458# a_n2129_44697# 0.035428f
C10960 a_15861_45028# a_15682_43940# 8.44e-19
C10961 a_9803_42558# a_526_44458# 2.85e-19
C10962 a_2437_43646# a_19123_46287# 7.12e-20
C10963 a_3357_43084# a_765_45546# 0.035297f
C10964 a_5691_45260# a_3090_45724# 1.29e-22
C10965 a_5883_43914# a_n881_46662# 2.63e-20
C10966 a_13163_45724# a_2324_44458# 7.36e-21
C10967 a_13249_42308# a_14275_46494# 8.84e-19
C10968 a_14495_45572# a_14493_46090# 0.00228f
C10969 a_10907_45822# a_9290_44172# 0.262972f
C10970 a_9159_45572# a_8199_44636# 0.049711f
C10971 a_10210_45822# a_11189_46129# 3.66e-19
C10972 a_7499_43078# a_6945_45028# 4.09e-22
C10973 a_18596_45572# a_11415_45002# 9.68e-19
C10974 a_5837_45028# a_5732_46660# 3.47e-21
C10975 a_10951_45334# a_10768_47026# 8.49e-21
C10976 a_742_44458# a_768_44030# 0.216263f
C10977 a_20205_45028# a_19321_45002# 5.38e-19
C10978 a_19721_31679# a_13747_46662# 0.001393f
C10979 a_5837_45348# a_5257_43370# 0.001158f
C10980 a_5342_30871# a_13070_42354# 2.82e-21
C10981 a_5534_30871# a_14456_42282# 4.39e-19
C10982 a_13635_43156# a_13657_42558# 4.38e-19
C10983 a_8128_46384# a_n2661_46634# 0.029397f
C10984 a_n1613_43370# a_n2312_38680# 4.23e-21
C10985 a_2747_46873# a_948_46660# 4.23e-19
C10986 a_n1435_47204# a_5257_43370# 2.43e-20
C10987 a_4915_47217# a_6969_46634# 1.7e-19
C10988 a_6151_47436# a_10554_47026# 1.71e-19
C10989 a_9067_47204# a_8667_46634# 0.005569f
C10990 a_9313_45822# a_7577_46660# 3.38e-19
C10991 a_2063_45854# a_10384_47026# 1.72e-19
C10992 a_17517_44484# a_19615_44636# 0.018532f
C10993 a_1307_43914# a_1568_43370# 0.182552f
C10994 a_10193_42453# a_12379_42858# 7.83e-20
C10995 a_5883_43914# a_7911_44260# 2.82e-19
C10996 a_6171_45002# a_6197_43396# 1.3e-20
C10997 a_2382_45260# a_3457_43396# 0.004922f
C10998 a_5205_44484# a_6031_43396# 9.87e-20
C10999 a_5111_44636# a_7112_43396# 0.041581f
C11000 a_n2017_45002# a_14579_43548# 0.003714f
C11001 a_3537_45260# a_6452_43396# 0.00408f
C11002 a_1606_42308# C9_P_btm 9.33e-20
C11003 a_n2661_44458# a_3483_46348# 1.44355f
C11004 a_949_44458# a_1208_46090# 2.47e-20
C11005 a_12883_44458# a_12741_44636# 0.073263f
C11006 a_15004_44636# a_11415_45002# 6.08e-19
C11007 a_11341_43940# a_12549_44172# 0.406618f
C11008 a_18079_43940# a_13661_43548# 0.028277f
C11009 a_1423_45028# a_8034_45724# 2.81e-21
C11010 a_2448_45028# a_526_44458# 7.21e-21
C11011 a_n1059_45260# a_n755_45592# 0.53237f
C11012 a_n967_45348# a_n863_45724# 4.28e-20
C11013 a_n37_45144# a_n2661_45546# 0.001732f
C11014 a_n913_45002# a_n357_42282# 0.309845f
C11015 a_n955_45028# a_n2293_45546# 0.002208f
C11016 a_2437_43646# a_2277_45546# 0.001212f
C11017 a_6031_43396# a_n971_45724# 4.44e-21
C11018 a_2982_43646# a_584_46384# 0.057754f
C11019 a_1568_43370# a_n443_46116# 0.584982f
C11020 a_n1630_35242# a_n2302_38778# 5.02e-20
C11021 a_14113_42308# a_18220_42308# 1.46e-20
C11022 a_5934_30871# a_n3565_39590# 6.35e-21
C11023 a_6851_47204# VDD 0.287724f
C11024 a_743_42282# CAL_N 4.51e-19
C11025 a_13467_32519# VDAC_N 3.73e-19
C11026 a_n2661_46634# a_n1641_46494# 6.71e-19
C11027 a_n2293_46634# a_n1853_46287# 0.014216f
C11028 a_n2312_38680# a_n2293_46098# 0.003636f
C11029 a_n2104_46634# a_n2157_46122# 0.013135f
C11030 a_3877_44458# a_765_45546# 0.001935f
C11031 a_6755_46942# a_15227_44166# 0.288173f
C11032 a_10428_46928# a_10425_46660# 2.36e-20
C11033 a_19386_47436# a_10809_44734# 9.09e-19
C11034 a_20894_47436# a_6945_45028# 0.016564f
C11035 a_13507_46334# a_19900_46494# 0.005187f
C11036 a_4883_46098# a_19335_46494# 0.007327f
C11037 a_12465_44636# a_18985_46122# 7.56e-21
C11038 a_11453_44696# a_17715_44484# 0.036977f
C11039 a_n881_46662# a_9569_46155# 2.93e-20
C11040 a_8128_46384# a_8199_44636# 3.12e-19
C11041 a_10037_47542# a_8016_46348# 3.96e-20
C11042 a_9804_47204# a_8349_46414# 3.47e-20
C11043 a_n2017_45002# a_20573_43172# 1.71e-20
C11044 a_n2472_43914# a_n4318_39304# 0.001031f
C11045 a_14539_43914# a_16664_43396# 0.001335f
C11046 a_n2661_43922# a_8685_43396# 4.82e-20
C11047 a_n356_44636# a_16137_43396# 0.001161f
C11048 a_13249_42308# a_13657_42308# 1.5e-19
C11049 a_7281_43914# a_7499_43940# 0.08213f
C11050 a_9672_43914# a_9895_44260# 0.011458f
C11051 a_9313_44734# a_14205_43396# 9.81e-20
C11052 a_10193_42453# a_18727_42674# 0.003839f
C11053 a_18326_43940# a_19478_44306# 3.31e-20
C11054 a_18451_43940# a_15493_43396# 2.04e-20
C11055 a_12429_44172# a_11341_43940# 0.001958f
C11056 a_18248_44752# a_18783_43370# 4.75e-20
C11057 a_18443_44721# a_18429_43548# 4.83e-19
C11058 a_3422_30871# VDD 1.12305f
C11059 a_11823_42460# a_13249_42308# 0.360411f
C11060 a_13163_45724# a_13527_45546# 0.124682f
C11061 a_9049_44484# a_10907_45822# 9.64e-21
C11062 a_2711_45572# a_8696_44636# 0.02621f
C11063 a_10053_45546# a_10210_45822# 0.18824f
C11064 a_8162_45546# a_8120_45572# 0.005491f
C11065 C2_N_btm C10_P_btm 3.9e-19
C11066 C0_dummy_P_btm C6_P_btm 0.1194f
C11067 C1_N_btm C9_P_btm 5.29e-19
C11068 C0_N_btm C8_P_btm 3.87e-19
C11069 C0_dummy_N_btm C7_P_btm 2.05e-19
C11070 C7_N_btm EN_VIN_BSTR_N 0.115875f
C11071 C0_P_btm C5_P_btm 0.138093f
C11072 C1_P_btm C4_P_btm 0.128167f
C11073 a_16241_44734# a_16375_45002# 1.69e-19
C11074 a_n2661_42834# a_n2293_45546# 4.84e-20
C11075 a_18204_44850# a_13259_45724# 1.43e-19
C11076 a_n2661_43922# a_n2956_38216# 2.48e-19
C11077 a_9028_43914# a_5937_45572# 2.88e-19
C11078 a_9672_43914# a_8199_44636# 0.043804f
C11079 a_10729_43914# a_8016_46348# 0.006537f
C11080 a_18083_42858# a_16327_47482# 0.591108f
C11081 a_15567_42826# a_10227_46804# 0.008041f
C11082 a_21356_42826# a_12861_44030# 1.38e-20
C11083 a_5193_43172# a_4791_45118# 8.86e-20
C11084 a_3080_42308# a_3090_45724# 0.002565f
C11085 a_13467_32519# a_21588_30879# 0.057457f
C11086 a_2698_46116# a_3699_46348# 6.47e-20
C11087 a_2804_46116# a_3483_46348# 4.05e-19
C11088 a_15227_44166# a_8049_45260# 0.036339f
C11089 a_12251_46660# a_12638_46436# 2.72e-19
C11090 a_11415_45002# a_13759_46122# 7.28e-21
C11091 a_1823_45246# a_5068_46348# 9.64e-20
C11092 a_20411_46873# a_6945_45028# 1.76e-19
C11093 a_17639_46660# a_17715_44484# 3.97e-19
C11094 a_20273_46660# a_21137_46414# 0.007288f
C11095 a_20841_46902# a_20708_46348# 3.45e-19
C11096 a_19551_46910# a_10809_44734# 0.006863f
C11097 a_5934_30871# a_3726_37500# 0.002188f
C11098 a_5932_42308# VDAC_P 0.009985f
C11099 a_11341_43940# a_21855_43396# 0.005468f
C11100 a_3499_42826# a_3681_42891# 0.033957f
C11101 a_9313_44734# a_22400_42852# 0.007141f
C11102 a_n356_44636# a_n784_42308# 0.084978f
C11103 a_15493_43940# a_13467_32519# 1.32e-20
C11104 a_n2109_47186# DATA[2] 0.05382f
C11105 SMPL_ON_P CLK_DATA 0.200962f
C11106 a_n1741_47186# DATA[0] 0.051737f
C11107 a_n2017_45002# a_n2956_37592# 2.81e-19
C11108 a_3357_43084# a_2382_45260# 0.219664f
C11109 a_20447_31679# a_413_45260# 0.226658f
C11110 a_n2109_45247# en_comp 0.108653f
C11111 a_n2293_45010# a_n967_45348# 0.018659f
C11112 a_n913_45002# a_n745_45366# 0.002509f
C11113 a_16211_45572# a_1307_43914# 1.74e-19
C11114 a_16147_45260# a_15415_45028# 6.7e-19
C11115 a_7499_43078# a_11827_44484# 0.104754f
C11116 a_6472_45840# a_n2661_44458# 1.35e-20
C11117 a_14209_32519# a_4185_45028# 0.091175f
C11118 a_4921_42308# a_n2293_46634# 4.37e-20
C11119 a_743_42282# a_8199_44636# 0.036554f
C11120 a_17324_43396# a_17715_44484# 0.002059f
C11121 a_17499_43370# a_18189_46348# 2.45e-20
C11122 a_18907_42674# a_13507_46334# 0.202065f
C11123 a_13258_32519# a_18479_47436# 1.35e-21
C11124 a_19511_42282# a_18597_46090# 0.156698f
C11125 a_21167_46155# VDD 8.63e-19
C11126 a_8162_45546# a_n881_46662# 1.32e-20
C11127 a_14495_45572# a_11453_44696# 7.3e-20
C11128 a_15765_45572# a_12861_44030# 0.026773f
C11129 a_8696_44636# a_9313_45822# 4.84e-20
C11130 a_n1925_42282# a_n755_45592# 0.020368f
C11131 a_n97_42460# a_15597_42852# 0.004581f
C11132 a_10807_43548# a_5742_30871# 0.020937f
C11133 a_14401_32519# a_14097_32519# 0.051264f
C11134 a_10341_43396# a_18083_42858# 5.86e-20
C11135 a_10249_46116# CLK 0.063525f
C11136 a_n2302_37984# a_n2216_37984# 0.011479f
C11137 a_18504_43218# VDD 0.077608f
C11138 a_9482_43914# a_13076_44458# 0.103066f
C11139 a_13348_45260# a_13720_44458# 2.46e-19
C11140 a_1423_45028# a_4743_44484# 0.022983f
C11141 a_1307_43914# a_5883_43914# 0.289388f
C11142 a_13556_45296# a_12883_44458# 8.08e-20
C11143 a_2711_45572# a_20365_43914# 7.09e-19
C11144 a_20841_45814# a_17517_44484# 4.23e-21
C11145 a_n2661_45010# a_n2661_42834# 0.01412f
C11146 a_15279_43071# a_n443_42852# 8.83e-21
C11147 a_20922_43172# a_n357_42282# 0.059485f
C11148 a_n2104_42282# a_n2956_38680# 2.5e-20
C11149 a_n3674_38216# a_n2956_39304# 0.023505f
C11150 VREF_GND VDD 0.482759f
C11151 a_11652_45724# a_11415_45002# 0.128811f
C11152 a_5907_45546# a_3483_46348# 6.03e-20
C11153 a_3775_45552# a_1823_45246# 0.070347f
C11154 a_4099_45572# a_4185_45028# 0.025863f
C11155 a_18479_45785# a_3090_45724# 0.259218f
C11156 a_5837_45348# a_5807_45002# 0.003033f
C11157 a_14797_45144# a_n743_46660# 2.35e-21
C11158 a_2382_45260# a_3877_44458# 0.395451f
C11159 a_2437_43646# a_6755_46942# 2.3e-19
C11160 a_413_45260# a_4817_46660# 1.37e-20
C11161 a_n2017_45002# a_5257_43370# 2.04e-19
C11162 a_2711_45572# a_4704_46090# 1.41e-19
C11163 a_n2661_43370# a_n1613_43370# 0.05744f
C11164 a_17719_45144# a_11453_44696# 0.105851f
C11165 a_18494_42460# a_4883_46098# 4.26e-20
C11166 a_20193_45348# a_18479_47436# 0.021013f
C11167 a_9838_44484# a_4791_45118# 1.34e-19
C11168 a_16977_43638# a_4958_30871# 7.21e-20
C11169 a_16409_43396# a_17303_42282# 7.54e-20
C11170 a_12379_42858# a_n784_42308# 1.29e-20
C11171 a_3681_42891# a_3318_42354# 0.001606f
C11172 a_4361_42308# a_11323_42473# 0.009186f
C11173 a_743_42282# a_13070_42354# 0.007989f
C11174 a_12281_43396# a_7174_31319# 4.88e-21
C11175 a_13467_32519# a_5742_30871# 0.004687f
C11176 a_18249_42858# a_19326_42852# 1.46e-19
C11177 a_19987_42826# a_20256_43172# 0.043356f
C11178 a_16137_43396# a_18727_42674# 0.007994f
C11179 a_8049_45260# EN_OFFSET_CAL 1.15e-20
C11180 a_n1741_47186# a_3524_46660# 1.63e-20
C11181 a_n237_47217# a_1799_45572# 0.417887f
C11182 a_2063_45854# a_948_46660# 4.3e-21
C11183 a_n1151_42308# a_171_46873# 6.23e-19
C11184 a_n746_45260# a_n2661_46098# 0.049386f
C11185 a_2124_47436# a_1983_46706# 5.47e-20
C11186 a_584_46384# a_2107_46812# 0.007756f
C11187 a_n971_45724# a_2443_46660# 0.004065f
C11188 a_3815_47204# a_n743_46660# 3.77e-20
C11189 a_4700_47436# a_n1925_46634# 7e-21
C11190 a_10227_46804# a_9804_47204# 4.77e-19
C11191 a_4915_47217# a_n2293_46634# 5.93e-19
C11192 a_6151_47436# a_n2661_46634# 0.140541f
C11193 a_n1435_47204# a_5807_45002# 3.71e-20
C11194 a_16327_47482# a_12549_44172# 0.123271f
C11195 a_15673_47210# a_15928_47570# 0.064178f
C11196 en_comp a_17538_32519# 8.81e-20
C11197 a_n1059_45260# a_n2129_43609# 0.005575f
C11198 a_n2661_45010# a_n1352_43396# 8.59e-22
C11199 a_n913_45002# a_n2433_43396# 5.3e-22
C11200 a_5111_44636# a_9801_43940# 2.57e-20
C11201 a_5205_44484# a_6671_43940# 0.049504f
C11202 a_n2017_45002# a_n2267_43396# 0.033995f
C11203 a_1307_43914# a_12495_44260# 3.12e-19
C11204 a_8783_44734# a_n2661_43922# 5.11e-21
C11205 a_13556_45296# a_15037_44260# 0.001318f
C11206 a_9313_44734# a_9159_44484# 0.056359f
C11207 a_16979_44734# a_17325_44484# 0.013377f
C11208 a_14537_43396# a_14021_43940# 0.048774f
C11209 a_n2661_44458# a_n2472_43914# 0.002397f
C11210 a_15004_44636# a_11967_42832# 3.52e-21
C11211 a_19963_31679# VDD 0.605279f
C11212 a_18175_45572# a_18051_46116# 2.57e-19
C11213 a_2437_43646# a_8049_45260# 0.041161f
C11214 a_n2810_45028# a_n1925_42282# 2.5e-20
C11215 a_13348_45260# a_13351_46090# 1.28e-19
C11216 a_1423_45028# a_8016_46348# 1.1e-20
C11217 a_13777_45326# a_10903_43370# 3.61e-19
C11218 a_9482_43914# a_12594_46348# 5.94e-21
C11219 a_8953_45002# a_2324_44458# 1.65784f
C11220 a_10405_44172# a_10227_46804# 0.011223f
C11221 a_19328_44172# a_12861_44030# 1.89e-19
C11222 a_13490_45067# a_11415_45002# 0.002913f
C11223 a_n2661_43370# a_n2293_46098# 0.027372f
C11224 a_21359_45002# a_20273_46660# 7.05e-22
C11225 a_10057_43914# a_3090_45724# 0.230475f
C11226 a_n984_44318# a_768_44030# 3.28e-20
C11227 a_19113_45348# a_19123_46287# 1.62e-19
C11228 a_20512_43084# a_19321_45002# 1.07e-19
C11229 a_22400_42852# a_22397_42558# 0.001581f
C11230 a_n1630_35242# a_4958_30871# 0.036823f
C11231 a_8325_42308# a_8791_42308# 0.173196f
C11232 C10_P_btm C8_P_btm 2.07867f
C11233 a_n743_46660# a_14976_45028# 0.024461f
C11234 a_5807_45002# a_13885_46660# 0.014137f
C11235 a_6540_46812# a_7577_46660# 3.44e-19
C11236 a_12549_44172# a_16434_46987# 6.15e-19
C11237 a_8128_46384# a_765_45546# 0.03129f
C11238 a_11453_44696# a_22365_46825# 0.001094f
C11239 a_21811_47423# a_12741_44636# 1.79e-20
C11240 a_13507_46334# a_21297_46660# 5.92e-19
C11241 a_21496_47436# a_21076_30879# 1.39e-19
C11242 a_4915_47217# a_9625_46129# 5.76e-20
C11243 a_6151_47436# a_8199_44636# 0.0013f
C11244 a_n1151_42308# a_10903_43370# 7.29e-19
C11245 a_20835_44721# a_14021_43940# 6.15e-21
C11246 a_22315_44484# a_15493_43940# 6.3e-21
C11247 a_20512_43084# a_20623_43914# 2.29e-20
C11248 a_n2661_44458# a_10695_43548# 9.47e-21
C11249 a_17719_45144# a_17324_43396# 1.66e-20
C11250 a_16922_45042# a_18783_43370# 1.97e-21
C11251 a_n356_44636# a_3080_42308# 0.072716f
C11252 a_3905_42865# a_n2661_42282# 3.49e-20
C11253 a_n913_45002# a_21356_42826# 7.3e-21
C11254 a_3232_43370# a_10341_42308# 2.53e-19
C11255 a_7640_43914# VDD 0.196713f
C11256 a_n4209_38502# C9_P_btm 3.26e-20
C11257 a_5907_45546# a_6472_45840# 0.041762f
C11258 a_5263_45724# a_6511_45714# 6.81e-21
C11259 a_2711_45572# a_7227_45028# 0.014767f
C11260 a_2998_44172# a_n2293_46098# 2.44e-19
C11261 a_17730_32519# a_4185_45028# 0.097949f
C11262 a_14021_43940# a_3090_45724# 0.049176f
C11263 a_10341_43396# a_12549_44172# 0.0385f
C11264 a_6452_43396# a_n2293_46634# 0.00445f
C11265 a_15682_43940# a_13059_46348# 9.48e-20
C11266 a_15004_44636# a_13259_45724# 6.12e-19
C11267 a_n2661_44458# a_n357_42282# 0.031616f
C11268 a_n1177_44458# a_n1079_45724# 6.5e-20
C11269 a_n1352_44484# a_n2293_45546# 1.39e-19
C11270 a_949_44458# a_n2661_45546# 1.19e-19
C11271 a_17517_44484# a_17957_46116# 2.11e-21
C11272 a_18204_44850# a_18189_46348# 2.34e-20
C11273 a_21259_43561# a_18597_46090# 0.005266f
C11274 a_5534_30871# w_1575_34946# 0.001804f
C11275 a_18909_45814# START 2.56e-21
C11276 a_19963_31679# a_22469_39537# 4.14e-20
C11277 a_n4209_39304# a_n3565_38216# 0.02945f
C11278 a_n3565_39304# a_n4209_38216# 0.02863f
C11279 a_4651_46660# VDD 0.457722f
C11280 a_14035_46660# a_3483_46348# 0.007996f
C11281 a_22000_46634# a_12741_44636# 0.044691f
C11282 a_21188_46660# a_22959_46660# 8.11e-21
C11283 a_4646_46812# a_8034_45724# 0.014576f
C11284 a_768_44030# a_3503_45724# 1.76e-21
C11285 a_5732_46660# a_5066_45546# 3.6e-22
C11286 a_5257_43370# a_526_44458# 0.003403f
C11287 a_n743_46660# a_18051_46116# 1.36e-19
C11288 a_14084_46812# a_10903_43370# 1.67e-21
C11289 a_12991_46634# a_13351_46090# 0.011685f
C11290 a_12816_46660# a_12594_46348# 1.63e-20
C11291 en_comp a_22465_38105# 0.533581f
C11292 a_n2810_45028# a_n4315_30879# 0.02588f
C11293 a_18114_32519# a_22400_42852# 1.47e-20
C11294 a_3737_43940# a_3626_43646# 7.51e-19
C11295 a_15493_43396# a_9145_43396# 1.4e-20
C11296 a_10807_43548# a_10849_43646# 0.003445f
C11297 a_9313_44734# a_22223_42860# 0.012144f
C11298 a_n4318_39304# a_n2433_43396# 6.19e-19
C11299 a_n2840_43370# a_n2129_43609# 0.001183f
C11300 a_14955_43940# a_14955_43396# 0.012141f
C11301 a_12429_44172# a_10341_43396# 9.54e-20
C11302 a_11322_45546# a_9482_43914# 8.92e-20
C11303 a_11823_42460# a_11787_45002# 0.217891f
C11304 a_11962_45724# a_13017_45260# 6.79e-20
C11305 a_18175_45572# a_19365_45572# 2.56e-19
C11306 a_6977_45572# a_6171_45002# 0.001188f
C11307 a_18451_43940# a_n357_42282# 4.34e-22
C11308 a_n2129_43609# a_n1925_42282# 5.05e-20
C11309 COMP_P a_n1613_43370# 0.001404f
C11310 VDAC_N VCM 11.7445f
C11311 a_9145_43396# a_3483_46348# 2.59e-19
C11312 a_16547_43609# a_12741_44636# 3.38e-20
C11313 a_20356_42852# a_12549_44172# 9.25e-21
C11314 VDAC_P VREF 0.008793f
C11315 a_n1379_46482# VDD 1.08e-19
C11316 a_2711_45572# a_15507_47210# 5.18e-21
C11317 a_11962_45724# a_2063_45854# 0.011034f
C11318 a_8746_45002# a_n1151_42308# 6.07e-20
C11319 a_8568_45546# a_4791_45118# 2.1e-20
C11320 a_1823_45246# a_3218_45724# 0.002867f
C11321 a_167_45260# a_1848_45724# 0.359783f
C11322 a_2698_46116# a_n755_45592# 1.12e-19
C11323 a_n2293_46098# a_2307_45899# 3.74e-19
C11324 a_22959_46124# a_8049_45260# 0.003236f
C11325 a_13759_46122# a_13259_45724# 7.02e-19
C11326 a_13925_46122# a_14383_46116# 0.027606f
C11327 a_5013_44260# a_5267_42460# 1.11e-21
C11328 a_18783_43370# a_15743_43084# 0.303966f
C11329 a_14955_43396# a_5649_42852# 3.11e-21
C11330 a_10341_43396# a_21855_43396# 0.011519f
C11331 a_n97_42460# a_18083_42858# 0.010531f
C11332 a_3626_43646# a_8387_43230# 3.45e-20
C11333 a_2982_43646# a_8952_43230# 9.76e-21
C11334 a_n2661_42282# a_n961_42308# 2.77e-19
C11335 a_22612_30879# VREF_GND 0.168163f
C11336 a_21588_30879# VCM 0.179761f
C11337 a_n1925_46634# DATA[2] 9.45e-20
C11338 a_n743_46660# DATA[0] 1.07e-19
C11339 a_16414_43172# VDD 0.201389f
C11340 a_n2810_45028# a_n3420_37440# 0.009781f
C11341 a_n2956_37592# a_n3690_37440# 0.015408f
C11342 en_comp a_19721_31679# 1.48e-19
C11343 a_n2293_45010# a_n1917_44484# 0.00169f
C11344 a_n2810_45028# a_n4318_40392# 0.026026f
C11345 a_3357_43084# a_5343_44458# 0.02588f
C11346 a_n2661_45010# a_n1352_44484# 0.051998f
C11347 a_n2956_37592# a_n2840_44458# 1.36e-20
C11348 a_n913_45002# a_n2433_44484# 1.25e-20
C11349 a_n745_45366# a_n2661_44458# 9.14e-19
C11350 a_n1059_45260# a_n2129_44697# 0.032443f
C11351 a_n2017_45002# a_n2267_44484# 0.034473f
C11352 a_8696_44636# a_9241_44734# 4.73e-19
C11353 a_13159_45002# a_13490_45067# 2.82e-19
C11354 a_14180_45002# a_14309_45348# 0.010132f
C11355 a_10193_42453# a_20679_44626# 1.62e-21
C11356 a_n1853_43023# a_n863_45724# 0.007839f
C11357 a_11136_42852# a_9290_44172# 0.001309f
C11358 a_10555_44260# CLK 9.69e-20
C11359 a_n2017_45002# a_5807_45002# 2.87e-20
C11360 a_19963_31679# a_22612_30879# 0.078731f
C11361 a_413_45260# a_11309_47204# 8.07e-21
C11362 a_3537_45260# a_n881_46662# 0.004983f
C11363 a_4574_45260# a_n1613_43370# 1.03e-20
C11364 a_11963_45334# a_11453_44696# 0.002899f
C11365 a_9482_43914# a_12465_44636# 0.069673f
C11366 a_13777_45326# a_4883_46098# 4.67e-21
C11367 a_n2661_43370# a_4791_45118# 0.408007f
C11368 a_14403_45348# a_n1151_42308# 1.39e-20
C11369 a_11823_42460# a_11813_46116# 6.35e-21
C11370 a_12427_45724# a_11901_46660# 1.11e-19
C11371 a_12791_45546# a_11735_46660# 4.28e-19
C11372 a_10180_45724# a_3090_45724# 4.56e-20
C11373 a_19987_42826# a_21195_42852# 4.49e-20
C11374 a_3626_43646# a_16522_42674# 0.002817f
C11375 a_13887_32519# a_22400_42852# 0.098244f
C11376 a_8605_42826# a_9061_43230# 4.2e-19
C11377 a_8387_43230# a_8649_43218# 0.001705f
C11378 a_n4318_39304# a_n4064_40160# 0.062069f
C11379 a_20922_43172# a_21356_42826# 0.017093f
C11380 a_4361_42308# a_20753_42852# 7.12e-19
C11381 a_5937_45572# CLK 1.52e-19
C11382 a_n2497_47436# a_n1613_43370# 0.402561f
C11383 a_n2109_47186# a_3094_47243# 0.003449f
C11384 a_n1741_47186# a_4842_47570# 2.25e-19
C11385 a_n237_47217# a_2747_46873# 5.93e-20
C11386 a_n971_45724# a_7_47243# 0.005756f
C11387 a_11459_47204# a_11599_46634# 0.019787f
C11388 a_13717_47436# a_13487_47204# 0.061247f
C11389 a_n1151_42308# a_4883_46098# 0.407909f
C11390 a_7174_31319# VDD 0.669838f
C11391 a_18587_45118# a_17517_44484# 5.57e-20
C11392 a_17767_44458# a_18248_44752# 0.041822f
C11393 a_1423_45028# a_1414_42308# 0.005518f
C11394 a_4743_44484# a_6109_44484# 2.06e-20
C11395 a_4223_44672# a_8375_44464# 0.001207f
C11396 a_16979_44734# a_18287_44626# 2.91e-20
C11397 a_1307_43914# a_2889_44172# 0.02756f
C11398 a_7499_43078# a_8147_43396# 0.227361f
C11399 a_5518_44484# a_5289_44734# 6.46e-20
C11400 a_11691_44458# a_15463_44811# 7.26e-19
C11401 a_14539_43914# a_18443_44721# 2.14e-20
C11402 a_626_44172# a_2127_44172# 3.19e-20
C11403 a_375_42282# a_895_43940# 5.29e-20
C11404 a_13249_42308# a_2982_43646# 1.48e-19
C11405 a_11827_44484# a_12189_44484# 1.28e-19
C11406 a_n2017_45002# a_19478_44306# 1.53e-20
C11407 a_3232_43370# a_3499_42826# 0.339727f
C11408 a_n1059_45260# a_15493_43396# 0.044794f
C11409 a_5147_45002# a_n2661_42282# 3.8e-19
C11410 a_8325_42308# a_n357_42282# 5.17e-20
C11411 a_n2302_40160# a_n1925_42282# 4.76e-20
C11412 a_8337_42558# a_n755_45592# 0.003302f
C11413 a_10306_45572# VDD 4.3e-19
C11414 a_n2661_43922# a_768_44030# 1.9176f
C11415 a_413_45260# a_472_46348# 1.26e-19
C11416 a_327_44734# a_376_46348# 8.78e-20
C11417 a_4574_45260# a_n2293_46098# 0.001761f
C11418 a_n356_44636# a_n2438_43548# 0.082195f
C11419 a_13213_44734# a_12891_46348# 0.052195f
C11420 a_9313_44734# a_13747_46662# 4.75e-21
C11421 a_6171_45002# a_12741_44636# 0.08387f
C11422 a_n2293_43922# a_12549_44172# 0.194293f
C11423 a_5343_44458# a_3877_44458# 3.14e-20
C11424 a_13163_45724# a_12839_46116# 5.88e-19
C11425 a_2711_45572# a_2957_45546# 0.056166f
C11426 a_8192_45572# a_8049_45260# 0.008707f
C11427 a_1990_45572# a_n2661_45546# 1.2e-19
C11428 a_19431_45546# a_18819_46122# 5.53e-19
C11429 a_18691_45572# a_18985_46122# 1.16e-19
C11430 a_18341_45572# a_19335_46494# 7.48e-19
C11431 a_2437_43646# a_8953_45546# 1.66e-19
C11432 a_20637_44484# a_16327_47482# 2.95e-19
C11433 a_2998_44172# a_4791_45118# 1.23e-19
C11434 a_2889_44172# a_n443_46116# 8.63e-19
C11435 a_1184_42692# a_2351_42308# 4.23e-20
C11436 a_n784_42308# a_3823_42558# 2.06e-20
C11437 a_14635_42282# a_14456_42282# 0.172313f
C11438 a_14097_32519# a_5934_30871# 2.14e-19
C11439 a_13291_42460# a_13249_42558# 0.002309f
C11440 a_22165_42308# a_22465_38105# 1.77e-19
C11441 a_1123_46634# a_1799_45572# 0.037438f
C11442 a_383_46660# a_n2661_46098# 0.002826f
C11443 a_9804_47204# a_10467_46802# 3.93e-21
C11444 a_n881_46662# a_6969_46634# 1.79e-19
C11445 a_n1613_43370# a_6682_46987# 1.74e-19
C11446 a_n2497_47436# a_n2293_46098# 0.039224f
C11447 a_13487_47204# a_14035_46660# 0.002982f
C11448 a_6151_47436# a_765_45546# 0.191559f
C11449 a_12861_44030# a_14180_46812# 0.238709f
C11450 a_13717_47436# a_14513_46634# 1.71e-20
C11451 a_18780_47178# a_15227_44166# 2.49e-19
C11452 a_14311_47204# a_13885_46660# 2.65e-19
C11453 a_18597_46090# a_18834_46812# 0.010699f
C11454 a_18479_47436# a_19333_46634# 5.75e-19
C11455 a_10227_46804# a_19692_46634# 0.239326f
C11456 a_4883_46098# a_14084_46812# 4.58e-20
C11457 a_13507_46334# a_3090_45724# 0.020036f
C11458 a_12465_44636# a_12816_46660# 4.51e-21
C11459 a_11453_44696# a_11901_46660# 2.64e-21
C11460 a_n2293_45010# a_n1853_43023# 4.48e-20
C11461 a_2382_45260# a_743_42282# 0.023665f
C11462 a_n2293_43922# a_12429_44172# 0.006182f
C11463 a_n2661_43370# a_8791_43396# 2.79e-21
C11464 a_9313_44734# a_20269_44172# 1.88e-20
C11465 a_7754_38636# VDD 0.036155f
C11466 a_4958_30871# a_11530_34132# 0.020719f
C11467 a_5742_30871# VCM 0.211981f
C11468 a_15890_42674# RST_Z 1.6e-20
C11469 a_3602_45348# a_3316_45546# 0.001923f
C11470 a_501_45348# a_n443_42852# 1.56e-19
C11471 a_16979_44734# a_15682_46116# 1.74e-20
C11472 a_7640_43914# a_7920_46348# 5.65e-22
C11473 a_4190_30871# w_1575_34946# 0.004947f
C11474 a_17517_44484# a_11415_45002# 0.006394f
C11475 a_14673_44172# a_12741_44636# 0.178572f
C11476 a_n2661_42834# a_1138_42852# 0.024191f
C11477 a_n97_42460# a_12549_44172# 1.69e-19
C11478 a_5013_44260# a_3090_45724# 0.009874f
C11479 a_20974_43370# a_13747_46662# 6.03e-20
C11480 a_21381_43940# a_19321_45002# 3e-20
C11481 a_11173_43940# a_n2293_46634# 2.54e-19
C11482 a_n4315_30879# a_n2302_40160# 0.407166f
C11483 a_n4334_40480# a_n4064_40160# 0.43652f
C11484 a_1606_42308# C0_N_btm 0.029189f
C11485 a_5342_30871# a_11206_38545# 2.16e-20
C11486 a_18834_46812# a_19123_46287# 0.039405f
C11487 a_15227_44166# a_18285_46348# 0.097182f
C11488 a_13885_46660# a_14226_46987# 0.003464f
C11489 a_19692_46634# a_17339_46660# 8.51e-21
C11490 a_n2472_46634# a_n2956_39304# 8.55e-19
C11491 a_9804_47204# a_8034_45724# 1.12e-19
C11492 a_4646_46812# a_8016_46348# 4.3e-21
C11493 a_5385_46902# a_5497_46414# 5.03e-20
C11494 a_5167_46660# a_5204_45822# 0.002145f
C11495 a_n2293_46634# a_10809_44734# 7.76e-20
C11496 a_4883_46098# a_19240_46482# 0.002371f
C11497 a_10227_46804# a_20692_30879# 1.56e-20
C11498 a_n443_46116# a_1990_45899# 0.002313f
C11499 a_5663_43940# a_6197_43396# 1.2e-19
C11500 a_6453_43914# a_6293_42852# 0.00419f
C11501 a_11967_42832# a_16759_43396# 0.001677f
C11502 a_15493_43940# a_19319_43548# 0.36082f
C11503 a_n2661_42282# a_4093_43548# 9.71e-22
C11504 a_21115_43940# a_21205_44306# 0.004764f
C11505 a_11173_44260# a_11257_43940# 0.002303f
C11506 a_20623_43914# a_21381_43940# 1.02e-19
C11507 a_2479_44172# a_2437_43396# 5.86e-20
C11508 a_19862_44208# a_17538_32519# 7.43e-20
C11509 a_11341_43940# a_19478_44056# 2.7e-20
C11510 a_3232_43370# a_3318_42354# 1.69e-19
C11511 a_n1059_45260# a_8791_42308# 8.01e-19
C11512 a_5111_44636# a_5379_42460# 0.118194f
C11513 a_n2017_45002# a_9223_42460# 0.003774f
C11514 a_n913_45002# a_8685_42308# 0.007967f
C11515 a_10729_43914# VDD 0.681371f
C11516 a_15599_45572# a_16333_45814# 0.053479f
C11517 a_15903_45785# a_15765_45572# 0.205788f
C11518 a_17538_32519# a_4185_45028# 0.043989f
C11519 a_13460_43230# a_n2293_46634# 4.99e-21
C11520 a_19339_43156# a_13661_43548# 2.81e-20
C11521 a_n1899_43946# a_n863_45724# 9.54e-20
C11522 a_n1331_43914# a_n1079_45724# 1.3e-20
C11523 a_n1549_44318# a_n2293_45546# 4.49e-19
C11524 a_8018_44260# a_8049_45260# 5.72e-20
C11525 a_9801_43940# a_9290_44172# 0.091547f
C11526 a_n327_42558# a_n1151_42308# 1.68e-19
C11527 a_1184_42692# a_584_46384# 3.73e-20
C11528 a_n3420_37984# C4_P_btm 1.42e-19
C11529 a_n4064_37984# C6_P_btm 1.01e-19
C11530 a_n1076_46494# VDD 0.294742f
C11531 C0_dummy_N_btm C2_N_btm 7.14548f
C11532 C0_N_btm C1_N_btm 11.2332f
C11533 C0_dummy_P_btm C3_N_btm 2.08e-19
C11534 C1_P_btm C5_N_btm 8.82e-20
C11535 C0_P_btm C4_N_btm 7.74e-20
C11536 a_13258_32519# CAL_N 0.020535f
C11537 a_3699_46348# a_526_44458# 0.00137f
C11538 a_3483_46348# a_n1925_42282# 0.536704f
C11539 a_1736_39587# a_3754_38802# 1.04e-19
C11540 a_n4064_40160# a_n2946_37690# 1.87e-20
C11541 a_n4209_39590# a_n4334_37440# 2.73e-19
C11542 a_2112_39137# a_2113_38308# 0.479143f
C11543 a_n4315_30879# a_n2302_37690# 1.98e-19
C11544 a_n3565_38502# a_n2302_37984# 2.07e-19
C11545 a_9823_46155# a_6945_45028# 1.27e-20
C11546 a_15015_46420# a_2324_44458# 0.027704f
C11547 a_n356_44636# a_15764_42576# 0.012586f
C11548 a_n2293_43922# a_7227_42308# 8.6e-20
C11549 a_n2661_42834# a_7963_42308# 2.63e-21
C11550 a_3626_43646# a_15743_43084# 2.37e-19
C11551 a_19478_44306# a_19164_43230# 4.47e-20
C11552 a_11341_43940# a_17701_42308# 7.35e-20
C11553 a_2982_43646# a_19700_43370# 3.31e-20
C11554 a_9145_43396# a_10695_43548# 0.053202f
C11555 a_8685_43396# a_14955_43396# 0.111211f
C11556 a_n2840_43370# a_n2840_42826# 0.026152f
C11557 a_21496_47436# SINGLE_ENDED 0.055146f
C11558 a_4883_46098# START 2.42e-19
C11559 a_21811_47423# RST_Z 5.42e-20
C11560 a_21487_43396# VDD 0.222231f
C11561 a_13249_42308# a_14539_43914# 0.032256f
C11562 a_1667_45002# a_1423_45028# 0.0017f
C11563 a_3537_45260# a_1307_43914# 0.290878f
C11564 a_6171_45002# a_13556_45296# 0.017156f
C11565 a_413_45260# a_2304_45348# 9.35e-20
C11566 a_9145_43396# a_n357_42282# 5.37e-19
C11567 a_8423_43396# a_n755_45592# 2.83e-20
C11568 a_2437_43396# a_n443_42852# 2.27e-19
C11569 a_12545_42858# a_9290_44172# 4.43e-19
C11570 a_19339_43156# a_4185_45028# 2.91e-21
C11571 a_n2293_42282# a_1138_42852# 1.83e-20
C11572 a_15037_45618# a_13747_46662# 0.009886f
C11573 a_2711_45572# a_7715_46873# 8.9e-19
C11574 a_4099_45572# a_5257_43370# 1.01e-19
C11575 a_16842_45938# a_n881_46662# 2.49e-19
C11576 a_3357_43084# a_10227_46804# 0.305304f
C11577 a_2437_43646# a_18780_47178# 0.008266f
C11578 a_21297_45572# a_16327_47482# 6.03e-19
C11579 a_21513_45002# a_18597_46090# 0.00344f
C11580 a_413_45260# a_7227_47204# 4.35e-19
C11581 a_n913_45002# a_12861_44030# 2.55e-20
C11582 a_4574_45260# a_4791_45118# 0.091783f
C11583 a_7229_43940# a_2063_45854# 0.003495f
C11584 a_3232_43370# a_n1151_42308# 0.003308f
C11585 a_3537_45260# a_n443_46116# 0.003861f
C11586 a_n863_45724# a_1848_45724# 5.68e-20
C11587 a_n2661_45546# a_n356_45724# 0.008001f
C11588 a_380_45546# a_n755_45592# 4.05e-19
C11589 a_n1099_45572# a_n357_42282# 0.013419f
C11590 a_3626_43646# a_1606_42308# 2.02e-20
C11591 a_8037_42858# a_8387_43230# 0.225358f
C11592 a_13887_32519# a_22223_42860# 0.013362f
C11593 a_n97_42460# a_7227_42308# 0.032716f
C11594 a_7871_42858# a_8952_43230# 0.102355f
C11595 a_20749_43396# a_20922_43172# 3.92e-19
C11596 a_3080_42308# a_3823_42558# 0.016209f
C11597 a_4905_42826# a_3318_42354# 4.93e-21
C11598 a_11341_43940# a_21613_42308# 4e-22
C11599 a_22000_46634# RST_Z 3.42e-20
C11600 a_21363_46634# SINGLE_ENDED 2.03e-20
C11601 a_7754_38636# a_8912_37509# 5.52e-19
C11602 a_n3420_37440# a_n2302_37690# 1.28e-19
C11603 a_n4209_37414# a_n3607_37440# 0.002294f
C11604 a_8530_39574# a_3726_37500# 1.35509f
C11605 a_n4334_37440# a_n4251_37440# 0.007692f
C11606 a_7754_38470# a_4338_37500# 0.208284f
C11607 a_3754_38470# a_5700_37509# 0.124176f
C11608 a_n2946_37690# a_n4064_37440# 0.053228f
C11609 a_5932_42308# VDD 0.534416f
C11610 a_1209_47178# a_1239_47204# 0.264529f
C11611 a_n971_45724# a_2952_47436# 0.019506f
C11612 a_n1605_47204# a_n1151_42308# 0.001389f
C11613 a_327_47204# a_1431_47204# 1.62e-20
C11614 a_n237_47217# a_2063_45854# 0.947844f
C11615 a_n1741_47186# a_3785_47178# 0.047034f
C11616 a_n2109_47186# a_4007_47204# 0.047269f
C11617 a_20193_45348# CAL_N 8.22e-19
C11618 a_413_45260# a_22315_44484# 1.08e-20
C11619 a_2437_43646# a_895_43940# 0.025092f
C11620 a_n2661_45010# a_n1549_44318# 2.9e-20
C11621 a_n2293_45010# a_n1899_43946# 0.18948f
C11622 a_n2017_45002# a_n2065_43946# 0.045593f
C11623 a_n2840_44458# a_n2267_44484# 4.89e-19
C11624 a_8696_44636# a_15682_43940# 0.001466f
C11625 a_13556_45296# a_14673_44172# 0.137701f
C11626 a_9482_43914# a_16241_44734# 9.38e-20
C11627 a_n4318_40392# a_n2129_44697# 4.04e-19
C11628 a_n2661_44458# a_n2433_44484# 0.039874f
C11629 a_16922_45042# a_17767_44458# 2.79e-19
C11630 a_17023_45118# a_16979_44734# 1.26e-19
C11631 a_22465_38105# a_4185_45028# 0.065539f
C11632 a_9223_42460# a_526_44458# 1.63e-20
C11633 a_10775_45002# a_10768_47026# 3.67e-22
C11634 a_16751_45260# a_6755_46942# 1.98e-19
C11635 a_19929_45028# a_19321_45002# 5.38e-19
C11636 a_18114_32519# a_13747_46662# 1.55e-19
C11637 a_4927_45028# a_3090_45724# 0.088804f
C11638 a_2437_43646# a_18285_46348# 6.42e-20
C11639 a_14495_45572# a_13925_46122# 2.46e-19
C11640 a_13249_42308# a_14493_46090# 6.35e-19
C11641 a_8791_45572# a_8199_44636# 0.003441f
C11642 a_5883_43914# a_n1613_43370# 0.352323f
C11643 a_n356_44636# a_13507_46334# 2.44e-20
C11644 a_19256_45572# a_11415_45002# 0.003224f
C11645 a_5534_30871# a_13575_42558# 0.002235f
C11646 a_14543_43071# a_14456_42282# 0.009977f
C11647 a_n881_46662# a_n2293_46634# 0.026189f
C11648 a_2747_46873# a_1123_46634# 2.46e-20
C11649 a_2266_47570# a_2107_46812# 2.38e-19
C11650 a_6575_47204# a_8667_46634# 0.01088f
C11651 a_4915_47217# a_6755_46942# 0.260675f
C11652 a_6151_47436# a_10623_46897# 4.99e-20
C11653 a_2063_45854# a_8270_45546# 0.017994f
C11654 a_20567_45036# a_14021_43940# 3.06e-22
C11655 a_17517_44484# a_11967_42832# 0.342031f
C11656 a_1307_43914# a_1049_43396# 0.001373f
C11657 a_10193_42453# a_10341_42308# 0.061874f
C11658 a_375_42282# a_458_43396# 0.014454f
C11659 a_5883_43914# a_7584_44260# 1.86e-20
C11660 a_3232_43370# a_6197_43396# 6.79e-20
C11661 a_5111_44636# a_7287_43370# 0.104641f
C11662 a_3537_45260# a_9396_43370# 5.47e-19
C11663 a_1423_45028# VDD 4.06861f
C11664 a_1606_42308# C10_P_btm 1.34e-19
C11665 a_n2661_44458# a_3147_46376# 7.41e-21
C11666 a_19721_31679# a_4185_45028# 0.004653f
C11667 a_12607_44458# a_12741_44636# 0.134974f
C11668 a_13720_44458# a_11415_45002# 0.001979f
C11669 a_5883_43914# a_n2293_46098# 0.069185f
C11670 a_11341_43940# a_12891_46348# 8.37e-19
C11671 a_21115_43940# a_12549_44172# 0.211261f
C11672 a_17973_43940# a_13661_43548# 0.031319f
C11673 a_15463_44811# a_15227_44166# 4.61e-19
C11674 a_2437_43646# a_1609_45822# 0.189329f
C11675 a_n143_45144# a_n2661_45546# 8.29e-19
C11676 a_6171_45002# a_16375_45002# 0.026914f
C11677 a_n2017_45002# a_n755_45592# 0.088948f
C11678 a_n1059_45260# a_n357_42282# 7.3759f
C11679 a_n967_45348# a_n1079_45724# 4.19e-20
C11680 a_n2661_43370# a_6945_45028# 0.006001f
C11681 a_2896_43646# a_584_46384# 0.00371f
C11682 a_1049_43396# a_n443_46116# 0.085877f
C11683 a_15890_42674# a_17303_42282# 1.66e-20
C11684 a_11551_42558# a_7174_31319# 4.88e-21
C11685 a_n4318_37592# a_n3565_38216# 5.63e-19
C11686 a_6491_46660# VDD 0.436756f
C11687 a_n1151_42308# a_11608_46482# 7.22e-19
C11688 a_n2312_38680# a_n2472_46090# 0.001445f
C11689 a_n2293_46634# a_n2157_46122# 0.04308f
C11690 a_n2104_46634# a_n2293_46098# 0.002261f
C11691 a_10150_46912# a_10425_46660# 0.007416f
C11692 a_19787_47423# a_6945_45028# 0.009959f
C11693 a_18597_46090# a_10809_44734# 0.036294f
C11694 a_20990_47178# a_20708_46348# 2.85e-21
C11695 a_13507_46334# a_20075_46420# 0.006404f
C11696 a_4883_46098# a_19553_46090# 0.005361f
C11697 a_4915_47217# a_8049_45260# 0.022494f
C11698 a_12465_44636# a_18819_46122# 2.8e-20
C11699 a_11453_44696# a_17583_46090# 1.99e-20
C11700 a_n881_46662# a_9625_46129# 3.67e-20
C11701 a_8128_46384# a_8349_46414# 0.101217f
C11702 a_9804_47204# a_8016_46348# 0.009763f
C11703 a_768_44030# a_5164_46348# 4.84e-20
C11704 a_n2017_45002# a_20256_43172# 3.49e-19
C11705 a_n1059_45260# a_18707_42852# 8.57e-19
C11706 a_n2661_42834# a_8685_43396# 9.54e-20
C11707 a_5343_44458# a_743_42282# 0.010119f
C11708 a_9672_43914# a_9801_44260# 0.010132f
C11709 a_10193_42453# a_18057_42282# 0.099046f
C11710 a_18287_44626# a_18429_43548# 8.45e-21
C11711 a_9313_44734# a_14358_43442# 5.8e-20
C11712 a_18079_43940# a_19478_44306# 2.26e-20
C11713 a_18326_43940# a_15493_43396# 3.68e-20
C11714 a_11750_44172# a_11341_43940# 0.002015f
C11715 a_18451_43940# a_19328_44172# 0.008311f
C11716 a_n2840_43914# a_n4318_39304# 0.002229f
C11717 a_21398_44850# VDD 0.077608f
C11718 a_11823_42460# a_13904_45546# 0.067334f
C11719 a_7499_43078# a_10907_45822# 5.14e-19
C11720 a_9049_44484# a_10210_45822# 1.6e-20
C11721 C1_N_btm C10_P_btm 9.71e-19
C11722 C0_dummy_P_btm C7_P_btm 0.119061f
C11723 C0_N_btm C9_P_btm 4.64e-19
C11724 C0_dummy_N_btm C8_P_btm 3.42e-19
C11725 C6_N_btm EN_VIN_BSTR_N 0.118916f
C11726 C1_P_btm C5_P_btm 0.127408f
C11727 C0_P_btm C6_P_btm 0.139059f
C11728 a_4699_43561# a_3090_45724# 1.16e-20
C11729 a_18533_44260# a_17339_46660# 0.002232f
C11730 a_17517_44484# a_13259_45724# 0.028602f
C11731 a_n2661_43922# a_n2472_45546# 2.25e-19
C11732 a_n89_44484# a_n755_45592# 3.83e-19
C11733 a_8333_44056# a_5937_45572# 7.94e-19
C11734 a_10405_44172# a_8016_46348# 0.098226f
C11735 a_17701_42308# a_16327_47482# 0.001161f
C11736 a_5342_30871# a_10227_46804# 0.163388f
C11737 a_14021_43940# a_21076_30879# 1.4e-20
C11738 a_n3420_38528# C1_P_btm 5.88e-20
C11739 a_5742_30871# VDAC_Ni 3.56e-19
C11740 a_2698_46116# a_3483_46348# 1.66e-19
C11741 a_2804_46116# a_3147_46376# 0.017019f
C11742 a_12251_46660# a_12379_46436# 4.35e-19
C11743 a_3090_45724# a_10586_45546# 0.002067f
C11744 a_12741_44636# a_10903_43370# 4.89e-19
C11745 a_11415_45002# a_13351_46090# 4.86e-21
C11746 a_1823_45246# a_4704_46090# 0.164557f
C11747 a_19123_46287# a_10809_44734# 0.009463f
C11748 a_17639_46660# a_17583_46090# 3.95e-19
C11749 a_20273_46660# a_20708_46348# 0.004461f
C11750 a_20107_46660# a_6945_45028# 0.024966f
C11751 a_20411_46873# a_21137_46414# 2.11e-20
C11752 a_11341_43940# a_4361_42308# 0.001978f
C11753 a_n2661_42282# a_685_42968# 1.62e-20
C11754 a_1427_43646# a_1512_43396# 1.48e-19
C11755 a_4905_42826# a_6197_43396# 1.53e-20
C11756 a_3626_43646# a_3539_42460# 0.017877f
C11757 a_3499_42826# a_2905_42968# 0.00265f
C11758 a_18494_42460# a_15803_42450# 1.58e-20
C11759 a_14021_43940# a_17486_43762# 1.72e-19
C11760 a_9313_44734# a_20836_43172# 9.15e-20
C11761 a_n1741_47186# CLK_DATA 8.62e-20
C11762 a_n1920_47178# DATA[0] 7.82e-20
C11763 a_n2109_47186# DATA[1] 0.049689f
C11764 a_n2109_45247# a_n2956_37592# 3.33e-19
C11765 a_n2017_45002# a_n2810_45028# 1.6e-19
C11766 a_n1059_45260# a_n745_45366# 0.0613f
C11767 a_n2293_45010# en_comp 0.066194f
C11768 a_22959_45572# a_413_45260# 0.021231f
C11769 a_16147_45260# a_14797_45144# 1.1e-19
C11770 a_10193_42453# a_18494_42460# 0.074751f
C11771 a_13249_42308# a_14309_45028# 0.008249f
C11772 a_22591_43396# a_4185_45028# 0.008398f
C11773 a_n97_42460# a_n2661_45546# 0.038952f
C11774 a_17499_43370# a_17715_44484# 0.001287f
C11775 a_18727_42674# a_13507_46334# 0.093566f
C11776 a_21613_42308# a_16327_47482# 1.68e-19
C11777 a_20850_46155# VDD 6.25e-20
C11778 a_2711_45572# a_13747_46662# 0.032065f
C11779 a_7230_45938# a_n881_46662# 8.9e-20
C11780 a_8162_45546# a_n1613_43370# 1.42e-20
C11781 a_13249_42308# a_11453_44696# 0.026348f
C11782 a_15037_45618# a_11599_46634# 1.12e-19
C11783 a_15903_45785# a_12861_44030# 0.156145f
C11784 a_526_44458# a_n755_45592# 0.065199f
C11785 a_n1925_42282# a_n357_42282# 0.023161f
C11786 a_14401_32519# a_22400_42852# 8.97e-20
C11787 a_21381_43940# a_14097_32519# 1.99e-20
C11788 a_10807_43548# a_11323_42473# 0.109765f
C11789 a_10341_43396# a_17701_42308# 2.12e-19
C11790 a_10554_47026# CLK 0.014924f
C11791 a_6755_46942# DATA[5] 2.62e-19
C11792 a_n4064_37984# a_n2216_37984# 0.005565f
C11793 a_13348_45260# a_13076_44458# 4.88e-20
C11794 a_1423_45028# a_n699_43396# 0.008455f
C11795 a_1307_43914# a_8701_44490# 7.15e-21
C11796 a_9482_43914# a_12883_44458# 7.92e-20
C11797 a_13556_45296# a_12607_44458# 0.01896f
C11798 a_7499_43078# a_n2661_42282# 5.53e-21
C11799 a_2711_45572# a_20269_44172# 8.26e-19
C11800 a_3065_45002# a_4181_44734# 3.66e-20
C11801 a_5534_30871# a_n443_42852# 8.98e-20
C11802 a_19987_42826# a_n357_42282# 0.016903f
C11803 a_n2293_42282# a_n2956_38216# 2.83e-20
C11804 a_n2104_42282# a_n2956_39304# 2.99e-20
C11805 a_n4318_38216# a_n2956_38680# 0.023189f
C11806 a_2711_45572# a_4419_46090# 0.026096f
C11807 VREF VDD 4.8299f
C11808 a_11525_45546# a_11415_45002# 1.34e-19
C11809 a_5263_45724# a_3483_46348# 9.89e-20
C11810 a_18175_45572# a_3090_45724# 0.130163f
C11811 a_14537_43396# a_n743_46660# 6.18e-20
C11812 a_1307_43914# a_n2293_46634# 0.184387f
C11813 a_16147_45260# a_14976_45028# 0.001993f
C11814 a_3357_43084# a_10467_46802# 1.38e-20
C11815 a_2437_43646# a_10249_46116# 1.78e-19
C11816 a_2274_45254# a_3877_44458# 7.27e-21
C11817 a_413_45260# a_4955_46873# 2.73e-20
C11818 a_17613_45144# a_11453_44696# 3.78e-19
C11819 a_18184_42460# a_4883_46098# 6.32e-21
C11820 a_20567_45036# a_13507_46334# 2.05e-21
C11821 a_16237_45028# a_10227_46804# 7.21e-19
C11822 a_n1243_44484# a_n2497_47436# 2.69e-19
C11823 a_5883_43914# a_4791_45118# 7.11e-19
C11824 a_16409_43396# a_4958_30871# 5.65e-20
C11825 a_10341_43396# a_21613_42308# 2.29e-20
C11826 a_10341_42308# a_n784_42308# 1.87e-21
C11827 a_19164_43230# a_20256_43172# 1.29e-19
C11828 a_4361_42308# a_10723_42308# 0.010334f
C11829 a_743_42282# a_12563_42308# 0.00803f
C11830 a_16137_43396# a_18057_42282# 0.01884f
C11831 a_3080_42308# a_1177_38525# 2.16e-19
C11832 a_n443_46116# a_n2293_46634# 0.050675f
C11833 a_n1741_47186# a_3699_46634# 1.51e-19
C11834 a_584_46384# a_948_46660# 0.002817f
C11835 a_n1151_42308# a_n133_46660# 0.002432f
C11836 a_2124_47436# a_2107_46812# 0.010665f
C11837 a_n971_45724# a_n2661_46098# 0.023255f
C11838 a_3785_47178# a_n743_46660# 2.74e-21
C11839 a_4007_47204# a_n1925_46634# 8.66e-20
C11840 a_n746_45260# a_1799_45572# 4.63e-22
C11841 a_13381_47204# a_5807_45002# 5.2e-20
C11842 a_5815_47464# a_n2661_46634# 1.29e-19
C11843 a_15673_47210# a_768_44030# 2.86e-20
C11844 a_15507_47210# a_16119_47582# 3.82e-19
C11845 a_15811_47375# a_15928_47570# 0.161235f
C11846 a_3422_30871# VDAC_N 0.480156f
C11847 a_3232_43370# a_8415_44056# 1.41e-19
C11848 a_n1059_45260# a_n2433_43396# 3.64e-21
C11849 a_n2017_45002# a_n2129_43609# 0.024338f
C11850 a_8333_44734# a_n2661_43922# 1.54e-35
C11851 a_14180_45002# a_14021_43940# 2.49e-20
C11852 a_14539_43914# a_17325_44484# 2.02e-20
C11853 a_18374_44850# a_18204_44850# 2.6e-19
C11854 a_16979_44734# a_17061_44484# 0.003935f
C11855 a_9313_44734# a_10617_44484# 0.006463f
C11856 a_9241_44734# a_9159_44484# 5.37e-19
C11857 a_18989_43940# a_17517_44484# 0.021791f
C11858 a_13720_44458# a_11967_42832# 1.06e-21
C11859 a_n2661_44458# a_n2840_43914# 0.002411f
C11860 a_n2946_39866# a_n2810_45572# 4.32e-20
C11861 a_n3565_39590# a_n2956_38216# 0.021271f
C11862 a_22591_45572# VDD 0.314172f
C11863 a_20567_45036# a_20623_46660# 3.11e-20
C11864 a_10440_44484# a_3090_45724# 1.35e-20
C11865 a_n809_44244# a_768_44030# 4.27e-19
C11866 a_18341_45572# a_19240_46482# 1.94e-19
C11867 a_16147_45260# a_18051_46116# 5.51e-19
C11868 a_21513_45002# a_8049_45260# 0.007177f
C11869 a_13017_45260# a_13759_46122# 9.47e-21
C11870 a_13348_45260# a_12594_46348# 7.19e-21
C11871 a_13556_45296# a_10903_43370# 2.71e-19
C11872 a_8191_45002# a_2324_44458# 0.120399f
C11873 a_9672_43914# a_10227_46804# 6.27e-19
C11874 a_18451_43940# a_12861_44030# 0.001042f
C11875 a_2448_45028# a_167_45260# 1.54e-19
C11876 a_15685_45394# a_11415_45002# 1.56e-19
C11877 a_5934_30871# a_9377_42558# 0.001873f
C11878 a_8325_42308# a_8685_42308# 0.141819f
C11879 C10_P_btm C9_P_btm 53.3168f
C11880 a_12549_44172# a_16721_46634# 0.013883f
C11881 a_n743_46660# a_3090_45724# 0.050883f
C11882 a_5732_46660# a_7577_46660# 3.52e-20
C11883 a_6540_46812# a_7715_46873# 1.3e-19
C11884 a_5807_45002# a_13170_46660# 3.81e-19
C11885 a_5159_47243# a_765_45546# 2e-19
C11886 a_4883_46098# a_12741_44636# 0.076276f
C11887 a_n1435_47204# a_3483_46348# 1.31e-20
C11888 a_6545_47178# a_8016_46348# 4.25e-20
C11889 a_4915_47217# a_8953_45546# 1.73e-19
C11890 a_6151_47436# a_8349_46414# 1.15e-19
C11891 a_n1151_42308# a_11387_46155# 0.195225f
C11892 a_17613_45144# a_17324_43396# 4.37e-19
C11893 a_6298_44484# a_6655_43762# 5.21e-20
C11894 a_20679_44626# a_14021_43940# 2.62e-20
C11895 a_3422_30871# a_15493_43940# 0.014587f
C11896 a_22315_44484# a_22223_43948# 0.012307f
C11897 a_20512_43084# a_20365_43914# 1.4e-19
C11898 a_n356_44636# a_4699_43561# 2.33e-21
C11899 a_5883_43914# a_8791_43396# 1.82e-19
C11900 a_n2661_44458# a_9803_43646# 6.14e-21
C11901 a_17719_45144# a_17499_43370# 2.73e-21
C11902 a_18494_42460# a_16137_43396# 0.115144f
C11903 a_n913_45002# a_20922_43172# 0.010679f
C11904 en_comp a_18599_43230# 9.77e-22
C11905 a_n2017_45002# a_21195_42852# 8.32e-21
C11906 a_6109_44484# VDD 0.243629f
C11907 a_n4209_38502# C10_P_btm 2.25e-20
C11908 a_n4064_39616# VCM 0.068103f
C11909 a_5907_45546# a_6194_45824# 0.233657f
C11910 a_2711_45572# a_6598_45938# 0.011792f
C11911 a_22591_44484# a_4185_45028# 0.013394f
C11912 a_14955_43940# a_13059_46348# 0.001717f
C11913 a_10341_43396# a_12891_46348# 7.46e-20
C11914 a_9396_43370# a_n2293_46634# 0.012588f
C11915 a_n1177_44458# a_n2293_45546# 3.48e-19
C11916 a_13720_44458# a_13259_45724# 0.016851f
C11917 a_11691_44458# a_n443_42852# 4.69e-20
C11918 a_n2661_44458# a_310_45028# 0.003131f
C11919 a_10809_44484# a_10809_44734# 0.009578f
C11920 a_17517_44484# a_18189_46348# 1.78e-19
C11921 a_4190_30871# a_18479_47436# 1.1e-19
C11922 a_4361_42308# a_16327_47482# 0.029635f
C11923 a_743_42282# a_10227_46804# 0.045325f
C11924 a_18341_45572# START 7.1e-21
C11925 a_20447_31679# a_22521_39511# 3.7e-20
C11926 a_4646_46812# VDD 2.53408f
C11927 a_13885_46660# a_3483_46348# 2.24e-19
C11928 a_21188_46660# a_12741_44636# 0.052893f
C11929 a_20841_46902# a_21297_46660# 4.2e-19
C11930 a_22000_46634# a_20820_30879# 0.001417f
C11931 a_5907_46634# a_5066_45546# 9.12e-19
C11932 a_768_44030# a_3316_45546# 5.1e-21
C11933 a_n743_46660# a_15002_46116# 1.44e-19
C11934 a_12991_46634# a_12594_46348# 7.99e-21
C11935 a_6755_46942# a_10809_44734# 0.042402f
C11936 a_n881_46662# a_2277_45546# 1.72e-20
C11937 a_10807_43548# a_10765_43646# 9.53e-19
C11938 a_453_43940# a_743_42282# 8.67e-23
C11939 a_9313_44734# a_22165_42308# 0.028818f
C11940 a_n2840_43370# a_n2433_43396# 0.039807f
C11941 a_11750_44172# a_10341_43396# 2.18e-21
C11942 a_14955_43940# a_15095_43370# 1.49e-19
C11943 a_19256_45572# a_20273_45572# 1.1e-19
C11944 a_11962_45724# a_11963_45334# 0.006674f
C11945 a_11823_42460# a_10951_45334# 8.18e-20
C11946 a_17568_45572# a_17668_45572# 0.005294f
C11947 a_11322_45546# a_13348_45260# 4.97e-20
C11948 a_11652_45724# a_13017_45260# 8.37e-21
C11949 a_18479_45785# a_20528_45572# 7.66e-21
C11950 a_6905_45572# a_6171_45002# 5.84e-19
C11951 a_743_42282# a_17339_46660# 4.84e-20
C11952 a_8333_44056# a_n443_42852# 3.11e-19
C11953 a_18326_43940# a_n357_42282# 6.84e-21
C11954 a_n2433_43396# a_n1925_42282# 0.001028f
C11955 a_6655_43762# a_5937_45572# 8.87e-19
C11956 VDAC_N VREF_GND 0.203821f
C11957 a_16243_43396# a_12741_44636# 5.87e-20
C11958 a_n1545_46494# VDD 1.74e-19
C11959 a_2711_45572# a_11599_46634# 0.018466f
C11960 a_4880_45572# a_6151_47436# 9.96e-20
C11961 a_10193_42453# a_n1151_42308# 0.238612f
C11962 a_11652_45724# a_2063_45854# 0.002983f
C11963 a_8162_45546# a_4791_45118# 3.59e-20
C11964 a_1823_45246# a_2957_45546# 0.009473f
C11965 a_167_45260# a_997_45618# 0.052039f
C11966 a_2521_46116# a_n755_45592# 3.63e-20
C11967 a_n2293_46098# a_1990_45899# 6.77e-19
C11968 a_10809_44734# a_8049_45260# 0.059599f
C11969 a_13759_46122# a_14383_46116# 9.73e-19
C11970 a_13351_46090# a_13259_45724# 7.81e-20
C11971 a_14275_46494# a_14537_46482# 0.001705f
C11972 a_14493_46090# a_14949_46494# 4.2e-19
C11973 a_5204_45822# a_n2661_45546# 5.48e-19
C11974 a_5244_44056# a_5267_42460# 1.4e-21
C11975 a_18525_43370# a_15743_43084# 0.058072f
C11976 a_10341_43396# a_4361_42308# 0.027045f
C11977 a_n97_42460# a_17701_42308# 0.001768f
C11978 a_2982_43646# a_9127_43156# 2.28e-19
C11979 a_3499_42826# a_n784_42308# 4.32e-21
C11980 a_3905_42865# a_5379_42460# 1.34e-20
C11981 a_3626_43646# a_8605_42826# 2.77e-20
C11982 a_n2661_42282# a_n1329_42308# 2.6e-19
C11983 a_16759_43396# a_16867_43762# 0.057222f
C11984 a_16137_43396# a_15940_43402# 4.65e-19
C11985 a_3422_30871# a_5742_30871# 0.029732f
C11986 a_20974_43370# a_22165_42308# 8.68e-20
C11987 a_14401_32519# a_22223_42860# 8.04e-20
C11988 a_21588_30879# VREF_GND 0.083908f
C11989 a_22612_30879# VREF 1.73216f
C11990 a_n1925_46634# DATA[1] 4.06e-21
C11991 a_n2661_46634# CLK 0.032279f
C11992 a_15567_42826# VDD 0.163583f
C11993 a_n2810_45028# a_n3690_37440# 5.77e-19
C11994 a_n2956_37592# a_n3565_37414# 0.304738f
C11995 en_comp a_18114_32519# 1.07e-19
C11996 a_n2293_45010# a_n1699_44726# 0.005129f
C11997 a_3357_43084# a_4743_44484# 2.98e-20
C11998 a_n1059_45260# a_n2433_44484# 3e-21
C11999 a_n2661_45010# a_n1177_44458# 0.052759f
C12000 a_n2810_45028# a_n2840_44458# 4.31e-19
C12001 a_n913_45002# a_n2661_44458# 0.024357f
C12002 a_n2017_45002# a_n2129_44697# 0.033299f
C12003 a_n2109_45247# a_n2267_44484# 3.19e-19
C12004 a_8696_44636# a_8855_44734# 2.74e-19
C12005 a_17668_45572# a_17767_44458# 7.33e-21
C12006 a_n4209_38216# a_n2312_38680# 2.66e-20
C12007 a_n2157_42858# a_n863_45724# 7.79e-21
C12008 a_13157_43218# a_9290_44172# 8.98e-21
C12009 a_11823_42460# a_11735_46660# 6.67e-20
C12010 a_11962_45724# a_11901_46660# 3.74e-20
C12011 a_19963_31679# a_21588_30879# 0.055898f
C12012 a_3429_45260# a_n881_46662# 1.13e-19
C12013 a_3537_45260# a_n1613_43370# 0.095192f
C12014 a_11787_45002# a_11453_44696# 0.005756f
C12015 a_13348_45260# a_12465_44636# 1.39e-21
C12016 a_14180_45002# a_13507_46334# 1.58e-22
C12017 a_8560_45348# a_6151_47436# 1.29e-20
C12018 a_5649_42852# a_14097_32519# 1.23e-20
C12019 a_n4318_39304# a_n4334_40480# 3.36e-19
C12020 a_8037_42858# a_9061_43230# 2.36e-20
C12021 a_8605_42826# a_8649_43218# 3.69e-19
C12022 a_2982_43646# a_17124_42282# 3.02e-19
C12023 a_19164_43230# a_21195_42852# 3.2e-21
C12024 a_7871_42858# a_8495_42852# 9.73e-19
C12025 a_22223_43396# a_22400_42852# 4.88e-19
C12026 a_13467_32519# a_20753_42852# 1.97e-19
C12027 a_8199_44636# CLK 0.231904f
C12028 a_20712_42282# VDD 0.282526f
C12029 a_n971_45724# a_n310_47243# 0.007307f
C12030 a_n452_47436# a_7_47243# 6.64e-19
C12031 a_6151_47436# a_10227_46804# 0.032659f
C12032 a_13717_47436# a_12861_44030# 0.319645f
C12033 a_n1435_47204# a_13487_47204# 0.135076f
C12034 a_3160_47472# a_4883_46098# 1.62e-19
C12035 a_2711_45572# a_14358_43442# 1.67e-21
C12036 a_17767_44458# a_17970_44736# 0.233657f
C12037 a_14539_43914# a_18287_44626# 3.64e-20
C12038 a_1307_43914# a_2675_43914# 0.453622f
C12039 a_626_44172# a_453_43940# 0.163589f
C12040 a_4223_44672# a_7640_43914# 0.002847f
C12041 a_7499_43078# a_7112_43396# 0.012965f
C12042 a_11827_44484# a_11909_44484# 0.00995f
C12043 a_n2661_44458# a_556_44484# 1.56e-19
C12044 a_5518_44484# a_5205_44734# 3.77e-20
C12045 a_11691_44458# a_15146_44811# 0.002578f
C12046 a_n2017_45002# a_15493_43396# 6.52e-20
C12047 a_5147_45002# a_6101_44260# 3.6e-20
C12048 a_4169_42308# a_n755_45592# 1.51e-19
C12049 a_10216_45572# VDD 4.83e-19
C12050 a_5534_30871# CAL_P 0.006743f
C12051 a_n2661_42834# a_768_44030# 4.99505f
C12052 a_n356_44636# a_n743_46660# 4.32e-20
C12053 a_413_45260# a_376_46348# 1.85e-19
C12054 a_3537_45260# a_n2293_46098# 0.019207f
C12055 a_n2661_43922# a_12549_44172# 0.061277f
C12056 a_9313_44734# a_13661_43548# 3.79e-19
C12057 a_3232_43370# a_12741_44636# 4.67e-19
C12058 a_n2293_43922# a_12891_46348# 8.04e-19
C12059 a_12791_45546# a_12839_46116# 2.39e-19
C12060 a_4099_45572# a_n755_45592# 0.001267f
C12061 a_8120_45572# a_8049_45260# 0.0028f
C12062 a_3733_45822# a_n2661_45546# 1.54e-35
C12063 a_18691_45572# a_18819_46122# 5.44e-20
C12064 a_3357_43084# a_8016_46348# 1.25e-21
C12065 a_2437_43646# a_5937_45572# 3.38e-20
C12066 a_17325_44484# a_11453_44696# 1.07e-19
C12067 a_18579_44172# a_18597_46090# 9.48e-21
C12068 a_20397_44484# a_16327_47482# 0.001966f
C12069 a_2675_43914# a_n443_46116# 0.011921f
C12070 a_1184_42692# a_2123_42473# 0.107417f
C12071 a_961_42354# a_1755_42282# 3.85e-19
C12072 a_n784_42308# a_3318_42354# 1.96e-20
C12073 a_13291_42460# a_14456_42282# 0.015899f
C12074 a_14635_42282# a_13575_42558# 5.53e-19
C12075 a_22165_42308# a_22397_42558# 8.87e-19
C12076 a_n743_46660# a_3699_46634# 1.08e-19
C12077 a_383_46660# a_1799_45572# 2.74e-20
C12078 a_601_46902# a_n2661_46098# 0.003957f
C12079 a_n1925_46634# a_2864_46660# 0.004284f
C12080 a_n2438_43548# a_2959_46660# 3.53e-20
C12081 a_9804_47204# a_10428_46928# 3.61e-20
C12082 a_n881_46662# a_6755_46942# 0.063288f
C12083 a_13487_47204# a_13885_46660# 0.002202f
C12084 a_5815_47464# a_765_45546# 0.01398f
C12085 a_13717_47436# a_14180_46812# 1e-20
C12086 a_12861_44030# a_14035_46660# 0.153051f
C12087 a_18780_47178# a_18834_46812# 0.010748f
C12088 a_18479_47436# a_15227_44166# 0.199537f
C12089 a_10227_46804# a_19466_46812# 1.18e-19
C12090 a_18597_46090# a_17609_46634# 8.28e-19
C12091 a_13507_46334# a_15009_46634# 7.3e-20
C12092 a_11453_44696# a_11813_46116# 5.74e-21
C12093 a_n1613_43370# a_6969_46634# 3.94e-19
C12094 a_n2661_45010# a_n1991_42858# 6.37e-20
C12095 en_comp a_13887_32519# 8.37e-20
C12096 a_n2293_45010# a_n2157_42858# 3.31e-20
C12097 a_9313_44734# a_19862_44208# 0.024263f
C12098 a_n2661_43922# a_12429_44172# 0.004259f
C12099 a_5742_30871# VREF_GND 0.191352f
C12100 a_15959_42545# RST_Z 3.5e-20
C12101 a_5244_44056# a_3090_45724# 0.002228f
C12102 a_10867_43940# a_n2293_46634# 7.16e-19
C12103 a_22959_45036# a_8049_45260# 0.002194f
C12104 a_375_42282# a_n443_42852# 0.075658f
C12105 a_3495_45348# a_3316_45546# 0.004904f
C12106 a_n2129_44697# a_526_44458# 4.74e-20
C12107 a_14539_43914# a_15682_46116# 2.11e-19
C12108 a_5883_43914# a_6945_45028# 1.46e-20
C12109 a_9145_43396# a_12861_44030# 1.84e-19
C12110 a_17517_44484# a_20202_43084# 0.021286f
C12111 a_9313_44734# a_4185_45028# 0.078424f
C12112 a_14581_44484# a_12741_44636# 2.79e-20
C12113 a_9804_47204# VDD 0.410522f
C12114 a_n4315_30879# a_n4064_40160# 0.363059f
C12115 a_n784_42308# C10_N_btm 1.34e-19
C12116 a_1606_42308# C0_dummy_N_btm 0.007541f
C12117 a_18834_46812# a_18285_46348# 0.144972f
C12118 a_13885_46660# a_14513_46634# 0.101344f
C12119 a_14035_46660# a_14180_46812# 0.00994f
C12120 a_15227_44166# a_17829_46910# 1.41e-19
C12121 a_17609_46634# a_19123_46287# 1.84e-20
C12122 a_19466_46812# a_17339_46660# 1.16e-20
C12123 a_768_44030# a_5066_45546# 2.81e-20
C12124 a_n2956_39768# a_n2956_38680# 0.043291f
C12125 a_n2661_46634# a_n2956_39304# 4.64e-19
C12126 a_9804_47204# a_8283_46482# 3.67e-21
C12127 a_n881_46662# a_8049_45260# 0.025172f
C12128 a_8128_46384# a_8034_45724# 0.003967f
C12129 a_4646_46812# a_7920_46348# 2.09e-20
C12130 a_4817_46660# a_5497_46414# 0.001967f
C12131 a_5167_46660# a_5164_46348# 0.003259f
C12132 a_5385_46902# a_5204_45822# 1.84e-20
C12133 a_4883_46098# a_16375_45002# 0.01007f
C12134 a_13507_46334# a_19431_46494# 0.001128f
C12135 a_18479_47436# a_21071_46482# 5.89e-19
C12136 a_n443_46116# a_2277_45546# 0.048113f
C12137 a_5534_30871# CAL_N 0.004303f
C12138 a_5342_30871# VDAC_P 0.007533f
C12139 a_5663_43940# a_6293_42852# 7.17e-19
C12140 a_6453_43914# a_6031_43396# 0.001451f
C12141 a_1414_42308# a_3457_43396# 0.094207f
C12142 a_11967_42832# a_16977_43638# 0.001333f
C12143 a_19862_44208# a_20974_43370# 0.026213f
C12144 a_n356_44636# a_1847_42826# 3.12e-20
C12145 a_3499_42826# a_3080_42308# 4.95e-19
C12146 a_11173_44260# a_11173_43940# 8.81e-19
C12147 a_11341_43940# a_18533_43940# 0.005886f
C12148 a_20365_43914# a_21381_43940# 3.94e-20
C12149 a_n2293_43922# a_4361_42308# 0.035634f
C12150 a_10057_43914# a_10341_42308# 2.07e-20
C12151 a_3065_45002# a_4921_42308# 4.26e-19
C12152 a_3537_45260# a_3905_42558# 1.27e-20
C12153 a_n1059_45260# a_8685_42308# 5.76e-19
C12154 a_5111_44636# a_5267_42460# 0.047489f
C12155 a_n913_45002# a_8325_42308# 0.233489f
C12156 a_n2017_45002# a_8791_42308# 0.004421f
C12157 a_10405_44172# VDD 0.408512f
C12158 a_2711_45572# en_comp 4.72e-20
C12159 a_15599_45572# a_15765_45572# 0.576512f
C12160 a_20974_43370# a_4185_45028# 0.184625f
C12161 a_8685_43396# a_13059_46348# 0.002513f
C12162 a_18599_43230# a_13661_43548# 0.001237f
C12163 a_n2293_42282# a_768_44030# 1.83e-20
C12164 a_9127_43156# a_2107_46812# 6e-20
C12165 a_13635_43156# a_n2293_46634# 1.15e-19
C12166 a_n1761_44111# a_n863_45724# 6.9e-20
C12167 a_n1899_43946# a_n1079_45724# 1.2e-21
C12168 a_n984_44318# a_n2661_45546# 1.23e-21
C12169 a_2455_43940# a_2324_44458# 1.69e-19
C12170 a_9420_43940# a_9290_44172# 0.002091f
C12171 a_16328_43172# a_10227_46804# 1.46e-21
C12172 a_n784_42308# a_n1151_42308# 0.154055f
C12173 a_1576_42282# a_584_46384# 6.73e-21
C12174 a_n3420_37984# C5_P_btm 1.22e-19
C12175 a_n4064_37984# C7_P_btm 4.26e-20
C12176 VDAC_Pi a_n923_35174# 0.001372f
C12177 a_10903_45394# CLK 0.001362f
C12178 a_n901_46420# VDD 0.518805f
C12179 a_19647_42308# CAL_N 0.001755f
C12180 a_n4064_40160# a_n3420_37440# 0.062634f
C12181 a_n4209_39590# a_n4209_37414# 0.031971f
C12182 a_7174_31319# VDAC_N 0.006576f
C12183 a_n4315_30879# a_n4064_37440# 0.035563f
C12184 a_n3565_38502# a_n4064_37984# 0.028083f
C12185 a_n3420_38528# a_n3420_37984# 0.113087f
C12186 a_1343_38525# a_3754_39134# 1.67e-19
C12187 C0_dummy_N_btm C1_N_btm 1.24905f
C12188 C0_dummy_P_btm C2_N_btm 2.79e-20
C12189 C0_P_btm C3_N_btm 3.06e-19
C12190 C1_P_btm C4_N_btm 8.82e-20
C12191 a_3483_46348# a_526_44458# 0.134907f
C12192 a_167_45260# a_1337_46116# 2.67e-20
C12193 a_15227_44166# a_n443_42852# 0.023429f
C12194 a_9569_46155# a_6945_45028# 3.28e-20
C12195 a_15015_46420# a_14840_46494# 0.233657f
C12196 a_14275_46494# a_2324_44458# 5.45e-20
C12197 a_n4318_40392# a_n4064_40160# 0.077948f
C12198 a_14539_43914# a_17124_42282# 3.94e-20
C12199 a_n356_44636# a_15486_42560# 1.56e-19
C12200 a_5891_43370# a_10723_42308# 2.6e-20
C12201 a_n2293_43922# a_6761_42308# 4.97e-20
C12202 a_n2661_42834# a_6123_31319# 3.51e-21
C12203 a_n97_42460# a_4361_42308# 0.15989f
C12204 a_11341_43940# a_17595_43084# 3.11e-20
C12205 a_15493_43940# a_16414_43172# 3.51e-21
C12206 a_3626_43646# a_18783_43370# 6.43e-21
C12207 a_2982_43646# a_19268_43646# 3.9e-21
C12208 a_8685_43396# a_15095_43370# 0.064911f
C12209 a_9145_43396# a_9803_43646# 0.055143f
C12210 a_19478_44306# a_19339_43156# 1.67e-19
C12211 a_15493_43396# a_19164_43230# 8.79e-19
C12212 a_13507_46334# SINGLE_ENDED 0.111959f
C12213 a_21496_47436# START 3e-20
C12214 a_4883_46098# RST_Z 1.25e-19
C12215 a_20556_43646# VDD 0.34939f
C12216 a_18691_45572# a_18911_45144# 0.006432f
C12217 a_18479_45785# a_18494_42460# 3.74e-20
C12218 a_6171_45002# a_9482_43914# 0.016128f
C12219 a_8423_43396# a_n357_42282# 1.68e-19
C12220 a_8317_43396# a_n755_45592# 0.007502f
C12221 a_12089_42308# a_9290_44172# 0.047614f
C12222 a_10991_42826# a_10903_43370# 9.88e-21
C12223 a_18599_43230# a_4185_45028# 1.09e-20
C12224 a_15037_45618# a_13661_43548# 0.001104f
C12225 a_6598_45938# a_6540_46812# 1.76e-21
C12226 a_17478_45572# a_12549_44172# 8.8e-20
C12227 a_2711_45572# a_7411_46660# 5.52e-20
C12228 a_14033_45822# a_13747_46662# 0.021007f
C12229 a_14127_45572# a_n881_46662# 7.26e-20
C12230 a_21188_45572# a_21496_47436# 1.76e-21
C12231 a_21363_45546# a_4883_46098# 2.24e-20
C12232 a_3357_43084# a_17591_47464# 5.7e-19
C12233 a_2437_43646# a_18479_47436# 0.041425f
C12234 a_20885_45572# a_18597_46090# 0.002608f
C12235 a_20447_31679# a_16327_47482# 2.78e-20
C12236 a_3232_43370# a_3160_47472# 2.79e-20
C12237 a_5691_45260# a_n1151_42308# 1.4e-20
C12238 a_3537_45260# a_4791_45118# 0.33264f
C12239 a_n1059_45260# a_12861_44030# 7.52e-20
C12240 a_413_45260# a_6851_47204# 9.63e-20
C12241 a_n2661_45546# a_3503_45724# 0.006856f
C12242 a_380_45546# a_n357_42282# 0.071576f
C12243 a_n452_45724# a_n755_45592# 0.03904f
C12244 a_n1099_45572# a_310_45028# 0.333219f
C12245 a_n863_45724# a_997_45618# 3.46e-19
C12246 a_22223_43396# a_22223_42860# 0.026152f
C12247 a_8037_42858# a_8605_42826# 0.178024f
C12248 a_7871_42858# a_9127_43156# 0.043633f
C12249 a_13887_32519# a_22165_42308# 0.002652f
C12250 a_3080_42308# a_3318_42354# 0.036372f
C12251 a_n97_42460# a_6761_42308# 0.012266f
C12252 a_11341_43940# a_21887_42336# 1.43e-20
C12253 a_7765_42852# a_8387_43230# 4.21e-19
C12254 a_15095_43370# a_15953_42852# 2.26e-19
C12255 a_2982_43646# a_1755_42282# 0.051666f
C12256 a_21188_46660# RST_Z 1.88e-21
C12257 a_765_45546# CLK 0.0309f
C12258 a_20623_46660# SINGLE_ENDED 2.87e-20
C12259 a_n3565_37414# a_n2860_37690# 2.96e-19
C12260 a_n4209_37414# a_n4251_37440# 0.00226f
C12261 a_7754_38470# a_3726_37500# 0.124796f
C12262 a_7754_38636# VDAC_N 9.38e-20
C12263 VDAC_Ni a_6886_37412# 0.178275f
C12264 a_3754_38470# a_5088_37509# 0.632585f
C12265 a_n3420_37440# a_n4064_37440# 8.19012f
C12266 a_6171_42473# VDD 0.184622f
C12267 a_n237_47217# a_584_46384# 0.645142f
C12268 a_n971_45724# a_2553_47502# 0.23907f
C12269 a_327_47204# a_1239_47204# 6.56e-19
C12270 a_n1741_47186# a_3381_47502# 0.011573f
C12271 a_n2109_47186# a_3815_47204# 0.045952f
C12272 a_n785_47204# a_1431_47204# 6.54e-19
C12273 SMPL_ON_P a_n1151_42308# 2.27e-19
C12274 a_n2293_45010# a_n1761_44111# 0.148418f
C12275 a_413_45260# a_3422_30871# 3.37e-19
C12276 a_3357_43084# a_1414_42308# 6.88e-19
C12277 a_2437_43646# a_2479_44172# 0.00389f
C12278 a_n2109_45247# a_n2065_43946# 7.64e-21
C12279 a_n2661_45010# a_n1331_43914# 4.98e-21
C12280 a_13556_45296# a_14581_44484# 2.18e-19
C12281 a_n2293_42834# a_7640_43914# 0.040893f
C12282 a_16680_45572# a_15682_43940# 1.27e-20
C12283 a_9482_43914# a_14673_44172# 0.42967f
C12284 a_n4318_40392# a_n2433_44484# 0.001155f
C12285 a_n2840_44458# a_n2129_44697# 6.34e-19
C12286 a_16922_45042# a_16979_44734# 7.83e-19
C12287 a_17023_45118# a_14539_43914# 7.91e-19
C12288 a_8791_42308# a_526_44458# 1.73e-21
C12289 a_14635_42282# a_n443_42852# 4.48e-20
C12290 a_4190_30871# CAL_P 0.007081f
C12291 a_18341_45572# a_12741_44636# 2.38e-20
C12292 a_19431_45546# a_11415_45002# 0.005163f
C12293 a_1307_43914# a_6755_46942# 0.076439f
C12294 a_18545_45144# a_19321_45002# 8.98e-21
C12295 a_11691_44458# a_n2661_46634# 8.5e-20
C12296 a_21188_45572# a_21363_46634# 9.99e-20
C12297 a_20731_45938# a_20841_46902# 1.09e-20
C12298 a_6171_45002# a_12816_46660# 6.34e-21
C12299 a_5111_44636# a_3090_45724# 0.063636f
C12300 a_11823_42460# a_2324_44458# 0.058835f
C12301 a_14495_45572# a_13759_46122# 2.94e-20
C12302 a_13249_42308# a_13925_46122# 0.001657f
C12303 a_10210_45822# a_10355_46116# 1.86e-19
C12304 a_8162_45546# a_6945_45028# 2.68e-20
C12305 a_8697_45572# a_8199_44636# 4.76e-19
C12306 a_8701_44490# a_n1613_43370# 2.9e-20
C12307 a_18287_44626# a_11453_44696# 0.001467f
C12308 a_5534_30871# a_13070_42354# 0.025818f
C12309 a_3080_42308# C10_N_btm 1.34e-19
C12310 a_12549_44172# a_19594_46812# 7.14e-20
C12311 a_n881_46662# a_n2442_46660# 1.71e-20
C12312 a_n1613_43370# a_n2293_46634# 0.103089f
C12313 a_9313_45822# a_7411_46660# 1.38e-19
C12314 a_6575_47204# a_7927_46660# 1.99e-19
C12315 a_6151_47436# a_10467_46802# 2.6e-19
C12316 a_4915_47217# a_10249_46116# 0.001348f
C12317 a_n1151_42308# a_8035_47026# 6.49e-20
C12318 a_4791_45118# a_6969_46634# 0.001756f
C12319 a_18494_42460# a_14021_43940# 0.026241f
C12320 a_1307_43914# a_1209_43370# 0.001241f
C12321 a_8746_45002# a_10991_42826# 2.47e-21
C12322 a_10193_42453# a_10922_42852# 3.71e-21
C12323 a_17517_44484# a_19006_44850# 0.016181f
C12324 a_17061_44734# a_11967_42832# 2.07e-20
C12325 a_5343_44458# a_9028_43914# 1.94e-20
C12326 a_6171_45002# a_6031_43396# 6.47e-22
C12327 a_3232_43370# a_6293_42852# 0.004069f
C12328 a_5111_44636# a_6547_43396# 0.035842f
C12329 a_3537_45260# a_8791_43396# 0.071369f
C12330 a_n1059_45260# a_9803_43646# 1.87e-20
C12331 a_n913_45002# a_9145_43396# 0.004598f
C12332 a_n2661_44458# a_2804_46116# 4.17e-21
C12333 a_18114_32519# a_4185_45028# 0.080343f
C12334 a_13076_44458# a_11415_45002# 3.9e-21
C12335 a_949_44458# a_472_46348# 7.78e-21
C12336 a_8975_43940# a_12741_44636# 3.01e-19
C12337 a_15682_43940# a_13747_46662# 3.79e-21
C12338 a_20935_43940# a_12549_44172# 0.110704f
C12339 a_n2661_42282# a_n2312_38680# 4.25e-20
C12340 a_17737_43940# a_13661_43548# 0.031811f
C12341 a_15146_44811# a_15227_44166# 1.56e-20
C12342 a_1307_43914# a_8049_45260# 1.63e-19
C12343 a_2437_43646# a_n443_42852# 0.006604f
C12344 a_n913_45002# a_n1099_45572# 2.98e-19
C12345 a_n467_45028# a_n2661_45546# 0.002796f
C12346 a_n2017_45002# a_n357_42282# 0.580077f
C12347 a_n967_45348# a_n2293_45546# 0.119714f
C12348 a_18533_43940# a_16327_47482# 0.001702f
C12349 a_15037_43940# a_10227_46804# 0.002378f
C12350 a_1987_43646# a_584_46384# 2.38e-19
C12351 a_1209_43370# a_n443_46116# 0.061682f
C12352 a_5742_30871# a_7174_31319# 0.34728f
C12353 a_15890_42674# a_4958_30871# 0.017137f
C12354 a_15803_42450# a_17531_42308# 6.07e-21
C12355 a_15959_42545# a_17303_42282# 6.6e-20
C12356 a_n4318_37592# a_n4334_38304# 7.52e-20
C12357 a_5934_30871# a_n4209_39590# 1.08e-21
C12358 a_6123_31319# a_n3565_39590# 5.77e-21
C12359 a_6545_47178# VDD 0.386368f
C12360 a_n1151_42308# a_11387_46482# 0.005536f
C12361 a_4190_30871# CAL_N 0.045535f
C12362 a_n2312_38680# a_n2840_46090# 0.003997f
C12363 a_n2661_46634# a_n1991_46122# 9.31e-19
C12364 a_n2293_46634# a_n2293_46098# 0.062583f
C12365 a_4883_46098# a_18985_46122# 0.027089f
C12366 a_13507_46334# a_19335_46494# 0.004216f
C12367 a_20894_47436# a_20708_46348# 1.02e-19
C12368 a_19386_47436# a_6945_45028# 0.008586f
C12369 a_18780_47178# a_10809_44734# 0.002996f
C12370 a_6151_47436# a_8034_45724# 9.18e-19
C12371 a_11453_44696# a_15682_46116# 1.17e-20
C12372 a_8128_46384# a_8016_46348# 0.09182f
C12373 a_n881_46662# a_8953_45546# 1.01e-19
C12374 a_n2017_45002# a_18707_42852# 0.026353f
C12375 a_11823_42460# a_16522_42674# 1.68e-21
C12376 a_1307_43914# a_3059_42968# 1.72e-19
C12377 a_10807_43548# a_11341_43940# 0.049779f
C12378 a_6453_43914# a_6671_43940# 0.08213f
C12379 a_10193_42453# a_17531_42308# 7.42e-19
C12380 a_9313_44734# a_14579_43548# 0.038528f
C12381 a_17973_43940# a_19478_44306# 0.001007f
C12382 a_18079_43940# a_15493_43396# 1.94e-19
C12383 a_5891_43370# a_10341_43396# 0.087957f
C12384 a_n2840_43914# a_n2840_43370# 0.025171f
C12385 a_18248_44752# a_18429_43548# 5.65e-19
C12386 a_16979_44734# a_15743_43084# 1.34e-20
C12387 a_20980_44850# VDD 0.132317f
C12388 a_11823_42460# a_13527_45546# 0.027805f
C12389 a_2711_45572# a_16855_45546# 2.31e-22
C12390 a_12791_45546# a_13163_45724# 1.53e-19
C12391 a_9049_44484# a_9241_45822# 3.68e-20
C12392 C0_N_btm C10_P_btm 8.52e-19
C12393 C0_dummy_P_btm C8_P_btm 0.234177f
C12394 C0_dummy_N_btm C9_P_btm 4.11e-19
C12395 C5_N_btm EN_VIN_BSTR_N 0.115337f
C12396 C0_P_btm C7_P_btm 0.140846f
C12397 C1_P_btm C6_P_btm 0.127656f
C12398 a_4235_43370# a_3090_45724# 1.99e-22
C12399 a_n310_44484# a_n755_45592# 0.001049f
C12400 a_n2661_43922# a_n2661_45546# 0.028803f
C12401 a_n2293_43922# a_n2810_45572# 2.93e-20
C12402 a_9672_43914# a_8016_46348# 0.074243f
C12403 a_8018_44260# a_5937_45572# 1.38e-20
C12404 a_8333_44056# a_8199_44636# 2.67e-19
C12405 a_n1533_42852# a_n1613_43370# 0.012196f
C12406 a_17595_43084# a_16327_47482# 0.007234f
C12407 a_15279_43071# a_10227_46804# 0.001583f
C12408 a_19987_42826# a_12861_44030# 1.24e-19
C12409 a_19692_46634# VDD 2.53528f
C12410 a_5932_42308# VDAC_N 0.007321f
C12411 a_6123_31319# a_3726_37500# 0.002503f
C12412 a_2698_46116# a_3147_46376# 0.003074f
C12413 a_2521_46116# a_3483_46348# 1.75e-19
C12414 a_167_45260# a_3699_46348# 4.42e-20
C12415 a_17609_46634# a_8049_45260# 1.64e-21
C12416 a_11901_46660# a_12638_46436# 4.56e-19
C12417 a_12469_46902# a_12379_46436# 5.5e-19
C12418 a_11415_45002# a_12594_46348# 1.51e-20
C12419 a_20411_46873# a_20708_46348# 0.081063f
C12420 a_20273_46660# a_19900_46494# 3.92e-19
C12421 a_20107_46660# a_21137_46414# 0.001469f
C12422 a_18285_46348# a_10809_44734# 0.014976f
C12423 a_1823_45246# a_4419_46090# 0.340207f
C12424 a_15493_43940# a_21487_43396# 1.34e-19
C12425 a_4223_44672# a_5932_42308# 1.08e-20
C12426 a_3080_42308# a_6197_43396# 3.94e-21
C12427 a_n1557_42282# a_1512_43396# 1.26e-20
C12428 a_3499_42826# a_2075_43172# 1.63e-19
C12429 a_n97_42460# a_7274_43762# 4.27e-20
C12430 a_11341_43940# a_13467_32519# 0.001199f
C12431 a_n1920_47178# CLK_DATA 3.9e-19
C12432 a_n2109_47186# DATA[0] 0.08202f
C12433 a_3457_43396# VDD 0.004013f
C12434 a_n2661_45010# a_n967_45348# 0.019427f
C12435 a_n2109_45247# a_n2810_45028# 4.84e-19
C12436 a_19963_31679# a_413_45260# 0.0432f
C12437 a_n2472_45002# en_comp 0.117861f
C12438 a_n2017_45002# a_n745_45366# 7.49e-21
C12439 a_n2293_45010# a_n2956_37592# 0.005894f
C12440 a_n1059_45260# a_n913_45002# 1.19505f
C12441 a_10193_42453# a_18184_42460# 0.216199f
C12442 a_16147_45260# a_14537_43396# 5.04e-19
C12443 a_10907_45822# a_n2661_43370# 0.057449f
C12444 a_5907_45546# a_n2661_44458# 6.68e-20
C12445 a_13887_32519# a_4185_45028# 0.044689f
C12446 a_n1917_43396# a_n2293_45546# 9.31e-20
C12447 a_743_42282# a_8016_46348# 1.7e-20
C12448 a_18057_42282# a_13507_46334# 6.56e-20
C12449 a_20692_30879# VDD 0.499615f
C12450 a_3775_45552# a_768_44030# 1.42e-21
C12451 a_2711_45572# a_13661_43548# 0.552383f
C12452 a_6812_45938# a_n881_46662# 1.43e-19
C12453 a_15037_45618# a_14955_47212# 4.91e-20
C12454 a_15599_45572# a_12861_44030# 0.025507f
C12455 a_8049_45260# a_19443_46116# 0.001302f
C12456 a_526_44458# a_n357_42282# 0.220537f
C12457 a_10729_43914# a_5742_30871# 1.45e-20
C12458 a_3422_30871# a_n4064_39616# 0.003743f
C12459 a_21381_43940# a_22400_42852# 1.44e-20
C12460 a_10807_43548# a_10723_42308# 8.52e-19
C12461 a_10341_43396# a_17595_43084# 3.94e-20
C12462 a_10623_46897# CLK 0.016177f
C12463 a_10249_46116# DATA[5] 3.81e-19
C12464 a_6755_46942# DATA[4] 4.06e-21
C12465 a_6969_46634# DATA[3] 6.68e-20
C12466 a_n4064_37984# a_n2860_37984# 0.003765f
C12467 a_19431_45546# a_11967_42832# 1.18e-20
C12468 a_20107_45572# a_17517_44484# 2.01e-21
C12469 a_13159_45002# a_13076_44458# 3.32e-19
C12470 a_9482_43914# a_12607_44458# 0.151452f
C12471 a_13017_45260# a_13720_44458# 2.63e-20
C12472 a_1423_45028# a_4223_44672# 0.013079f
C12473 a_2711_45572# a_19862_44208# 0.002631f
C12474 a_5111_44636# a_n356_44636# 1.45e-19
C12475 a_8515_42308# a_4185_45028# 6.87e-20
C12476 a_14543_43071# a_n443_42852# 6.35e-20
C12477 a_19164_43230# a_n357_42282# 0.011328f
C12478 a_n2472_42282# a_n2956_38680# 2.5e-20
C12479 a_n4318_38216# a_n2956_39304# 0.023331f
C12480 VIN_N VDD 1.46155f
C12481 a_11322_45546# a_11415_45002# 0.527707f
C12482 a_4099_45572# a_3483_46348# 0.15767f
C12483 a_2711_45572# a_4185_45028# 0.102913f
C12484 a_10193_42453# a_12741_44636# 0.078619f
C12485 a_16147_45260# a_3090_45724# 0.076341f
C12486 a_14180_45002# a_n743_46660# 7.43e-22
C12487 a_5093_45028# a_768_44030# 1.51e-19
C12488 a_3357_43084# a_10428_46928# 1.41e-20
C12489 a_413_45260# a_4651_46660# 3.36e-20
C12490 a_17023_45118# a_11453_44696# 1.62e-19
C12491 a_19778_44110# a_4883_46098# 3.83e-22
C12492 a_18494_42460# a_13507_46334# 0.234442f
C12493 a_8701_44490# a_4791_45118# 0.138973f
C12494 a_16547_43609# a_4958_30871# 6.55e-19
C12495 a_16243_43396# a_17303_42282# 2.6e-19
C12496 a_10922_42852# a_n784_42308# 4.32e-21
C12497 a_2905_42968# a_2903_42308# 1.75e-19
C12498 a_4361_42308# a_10533_42308# 0.017218f
C12499 a_16137_43396# a_17531_42308# 0.001298f
C12500 a_10341_43396# a_21887_42336# 2.25e-20
C12501 a_743_42282# a_11633_42558# 0.005183f
C12502 a_1847_42826# a_3823_42558# 1.7e-20
C12503 a_20692_30879# a_22469_39537# 6.23e-20
C12504 a_n2109_47186# a_3524_46660# 6.67e-20
C12505 a_n1741_47186# a_2959_46660# 3.8e-20
C12506 a_n971_45724# a_1799_45572# 2.58e-19
C12507 a_584_46384# a_1123_46634# 0.370049f
C12508 a_n1151_42308# a_n2438_43548# 0.093859f
C12509 a_327_47204# a_491_47026# 0.001941f
C12510 a_3815_47204# a_n1925_46634# 2.59e-20
C12511 a_4791_45118# a_n2293_46634# 0.030843f
C12512 a_n746_45260# a_645_46660# 4.3e-19
C12513 a_n2312_40392# a_n2312_39304# 0.057374f
C12514 a_13487_47204# a_13759_47204# 0.001672f
C12515 a_11459_47204# a_5807_45002# 5.3e-20
C12516 a_5129_47502# a_n2661_46634# 5.07e-21
C12517 a_15811_47375# a_768_44030# 9.22e-21
C12518 a_15673_47210# a_12549_44172# 3.81e-20
C12519 a_15507_47210# a_15928_47570# 0.089677f
C12520 en_comp a_14401_32519# 7.39e-20
C12521 a_n2661_45010# a_n1917_43396# 3.02e-20
C12522 a_5111_44636# a_9165_43940# 1.1e-19
C12523 a_n2017_45002# a_n2433_43396# 0.035979f
C12524 a_8238_44734# a_n2661_43922# 7.85e-20
C12525 a_n2661_43370# a_n2661_42282# 1.08e-20
C12526 a_11823_42460# a_15743_43084# 1.48e-19
C12527 a_1307_43914# a_11173_44260# 1.43e-19
C12528 a_14539_43914# a_17061_44484# 0.003953f
C12529 a_484_44484# a_556_44484# 0.003395f
C12530 a_5891_43370# a_n2293_43922# 1.56e-19
C12531 a_n4318_40392# a_n2840_43914# 4.88e-19
C12532 a_18374_44850# a_17517_44484# 0.019155f
C12533 a_8696_44636# a_8685_43396# 2.24e-19
C12534 a_n3420_39616# a_n2810_45572# 1.68e-19
C12535 a_3357_43084# VDD 1.66202f
C12536 a_2809_45028# a_1823_45246# 0.076288f
C12537 a_117_45144# a_167_45260# 0.003885f
C12538 a_15060_45348# a_11415_45002# 0.001314f
C12539 a_20512_43084# a_13747_46662# 5.53e-21
C12540 a_18341_45572# a_16375_45002# 9.37e-19
C12541 a_n913_45002# a_n1925_42282# 0.017956f
C12542 a_20885_45572# a_8049_45260# 3.49e-19
C12543 a_9482_43914# a_10903_43370# 1.20611f
C12544 a_13017_45260# a_13351_46090# 1.33e-20
C12545 a_1423_45028# a_6419_46155# 3.69e-22
C12546 a_13159_45002# a_12594_46348# 2.01e-20
C12547 a_1307_43914# a_8953_45546# 0.022061f
C12548 a_14537_43396# a_9290_44172# 3.99e-19
C12549 a_7705_45326# a_2324_44458# 0.029419f
C12550 a_3537_45260# a_6945_45028# 9.87e-21
C12551 a_1241_43940# a_584_46384# 0.007526f
C12552 a_5934_30871# a_9293_42558# 0.001273f
C12553 a_8337_42558# a_8685_42308# 4.27e-19
C12554 a_5932_42308# a_5742_30871# 1.14154f
C12555 EN_VIN_BSTR_P C2_P_btm 0.118072f
C12556 a_n923_35174# RST_Z 0.001488f
C12557 a_22469_39537# VIN_N 2.79e-20
C12558 a_n743_46660# a_15009_46634# 1.24e-21
C12559 a_12549_44172# a_16388_46812# 0.03419f
C12560 a_6540_46812# a_7411_46660# 5.06e-21
C12561 a_5732_46660# a_7715_46873# 1.03e-20
C12562 a_768_44030# a_13059_46348# 0.062321f
C12563 a_5907_46634# a_7577_46660# 5.36e-20
C12564 a_5072_46660# a_5257_43370# 1.51e-20
C12565 a_5807_45002# a_12925_46660# 9.54e-20
C12566 a_4842_47243# a_765_45546# 4.26e-19
C12567 a_22223_47212# a_20202_43084# 1.25e-19
C12568 a_12465_44636# a_11415_45002# 0.375509f
C12569 a_21496_47436# a_12741_44636# 4.23e-20
C12570 a_4883_46098# a_20820_30879# 1.84e-19
C12571 a_n1435_47204# a_3147_46376# 6.37e-21
C12572 a_4915_47217# a_5937_45572# 2.78e-20
C12573 a_6151_47436# a_8016_46348# 1.03e-19
C12574 a_n1151_42308# a_11133_46155# 0.162011f
C12575 a_17613_45144# a_17499_43370# 5.51e-21
C12576 a_8701_44490# a_8791_43396# 1.69e-20
C12577 a_20640_44752# a_14021_43940# 8.61e-21
C12578 a_3422_30871# a_22223_43948# 0.011616f
C12579 a_n356_44636# a_4235_43370# 5.73e-21
C12580 a_5883_43914# a_8147_43396# 3.36e-20
C12581 a_5891_43370# a_n97_42460# 0.957548f
C12582 a_20512_43084# a_20269_44172# 2.47e-20
C12583 a_11823_42460# a_1606_42308# 4.73e-20
C12584 a_18184_42460# a_16137_43396# 0.029846f
C12585 a_n2661_44458# a_9145_43396# 2.4e-20
C12586 a_n913_45002# a_19987_42826# 4.56e-20
C12587 en_comp a_18817_42826# 4.89e-21
C12588 a_n2017_45002# a_21356_42826# 1.31e-20
C12589 a_5826_44734# VDD 0.007376f
C12590 a_n4064_39616# VREF_GND 0.241027f
C12591 a_5263_45724# a_6194_45824# 1.4e-19
C12592 a_2711_45572# a_6667_45809# 0.010894f
C12593 a_22485_44484# a_4185_45028# 0.080982f
C12594 a_13483_43940# a_13059_46348# 0.124566f
C12595 a_8791_43396# a_n2293_46634# 0.010288f
C12596 a_14955_43396# a_12549_44172# 4.21e-19
C12597 a_22959_43948# a_19692_46634# 8.6e-20
C12598 a_13076_44458# a_13259_45724# 0.188498f
C12599 a_n2661_44458# a_n1099_45572# 9.19e-21
C12600 a_3363_44484# a_526_44458# 0.119556f
C12601 a_n1917_44484# a_n2293_45546# 6.29e-19
C12602 a_17517_44484# a_17715_44484# 0.163303f
C12603 a_15367_44484# a_2324_44458# 3.72e-19
C12604 a_13467_32519# a_16327_47482# 0.004353f
C12605 a_n2302_39072# a_n2302_38778# 0.050477f
C12606 a_n4209_39304# a_n4209_38216# 0.029694f
C12607 a_3877_44458# VDD 0.786903f
C12608 a_21188_46660# a_20820_30879# 3.56e-19
C12609 a_21363_46634# a_12741_44636# 0.053741f
C12610 a_20273_46660# a_21297_46660# 2.36e-20
C12611 a_768_44030# a_3218_45724# 3.61e-19
C12612 a_5167_46660# a_5066_45546# 1.61e-20
C12613 a_22612_30879# a_20692_30879# 0.07827f
C12614 a_n1613_43370# a_2277_45546# 3.18e-21
C12615 a_10249_46116# a_10809_44734# 4.78e-19
C12616 a_3090_45724# a_9290_44172# 0.196232f
C12617 a_6969_46634# a_6945_45028# 0.017662f
C12618 a_12251_46660# a_12594_46348# 0.011817f
C12619 a_12816_46660# a_10903_43370# 3.28e-19
C12620 a_10057_43914# a_10752_42852# 1.23e-20
C12621 a_19237_31679# a_17364_32525# 0.054573f
C12622 a_n2293_42834# a_5932_42308# 2.23e-19
C12623 a_9313_44734# a_21671_42860# 0.012466f
C12624 a_14955_43940# a_14205_43396# 4.77e-19
C12625 a_1414_42308# a_743_42282# 0.004767f
C12626 a_n2840_43370# a_n4318_39304# 0.158695f
C12627 a_14537_43396# a_15051_42282# 7.92e-20
C12628 a_10807_43548# a_10341_43396# 0.042318f
C12629 a_11962_45724# a_11787_45002# 4.92e-19
C12630 a_19256_45572# a_20107_45572# 4.08e-19
C12631 a_8746_45002# a_9482_43914# 0.002141f
C12632 a_11322_45546# a_13159_45002# 4.52e-20
C12633 a_11652_45724# a_11963_45334# 8.93e-19
C12634 a_11823_42460# a_10775_45002# 2.94e-20
C12635 a_18175_45572# a_20528_45572# 2.64e-21
C12636 a_6469_45572# a_6171_45002# 4.62e-19
C12637 a_16137_43396# a_12741_44636# 3.03e-20
C12638 a_8952_43230# a_8270_45546# 1.53e-20
C12639 a_18079_43940# a_n357_42282# 1.54e-20
C12640 a_9396_43370# a_8953_45546# 0.007396f
C12641 a_n1736_42282# a_n1613_43370# 1.08e-20
C12642 VDAC_N VREF 0.008793f
C12643 VDAC_P VIN_P 0.255243f
C12644 a_n1736_46482# VDD 0.083417f
C12645 a_2711_45572# a_14955_47212# 1.19e-21
C12646 a_7230_45938# a_4791_45118# 0.010716f
C12647 a_11525_45546# a_2063_45854# 0.001514f
C12648 a_10180_45724# a_n1151_42308# 6.68e-20
C12649 a_4808_45572# a_6151_47436# 2.53e-20
C12650 a_n2293_46098# a_2277_45546# 0.005746f
C12651 a_n1853_46287# a_n443_42852# 0.003661f
C12652 a_167_45260# a_n755_45592# 1.02724f
C12653 a_1823_45246# a_1848_45724# 0.028459f
C12654 a_1431_46436# a_1337_46116# 1.26e-19
C12655 a_12594_46348# a_13259_45724# 0.012487f
C12656 a_22223_46124# a_8049_45260# 0.007569f
C12657 a_14493_46090# a_14537_46482# 3.69e-19
C12658 a_13925_46122# a_14949_46494# 2.36e-20
C12659 a_5164_46348# a_n2661_45546# 8.06e-20
C12660 a_18525_43370# a_18783_43370# 0.22264f
C12661 a_16977_43638# a_16867_43762# 0.097745f
C12662 a_14205_43396# a_5649_42852# 4.06e-21
C12663 a_18429_43548# a_15743_43084# 0.053516f
C12664 a_10341_43396# a_13467_32519# 0.007243f
C12665 a_n97_42460# a_17595_43084# 0.0027f
C12666 a_20974_43370# a_21671_42860# 8.3e-20
C12667 a_3626_43646# a_8037_42858# 5.94e-20
C12668 a_2982_43646# a_8387_43230# 3.53e-20
C12669 a_n2661_42282# COMP_P 0.02767f
C12670 a_3905_42865# a_5267_42460# 9.02e-20
C12671 a_12281_43396# a_743_42282# 0.036414f
C12672 a_16759_43396# a_16664_43396# 0.049827f
C12673 a_16137_43396# a_15868_43402# 5.04e-20
C12674 a_21588_30879# VREF 0.860047f
C12675 a_22612_30879# VIN_N 0.19035f
C12676 a_n1925_46634# DATA[0] 2.87e-19
C12677 a_5342_30871# VDD 0.496295f
C12678 a_n2810_45028# a_n3565_37414# 0.135518f
C12679 a_3357_43084# a_n699_43396# 0.004379f
C12680 a_n2661_45010# a_n1917_44484# 0.015623f
C12681 a_n1059_45260# a_n2661_44458# 0.028647f
C12682 a_n2017_45002# a_n2433_44484# 0.039498f
C12683 a_n2109_45247# a_n2129_44697# 0.003166f
C12684 a_n2293_45010# a_n2267_44484# 0.0118f
C12685 a_8696_44636# a_8783_44734# 7.48e-19
C12686 a_1423_45028# a_n2293_42834# 0.033636f
C12687 a_18596_45572# a_18443_44721# 1.58e-20
C12688 a_18799_45938# a_18287_44626# 2.22e-20
C12689 a_15051_42282# a_3090_45724# 1.14e-20
C12690 a_12991_43230# a_9290_44172# 1.31e-20
C12691 a_11962_45724# a_11813_46116# 1.15e-19
C12692 a_2437_43646# a_n2661_46634# 0.02989f
C12693 a_3065_45002# a_n881_46662# 1.23e-20
C12694 a_3429_45260# a_n1613_43370# 2.46e-21
C12695 a_13159_45002# a_12465_44636# 6.58e-20
C12696 a_10951_45334# a_11453_44696# 5.15e-19
C12697 a_9482_43914# a_4883_46098# 0.025151f
C12698 a_3626_43646# a_13921_42308# 5.3e-19
C12699 a_5649_42852# a_22400_42852# 6.16e-20
C12700 a_19987_42826# a_20922_43172# 0.001853f
C12701 a_13678_32519# a_14097_32519# 0.04945f
C12702 a_13467_32519# a_20356_42852# 1.53e-20
C12703 a_8953_45546# DATA[4] 7.93e-19
C12704 a_20107_42308# VDD 0.284252f
C12705 a_n971_45724# a_2747_46873# 0.047519f
C12706 a_n452_47436# a_n310_47243# 0.005572f
C12707 a_n1435_47204# a_12861_44030# 0.036547f
C12708 a_13381_47204# a_13487_47204# 0.152045f
C12709 a_2905_45572# a_4883_46098# 3.03e-20
C12710 a_n1151_42308# a_13507_46334# 0.001912f
C12711 a_17719_45144# a_17517_44484# 1.47e-19
C12712 a_11691_44458# a_15433_44458# 0.110923f
C12713 a_16979_44734# a_17970_44736# 5.21e-19
C12714 a_1307_43914# a_895_43940# 0.754684f
C12715 a_4223_44672# a_6109_44484# 0.003455f
C12716 a_7499_43078# a_7287_43370# 0.057949f
C12717 a_n2129_44697# a_n310_44484# 2.88e-19
C12718 a_11827_44484# a_11541_44484# 0.0442f
C12719 a_14539_43914# a_18248_44752# 5.77e-20
C12720 a_626_44172# a_1414_42308# 0.002821f
C12721 a_1423_45028# a_1115_44172# 3.06e-20
C12722 a_n1059_45260# a_18451_43940# 2.97e-21
C12723 a_5147_45002# a_5841_44260# 1.74e-19
C12724 a_4921_42308# a_n443_42852# 4.12e-19
C12725 a_3905_42308# a_n755_45592# 6.37e-19
C12726 a_9159_45572# VDD 0.004886f
C12727 a_3429_45260# a_n2293_46098# 2.13e-20
C12728 a_n699_43396# a_3877_44458# 0.061672f
C12729 a_9313_44734# a_5807_45002# 7.63e-20
C12730 a_4223_44672# a_4646_46812# 0.018453f
C12731 a_n2661_43922# a_12891_46348# 1.94e-19
C12732 a_n2661_42834# a_12549_44172# 0.04571f
C12733 a_3175_45822# a_n755_45592# 0.046968f
C12734 a_10193_42453# a_16375_45002# 0.125364f
C12735 a_11682_45822# a_8049_45260# 0.011453f
C12736 a_11322_45546# a_13259_45724# 5.48e-21
C12737 a_11823_42460# a_12839_46116# 2.9e-19
C12738 a_3638_45822# a_n2661_45546# 2.27e-21
C12739 a_18341_45572# a_18985_46122# 7.1e-19
C12740 a_18909_45814# a_18819_46122# 0.003441f
C12741 a_18175_45572# a_19335_46494# 1.2e-19
C12742 a_2437_43646# a_8199_44636# 3.38e-20
C12743 a_11967_42832# a_12465_44636# 1.63e-20
C12744 a_17061_44484# a_11453_44696# 3.88e-19
C12745 a_20159_44458# a_4883_46098# 4.39e-22
C12746 a_20640_44752# a_13507_46334# 8.68e-20
C12747 a_n822_43940# a_n971_45724# 1.37e-19
C12748 a_n2661_42282# a_n2497_47436# 4.56e-21
C12749 a_261_44278# a_n746_45260# 5.72e-19
C12750 a_895_43940# a_n443_46116# 0.163929f
C12751 a_1576_42282# a_2123_42473# 4.32e-19
C12752 a_1184_42692# a_1755_42282# 0.016329f
C12753 a_n784_42308# a_2903_42308# 3.86e-20
C12754 a_13291_42460# a_13575_42558# 0.074792f
C12755 a_14635_42282# a_13070_42354# 2.81e-20
C12756 a_14097_32519# a_6123_31319# 0.003315f
C12757 a_3080_42308# VDAC_Pi 3.65e-19
C12758 a_n1925_46634# a_3524_46660# 0.008296f
C12759 a_n743_46660# a_2959_46660# 1.5e-20
C12760 a_601_46902# a_1799_45572# 1.3e-20
C12761 a_n133_46660# a_2609_46660# 1.38e-21
C12762 a_33_46660# a_n2661_46098# 0.007289f
C12763 a_948_46660# a_1110_47026# 0.006453f
C12764 a_383_46660# a_645_46660# 0.001705f
C12765 a_n2438_43548# a_3177_46902# 2.59e-20
C12766 a_n2661_46634# a_3686_47026# 1.44e-19
C12767 a_5807_45002# a_5072_46660# 7.94e-20
C12768 a_9804_47204# a_10150_46912# 3.14e-19
C12769 a_13717_47436# a_14035_46660# 2.07e-20
C12770 a_5129_47502# a_765_45546# 0.004549f
C12771 a_12861_44030# a_13885_46660# 0.042236f
C12772 a_18143_47464# a_15227_44166# 1.06e-19
C12773 a_10227_46804# a_19333_46634# 8.89e-20
C12774 a_4883_46098# a_12816_46660# 3.12e-20
C12775 a_13507_46334# a_14084_46812# 4.22e-20
C12776 a_11453_44696# a_11735_46660# 5.11e-21
C12777 a_n1613_43370# a_6755_46942# 0.006199f
C12778 a_n881_46662# a_10249_46116# 3.58e-19
C12779 a_n2661_45010# a_n1853_43023# 1.08e-20
C12780 a_n2293_43922# a_10807_43548# 1.85e-21
C12781 a_n4318_40392# a_n4318_39304# 0.024428f
C12782 a_16922_45042# a_2982_43646# 0.010868f
C12783 a_9313_44734# a_19478_44306# 5.64e-21
C12784 a_n2661_42834# a_12429_44172# 0.002835f
C12785 a_n2661_43922# a_11750_44172# 3.46e-20
C12786 a_9838_44484# a_9801_43940# 2.53e-21
C12787 a_16237_45028# VDD 0.248452f
C12788 a_4958_30871# EN_VIN_BSTR_P 0.021638f
C12789 a_15803_42450# RST_Z 1.82e-19
C12790 a_3905_42865# a_3090_45724# 0.025179f
C12791 a_21381_43940# a_13747_46662# 0.030122f
C12792 a_10651_43940# a_n2293_46634# 6.07e-19
C12793 a_117_45144# a_n863_45724# 2.14e-19
C12794 a_2809_45028# a_n2293_45546# 5.9e-20
C12795 a_n2661_44458# a_n1925_42282# 0.029506f
C12796 a_15060_45348# a_13259_45724# 4.35e-19
C12797 a_16112_44458# a_15682_46116# 2.03e-21
C12798 a_14539_43914# a_2324_44458# 0.028976f
C12799 a_n356_44636# a_9290_44172# 8.05e-19
C12800 a_6109_44484# a_6419_46155# 1.19e-21
C12801 a_10193_42453# RST_Z 4.5e-19
C12802 a_8128_46384# VDD 0.403575f
C12803 a_n4315_30879# a_n4334_40480# 0.253307f
C12804 a_n784_42308# C9_N_btm 9.31e-20
C12805 a_1606_42308# C0_dummy_P_btm 0.007541f
C12806 a_5534_30871# a_11206_38545# 2.6e-20
C12807 a_13885_46660# a_14180_46812# 0.150851f
C12808 a_17609_46634# a_18285_46348# 0.115413f
C12809 a_15227_44166# a_765_45546# 3.46e-20
C12810 a_n2956_39768# a_n2956_39304# 0.098523f
C12811 a_8128_46384# a_8283_46482# 0.007532f
C12812 a_4646_46812# a_6419_46155# 6.54e-20
C12813 a_5385_46902# a_5164_46348# 0.001231f
C12814 a_4817_46660# a_5204_45822# 0.001084f
C12815 a_2107_46812# a_2324_44458# 0.051531f
C12816 a_n1613_43370# a_8049_45260# 2.61e-20
C12817 a_12465_44636# a_13259_45724# 0.096616f
C12818 a_13507_46334# a_19240_46482# 0.002125f
C12819 a_4883_46098# a_18243_46436# 1.03e-19
C12820 a_18597_46090# a_20254_46482# 0.002021f
C12821 a_18479_47436# a_20850_46482# 7.88e-19
C12822 a_4915_47217# a_n443_42852# 1.15e-20
C12823 a_n443_46116# a_1609_45822# 0.096281f
C12824 a_22315_44484# a_10341_43396# 7.96e-19
C12825 a_1414_42308# a_2813_43396# 0.00815f
C12826 a_5663_43940# a_6031_43396# 1.67e-19
C12827 a_20365_43914# a_19741_43940# 8.59e-20
C12828 a_3499_42826# a_4699_43561# 4.46e-21
C12829 a_n2661_42282# a_1568_43370# 1.94e-21
C12830 a_11967_42832# a_16409_43396# 0.004815f
C12831 a_11341_43940# a_19319_43548# 0.042701f
C12832 a_n356_44636# a_791_42968# 0.003419f
C12833 a_20269_44172# a_21381_43940# 1.62e-20
C12834 a_10807_43548# a_n97_42460# 5.41e-19
C12835 a_19862_44208# a_14401_32519# 2.61e-20
C12836 a_n1059_45260# a_8325_42308# 6.3e-20
C12837 a_n2017_45002# a_8685_42308# 0.016058f
C12838 en_comp a_5934_30871# 0.028694f
C12839 a_n913_45002# a_8337_42558# 5.84e-19
C12840 a_9672_43914# VDD 0.150499f
C12841 a_15297_45822# a_15765_45572# 3.14e-20
C12842 a_15599_45572# a_15903_45785# 0.161702f
C12843 a_n3420_37984# C6_P_btm 1.22e-19
C12844 a_7754_39964# a_n923_35174# 3.06e-20
C12845 a_14401_32519# a_4185_45028# 0.040395f
C12846 a_n809_44244# a_n2661_45546# 2.15e-20
C12847 a_n2065_43946# a_n863_45724# 4.6e-21
C12848 a_n1899_43946# a_n2293_45546# 2.4e-20
C12849 a_2253_43940# a_2324_44458# 2.21e-19
C12850 a_9165_43940# a_9290_44172# 0.01396f
C12851 a_10555_44260# a_10809_44734# 6.94e-19
C12852 a_18695_43230# a_16327_47482# 0.003378f
C12853 a_15785_43172# a_10227_46804# 4.06e-19
C12854 a_1067_42314# a_584_46384# 4.65e-21
C12855 a_196_42282# a_n1151_42308# 1.47e-19
C12856 a_n327_42308# a_n971_45724# 0.001391f
C12857 a_n1641_46494# VDD 0.226065f
C12858 C0_dummy_N_btm C0_N_btm 7.97415f
C12859 C0_dummy_P_btm C1_N_btm 1.59e-19
C12860 C1_P_btm C3_N_btm 5.17e-19
C12861 C0_P_btm C2_N_btm 2.79e-20
C12862 a_19511_42282# CAL_N 0.001217f
C12863 a_n4064_40160# a_n3690_37440# 2.54e-19
C12864 a_7174_31319# a_6886_37412# 4.9e-19
C12865 a_n4315_30879# a_n2946_37690# 1.33e-19
C12866 a_n3565_38502# a_n2946_37984# 0.001251f
C12867 a_n3420_38528# a_n3690_38304# 0.018295f
C12868 a_n4209_38502# a_n2302_37984# 0.001417f
C12869 a_n3690_38528# a_n3420_37984# 8.87e-19
C12870 a_n4334_38528# a_n4064_37984# 7.91e-19
C12871 a_3147_46376# a_526_44458# 0.352f
C12872 a_3483_46348# a_2981_46116# 2.44e-19
C12873 a_5937_45572# a_10809_44734# 0.001476f
C12874 a_14275_46494# a_14840_46494# 7.99e-20
C12875 a_9625_46129# a_6945_45028# 1.2e-19
C12876 a_14493_46090# a_2324_44458# 6.29e-20
C12877 a_20512_43084# a_20836_43172# 8.79e-20
C12878 a_3422_30871# a_20753_42852# 0.048434f
C12879 a_n4318_40392# a_n4334_40480# 0.089305f
C12880 a_n356_44636# a_15051_42282# 8.17e-19
C12881 a_19328_44172# a_19164_43230# 2.78e-20
C12882 a_15493_43940# a_15567_42826# 6.99e-20
C12883 a_2982_43646# a_15743_43084# 0.023587f
C12884 a_8685_43396# a_14205_43396# 0.011249f
C12885 a_15493_43396# a_19339_43156# 3.83e-19
C12886 a_5891_43370# a_10533_42308# 5.45e-19
C12887 a_21177_47436# SINGLE_ENDED 0.057266f
C12888 a_13507_46334# START 4.08e-19
C12889 a_10227_46804# CLK 0.207445f
C12890 a_21496_47436# RST_Z 5.48e-20
C12891 a_743_42282# VDD 0.597869f
C12892 a_18909_45814# a_18911_45144# 0.0027f
C12893 a_18479_45785# a_18184_42460# 3.17e-20
C12894 a_1667_45002# a_626_44172# 1.79e-19
C12895 a_3065_45002# a_1307_43914# 0.033168f
C12896 a_6171_45002# a_13348_45260# 0.009869f
C12897 a_413_45260# a_1423_45028# 0.194002f
C12898 a_3232_43370# a_9482_43914# 0.129525f
C12899 a_n2293_45010# a_117_45144# 2.83e-21
C12900 a_8191_45002# a_8953_45002# 1.72e-19
C12901 a_18817_42826# a_4185_45028# 1.72e-20
C12902 a_8229_43396# a_n755_45592# 0.002439f
C12903 a_16409_43396# a_13259_45724# 7.07e-20
C12904 a_6452_43396# a_n443_42852# 0.001812f
C12905 a_10796_42968# a_10903_43370# 0.001425f
C12906 a_12379_42858# a_9290_44172# 0.001587f
C12907 a_15037_45618# a_5807_45002# 4.32e-21
C12908 a_6667_45809# a_6540_46812# 2.06e-20
C12909 a_2711_45572# a_5257_43370# 0.082068f
C12910 a_15861_45028# a_12549_44172# 7.24e-20
C12911 a_8696_44636# a_768_44030# 0.031444f
C12912 a_14033_45572# a_n881_46662# 5.52e-20
C12913 a_21363_45546# a_21496_47436# 4.09e-21
C12914 a_20623_45572# a_4883_46098# 2.03e-20
C12915 a_21188_45572# a_13507_46334# 8.13e-19
C12916 a_3429_45260# a_4791_45118# 6.17e-21
C12917 a_5205_44484# a_2063_45854# 1.89e-20
C12918 a_3065_45002# a_n443_46116# 1.4e-20
C12919 a_4927_45028# a_n1151_42308# 9.34e-21
C12920 a_n2017_45002# a_12861_44030# 6.5e-19
C12921 a_413_45260# a_6491_46660# 3.19e-19
C12922 a_21513_45002# a_18479_47436# 4.09e-20
C12923 a_22959_45572# a_16327_47482# 5.96e-20
C12924 a_20719_45572# a_18597_46090# 0.005294f
C12925 a_2437_43646# a_18143_47464# 0.013364f
C12926 a_3357_43084# a_16588_47582# 1.09e-19
C12927 a_n2661_45546# a_3316_45546# 0.027868f
C12928 a_380_45546# a_310_45028# 0.057269f
C12929 a_n863_45724# a_n755_45592# 1.76733f
C12930 a_21363_46634# RST_Z 2.85e-20
C12931 a_2982_43646# a_1606_42308# 0.021878f
C12932 a_13887_32519# a_21671_42860# 5.19e-19
C12933 a_4235_43370# a_3823_42558# 3.1e-19
C12934 a_5649_42852# a_22223_42860# 5.33e-19
C12935 a_7871_42858# a_8387_43230# 0.106107f
C12936 a_22223_43396# a_22165_42308# 0.00197f
C12937 a_13678_32519# a_22959_42860# 4.44e-20
C12938 a_648_43396# a_564_42282# 1.99e-20
C12939 a_3080_42308# a_2903_42308# 0.154008f
C12940 a_14021_43940# a_17531_42308# 1.76e-21
C12941 a_15095_43370# a_15597_42852# 0.071983f
C12942 a_7765_42852# a_8605_42826# 6.55e-19
C12943 a_14579_43548# a_16877_42852# 2.78e-22
C12944 a_n97_42460# a_6773_42558# 6.7e-19
C12945 a_20841_46902# SINGLE_ENDED 3.74e-21
C12946 a_n4209_37414# a_n2216_37690# 0.001361f
C12947 VDAC_Ni a_5700_37509# 0.079762f
C12948 a_3754_38470# a_4338_37500# 0.473597f
C12949 a_n3565_37414# a_n2302_37690# 0.046906f
C12950 a_n3690_37440# a_n4064_37440# 0.085414f
C12951 a_n3420_37440# a_n2946_37690# 0.236674f
C12952 a_5755_42308# VDD 0.229304f
C12953 a_n1741_47186# a_n1151_42308# 2.98024f
C12954 a_n237_47217# a_2124_47436# 0.001177f
C12955 a_n971_45724# a_2063_45854# 0.164981f
C12956 a_n2109_47186# a_3785_47178# 0.190973f
C12957 a_n746_45260# a_584_46384# 0.491308f
C12958 a_n785_47204# a_1239_47204# 4.16e-19
C12959 en_comp a_20512_43084# 4.89e-21
C12960 a_n2661_45010# a_n1899_43946# 2.77e-19
C12961 a_n2293_45010# a_n2065_43946# 0.023134f
C12962 a_2437_43646# a_2127_44172# 0.017247f
C12963 a_n2661_43370# a_n310_44811# 3.23e-19
C12964 a_7639_45394# a_7640_43914# 2.67e-20
C12965 a_13556_45296# a_13940_44484# 8.88e-19
C12966 a_8696_44636# a_13483_43940# 9.44e-22
C12967 a_16855_45546# a_15682_43940# 4.92e-20
C12968 a_n2840_44458# a_n2433_44484# 0.039807f
C12969 a_n4318_40392# a_n2661_44458# 0.026979f
C12970 a_16922_45042# a_14539_43914# 0.001347f
C12971 a_8685_42308# a_526_44458# 6.82e-21
C12972 a_13291_42460# a_n443_42852# 1.19e-21
C12973 a_17749_42852# a_n357_42282# 0.001128f
C12974 a_16137_43396# RST_Z 1.66e-20
C12975 a_20273_45572# a_20528_46660# 9.08e-22
C12976 a_18479_45785# a_12741_44636# 0.035678f
C12977 a_18691_45572# a_11415_45002# 0.002376f
C12978 a_16019_45002# a_6755_46942# 0.005906f
C12979 a_n2293_42834# a_4646_46812# 0.152973f
C12980 a_11827_44484# a_n2293_46634# 0.002225f
C12981 a_6194_45824# a_526_44458# 7.16e-21
C12982 a_2437_43646# a_765_45546# 0.030322f
C12983 a_21363_45546# a_21363_46634# 0.001846f
C12984 a_5147_45002# a_3090_45724# 0.023629f
C12985 a_6298_44484# a_n881_46662# 0.002351f
C12986 a_12427_45724# a_2324_44458# 0.001185f
C12987 a_8192_45572# a_8199_44636# 0.04905f
C12988 a_11823_42460# a_14840_46494# 0.004799f
C12989 a_13249_42308# a_13759_46122# 0.001706f
C12990 a_13904_45546# a_13925_46122# 5.43e-19
C12991 a_10210_45822# a_9823_46155# 0.001193f
C12992 a_7230_45938# a_6945_45028# 5.3e-19
C12993 a_18248_44752# a_11453_44696# 0.004115f
C12994 a_5534_30871# a_12563_42308# 0.179331f
C12995 a_13460_43230# a_13575_42558# 1.38e-19
C12996 a_3080_42308# C9_N_btm 9.33e-20
C12997 a_12549_44172# a_19321_45002# 0.238866f
C12998 a_n1613_43370# a_n2442_46660# 4.46e-21
C12999 a_6151_47436# a_10428_46928# 0.001405f
C13000 a_6575_47204# a_8145_46902# 0.001541f
C13001 a_7903_47542# a_7927_46660# 1.47e-20
C13002 a_n2109_47186# a_3090_45724# 2.79e-20
C13003 a_4791_45118# a_6755_46942# 2.99e-19
C13004 a_18184_42460# a_14021_43940# 0.029776f
C13005 a_5343_44458# a_8333_44056# 0.092296f
C13006 a_1307_43914# a_458_43396# 3.65e-20
C13007 a_n356_44636# a_3905_42865# 3.95e-20
C13008 a_10193_42453# a_10991_42826# 5.97e-20
C13009 a_17517_44484# a_18588_44850# 0.026595f
C13010 a_5883_43914# a_n2661_42282# 0.107496f
C13011 a_7499_43078# a_12089_42308# 9.57e-21
C13012 a_3232_43370# a_6031_43396# 4.81e-20
C13013 a_3537_45260# a_8147_43396# 0.088185f
C13014 a_5111_44636# a_6765_43638# 0.022146f
C13015 a_n1059_45260# a_9145_43396# 0.016142f
C13016 a_5147_45002# a_6547_43396# 2e-19
C13017 a_n913_45002# a_8423_43396# 7.65e-20
C13018 a_626_44172# VDD 0.621601f
C13019 a_n784_42308# RST_Z 0.033698f
C13020 a_n2661_44458# a_2698_46116# 1.03e-21
C13021 a_15433_44458# a_15227_44166# 0.026124f
C13022 a_15682_43940# a_13661_43548# 0.055235f
C13023 a_20623_43914# a_12549_44172# 0.033887f
C13024 a_16019_45002# a_8049_45260# 2.24e-21
C13025 a_n745_45366# a_n452_45724# 0.00143f
C13026 a_n1059_45260# a_n1099_45572# 2.72e-19
C13027 a_n2293_45010# a_n755_45592# 0.159033f
C13028 en_comp a_n2293_45546# 2.1e-19
C13029 a_458_43396# a_n443_46116# 1.87e-21
C13030 a_1891_43646# a_584_46384# 4.57e-19
C13031 a_13565_43940# a_10227_46804# 5.26e-19
C13032 a_19319_43548# a_16327_47482# 0.021453f
C13033 a_15959_42545# a_4958_30871# 0.043235f
C13034 a_15803_42450# a_17303_42282# 0.00508f
C13035 a_11323_42473# a_7174_31319# 4.88e-21
C13036 a_n3674_38216# a_n3565_38216# 0.128699f
C13037 a_n4318_37592# a_n4209_38216# 1.11e-19
C13038 a_15890_42674# a_16269_42308# 3.16e-19
C13039 a_n3674_37592# a_n4064_38528# 0.019942f
C13040 a_6151_47436# VDD 4.39915f
C13041 a_4190_30871# a_11206_38545# 1.56e-20
C13042 a_n1151_42308# a_10586_45546# 0.02493f
C13043 a_4791_45118# a_8049_45260# 3.69e-19
C13044 a_n2661_46634# a_n1853_46287# 2.3e-19
C13045 a_n2293_46634# a_n2472_46090# 3.35e-19
C13046 a_9863_46634# a_10185_46660# 0.007399f
C13047 a_3686_47026# a_765_45546# 1.39e-19
C13048 a_11453_44696# a_2324_44458# 0.023884f
C13049 a_12465_44636# a_18189_46348# 1.08e-20
C13050 a_6575_47204# a_5066_45546# 2.37e-20
C13051 a_4883_46098# a_18819_46122# 0.054304f
C13052 a_13507_46334# a_19553_46090# 0.002559f
C13053 a_18597_46090# a_6945_45028# 0.049383f
C13054 a_18479_47436# a_10809_44734# 0.04504f
C13055 a_n1613_43370# a_8953_45546# 0.024821f
C13056 a_n881_46662# a_5937_45572# 0.195456f
C13057 a_8128_46384# a_7920_46348# 0.197919f
C13058 a_1307_43914# a_2987_42968# 3.55e-20
C13059 a_5891_43370# a_9885_43646# 0.004104f
C13060 a_10949_43914# a_11341_43940# 0.0383f
C13061 a_9028_43914# a_9248_44260# 0.009965f
C13062 a_n699_43396# a_743_42282# 3.69e-20
C13063 a_10193_42453# a_17303_42282# 0.028322f
C13064 a_14539_43914# a_15743_43084# 0.024623f
C13065 a_9313_44734# a_13667_43396# 2.37e-20
C13066 a_18326_43940# a_18451_43940# 0.145292f
C13067 a_17973_43940# a_15493_43396# 8.43e-20
C13068 a_11823_42460# a_13163_45724# 0.038493f
C13069 a_2711_45572# a_16115_45572# 0.00431f
C13070 a_9049_44484# a_8697_45822# 7.16e-20
C13071 C0_dummy_N_btm C10_P_btm 7.53e-19
C13072 C0_P_btm C8_P_btm 0.146541f
C13073 C1_P_btm C7_P_btm 0.128479f
C13074 C4_N_btm EN_VIN_BSTR_N 0.116925f
C13075 C0_dummy_P_btm C9_P_btm 0.111645f
C13076 a_14021_43940# a_12741_44636# 2.11e-19
C13077 a_4093_43548# a_3090_45724# 0.00131f
C13078 a_n2661_42834# a_n2661_45546# 0.029567f
C13079 a_7911_44260# a_5937_45572# 2.23e-20
C13080 a_n722_43218# a_n1613_43370# 0.00237f
C13081 a_16795_42852# a_16327_47482# 6.73e-19
C13082 a_5534_30871# a_10227_46804# 0.304847f
C13083 a_19164_43230# a_12861_44030# 5.09e-21
C13084 a_19466_46812# VDD 0.664497f
C13085 a_1823_45246# a_4185_45028# 0.081652f
C13086 a_2698_46116# a_2804_46116# 0.313533f
C13087 a_167_45260# a_3483_46348# 1.26e-19
C13088 a_11813_46116# a_12638_46436# 3.97e-19
C13089 a_11415_45002# a_12005_46116# 1.53e-20
C13090 a_20411_46873# a_19900_46494# 6.79e-19
C13091 a_20107_46660# a_20708_46348# 2.61e-20
C13092 a_20273_46660# a_20075_46420# 5.46e-21
C13093 a_19123_46287# a_6945_45028# 1.85e-19
C13094 a_17829_46910# a_10809_44734# 0.02024f
C13095 a_5932_42308# a_6886_37412# 5.75e-19
C13096 a_19319_43548# a_10341_43396# 0.027205f
C13097 a_2982_43646# a_3539_42460# 0.01563f
C13098 a_3540_43646# a_3626_43646# 0.100706f
C13099 a_n1557_42282# a_648_43396# 0.048175f
C13100 a_9313_44734# a_20256_43172# 0.0039f
C13101 a_4699_43561# a_6197_43396# 9.72e-21
C13102 a_n97_42460# a_5837_43396# 6.05e-19
C13103 a_3499_42826# a_1847_42826# 0.006199f
C13104 a_n2109_47186# CLK_DATA 6.42e-19
C13105 a_2813_43396# VDD 0.004385f
C13106 a_2437_43646# a_2382_45260# 0.005858f
C13107 a_n2293_45010# a_n2810_45028# 7.12e-19
C13108 a_n2661_45010# en_comp 0.10363f
C13109 a_n2017_45002# a_n913_45002# 0.275686f
C13110 a_n2472_45002# a_n2956_37592# 0.152938f
C13111 a_22591_45572# a_413_45260# 0.003236f
C13112 a_10907_45822# a_11361_45348# 1.86e-19
C13113 a_10193_42453# a_19778_44110# 8.12e-21
C13114 a_16147_45260# a_14180_45002# 4.1e-21
C13115 a_22223_43396# a_4185_45028# 3.93e-19
C13116 a_9803_43646# a_526_44458# 0.170855f
C13117 a_n2129_43609# a_n863_45724# 0.003134f
C13118 a_n1699_43638# a_n2293_45546# 6.05e-20
C13119 a_17531_42308# a_13507_46334# 1.18e-20
C13120 a_21335_42336# a_16327_47482# 0.081786f
C13121 a_20205_31679# VDD 0.737305f
C13122 a_2711_45572# a_5807_45002# 0.065611f
C13123 a_5437_45600# a_n881_46662# 0.001471f
C13124 a_6812_45938# a_n1613_43370# 0.00201f
C13125 a_13527_45546# a_11453_44696# 4.99e-21
C13126 a_10809_44734# a_n443_42852# 3.02e-20
C13127 a_5066_45546# a_n2661_45546# 9.86e-19
C13128 a_526_44458# a_310_45028# 1.77e-21
C13129 a_n97_42460# a_18695_43230# 0.001854f
C13130 a_10807_43548# a_10533_42308# 4.25e-19
C13131 a_10341_43396# a_16795_42852# 1.46e-20
C13132 a_22959_43396# a_17364_32525# 0.156288f
C13133 a_10467_46802# CLK 0.028547f
C13134 a_6755_46942# DATA[3] 6.6e-21
C13135 a_n2946_37984# a_n2860_37984# 0.011479f
C13136 a_n3420_37984# a_n2216_37984# 5.9e-20
C13137 a_13348_45260# a_12607_44458# 5.28e-21
C13138 a_13017_45260# a_13076_44458# 0.011055f
C13139 a_1423_45028# a_2779_44458# 0.246285f
C13140 a_1307_43914# a_6298_44484# 4.3e-19
C13141 a_9482_43914# a_8975_43940# 0.186623f
C13142 a_18479_45785# a_20362_44736# 2.03e-36
C13143 a_626_44172# a_n699_43396# 0.042617f
C13144 a_2711_45572# a_19478_44306# 0.006321f
C13145 a_2382_45260# a_4181_44734# 7.54e-21
C13146 a_5934_30871# a_4185_45028# 0.060401f
C13147 a_19339_43156# a_n357_42282# 0.008506f
C13148 a_n2472_42282# a_n2956_39304# 2.99e-20
C13149 a_n3674_38680# a_n2956_38680# 0.023107f
C13150 a_3080_42308# RST_Z 0.00595f
C13151 VIN_P VDD 1.47957f
C13152 a_2711_45572# a_3699_46348# 2.78e-20
C13153 a_10490_45724# a_11415_45002# 1.25e-19
C13154 a_13777_45326# a_n743_46660# 1.09e-20
C13155 a_17786_45822# a_3090_45724# 0.003629f
C13156 a_3357_43084# a_10150_46912# 1.08e-20
C13157 a_413_45260# a_4646_46812# 3.52e-20
C13158 a_16922_45042# a_11453_44696# 0.07136f
C13159 a_18184_42460# a_13507_46334# 0.505552f
C13160 a_18911_45144# a_4883_46098# 8.04e-21
C13161 a_8103_44636# a_4791_45118# 0.048713f
C13162 a_11827_44484# a_18597_46090# 0.039373f
C13163 a_11691_44458# a_10227_46804# 0.012084f
C13164 a_16243_43396# a_4958_30871# 2.01e-19
C13165 a_10991_42826# a_n784_42308# 4.32e-21
C13166 a_2905_42968# a_2713_42308# 1.96e-19
C13167 a_743_42282# a_11551_42558# 0.014689f
C13168 a_16137_43396# a_17303_42282# 8.65e-19
C13169 a_1847_42826# a_3318_42354# 9.4e-21
C13170 a_20692_30879# a_22821_38993# 8.99e-20
C13171 a_20205_31679# a_22469_39537# 4.7e-20
C13172 a_n1151_42308# a_n743_46660# 0.195953f
C13173 a_n2109_47186# a_3699_46634# 6.42e-20
C13174 a_584_46384# a_383_46660# 0.001651f
C13175 a_n815_47178# a_n2661_46098# 3.57e-20
C13176 a_3785_47178# a_n1925_46634# 3.96e-20
C13177 a_3160_47472# a_n2438_43548# 3.61e-21
C13178 a_n746_45260# a_479_46660# 0.001012f
C13179 a_4915_47217# a_n2661_46634# 9.46e-19
C13180 a_9313_45822# a_5807_45002# 0.031627f
C13181 a_13487_47204# a_13675_47204# 0.001217f
C13182 a_12861_44030# a_13759_47204# 0.001988f
C13183 a_15507_47210# a_768_44030# 5.43e-20
C13184 a_15811_47375# a_12549_44172# 0.024519f
C13185 a_n2293_45010# a_n2129_43609# 8.68e-20
C13186 a_n2661_45010# a_n1699_43638# 6.02e-20
C13187 a_n2017_45002# a_n4318_39304# 9.41e-20
C13188 a_5111_44636# a_8487_44056# 0.004423f
C13189 en_comp a_21381_43940# 3.87e-21
C13190 a_14539_43914# a_16789_44484# 3.44e-19
C13191 a_1307_43914# a_10555_44260# 5.81e-19
C13192 a_18443_44721# a_17517_44484# 0.029904f
C13193 a_13556_45296# a_14021_43940# 1.12e-19
C13194 a_5891_43370# a_n2661_43922# 0.042536f
C13195 a_n2840_44458# a_n2840_43914# 0.026152f
C13196 a_n4209_39590# a_n2956_38216# 0.021267f
C13197 a_19479_31679# VDD 0.579914f
C13198 a_45_45144# a_167_45260# 0.002149f
C13199 a_4185_45348# a_4185_45028# 0.009825f
C13200 a_2448_45028# a_1823_45246# 7.38e-19
C13201 a_14976_45348# a_11415_45002# 7.17e-19
C13202 a_20567_45036# a_20273_46660# 4.15e-22
C13203 a_10157_44484# a_3090_45724# 5.31e-20
C13204 a_11691_44458# a_17339_46660# 0.018074f
C13205 a_20512_43084# a_13661_43548# 0.00101f
C13206 a_20637_44484# a_19321_45002# 1.7e-20
C13207 a_21145_44484# a_13747_46662# 8.01e-19
C13208 a_18479_45785# a_16375_45002# 1.81e-19
C13209 a_n913_45002# a_526_44458# 0.250864f
C13210 a_n1059_45260# a_n1925_42282# 0.023119f
C13211 a_20719_45572# a_8049_45260# 6.29e-19
C13212 a_13348_45260# a_10903_43370# 0.011259f
C13213 a_1423_45028# a_6165_46155# 4.27e-22
C13214 a_13017_45260# a_12594_46348# 4.35e-20
C13215 a_1307_43914# a_5937_45572# 0.101589f
C13216 a_895_43940# a_n1613_43370# 8.02e-21
C13217 a_6709_45028# a_2324_44458# 0.076559f
C13218 a_5934_30871# a_9803_42558# 0.001422f
C13219 a_8337_42558# a_8325_42308# 0.01416f
C13220 a_14097_32519# a_22775_42308# 0.001341f
C13221 a_6171_42473# a_5742_30871# 1.16e-20
C13222 EN_VIN_BSTR_P C3_P_btm 0.100325f
C13223 a_n1925_46634# a_3090_45724# 8.91e-20
C13224 a_5907_46634# a_7715_46873# 8.55e-21
C13225 a_6540_46812# a_5257_43370# 0.00507f
C13226 a_5732_46660# a_7411_46660# 1.96e-20
C13227 a_12549_44172# a_13059_46348# 0.808395f
C13228 a_5807_45002# a_12513_46660# 7.17e-19
C13229 a_12465_44636# a_20202_43084# 8.04e-20
C13230 a_22223_47212# a_22365_46825# 0.011422f
C13231 a_13507_46334# a_12741_44636# 0.137731f
C13232 a_11453_44696# a_21350_47026# 3.86e-19
C13233 a_6545_47178# a_6419_46155# 0.080336f
C13234 a_4915_47217# a_8199_44636# 2.73e-20
C13235 a_n1151_42308# a_11189_46129# 0.12414f
C13236 a_4791_45118# a_8953_45546# 1.45e-19
C13237 a_n443_46116# a_5937_45572# 4.89e-20
C13238 a_3422_30871# a_11341_43940# 0.030182f
C13239 a_5883_43914# a_7112_43396# 2.7e-20
C13240 a_n356_44636# a_4093_43548# 1.07e-21
C13241 a_20512_43084# a_19862_44208# 0.023947f
C13242 a_n699_43396# a_2813_43396# 0.001609f
C13243 a_3232_43370# a_10796_42968# 1.9e-20
C13244 en_comp a_18249_42858# 8.38e-21
C13245 a_n913_45002# a_19164_43230# 8.4e-21
C13246 a_n2017_45002# a_20922_43172# 1.61e-20
C13247 a_5289_44734# VDD 5.21e-19
C13248 a_n4064_39616# VREF 1.53e-20
C13249 a_n4064_39072# C2_P_btm 1.14e-20
C13250 a_n3420_39616# VCM 0.0424f
C13251 a_n4064_38528# EN_VIN_BSTR_P 0.032853f
C13252 a_5263_45724# a_5907_45546# 0.001537f
C13253 a_2711_45572# a_6511_45714# 0.04109f
C13254 VDAC_N a_20692_30879# 9.25e-19
C13255 a_20512_43084# a_4185_45028# 2.96e-20
C13256 a_8147_43396# a_n2293_46634# 0.011922f
C13257 a_15493_43940# a_19692_46634# 0.16692f
C13258 a_12429_44172# a_13059_46348# 8.69e-20
C13259 a_n2661_44458# a_380_45546# 2.29e-20
C13260 a_n2129_44697# a_n863_45724# 2.81e-19
C13261 a_556_44484# a_526_44458# 0.077901f
C13262 a_12883_44458# a_13259_45724# 0.003043f
C13263 a_n1699_44726# a_n2293_45546# 0.001074f
C13264 a_17517_44484# a_17583_46090# 5.71e-21
C13265 a_15743_43084# a_11453_44696# 9.67e-22
C13266 a_19095_43396# a_16327_47482# 6.39e-19
C13267 a_4190_30871# a_10227_46804# 6.29e-20
C13268 a_20447_31679# a_22459_39145# 2.66e-20
C13269 a_19963_31679# a_22521_39511# 2.93e-20
C13270 a_19479_31679# a_22469_39537# 3.29e-20
C13271 a_n4064_39072# a_n2302_38778# 2.59e-20
C13272 a_n2302_39072# a_n4064_38528# 2.59e-20
C13273 a_22000_46634# a_11415_45002# 1.58e-19
C13274 a_21188_46660# a_22591_46660# 1.52e-20
C13275 a_20623_46660# a_12741_44636# 0.034292f
C13276 a_21363_46634# a_20820_30879# 2.73e-19
C13277 a_12991_46634# a_10903_43370# 1.94e-19
C13278 a_6755_46942# a_6945_45028# 0.024014f
C13279 a_12251_46660# a_12005_46116# 8.94e-19
C13280 a_12469_46902# a_12594_46348# 4.31e-19
C13281 a_n881_46662# a_n443_42852# 0.005862f
C13282 a_21588_30879# a_20692_30879# 0.056225f
C13283 a_22612_30879# a_20205_31679# 0.111294f
C13284 a_768_44030# a_2957_45546# 0.027276f
C13285 a_10807_43548# a_9885_43646# 1.34e-20
C13286 a_n2293_42834# a_6171_42473# 2.63e-20
C13287 a_9313_44734# a_21195_42852# 0.02195f
C13288 a_19319_43548# a_n97_42460# 0.029676f
C13289 a_1467_44172# a_743_42282# 3.61e-22
C13290 a_10949_43914# a_10341_43396# 4.22e-20
C13291 a_15037_43940# VDD 0.190221f
C13292 a_10193_42453# a_9482_43914# 0.029531f
C13293 a_19431_45546# a_20107_45572# 0.001119f
C13294 a_11652_45724# a_11787_45002# 0.077604f
C13295 a_11525_45546# a_11963_45334# 2.67e-19
C13296 a_18596_45572# a_18787_45572# 4.61e-19
C13297 a_11322_45546# a_13017_45260# 0.003434f
C13298 a_11823_42460# a_8953_45002# 1.65e-20
C13299 a_9127_43156# a_8270_45546# 0.002724f
C13300 a_4190_30871# a_17339_46660# 0.005828f
C13301 a_15493_43940# a_20692_30879# 1.18e-20
C13302 a_15037_44260# a_13259_45724# 3.72e-21
C13303 a_14021_43940# a_16375_45002# 3.38e-20
C13304 a_8791_43396# a_8953_45546# 0.012124f
C13305 VDAC_N VIN_N 0.256435f
C13306 a_n2956_38680# VDD 0.871805f
C13307 a_11322_45546# a_2063_45854# 0.105268f
C13308 a_10053_45546# a_n1151_42308# 2.02e-20
C13309 a_2711_45572# a_14311_47204# 3.64e-21
C13310 a_167_45260# a_n357_42282# 0.148401f
C13311 a_2202_46116# a_n755_45592# 2.03e-20
C13312 a_376_46348# a_n356_45724# 7.46e-20
C13313 a_n2293_46098# a_1609_45822# 0.002761f
C13314 a_1337_46436# a_1337_46116# 6.96e-20
C13315 a_6945_45028# a_8049_45260# 0.009745f
C13316 a_13759_46122# a_14949_46494# 2.56e-19
C13317 a_14955_43396# a_4361_42308# 3.74e-21
C13318 a_11967_42832# a_15890_42674# 0.001386f
C13319 a_17324_43396# a_15743_43084# 0.050725f
C13320 a_18429_43548# a_18783_43370# 0.001885f
C13321 a_n97_42460# a_16795_42852# 0.126591f
C13322 a_20974_43370# a_21195_42852# 1.06e-20
C13323 a_3905_42865# a_3823_42558# 1.35e-19
C13324 a_3626_43646# a_7765_42852# 3.92e-20
C13325 a_2982_43646# a_8605_42826# 2.81e-20
C13326 a_n2661_42282# a_n4318_37592# 0.03806f
C13327 a_16409_43396# a_16867_43762# 0.027606f
C13328 a_10341_43396# a_19095_43396# 0.004123f
C13329 a_21381_43940# a_22165_42308# 1.75e-19
C13330 a_n2661_46634# DATA[5] 6.56e-19
C13331 a_21588_30879# VIN_N 0.106594f
C13332 a_15279_43071# VDD 0.189193f
C13333 a_n2810_45028# a_n4334_37440# 6.16e-20
C13334 a_n2956_37592# a_n4209_37414# 0.145558f
C13335 a_3357_43084# a_4223_44672# 0.029613f
C13336 a_n2109_45247# a_n2433_44484# 1.13e-19
C13337 a_n2661_45010# a_n1699_44726# 0.04137f
C13338 a_n2293_45010# a_n2129_44697# 0.021404f
C13339 a_n2017_45002# a_n2661_44458# 0.034362f
C13340 a_18691_45572# a_18989_43940# 1.88e-19
C13341 a_13017_45260# a_15060_45348# 7e-21
C13342 a_13556_45296# a_13711_45394# 0.005081f
C13343 a_18799_45938# a_18248_44752# 5.06e-22
C13344 a_14113_42308# a_3090_45724# 2.41e-20
C13345 a_12800_43218# a_9290_44172# 1.74e-20
C13346 a_14021_43940# RST_Z 0.007254f
C13347 a_11962_45724# a_11735_46660# 4.42e-20
C13348 a_7499_43078# a_3090_45724# 0.23734f
C13349 a_2711_45572# a_14226_46987# 3.21e-22
C13350 a_19479_31679# a_22612_30879# 0.064572f
C13351 a_413_45260# a_9804_47204# 6.79e-20
C13352 a_3065_45002# a_n1613_43370# 1.12e-20
C13353 a_13017_45260# a_12465_44636# 1.71e-20
C13354 a_10775_45002# a_11453_44696# 6.82e-19
C13355 a_8016_46348# CLK 0.001431f
C13356 a_5937_45572# DATA[4] 8.55e-21
C13357 a_3626_43646# a_13657_42308# 0.00116f
C13358 a_13678_32519# a_22400_42852# 0.035124f
C13359 a_7871_42858# a_9061_43230# 2.56e-19
C13360 a_19164_43230# a_20922_43172# 8.1e-20
C13361 a_13467_32519# a_20256_42852# 2.92e-20
C13362 a_13258_32519# VDD 3.19231f
C13363 a_n2109_47186# a_2583_47243# 8.31e-19
C13364 a_n971_45724# a_2487_47570# 6.45e-19
C13365 a_n1741_47186# a_3315_47570# 2.13e-19
C13366 a_n1435_47204# a_13717_47436# 0.196889f
C13367 a_13381_47204# a_12861_44030# 4.15e-20
C13368 a_n237_47217# a_n89_47570# 0.005668f
C13369 a_n785_47204# a_n2312_39304# 9.48e-20
C13370 a_17613_45144# a_17517_44484# 1.32e-20
C13371 a_16979_44734# a_17767_44458# 0.011457f
C13372 a_14539_43914# a_17970_44736# 2.85e-19
C13373 a_1307_43914# a_2479_44172# 0.300587f
C13374 a_11691_44458# a_14815_43914# 0.018499f
C13375 a_11823_42460# a_3626_43646# 0.011402f
C13376 a_375_42282# a_453_43940# 0.021162f
C13377 a_626_44172# a_1467_44172# 4.19e-19
C13378 a_7499_43078# a_6547_43396# 1.37e-19
C13379 a_11827_44484# a_10809_44484# 2.9e-20
C13380 a_n2017_45002# a_18451_43940# 4.02e-22
C13381 a_3537_45260# a_n2661_42282# 0.105917f
C13382 a_n1059_45260# a_18326_43940# 7.46e-21
C13383 a_8515_42308# a_n755_45592# 0.003799f
C13384 a_n4315_30879# a_n1925_42282# 3.26e-20
C13385 a_15890_42674# a_13259_45724# 8.67e-20
C13386 a_3065_45002# a_n2293_46098# 2.43e-19
C13387 a_4223_44672# a_3877_44458# 0.007855f
C13388 a_6171_45002# a_11415_45002# 1.05801f
C13389 a_11827_44484# a_6755_46942# 0.529579f
C13390 a_9159_44484# a_768_44030# 0.003496f
C13391 a_n745_45366# a_167_45260# 7.9e-20
C13392 a_n2661_42834# a_12891_46348# 9.68e-21
C13393 a_3775_45552# a_n2661_45546# 0.006201f
C13394 a_2711_45572# a_n755_45592# 0.168218f
C13395 a_11280_45822# a_8049_45260# 1.62e-19
C13396 a_10490_45724# a_13259_45724# 1.48e-19
C13397 a_n2661_43922# a_11309_47204# 1.06e-21
C13398 a_18479_45785# a_18985_46122# 1.04e-21
C13399 a_18341_45572# a_18819_46122# 0.00524f
C13400 a_20362_44736# a_13507_46334# 5.2e-22
C13401 a_2479_44172# a_n443_46116# 0.732848f
C13402 a_18579_44172# a_18479_47436# 1.01e-20
C13403 a_3422_30871# a_16327_47482# 0.220296f
C13404 a_22959_42860# a_22775_42308# 0.019713f
C13405 a_1576_42282# a_1755_42282# 0.168925f
C13406 a_1184_42692# a_1606_42308# 0.125247f
C13407 a_n784_42308# a_2713_42308# 2.26e-20
C13408 a_13291_42460# a_13070_42354# 0.155164f
C13409 a_n3674_37592# a_n39_42308# 0.003612f
C13410 a_n2833_47464# a_n2840_46090# 2.94e-20
C13411 a_5807_45002# a_6540_46812# 0.007069f
C13412 a_n1925_46634# a_3699_46634# 0.014429f
C13413 a_n133_46660# a_2443_46660# 4.17e-21
C13414 a_171_46873# a_n2661_46098# 0.168482f
C13415 a_383_46660# a_479_46660# 0.013793f
C13416 a_601_46902# a_645_46660# 3.69e-19
C13417 a_n2438_43548# a_2609_46660# 8.62e-19
C13418 a_33_46660# a_1799_45572# 3.91e-21
C13419 a_13717_47436# a_13885_46660# 0.003475f
C13420 a_4915_47217# a_765_45546# 0.169406f
C13421 a_12861_44030# a_13170_46660# 9.11e-20
C13422 a_18479_47436# a_17609_46634# 3.14e-19
C13423 a_10227_46804# a_15227_44166# 0.013242f
C13424 a_4883_46098# a_12991_46634# 8.79e-20
C13425 a_9804_47204# a_9863_46634# 0.017882f
C13426 a_n2661_45010# a_n2157_42858# 4.56e-21
C13427 en_comp a_5649_42852# 2.63e-19
C13428 a_n2293_43922# a_10949_43914# 0.008394f
C13429 a_n2661_43370# a_7287_43370# 3.73e-21
C13430 a_9313_44734# a_15493_43396# 0.001749f
C13431 a_n2661_42834# a_11750_44172# 0.006203f
C13432 a_n2661_43922# a_10807_43548# 2.2e-19
C13433 a_22959_44484# a_19237_31679# 0.155744f
C13434 a_3754_38802# VDD 0.002173f
C13435 a_20193_45348# VDD 0.793111f
C13436 a_4958_30871# a_n923_35174# 0.015856f
C13437 a_15764_42576# RST_Z 1.86e-19
C13438 a_5742_30871# VIN_N 0.042613f
C13439 a_9313_44734# a_3483_46348# 0.015646f
C13440 a_14673_44172# a_11415_45002# 0.229077f
C13441 a_5708_44484# a_1823_45246# 5.34e-19
C13442 a_3600_43914# a_3090_45724# 3.95e-19
C13443 a_19478_44056# a_19321_45002# 1.84e-21
C13444 a_n2661_44458# a_526_44458# 0.087308f
C13445 a_1307_43914# a_n443_42852# 0.05746f
C13446 a_2448_45028# a_n2293_45546# 9.06e-19
C13447 a_45_45144# a_n863_45724# 2.41e-19
C13448 a_11827_44484# a_8049_45260# 1.09e-19
C13449 a_458_43396# a_n1613_43370# 4.14e-20
C13450 a_5159_47243# VDD 2.18e-20
C13451 a_n784_42308# C8_N_btm 6.79e-20
C13452 a_1606_42308# C0_P_btm 0.029189f
C13453 a_5534_30871# VDAC_P 0.004862f
C13454 a_5342_30871# VDAC_N 0.011631f
C13455 a_5257_43370# a_1823_45246# 0.003231f
C13456 a_15227_44166# a_17339_46660# 0.524034f
C13457 a_13885_46660# a_14035_46660# 0.25868f
C13458 a_17609_46634# a_17829_46910# 0.111805f
C13459 a_n2840_46634# a_n2956_39304# 0.001899f
C13460 a_8128_46384# a_8062_46482# 7.91e-19
C13461 a_n881_46662# a_6633_46155# 8.73e-19
C13462 a_4646_46812# a_6165_46155# 3.41e-20
C13463 a_3877_44458# a_6419_46155# 0.002843f
C13464 a_4651_46660# a_5497_46414# 2.21e-19
C13465 a_4817_46660# a_5164_46348# 5.41e-19
C13466 a_n2661_46634# a_10809_44734# 0.023983f
C13467 a_4955_46873# a_5204_45822# 3.57e-19
C13468 a_12465_44636# a_14383_46116# 0.00348f
C13469 a_13507_46334# a_16375_45002# 0.002576f
C13470 a_4883_46098# a_18147_46436# 2.8e-19
C13471 a_18479_47436# a_19443_46116# 3.9e-22
C13472 a_18597_46090# a_20009_46494# 8.96e-19
C13473 a_n443_46116# a_n443_42852# 0.145452f
C13474 a_3422_30871# a_10341_43396# 0.029183f
C13475 a_11967_42832# a_16547_43609# 0.176385f
C13476 a_n356_44636# a_685_42968# 3.75e-19
C13477 a_19862_44208# a_21381_43940# 0.113704f
C13478 a_3499_42826# a_4235_43370# 4.6e-20
C13479 a_15493_43396# a_20974_43370# 1.15e-20
C13480 a_18479_45785# a_17303_42282# 1.31e-20
C13481 a_3065_45002# a_3905_42558# 0.044632f
C13482 a_n2017_45002# a_8325_42308# 0.009217f
C13483 a_9028_43914# VDD 0.17194f
C13484 a_15225_45822# a_15765_45572# 2.89e-20
C13485 a_n3420_37984# C7_P_btm 2.68e-20
C13486 a_21381_43940# a_4185_45028# 1.24e-20
C13487 a_18249_42858# a_13661_43548# 2.04e-19
C13488 a_15781_43660# a_3090_45724# 5.85e-20
C13489 a_n2065_43946# a_n1079_45724# 5.59e-22
C13490 a_n1549_44318# a_n2661_45546# 1.94e-21
C13491 a_n1761_44111# a_n2293_45546# 2.91e-20
C13492 a_n473_42460# a_n1151_42308# 0.006908f
C13493 a_18504_43218# a_16327_47482# 0.002118f
C13494 a_14635_42282# a_10227_46804# 0.008414f
C13495 a_n1423_46090# VDD 0.227012f
C13496 C0_dummy_P_btm C0_N_btm 1.3e-19
C13497 C0_P_btm C1_N_btm 2.15e-19
C13498 C1_P_btm C2_N_btm 2.79e-20
C13499 a_2698_46116# a_n1925_42282# 1.04e-20
C13500 a_1823_45246# a_1337_46116# 1.69e-19
C13501 a_3147_46376# a_2981_46116# 0.003565f
C13502 a_2804_46116# a_526_44458# 0.00297f
C13503 a_n4064_40160# a_n3565_37414# 4.29714f
C13504 a_n4315_30879# a_n3420_37440# 0.039346f
C13505 a_n4209_38502# a_n4064_37984# 0.028133f
C13506 a_n3565_38502# a_n3420_37984# 0.028236f
C13507 a_n3690_38528# a_n3690_38304# 0.052468f
C13508 a_14493_46090# a_14840_46494# 0.051162f
C13509 a_8199_44636# a_10809_44734# 0.022266f
C13510 a_8953_45546# a_6945_45028# 2.77e-19
C13511 a_13925_46122# a_2324_44458# 4.65e-20
C13512 a_13759_46122# a_15682_46116# 1.44e-20
C13513 a_n97_42460# a_19095_43396# 0.003217f
C13514 a_5891_43370# a_10545_42558# 1.64e-20
C13515 a_3422_30871# a_20356_42852# 3.72e-19
C13516 a_20512_43084# a_20573_43172# 0.00112f
C13517 a_9396_43370# a_9885_43396# 4.89e-20
C13518 a_n4318_40392# a_n4315_30879# 0.151169f
C13519 a_n356_44636# a_14113_42308# 0.019853f
C13520 a_15493_43396# a_18599_43230# 5.54e-20
C13521 a_11341_43940# a_16414_43172# 3.69e-21
C13522 a_2982_43646# a_18783_43370# 4.48e-21
C13523 a_8685_43396# a_14358_43442# 0.002184f
C13524 a_19328_44172# a_19339_43156# 1.37e-19
C13525 a_13507_46334# RST_Z 0.004909f
C13526 a_20990_47178# SINGLE_ENDED 0.067698f
C13527 a_21177_47436# START 7.35e-20
C13528 a_20301_43646# VDD 0.296691f
C13529 a_18341_45572# a_18911_45144# 0.006584f
C13530 a_13249_42308# a_13720_44458# 1.19e-19
C13531 a_8192_45572# a_5343_44458# 6.07e-21
C13532 a_7499_43078# a_n356_44636# 4.62e-19
C13533 a_18479_45785# a_19778_44110# 0.009f
C13534 a_327_44734# a_626_44172# 0.120093f
C13535 a_2680_45002# a_1307_43914# 9.4e-20
C13536 a_6171_45002# a_13159_45002# 0.012283f
C13537 a_3357_43084# a_n2293_42834# 0.045124f
C13538 a_n2293_45010# a_45_45144# 3.59e-21
C13539 a_7705_45326# a_8953_45002# 1.82e-20
C13540 a_18249_42858# a_4185_45028# 3.07e-20
C13541 a_13258_32519# a_22612_30879# 0.065697f
C13542 a_9396_43370# a_n443_42852# 0.039136f
C13543 a_16547_43609# a_13259_45724# 3.22e-20
C13544 a_n4318_38680# a_n2956_38680# 0.023283f
C13545 a_10835_43094# a_10903_43370# 0.001283f
C13546 a_10341_42308# a_9290_44172# 0.051084f
C13547 a_8696_44636# a_12549_44172# 0.035105f
C13548 a_3065_45002# a_4791_45118# 0.006346f
C13549 a_2680_45002# a_n443_46116# 0.009148f
C13550 a_5111_44636# a_n1151_42308# 8.63e-19
C13551 a_413_45260# a_6545_47178# 3.66e-19
C13552 a_20885_45572# a_18479_47436# 6.01e-19
C13553 a_19963_31679# a_16327_47482# 1.05e-19
C13554 a_2437_43646# a_10227_46804# 0.150025f
C13555 a_3357_43084# a_16763_47508# 4.84e-19
C13556 a_21363_45546# a_13507_46334# 3.97e-19
C13557 a_20841_45814# a_4883_46098# 5.36e-20
C13558 a_20731_45938# a_20894_47436# 3.6e-21
C13559 a_n2661_45546# a_3218_45724# 0.010947f
C13560 a_n863_45724# a_n357_42282# 0.172013f
C13561 a_n1079_45724# a_n755_45592# 0.109544f
C13562 a_380_45546# a_n1099_45572# 0.148825f
C13563 a_n452_45724# a_310_45028# 5.77e-21
C13564 a_4361_42308# a_n2293_42282# 2.71e-21
C13565 a_4093_43548# a_3823_42558# 1.14e-20
C13566 a_5649_42852# a_22165_42308# 0.077779f
C13567 a_7765_42852# a_8037_42858# 0.309282f
C13568 a_7871_42858# a_8605_42826# 0.06628f
C13569 a_13678_32519# a_22223_42860# 0.002285f
C13570 a_3080_42308# a_2713_42308# 0.004874f
C13571 a_14021_43940# a_17303_42282# 3.16e-21
C13572 a_15493_43940# a_20107_42308# 7.88e-22
C13573 a_15095_43370# a_14853_42852# 6.13e-21
C13574 a_14579_43548# a_16245_42852# 6.32e-20
C13575 a_13887_32519# a_21195_42852# 9.75e-21
C13576 a_765_45546# DATA[5] 0.027477f
C13577 a_20623_46660# RST_Z 2.19e-20
C13578 a_20273_46660# SINGLE_ENDED 1.13e-20
C13579 VDAC_Ni a_5088_37509# 1.70462f
C13580 a_3754_38470# a_3726_37500# 0.554457f
C13581 a_n3565_37414# a_n4064_37440# 0.230258f
C13582 a_5421_42558# VDD 0.007373f
C13583 a_n971_45724# a_584_46384# 0.152617f
C13584 a_n237_47217# a_1431_47204# 0.045044f
C13585 a_n1741_47186# a_3160_47472# 0.012286f
C13586 a_n2109_47186# a_3381_47502# 0.035813f
C13587 a_n23_47502# a_1239_47204# 8.7e-21
C13588 a_n785_47204# a_1209_47178# 3.43e-19
C13589 a_n1920_47178# a_n1151_42308# 8.17e-19
C13590 a_6171_45002# a_11967_42832# 5.32e-19
C13591 a_n2661_45010# a_n1761_44111# 8.36e-20
C13592 a_2437_43646# a_453_43940# 1.7e-19
C13593 a_n2293_45010# a_n2472_43914# 1.49e-19
C13594 a_5837_45028# a_5891_43370# 6.5e-21
C13595 a_8696_44636# a_12429_44172# 2.76e-20
C13596 a_n2661_43370# a_n23_44458# 9.21e-19
C13597 a_n2840_44458# a_n2661_44458# 0.179135f
C13598 a_16115_45572# a_15682_43940# 2.15e-19
C13599 a_13003_42852# a_n443_42852# 1.06e-19
C13600 a_17665_42852# a_n357_42282# 8.95e-19
C13601 a_15037_45618# a_3483_46348# 1.96e-21
C13602 a_18909_45814# a_11415_45002# 0.002265f
C13603 a_18175_45572# a_12741_44636# 7.5e-20
C13604 a_20107_45572# a_20528_46660# 5.09e-21
C13605 a_15595_45028# a_6755_46942# 0.012879f
C13606 a_n2293_42834# a_3877_44458# 3.47e-22
C13607 a_5907_45546# a_526_44458# 3.52e-20
C13608 a_413_45260# a_19692_46634# 6.26e-20
C13609 a_4558_45348# a_3090_45724# 0.147318f
C13610 a_2437_43646# a_17339_46660# 3.78e-20
C13611 a_11962_45724# a_2324_44458# 0.004603f
C13612 a_11823_42460# a_15015_46420# 0.001494f
C13613 a_13904_45546# a_13759_46122# 0.008324f
C13614 a_8192_45572# a_8349_46414# 2.67e-20
C13615 a_10907_45822# a_9625_46129# 2.68e-19
C13616 a_14495_45572# a_12594_46348# 5.14e-20
C13617 a_6812_45938# a_6945_45028# 0.002475f
C13618 a_6298_44484# a_n1613_43370# 0.02075f
C13619 a_17970_44736# a_11453_44696# 0.008957f
C13620 a_15433_44458# a_4915_47217# 3.72e-20
C13621 a_5342_30871# a_5742_30871# 0.031909f
C13622 a_13635_43156# a_13575_42558# 0.00691f
C13623 a_3080_42308# C8_N_btm 0.006767f
C13624 a_768_44030# a_13747_46662# 0.434325f
C13625 a_n881_46662# a_n2661_46634# 0.035376f
C13626 a_6151_47436# a_10150_46912# 0.006237f
C13627 a_6575_47204# a_7577_46660# 3.98e-19
C13628 a_7903_47542# a_8145_46902# 0.010369f
C13629 a_4915_47217# a_10623_46897# 0.002626f
C13630 a_2063_45854# a_8654_47026# 1.72e-19
C13631 a_19778_44110# a_14021_43940# 4.06e-19
C13632 a_4223_44672# a_9672_43914# 4.35e-21
C13633 a_14673_44172# a_11967_42832# 3.97e-20
C13634 a_10193_42453# a_10796_42968# 0.015009f
C13635 a_17517_44484# a_17325_44484# 1.97e-19
C13636 a_5883_43914# a_6101_44260# 0.001046f
C13637 a_5343_44458# a_8018_44260# 0.003899f
C13638 a_20193_45348# a_22959_43948# 2.96e-19
C13639 a_5691_45260# a_6031_43396# 1.62e-21
C13640 a_5111_44636# a_6197_43396# 0.025934f
C13641 a_3537_45260# a_7112_43396# 0.046531f
C13642 a_n2017_45002# a_9145_43396# 2.64e-19
C13643 a_n784_42308# C2_P_btm 0.005178f
C13644 a_12607_44458# a_11415_45002# 1.53e-19
C13645 a_14955_43940# a_13661_43548# 0.010124f
C13646 a_20365_43914# a_12549_44172# 0.069119f
C13647 a_14815_43914# a_15227_44166# 4.45e-19
C13648 a_n2661_42282# a_n2293_46634# 0.039408f
C13649 a_15595_45028# a_8049_45260# 2.98e-20
C13650 a_6171_45002# a_13259_45724# 0.068737f
C13651 a_n745_45366# a_n863_45724# 7.61e-20
C13652 a_413_45260# a_20692_30879# 0.111034f
C13653 a_n2293_45010# a_n357_42282# 0.020718f
C13654 en_comp a_n2956_38216# 1.61e-19
C13655 a_n659_45366# a_n2661_45546# 5.25e-19
C13656 a_1427_43646# a_584_46384# 0.003548f
C13657 a_n144_43396# a_n971_45724# 0.010576f
C13658 a_17538_32519# a_12861_44030# 4.84e-19
C13659 a_19808_44306# a_16327_47482# 3.3e-21
C13660 a_15803_42450# a_4958_30871# 0.093396f
C13661 a_15764_42576# a_17303_42282# 1.02e-19
C13662 a_10723_42308# a_7174_31319# 9.76e-21
C13663 a_n3674_38216# a_n4334_38304# 0.059852f
C13664 a_15959_42545# a_16269_42308# 0.013793f
C13665 a_15890_42674# a_16197_42308# 3.69e-19
C13666 a_6123_31319# a_n4209_39590# 9.76e-22
C13667 a_5815_47464# VDD 0.399354f
C13668 a_4190_30871# VDAC_P 0.044618f
C13669 a_768_44030# a_4419_46090# 2.08e-20
C13670 a_n2661_46634# a_n2157_46122# 1.89e-19
C13671 a_n2472_46634# a_n2293_46098# 0.00197f
C13672 a_n2442_46660# a_n2472_46090# 6.07e-19
C13673 a_n743_46660# a_12741_44636# 9.6e-19
C13674 a_11453_44696# a_14840_46494# 7.84e-22
C13675 a_12465_44636# a_17715_44484# 1.19e-20
C13676 a_n1435_47204# a_n1925_42282# 4.56e-21
C13677 a_4883_46098# a_17957_46116# 0.013641f
C13678 a_13507_46334# a_18985_46122# 0.002665f
C13679 a_18143_47464# a_10809_44734# 0.006426f
C13680 a_18780_47178# a_6945_45028# 0.013003f
C13681 a_18479_47436# a_22223_46124# 5.82e-20
C13682 a_n1613_43370# a_5937_45572# 0.117604f
C13683 a_n881_46662# a_8199_44636# 2.26e-20
C13684 a_6755_46942# a_15559_46634# 1.64e-19
C13685 a_11823_42460# a_13921_42308# 3.14e-20
C13686 a_5663_43940# a_5829_43940# 0.143754f
C13687 a_10193_42453# a_4958_30871# 0.108497f
C13688 a_3422_30871# a_n97_42460# 3.53e-20
C13689 a_n356_44636# a_15781_43660# 6.74e-21
C13690 a_9313_44734# a_10695_43548# 2.41e-19
C13691 a_17737_43940# a_15493_43396# 1.12e-19
C13692 a_18079_43940# a_18451_43940# 9.65e-20
C13693 a_17973_43940# a_19328_44172# 4.29e-20
C13694 a_10729_43914# a_11341_43940# 0.243062f
C13695 a_20596_44850# VDD 4.6e-19
C13696 a_11823_42460# a_12791_45546# 0.030093f
C13697 a_7499_43078# a_8697_45822# 0.038073f
C13698 a_2711_45572# a_16333_45814# 9.94e-19
C13699 a_8568_45546# a_9241_45822# 7.63e-21
C13700 a_11962_45724# a_13527_45546# 1.48e-19
C13701 C0_dummy_P_btm C10_P_btm 0.749362f
C13702 C1_P_btm C8_P_btm 0.129306f
C13703 C0_P_btm C9_P_btm 0.146135f
C13704 C3_N_btm EN_VIN_BSTR_N 0.100325f
C13705 a_14021_43940# a_20820_30879# 1.28e-20
C13706 a_17737_43940# a_3483_46348# 8.22e-21
C13707 a_14761_44260# a_11415_45002# 1.35e-19
C13708 a_5649_42852# a_13661_43548# 3.72e-21
C13709 a_14673_44172# a_13259_45724# 0.006759f
C13710 a_9313_44734# a_n357_42282# 5.02008f
C13711 a_7584_44260# a_5937_45572# 2.31e-20
C13712 a_n967_43230# a_n1613_43370# 2.95e-19
C13713 a_14543_43071# a_10227_46804# 0.00196f
C13714 a_19339_43156# a_12861_44030# 1.64e-21
C13715 a_19333_46634# VDD 0.199048f
C13716 a_1823_45246# a_3699_46348# 2.62e-19
C13717 a_2202_46116# a_3483_46348# 9.66e-20
C13718 a_167_45260# a_3147_46376# 3.32e-19
C13719 a_15559_46634# a_8049_45260# 3.55e-20
C13720 a_11735_46660# a_12638_46436# 1.61e-19
C13721 a_11813_46116# a_12379_46436# 0.001157f
C13722 a_11415_45002# a_10903_43370# 0.085164f
C13723 a_n2293_46098# a_5937_45572# 0.078393f
C13724 a_765_45546# a_10809_44734# 2.52248f
C13725 a_20107_46660# a_19900_46494# 1.04e-19
C13726 a_20411_46873# a_20075_46420# 0.007002f
C13727 a_18285_46348# a_6945_45028# 1.31e-19
C13728 a_14815_43914# a_14635_42282# 1.04e-19
C13729 a_20623_43914# a_4361_42308# 3.31e-21
C13730 a_3080_42308# a_6031_43396# 9.6e-22
C13731 a_4699_43561# a_6293_42852# 5.22e-21
C13732 a_11341_43940# a_21487_43396# 0.005254f
C13733 a_20512_43084# a_21671_42860# 2.28e-19
C13734 a_19862_44208# a_5649_42852# 1.34e-20
C13735 a_4223_44672# a_5755_42308# 7.11e-21
C13736 a_2982_43646# a_3626_43646# 6.553431f
C13737 a_766_43646# a_648_43396# 1.98e-20
C13738 a_n1557_42282# a_548_43396# 0.005988f
C13739 a_15493_43940# a_743_42282# 5.64e-20
C13740 a_n1741_47186# RST_Z 7.39e-20
C13741 a_n2288_47178# CLK_DATA 6.87e-19
C13742 a_n2497_47436# DATA[0] 0.008757f
C13743 a_n2661_45010# a_n2956_37592# 0.163638f
C13744 a_n2293_45010# a_n745_45366# 5.55e-20
C13745 a_n2017_45002# a_n1059_45260# 6.27837f
C13746 a_2437_43646# a_2274_45254# 0.01398f
C13747 a_3357_43084# a_413_45260# 7.24598f
C13748 a_n2472_45002# a_n2810_45028# 0.002586f
C13749 a_n2840_45002# en_comp 8.04e-20
C13750 a_4099_45572# a_n2661_44458# 2.29e-20
C13751 a_5649_42852# a_4185_45028# 8.049951f
C13752 a_n2433_43396# a_n863_45724# 3.43e-22
C13753 a_9145_43396# a_526_44458# 0.004932f
C13754 a_20974_43370# a_n357_42282# 7.13e-19
C13755 a_n2267_43396# a_n2293_45546# 1.47e-20
C13756 a_n2302_38778# SMPL_ON_P 5.6e-20
C13757 a_7174_31319# a_16327_47482# 4.51e-19
C13758 a_17303_42282# a_13507_46334# 1.68549f
C13759 a_20062_46116# VDD 4.6e-19
C13760 a_6428_45938# a_n881_46662# 4.11e-19
C13761 a_14495_45572# a_12465_44636# 0.019417f
C13762 a_526_44458# a_n1099_45572# 1.36e-19
C13763 a_3422_30871# a_n3420_39616# 0.005543f
C13764 a_n97_42460# a_18504_43218# 0.002932f
C13765 a_6293_42852# a_6101_43172# 9.07e-19
C13766 a_14209_32519# a_17364_32525# 0.056697f
C13767 a_12281_43396# a_5534_30871# 0.012136f
C13768 a_10341_43396# a_16414_43172# 8.63e-20
C13769 a_10428_46928# CLK 0.032943f
C13770 a_n4064_37984# a_n3607_38304# 4.68e-19
C13771 a_n3420_37984# a_n2860_37984# 0.003211f
C13772 a_18909_45814# a_11967_42832# 4.13e-21
C13773 a_13017_45260# a_12883_44458# 7.59e-19
C13774 a_13159_45002# a_12607_44458# 4.65e-20
C13775 a_1423_45028# a_949_44458# 0.06121f
C13776 a_1307_43914# a_5518_44484# 0.01058f
C13777 a_9482_43914# a_10057_43914# 0.401746f
C13778 a_2711_45572# a_15493_43396# 0.054674f
C13779 a_7963_42308# a_4185_45028# 6.87e-20
C13780 a_13635_43156# a_n443_42852# 1.86e-19
C13781 a_18599_43230# a_n357_42282# 0.006999f
C13782 a_n2840_42282# a_n2956_38680# 2.5e-20
C13783 a_n2293_42282# a_n2810_45572# 3.09e-20
C13784 a_n3674_38680# a_n2956_39304# 0.023226f
C13785 a_3080_42308# C2_P_btm 0.108823f
C13786 a_2711_45572# a_3483_46348# 0.167588f
C13787 a_3175_45822# a_3147_46376# 0.001132f
C13788 a_5437_45600# a_n2293_46098# 4.86e-19
C13789 a_13556_45296# a_n743_46660# 3.23e-21
C13790 a_2809_45028# a_768_44030# 0.005501f
C13791 a_16377_45572# a_3090_45724# 3.99e-19
C13792 a_2437_43646# a_10467_46802# 1.48e-20
C13793 a_413_45260# a_3877_44458# 3.15e-19
C13794 a_3357_43084# a_9863_46634# 1.66e-20
C13795 a_8953_45002# a_2107_46812# 0.016508f
C13796 CLK VDD 0.49309f
C13797 a_n23_44458# a_n2497_47436# 4.12e-19
C13798 a_6298_44484# a_4791_45118# 0.033887f
C13799 a_21359_45002# a_18597_46090# 0.008859f
C13800 a_19778_44110# a_13507_46334# 1.08e-20
C13801 a_16759_43396# a_17124_42282# 7.27e-19
C13802 a_1847_42826# a_2903_42308# 4.53e-19
C13803 a_5755_42852# a_1755_42282# 7.33e-21
C13804 a_10796_42968# a_n784_42308# 8.64e-21
C13805 a_16137_43396# a_4958_30871# 0.008832f
C13806 a_743_42282# a_5742_30871# 0.02341f
C13807 a_5649_42852# a_9803_42558# 6.94e-20
C13808 a_19164_43230# a_19273_43230# 0.007416f
C13809 a_19339_43156# a_19518_43218# 0.007399f
C13810 a_18599_43230# a_18707_42852# 0.057222f
C13811 a_10341_43396# a_7174_31319# 4.2e-20
C13812 a_20205_31679# a_22821_38993# 5.5e-20
C13813 a_1209_47178# a_2107_46812# 2.05e-19
C13814 a_n2109_47186# a_2959_46660# 1.8e-19
C13815 a_n1741_47186# a_2609_46660# 8.05e-20
C13816 a_584_46384# a_601_46902# 0.00376f
C13817 a_1239_47204# a_948_46660# 1.6e-20
C13818 a_n1151_42308# a_n1021_46688# 0.105326f
C13819 a_1431_47204# a_1123_46634# 0.012069f
C13820 a_3381_47502# a_n1925_46634# 2.29e-21
C13821 a_n443_46116# a_n2661_46634# 0.121882f
C13822 a_3160_47472# a_n743_46660# 0.011563f
C13823 a_2905_45572# a_n2438_43548# 2.97e-21
C13824 a_n746_45260# a_1110_47026# 5.54e-20
C13825 a_15507_47210# a_12549_44172# 7.15e-20
C13826 a_11599_46634# a_768_44030# 0.018831f
C13827 a_13487_47204# a_13569_47204# 0.014524f
C13828 a_13717_47436# a_13759_47204# 0.013673f
C13829 a_12861_44030# a_13675_47204# 0.001416f
C13830 a_5111_44636# a_8415_44056# 0.003443f
C13831 a_n2661_45010# a_n2267_43396# 2.61e-20
C13832 a_3232_43370# a_5829_43940# 5.72e-19
C13833 a_18248_44752# a_18204_44850# 1.46e-19
C13834 a_18287_44626# a_17517_44484# 0.031756f
C13835 a_9482_43914# a_14021_43940# 3.32e-19
C13836 a_5891_43370# a_n2661_42834# 0.091553f
C13837 a_8375_44464# a_n2661_43922# 0.007585f
C13838 a_n3565_39590# a_n2810_45572# 0.020853f
C13839 a_22223_45572# VDD 0.287831f
C13840 a_14403_45348# a_11415_45002# 3.58e-19
C13841 a_4640_45348# a_3483_46348# 3.32e-19
C13842 a_18494_42460# a_20273_46660# 1.49e-19
C13843 a_9838_44484# a_3090_45724# 2.74e-22
C13844 a_20567_45036# a_20411_46873# 1.28e-19
C13845 a_18175_45572# a_16375_45002# 0.001125f
C13846 a_n1059_45260# a_526_44458# 0.097646f
C13847 a_n2017_45002# a_n1925_42282# 0.041988f
C13848 a_21350_45938# a_8049_45260# 1.72e-19
C13849 a_1307_43914# a_8199_44636# 0.044343f
C13850 a_1423_45028# a_5497_46414# 2.85e-22
C13851 a_13159_45002# a_10903_43370# 2.53e-19
C13852 a_13777_45326# a_9290_44172# 1.57e-20
C13853 a_7229_43940# a_2324_44458# 0.008305f
C13854 a_6171_45002# a_18189_46348# 2.69e-20
C13855 a_n3674_39768# a_n2312_39304# 0.023328f
C13856 a_n784_42308# a_4958_30871# 0.020733f
C13857 a_22400_42852# a_22775_42308# 0.003696f
C13858 a_20753_42852# a_20712_42282# 5.65e-19
C13859 a_5934_30871# a_9223_42460# 0.051891f
C13860 a_8515_42308# a_8791_42308# 0.001038f
C13861 a_5755_42308# a_5742_30871# 2.87e-20
C13862 EN_VIN_BSTR_P C4_P_btm 0.116925f
C13863 a_20916_46384# a_19692_46634# 0.117693f
C13864 a_12891_46348# a_13059_46348# 0.372745f
C13865 a_5732_46660# a_5257_43370# 0.001523f
C13866 a_5072_46660# a_5263_46660# 4.61e-19
C13867 a_12549_44172# a_15227_46910# 0.008471f
C13868 a_4646_46812# a_8492_46660# 2.79e-21
C13869 a_5807_45002# a_12347_46660# 0.001248f
C13870 a_n881_46662# a_765_45546# 0.333008f
C13871 a_21811_47423# a_20202_43084# 1.66e-20
C13872 a_21177_47436# a_12741_44636# 4.05e-21
C13873 a_4883_46098# a_11415_45002# 1.14e-19
C13874 a_13507_46334# a_20820_30879# 3.67e-19
C13875 a_n1435_47204# a_2698_46116# 2.19e-21
C13876 a_9313_45822# a_3483_46348# 0.087132f
C13877 a_6151_47436# a_6419_46155# 0.004367f
C13878 a_2063_45854# a_12005_46116# 0.051126f
C13879 a_n1151_42308# a_9290_44172# 0.10853f
C13880 a_4791_45118# a_5937_45572# 0.151145f
C13881 a_n237_47217# a_2324_44458# 1.65e-19
C13882 a_16922_45042# a_17499_43370# 4.92e-21
C13883 a_20159_44458# a_14021_43940# 7.12e-20
C13884 a_3422_30871# a_21115_43940# 1.12e-21
C13885 a_5883_43914# a_7287_43370# 2.97e-19
C13886 a_n2293_42834# a_743_42282# 2.24e-19
C13887 a_3600_43914# a_3820_44260# 0.009965f
C13888 a_n1644_44306# a_n1453_44318# 4.61e-19
C13889 a_3905_42865# a_3499_42826# 6.78e-19
C13890 a_3232_43370# a_10835_43094# 2.81e-20
C13891 a_n913_45002# a_19339_43156# 3.67e-21
C13892 a_n2017_45002# a_19987_42826# 0.142839f
C13893 en_comp a_17333_42852# 1.3e-21
C13894 a_n1059_45260# a_19164_43230# 8.48e-22
C13895 a_5205_44734# VDD 0.001314f
C13896 a_n3420_39616# VREF_GND 0.117023f
C13897 a_n4064_38528# a_n923_35174# 0.004282f
C13898 a_n4064_39072# C3_P_btm 1.38e-20
C13899 a_2711_45572# a_6472_45840# 0.049759f
C13900 a_15493_43940# a_19466_46812# 4.43e-22
C13901 a_8685_43396# a_13661_43548# 8.18e-19
C13902 a_22223_43948# a_19692_46634# 0.003538f
C13903 a_7112_43396# a_n2293_46634# 0.012325f
C13904 a_14205_43396# a_12549_44172# 9.74e-21
C13905 a_12607_44458# a_13259_45724# 0.132105f
C13906 a_n2661_44458# a_n452_45724# 5.67e-21
C13907 a_n2129_44697# a_n1079_45724# 4.42e-21
C13908 a_n2267_44484# a_n2293_45546# 3.38e-19
C13909 a_n1177_44458# a_n2661_45546# 3.02e-20
C13910 a_n2433_44484# a_n863_45724# 1.5e-21
C13911 a_484_44484# a_526_44458# 0.003617f
C13912 a_11967_42832# a_10903_43370# 0.02192f
C13913 a_15743_43084# SMPL_ON_N 4.69e-20
C13914 a_4520_42826# a_584_46384# 0.001248f
C13915 a_20447_31679# a_22521_40055# 9.79e-21
C13916 a_n4064_39072# a_n4064_38528# 0.05966f
C13917 a_22000_46634# a_20202_43084# 0.154237f
C13918 a_20841_46902# a_12741_44636# 0.043075f
C13919 a_20107_46660# a_21297_46660# 2.56e-19
C13920 a_20623_46660# a_20820_30879# 8.87e-21
C13921 a_n1613_43370# a_n443_42852# 0.062474f
C13922 a_10249_46116# a_6945_45028# 6.69e-19
C13923 a_12469_46902# a_12005_46116# 0.003112f
C13924 a_12251_46660# a_10903_43370# 5.76e-22
C13925 a_11901_46660# a_12594_46348# 1.15e-19
C13926 a_11813_46116# a_13351_46090# 7.95e-20
C13927 a_8270_45546# a_2324_44458# 0.039817f
C13928 a_n881_46662# a_509_45822# 0.001201f
C13929 a_21588_30879# a_20205_31679# 0.058932f
C13930 a_20916_46384# a_20692_30879# 0.001701f
C13931 a_n743_46660# a_16375_45002# 0.03035f
C13932 a_4817_46660# a_5066_45546# 7.24e-20
C13933 a_768_44030# a_1848_45724# 5.61e-19
C13934 a_n913_45002# a_22465_38105# 2.35e-19
C13935 a_19237_31679# a_14209_32519# 0.052426f
C13936 a_17730_32519# a_17364_32525# 0.054843f
C13937 a_n2293_42834# a_5755_42308# 7.41e-20
C13938 a_9313_44734# a_21356_42826# 0.009873f
C13939 a_10729_43914# a_10341_43396# 2.83e-20
C13940 a_13565_43940# VDD 0.175245f
C13941 a_11322_45546# a_11963_45334# 0.028732f
C13942 a_11525_45546# a_11787_45002# 5.53e-19
C13943 a_10180_45724# a_9482_43914# 0.001194f
C13944 a_11652_45724# a_10951_45334# 1.16e-21
C13945 a_8685_43396# a_4185_45028# 2.24e-20
C13946 a_15493_43940# a_20205_31679# 1.01e-20
C13947 a_17737_43940# a_n357_42282# 1.35e-20
C13948 a_8791_43396# a_5937_45572# 2.23e-21
C13949 a_9396_43370# a_8199_44636# 0.004302f
C13950 a_n2956_39304# VDD 0.455981f
C13951 a_5437_45600# a_4791_45118# 0.001854f
C13952 a_10490_45724# a_2063_45854# 0.082703f
C13953 a_9049_44484# a_n1151_42308# 1.64e-19
C13954 a_7227_45028# a_6575_47204# 9.87e-21
C13955 a_167_45260# a_310_45028# 0.035247f
C13956 a_n2293_46098# a_n443_42852# 0.086171f
C13957 a_1138_42852# a_997_45618# 0.005258f
C13958 a_1823_45246# a_n755_45592# 0.390511f
C13959 a_526_44458# a_n1925_42282# 0.213917f
C13960 a_10903_43370# a_13259_45724# 0.600111f
C13961 a_21137_46414# a_8049_45260# 0.004656f
C13962 a_18429_43548# a_18525_43370# 0.419086f
C13963 a_16409_43396# a_16664_43396# 0.056391f
C13964 a_14579_43548# a_5649_42852# 3.24e-21
C13965 a_17499_43370# a_15743_43084# 0.049383f
C13966 a_10341_43396# a_21487_43396# 0.010314f
C13967 a_n97_42460# a_16414_43172# 0.044625f
C13968 a_20974_43370# a_21356_42826# 8.97e-20
C13969 a_3626_43646# a_7871_42858# 3.84e-20
C13970 a_2982_43646# a_8037_42858# 5.75e-20
C13971 a_21381_43940# a_21671_42860# 0.001657f
C13972 a_n2661_42282# a_n1736_42282# 3.68e-19
C13973 a_11967_42832# a_15959_42545# 6.6e-19
C13974 a_15095_43370# a_4361_42308# 1.65e-19
C13975 a_n2661_46634# DATA[4] 7.86e-20
C13976 a_n743_46660# RST_Z 1.57e-20
C13977 a_n2312_38680# CLK_DATA 1.56e-20
C13978 a_5534_30871# VDD 0.513761f
C13979 a_n2810_45028# a_n4209_37414# 0.09606f
C13980 a_6171_45002# a_18315_45260# 5.25e-20
C13981 a_n2017_45002# a_n4318_40392# 2.16e-20
C13982 a_n2661_45010# a_n2267_44484# 0.260289f
C13983 a_n2109_45247# a_n2661_44458# 0.001495f
C13984 a_n2293_45010# a_n2433_44484# 0.016908f
C13985 a_18909_45814# a_18989_43940# 4.16e-19
C13986 a_13017_45260# a_14976_45348# 5.79e-21
C13987 a_626_44172# a_n2293_42834# 2.37e-20
C13988 a_18691_45572# a_18374_44850# 2.44e-20
C13989 a_13887_32519# a_n357_42282# 3.9e-20
C13990 a_2711_45572# a_14513_46634# 3.9e-21
C13991 a_11322_45546# a_11901_46660# 8.73e-20
C13992 a_11525_45546# a_11813_46116# 6.46e-19
C13993 a_3357_43084# a_20916_46384# 7.98e-19
C13994 a_19479_31679# a_21588_30879# 0.055797f
C13995 a_2382_45260# a_n881_46662# 6.99e-22
C13996 a_413_45260# a_8128_46384# 4.76e-20
C13997 a_9482_43914# a_13507_46334# 2.01e-19
C13998 a_13159_45002# a_4883_46098# 2.87e-21
C13999 a_8953_45002# a_11453_44696# 6.78e-19
C14000 a_3080_42308# a_4958_30871# 0.01856f
C14001 a_19164_43230# a_19987_42826# 3.85e-19
C14002 a_n97_42460# a_7174_31319# 6.58e-20
C14003 a_7765_42852# a_7309_42852# 0.00456f
C14004 a_3626_43646# a_11897_42308# 3.42e-19
C14005 a_19647_42308# VDD 0.227331f
C14006 a_n2109_47186# a_2266_47243# 0.001164f
C14007 a_n971_45724# a_2266_47570# 4.39e-19
C14008 a_n1741_47186# a_3094_47570# 2.25e-19
C14009 a_4915_47217# a_10227_46804# 0.062269f
C14010 a_13381_47204# a_13717_47436# 4.77e-21
C14011 a_n746_45260# a_n89_47570# 0.004982f
C14012 a_n237_47217# a_n310_47570# 6.1e-19
C14013 a_n785_47204# a_n2312_40392# 2.56e-20
C14014 a_16112_44458# a_17970_44736# 6.26e-20
C14015 a_626_44172# a_1115_44172# 0.00354f
C14016 a_1307_43914# a_2127_44172# 0.127867f
C14017 a_4223_44672# a_5289_44734# 0.009506f
C14018 a_11691_44458# a_14112_44734# 0.005155f
C14019 a_14539_43914# a_17767_44458# 3.19e-19
C14020 a_375_42282# a_1414_42308# 6.78e-21
C14021 a_7499_43078# a_6765_43638# 3.15e-19
C14022 a_n1059_45260# a_18079_43940# 5.09e-19
C14023 a_5934_30871# a_n755_45592# 0.040823f
C14024 a_8515_42308# a_n357_42282# 2.87e-20
C14025 a_n2302_39866# a_n2956_38680# 2.07e-19
C14026 a_15959_42545# a_13259_45724# 1.16e-19
C14027 a_n2661_43370# a_3090_45724# 0.101361f
C14028 a_3232_43370# a_11415_45002# 4.11e-19
C14029 a_10617_44484# a_768_44030# 0.001771f
C14030 a_10907_45822# a_8049_45260# 0.010337f
C14031 a_2711_45572# a_n357_42282# 0.039058f
C14032 a_1260_45572# a_997_45618# 0.010598f
C14033 a_8192_45572# a_8034_45724# 0.002594f
C14034 a_1609_45572# a_n755_45592# 5.85e-19
C14035 a_15433_44458# a_n881_46662# 3.48e-21
C14036 a_18175_45572# a_18985_46122# 0.009338f
C14037 a_18479_45785# a_18819_46122# 2.67e-20
C14038 a_18341_45572# a_17957_46116# 1.43e-19
C14039 a_2437_43646# a_8016_46348# 3.18e-20
C14040 a_3357_43084# a_6165_46155# 0.009006f
C14041 a_n1441_43940# a_n971_45724# 7.56e-19
C14042 a_2127_44172# a_n443_46116# 0.196411f
C14043 a_19279_43940# a_18597_46090# 0.021978f
C14044 a_21398_44850# a_16327_47482# 2.55e-19
C14045 a_11967_42832# a_4883_46098# 5.15e-22
C14046 a_1576_42282# a_1606_42308# 0.176925f
C14047 a_1067_42314# a_1755_42282# 8.86e-19
C14048 a_961_42354# a_1149_42558# 7.47e-21
C14049 a_n3674_37592# a_n327_42308# 0.002227f
C14050 a_1184_42692# a_1221_42558# 3.52e-19
C14051 a_n443_46116# a_765_45546# 0.297346f
C14052 a_10227_46804# a_18834_46812# 2.09e-20
C14053 a_18143_47464# a_17609_46634# 0.001435f
C14054 a_4883_46098# a_12251_46660# 1.41e-19
C14055 a_9804_47204# a_8492_46660# 8.56e-22
C14056 a_171_46873# a_1799_45572# 2.16e-21
C14057 a_601_46902# a_479_46660# 3.16e-19
C14058 a_n133_46660# a_n2661_46098# 0.005588f
C14059 a_n2438_43548# a_2443_46660# 0.237765f
C14060 a_n743_46660# a_2609_46660# 6.69e-20
C14061 a_n1925_46634# a_2959_46660# 0.009513f
C14062 a_5807_45002# a_5732_46660# 9.62e-19
C14063 en_comp a_13678_32519# 1.37e-19
C14064 a_2711_45572# a_18707_42852# 2.52e-19
C14065 a_n2293_43922# a_10729_43914# 1.27e-20
C14066 a_5883_43914# a_9420_43940# 0.001123f
C14067 a_17730_32519# a_19237_31679# 0.058836f
C14068 a_14537_43396# a_15681_43442# 2.41e-19
C14069 a_n2661_42834# a_10807_43548# 0.003836f
C14070 a_n2661_43922# a_10949_43914# 9.62e-19
C14071 a_7754_38968# VDD 0.041093f
C14072 a_11691_44458# VDD 3.25709f
C14073 a_15486_42560# RST_Z 5.88e-19
C14074 a_5742_30871# VIN_P 0.042613f
C14075 a_n2661_43922# a_376_46348# 2.93e-22
C14076 a_14581_44484# a_11415_45002# 0.009374f
C14077 a_5608_44484# a_1823_45246# 3.64e-19
C14078 a_2998_44172# a_3090_45724# 0.001518f
C14079 a_18681_44484# a_17339_46660# 5.66e-19
C14080 a_21205_44306# a_13747_46662# 5.28e-19
C14081 a_21359_45002# a_8049_45260# 2.51e-22
C14082 a_14403_45348# a_13259_45724# 0.001862f
C14083 a_117_45144# a_n2293_45546# 6.33e-19
C14084 a_6298_44484# a_6945_45028# 0.00332f
C14085 a_15004_44636# a_2324_44458# 2.94e-20
C14086 a_n229_43646# a_n1613_43370# 3.21e-19
C14087 a_4842_47243# VDD 6.34e-20
C14088 a_n784_42308# C7_N_btm 0.002308f
C14089 a_1606_42308# C1_P_btm 0.096405f
C14090 a_5534_30871# a_8912_37509# 3.98e-19
C14091 a_17609_46634# a_765_45546# 0.256159f
C14092 a_16292_46812# a_17829_46910# 1.46e-19
C14093 a_4955_46873# a_5164_46348# 0.009022f
C14094 a_3877_44458# a_6165_46155# 1.87e-19
C14095 a_4646_46812# a_5497_46414# 2.5e-20
C14096 a_4651_46660# a_5204_45822# 2.21e-19
C14097 a_4817_46660# a_5068_46348# 0.001467f
C14098 a_4883_46098# a_13259_45724# 0.011246f
C14099 a_13507_46334# a_18243_46436# 6.14e-19
C14100 a_18597_46090# a_19597_46482# 0.002198f
C14101 a_10227_46804# a_20850_46482# 6.4e-19
C14102 a_16327_47482# a_20850_46155# 2.49e-19
C14103 a_4791_45118# a_n443_42852# 0.02747f
C14104 a_n443_46116# a_509_45822# 0.006202f
C14105 a_10057_43914# a_10796_42968# 1.53e-19
C14106 a_19862_44208# a_19741_43940# 0.038152f
C14107 a_n2661_42282# a_1209_43370# 2.03e-21
C14108 a_11967_42832# a_16243_43396# 0.269605f
C14109 a_17517_44484# a_19268_43646# 3.12e-21
C14110 a_10555_44260# a_10651_43940# 0.001863f
C14111 a_15493_43940# a_15037_43940# 0.004121f
C14112 a_3905_42865# a_6197_43396# 1.51e-20
C14113 a_10729_43914# a_n97_42460# 2.13e-20
C14114 a_3537_45260# a_5379_42460# 6.86e-20
C14115 en_comp a_6123_31319# 0.028738f
C14116 a_3065_45002# a_3581_42558# 0.003532f
C14117 a_n2017_45002# a_8337_42558# 4.83e-19
C14118 a_8333_44056# VDD 0.124235f
C14119 a_15037_45618# a_15765_45572# 3.63e-20
C14120 a_5649_42852# a_5257_43370# 8.9e-19
C14121 a_15681_43442# a_3090_45724# 3.44e-19
C14122 a_17333_42852# a_13661_43548# 1.34e-20
C14123 a_12545_42858# a_n2293_46634# 3.58e-20
C14124 a_16823_43084# a_6755_46942# 1.01e-19
C14125 a_n2065_43946# a_n2293_45546# 2.73e-20
C14126 a_564_42282# a_584_46384# 7.22e-21
C14127 a_n961_42308# a_n1151_42308# 0.109068f
C14128 a_13291_42460# a_10227_46804# 0.002348f
C14129 a_n1991_46122# VDD 0.581018f
C14130 C0_dummy_P_btm C0_dummy_N_btm 0.033338f
C14131 C1_P_btm C1_N_btm 0.065833f
C14132 C0_P_btm C0_N_btm 0.044249f
C14133 a_n4064_40160# a_n4334_37440# 0.007725f
C14134 a_n4315_30879# a_n3690_37440# 1.35e-19
C14135 a_n4209_38502# a_n2946_37984# 5.32e-20
C14136 a_n3565_38502# a_n3690_38304# 7.97e-20
C14137 a_1736_39043# a_2113_38308# 0.088667f
C14138 a_13258_32519# VDAC_N 4.18e-19
C14139 a_13759_46122# a_2324_44458# 8.3e-20
C14140 a_13925_46122# a_14840_46494# 0.118759f
C14141 a_5937_45572# a_6945_45028# 0.22046f
C14142 a_2698_46116# a_526_44458# 0.002083f
C14143 a_2804_46116# a_2981_46116# 0.134298f
C14144 a_1138_42852# a_1337_46116# 0.039951f
C14145 a_21177_47436# RST_Z 5.48e-20
C14146 a_20894_47436# SINGLE_ENDED 0.044283f
C14147 a_20990_47178# START 4.18e-19
C14148 a_3422_30871# a_20256_42852# 1.38e-20
C14149 a_17538_32519# a_17364_32525# 9.64512f
C14150 a_5891_43370# a_9885_42558# 0.001022f
C14151 a_n2293_43922# a_5932_42308# 0.178011f
C14152 a_20512_43084# a_20256_43172# 0.047194f
C14153 a_11341_43940# a_15567_42826# 3.04e-20
C14154 a_20974_43370# a_20749_43396# 0.0837f
C14155 a_3626_43646# a_17324_43396# 4.75e-21
C14156 a_8685_43396# a_14579_43548# 0.03481f
C14157 a_10227_46804# DATA[5] 2.13e-20
C14158 a_4190_30871# VDD 1.36846f
C14159 a_13904_45546# a_13720_44458# 2.89e-21
C14160 a_18341_45572# a_18587_45118# 8.86e-19
C14161 a_18479_45785# a_18911_45144# 0.00112f
C14162 a_13249_42308# a_13076_44458# 1.5e-19
C14163 a_1667_45002# a_375_42282# 2.16e-20
C14164 a_6171_45002# a_13017_45260# 0.045098f
C14165 a_413_45260# a_626_44172# 0.032584f
C14166 a_2382_45260# a_1307_43914# 0.53878f
C14167 a_7705_45326# a_8191_45002# 5.55e-19
C14168 a_17333_42852# a_4185_45028# 1.67e-20
C14169 a_13258_32519# a_21588_30879# 0.062822f
C14170 a_8791_43396# a_n443_42852# 0.053902f
C14171 a_16243_43396# a_13259_45724# 1.45e-20
C14172 a_n3674_39304# a_n2956_38680# 0.023431f
C14173 a_n4318_38680# a_n2956_39304# 0.023405f
C14174 a_5755_42852# a_2324_44458# 3.34e-19
C14175 a_10518_42984# a_10903_43370# 8.08e-19
C14176 a_10922_42852# a_9290_44172# 0.028552f
C14177 a_6472_45840# a_6540_46812# 3.24e-21
C14178 a_8696_44636# a_12891_46348# 0.028033f
C14179 a_8336_45822# a_n1925_46634# 0.003059f
C14180 a_11682_45822# a_n2661_46634# 0.010865f
C14181 a_20273_45572# a_4883_46098# 9.32e-20
C14182 a_2382_45260# a_n443_46116# 0.027844f
C14183 a_5147_45002# a_n1151_42308# 4.06e-20
C14184 a_6171_45002# a_2063_45854# 0.029207f
C14185 a_413_45260# a_6151_47436# 3.16e-19
C14186 a_19610_45572# a_18597_46090# 4.96e-19
C14187 a_22591_45572# a_16327_47482# 1.29e-19
C14188 a_2437_43646# a_17591_47464# 0.013209f
C14189 a_3357_43084# a_16023_47582# 2.06e-19
C14190 a_20623_45572# a_13507_46334# 1.7e-20
C14191 a_n2661_45546# a_2957_45546# 0.008098f
C14192 a_n863_45724# a_310_45028# 0.033427f
C14193 a_n2293_45546# a_n755_45592# 0.061822f
C14194 a_n452_45724# a_n1099_45572# 0.053931f
C14195 a_7871_42858# a_8037_42858# 0.772842f
C14196 a_5649_42852# a_21671_42860# 0.003655f
C14197 a_n97_42460# a_5932_42308# 2.52e-19
C14198 a_13678_32519# a_22165_42308# 0.018986f
C14199 a_14579_43548# a_15953_42852# 1.82e-19
C14200 a_1987_43646# a_1606_42308# 3.6e-36
C14201 a_14021_43940# a_4958_30871# 2.74e-20
C14202 a_765_45546# DATA[4] 0.006502f
C14203 a_20841_46902# RST_Z 1.47e-20
C14204 a_7754_38968# a_8912_37509# 6.06e-19
C14205 a_7754_38636# a_5088_37509# 0.288061f
C14206 VDAC_Ni a_4338_37500# 0.640521f
C14207 a_n4209_37414# a_n2302_37690# 0.407594f
C14208 a_n3565_37414# a_n2946_37690# 0.407439f
C14209 a_n3690_37440# a_n3420_37440# 0.431074f
C14210 a_n4334_37440# a_n4064_37440# 0.448688f
C14211 a_5337_42558# VDD 0.008564f
C14212 a_n785_47204# a_327_47204# 0.237391f
C14213 a_n971_45724# a_2124_47436# 0.352461f
C14214 a_n237_47217# a_1239_47204# 0.203126f
C14215 a_n1741_47186# a_2905_45572# 0.012244f
C14216 a_n2109_47186# a_n1151_42308# 0.235661f
C14217 a_n746_45260# a_1431_47204# 2.26e-19
C14218 a_n2293_45010# a_n2840_43914# 4.9e-20
C14219 a_2437_43646# a_1414_42308# 0.023872f
C14220 a_n2661_45010# a_n2065_43946# 0.001138f
C14221 a_n2472_45002# a_n2472_43914# 0.001034f
C14222 a_8696_44636# a_11750_44172# 3.79e-20
C14223 a_1307_43914# a_15433_44458# 2.11e-20
C14224 a_n2661_43370# a_n356_44636# 0.002184f
C14225 a_n2840_44458# a_n4318_40392# 0.161548f
C14226 a_10907_45822# a_11173_44260# 7.74e-20
C14227 a_16333_45814# a_15682_43940# 2.17e-19
C14228 a_16877_42852# a_n357_42282# 0.016936f
C14229 a_4169_42308# a_n1925_42282# 2.9e-19
C14230 a_5742_30871# a_n2956_38680# 4.45e-21
C14231 a_20273_45572# a_21188_46660# 3.8e-20
C14232 a_14033_45822# a_3483_46348# 0.030627f
C14233 a_18341_45572# a_11415_45002# 0.002269f
C14234 a_16147_45260# a_12741_44636# 0.023061f
C14235 a_5093_45028# a_4817_46660# 5.47e-21
C14236 a_15415_45028# a_6755_46942# 5.84e-21
C14237 a_7418_45394# a_4646_46812# 0.001071f
C14238 a_4099_45572# a_n1925_42282# 0.009682f
C14239 a_5263_45724# a_526_44458# 5.01e-19
C14240 a_21188_45572# a_20273_46660# 6.41e-21
C14241 a_20623_45572# a_20623_46660# 2.72e-19
C14242 a_20528_45572# a_20411_46873# 3.25e-21
C14243 a_413_45260# a_19466_46812# 2.56e-20
C14244 a_4574_45260# a_3090_45724# 0.002261f
C14245 a_5343_44458# a_n881_46662# 6.79e-19
C14246 a_11652_45724# a_2324_44458# 0.034041f
C14247 a_11823_42460# a_14275_46494# 1.34e-19
C14248 a_10210_45822# a_9625_46129# 0.002126f
C14249 a_13249_42308# a_12594_46348# 4.26e-20
C14250 a_17767_44458# a_11453_44696# 0.010225f
C14251 a_14815_43914# a_4915_47217# 0.006248f
C14252 a_9313_44734# a_12861_44030# 0.001011f
C14253 a_17364_32525# a_22465_38105# 2.07e-19
C14254 a_12089_42308# a_13333_42558# 2.22e-19
C14255 a_5534_30871# a_11551_42558# 5.08e-19
C14256 a_3080_42308# C7_N_btm 0.002948f
C14257 a_12549_44172# a_13747_46662# 0.072812f
C14258 a_768_44030# a_13661_43548# 0.175469f
C14259 a_15928_47570# a_5807_45002# 1.22e-19
C14260 a_n1613_43370# a_n2661_46634# 0.279652f
C14261 a_6151_47436# a_9863_46634# 0.0481f
C14262 a_6575_47204# a_7715_46873# 4.64e-19
C14263 a_7903_47542# a_7577_46660# 4e-20
C14264 a_4915_47217# a_10467_46802# 0.003258f
C14265 a_n2497_47436# a_3090_45724# 0.16041f
C14266 a_18911_45144# a_14021_43940# 1.04e-20
C14267 a_7499_43078# a_10341_42308# 0.42152f
C14268 a_4223_44672# a_9028_43914# 5.03e-20
C14269 a_20193_45348# a_15493_43940# 0.10893f
C14270 a_10193_42453# a_10835_43094# 0.041273f
C14271 a_5343_44458# a_7911_44260# 0.005844f
C14272 a_5883_43914# a_5841_44260# 2.9e-21
C14273 a_5111_44636# a_6293_42852# 0.072755f
C14274 a_3537_45260# a_7287_43370# 0.400907f
C14275 a_5147_45002# a_6197_43396# 9.61e-19
C14276 a_413_45260# a_2813_43396# 6.05e-21
C14277 a_375_42282# VDD 0.591443f
C14278 a_n784_42308# C3_P_btm 0.001962f
C14279 a_n2661_44458# a_167_45260# 4.36e-19
C14280 a_8975_43940# a_11415_45002# 6.59e-20
C14281 a_13483_43940# a_13661_43548# 0.057042f
C14282 a_20269_44172# a_12549_44172# 0.049822f
C14283 a_n2661_42282# a_n2442_46660# 7.91e-20
C14284 a_15415_45028# a_8049_45260# 2.92e-20
C14285 a_9482_43914# a_10586_45546# 1.67e-20
C14286 a_n2661_45010# a_n755_45592# 0.01648f
C14287 a_n1059_45260# a_n452_45724# 2.74e-19
C14288 a_n913_45002# a_n863_45724# 0.565852f
C14289 a_413_45260# a_20205_31679# 0.034773f
C14290 a_n2956_37592# a_n2956_38216# 0.103811f
C14291 a_n2810_45028# a_n2293_45546# 8.06e-21
C14292 a_n2293_45010# a_310_45028# 2.43e-21
C14293 en_comp a_n2472_45546# 5.76e-19
C14294 a_n967_45348# a_n2661_45546# 0.001666f
C14295 a_n998_43396# a_n971_45724# 1.52e-19
C14296 a_n1557_42282# a_584_46384# 0.032459f
C14297 a_20974_43370# a_12861_44030# 1.38e-19
C14298 a_18797_44260# a_16327_47482# 1.19e-19
C14299 a_15764_42576# a_4958_30871# 0.413236f
C14300 a_15486_42560# a_17303_42282# 3.91e-21
C14301 a_10533_42308# a_7174_31319# 4.88e-21
C14302 a_1606_42308# a_1736_39043# 7.77e-20
C14303 a_n3674_38216# a_n4209_38216# 0.059407f
C14304 a_n1630_35242# a_n3565_38502# 1.85e-19
C14305 a_5742_30871# a_13258_32519# 0.004591f
C14306 a_15890_42674# a_15761_42308# 4.2e-19
C14307 a_15959_42545# a_16197_42308# 0.001705f
C14308 a_15803_42450# a_16269_42308# 3.82e-19
C14309 a_14113_42308# a_18057_42282# 2.13e-20
C14310 a_n3674_37592# a_n3420_38528# 0.020112f
C14311 a_n784_42308# a_n4064_38528# 0.004411f
C14312 a_n4318_38216# a_n3565_38216# 3.9e-19
C14313 a_5129_47502# VDD 0.20906f
C14314 a_18597_46090# a_20708_46348# 0.003878f
C14315 a_10227_46804# a_10809_44734# 0.17883f
C14316 a_18479_47436# a_6945_45028# 0.348097f
C14317 a_4791_45118# a_6633_46155# 0.006879f
C14318 a_12465_44636# a_17583_46090# 1.75e-21
C14319 a_4915_47217# a_8034_45724# 7.21e-21
C14320 a_n1435_47204# a_526_44458# 4.56e-21
C14321 a_4883_46098# a_18189_46348# 0.012818f
C14322 a_13507_46334# a_18819_46122# 0.004962f
C14323 a_n1613_43370# a_8199_44636# 5.93e-20
C14324 a_n881_46662# a_8349_46414# 7.22e-20
C14325 a_6755_46942# a_15368_46634# 0.033754f
C14326 a_768_44030# a_4185_45028# 0.022613f
C14327 a_n2661_46634# a_n2293_46098# 2.67e-19
C14328 a_n2472_46634# a_n2472_46090# 0.026152f
C14329 a_20447_31679# a_14097_32519# 0.05131f
C14330 a_n1059_45260# a_17749_42852# 8.24e-19
C14331 a_11823_42460# a_13657_42308# 4.58e-19
C14332 a_10405_44172# a_11341_43940# 0.001372f
C14333 a_5663_43940# a_5745_43940# 0.096132f
C14334 a_19721_31679# a_17364_32525# 0.053872f
C14335 a_19237_31679# a_17538_32519# 0.060188f
C14336 a_9313_44734# a_9803_43646# 2.3e-19
C14337 a_17973_43940# a_18451_43940# 0.0015f
C14338 a_15682_43940# a_15493_43396# 9.79e-19
C14339 a_5495_43940# a_5829_43940# 0.001349f
C14340 a_18079_43940# a_18326_43940# 0.152347f
C14341 a_17970_44736# a_17499_43370# 9.31e-19
C14342 a_2711_45572# a_15765_45572# 0.005291f
C14343 a_11962_45724# a_13163_45724# 0.113317f
C14344 a_12427_45724# a_12791_45546# 0.124682f
C14345 a_8568_45546# a_8697_45822# 0.062574f
C14346 C1_P_btm C9_P_btm 0.132506f
C14347 C0_P_btm C10_P_btm 0.365593f
C14348 C2_N_btm EN_VIN_BSTR_N 0.118072f
C14349 a_15682_43940# a_3483_46348# 0.261013f
C14350 a_19279_43940# a_8049_45260# 2.89e-20
C14351 a_556_44484# a_n863_45724# 0.002594f
C14352 a_6756_44260# a_5937_45572# 0.010335f
C14353 a_n1379_43218# a_n1613_43370# 0.001903f
C14354 a_13460_43230# a_10227_46804# 0.243111f
C14355 a_18599_43230# a_12861_44030# 7.75e-20
C14356 a_8495_42852# a_n971_45724# 1.66e-19
C14357 a_15227_44166# VDD 2.69945f
C14358 a_1823_45246# a_3483_46348# 0.070929f
C14359 a_167_45260# a_2804_46116# 0.003847f
C14360 a_2521_46116# a_2698_46116# 0.159555f
C14361 a_15368_46634# a_8049_45260# 0.032468f
C14362 a_11813_46116# a_12005_46436# 6.29e-19
C14363 a_11415_45002# a_11387_46155# 3.86e-20
C14364 a_12741_44636# a_9290_44172# 0.004434f
C14365 a_20107_46660# a_20075_46420# 0.001101f
C14366 a_17339_46660# a_10809_44734# 0.003677f
C14367 a_9313_44734# a_19518_43218# 1.42e-19
C14368 a_20512_43084# a_21195_42852# 2.47e-19
C14369 a_11341_43940# a_20556_43646# 0.004978f
C14370 a_n2497_47436# CLK_DATA 0.026654f
C14371 a_6655_43762# VDD 0.132357f
C14372 a_n2661_45010# a_n2810_45028# 0.009249f
C14373 a_n2840_45002# a_n2956_37592# 0.035532f
C14374 a_n2293_45010# a_n913_45002# 0.015951f
C14375 a_19479_31679# a_413_45260# 0.055869f
C14376 a_n2109_45247# a_n1059_45260# 1.05e-19
C14377 a_2437_43646# a_1667_45002# 0.005688f
C14378 a_10193_42453# a_18587_45118# 7.6e-21
C14379 a_13678_32519# a_4185_45028# 0.037732f
C14380 a_n4064_38528# SMPL_ON_P 9.15e-21
C14381 a_20712_42282# a_16327_47482# 0.030215f
C14382 a_4958_30871# a_13507_46334# 6.72e-21
C14383 a_4880_45572# a_n881_46662# 2.99e-19
C14384 a_13249_42308# a_12465_44636# 0.541909f
C14385 a_15143_45578# a_4883_46098# 5.67e-21
C14386 a_15037_45618# a_12861_44030# 1.43e-20
C14387 a_14033_45822# a_13487_47204# 1.36e-20
C14388 a_12638_46436# a_12839_46116# 0.005425f
C14389 a_526_44458# a_380_45546# 8.89e-21
C14390 a_n97_42460# a_17141_43172# 3.1e-19
C14391 a_19237_31679# a_22465_38105# 2.6e-19
C14392 a_22591_43396# a_17364_32525# 7.75e-19
C14393 a_3539_42460# a_4649_42852# 0.006668f
C14394 a_21381_43940# a_20256_43172# 6.27e-20
C14395 a_10341_43396# a_15567_42826# 0.004039f
C14396 a_14209_32519# a_22959_43396# 0.015679f
C14397 a_10729_43914# a_10533_42308# 2.31e-20
C14398 a_10150_46912# CLK 0.004688f
C14399 a_10467_46802# DATA[5] 1.05e-19
C14400 a_n4064_37984# a_n4251_38304# 4.37e-19
C14401 a_14635_42282# VDD 0.369964f
C14402 a_18341_45572# a_11967_42832# 6.68e-21
C14403 a_1307_43914# a_5343_44458# 0.02568f
C14404 a_9482_43914# a_10440_44484# 0.001083f
C14405 a_18479_45785# a_19615_44636# 0.006445f
C14406 a_2711_45572# a_19328_44172# 0.010017f
C14407 a_375_42282# a_n699_43396# 0.127058f
C14408 a_1423_45028# a_742_44458# 0.019572f
C14409 a_n913_45002# a_9313_44734# 0.055701f
C14410 a_6123_31319# a_4185_45028# 0.068372f
C14411 a_18548_42308# a_17339_46660# 1.37e-19
C14412 a_18817_42826# a_n357_42282# 0.008235f
C14413 a_n2840_42282# a_n2956_39304# 2.99e-20
C14414 a_12895_43230# a_n443_42852# 1.14e-19
C14415 a_3080_42308# C3_P_btm 0.027071f
C14416 a_10193_42453# a_11415_45002# 0.024787f
C14417 a_2711_45572# a_3147_46376# 7.31e-20
C14418 a_6428_45938# a_n2293_46098# 5.88e-21
C14419 a_9482_43914# a_n743_46660# 7.74e-21
C14420 a_16211_45572# a_3090_45724# 7.88e-19
C14421 a_2437_43646# a_10428_46928# 3.53e-20
C14422 a_3537_45260# a_3524_46660# 1.28e-20
C14423 a_413_45260# a_3221_46660# 9.19e-19
C14424 EN_OFFSET_CAL VDD 0.489629f
C14425 a_5518_44484# a_4791_45118# 2.27e-19
C14426 a_n356_44636# a_n2497_47436# 0.019387f
C14427 a_11827_44484# a_18479_47436# 0.035345f
C14428 a_21101_45002# a_18597_46090# 0.033595f
C14429 a_18911_45144# a_13507_46334# 1.16e-20
C14430 a_18315_45260# a_4883_46098# 1.48e-20
C14431 a_4361_42308# a_9377_42558# 8.36e-20
C14432 a_1847_42826# a_2713_42308# 0.015903f
C14433 a_5111_42852# a_1755_42282# 2.49e-20
C14434 a_10835_43094# a_n784_42308# 1.43e-21
C14435 a_18817_42826# a_18707_42852# 0.097745f
C14436 a_5649_42852# a_9223_42460# 6.66e-20
C14437 a_743_42282# a_11323_42473# 0.008466f
C14438 a_16977_43638# a_17124_42282# 4.32e-20
C14439 a_10341_43396# a_20712_42282# 2.59e-20
C14440 a_3080_42308# a_n4064_38528# 0.001913f
C14441 a_20692_30879# a_22521_39511# 5.01e-20
C14442 a_10227_46804# a_n881_46662# 0.146883f
C14443 SMPL_ON_P a_n2661_46098# 0.004205f
C14444 a_n2109_47186# a_3177_46902# 1.13e-19
C14445 a_n1741_47186# a_2443_46660# 1.18e-19
C14446 a_584_46384# a_33_46660# 8.87e-19
C14447 a_1209_47178# a_948_46660# 0.002172f
C14448 a_1239_47204# a_1123_46634# 2.42e-19
C14449 a_n1151_42308# a_n1925_46634# 0.105874f
C14450 a_2905_45572# a_n743_46660# 0.03492f
C14451 a_4791_45118# a_n2661_46634# 0.026643f
C14452 a_11599_46634# a_12549_44172# 0.075725f
C14453 a_14955_47212# a_768_44030# 1.84e-19
C14454 a_13717_47436# a_13675_47204# 0.006407f
C14455 a_12861_44030# a_13569_47204# 6.43e-19
C14456 a_n1435_47204# a_13759_47204# 5.48e-19
C14457 a_n913_45002# a_20974_43370# 2.82e-20
C14458 a_3232_43370# a_5745_43940# 1.59e-19
C14459 a_n2661_45010# a_n2129_43609# 1.46e-20
C14460 a_17970_44736# a_18204_44850# 0.006453f
C14461 a_16112_44458# a_16335_44484# 0.011458f
C14462 a_19721_31679# a_19237_31679# 0.071506f
C14463 a_7640_43914# a_n2661_43922# 0.019048f
C14464 a_18248_44752# a_17517_44484# 0.561898f
C14465 a_8975_43940# a_11967_42832# 1.12e-20
C14466 a_8375_44464# a_n2661_42834# 3.77e-20
C14467 a_2437_43646# VDD 1.17411f
C14468 a_20567_45036# a_20107_46660# 5.96e-22
C14469 a_5883_43914# a_3090_45724# 0.132458f
C14470 a_n2293_43922# a_4646_46812# 8.64e-21
C14471 a_n1761_44111# a_768_44030# 2.61e-20
C14472 a_18341_45572# a_13259_45724# 1.51e-19
C14473 a_16147_45260# a_16375_45002# 1.01554f
C14474 a_n2017_45002# a_526_44458# 0.028467f
C14475 a_13017_45260# a_10903_43370# 2.86e-19
C14476 a_1423_45028# a_5204_45822# 3.01e-21
C14477 a_11963_45334# a_12005_46116# 1.6e-19
C14478 a_13556_45296# a_9290_44172# 2.5e-20
C14479 a_7276_45260# a_2324_44458# 0.049304f
C14480 a_6171_45002# a_17715_44484# 5.11e-20
C14481 a_n3674_39768# a_n2312_40392# 0.025146f
C14482 a_n4318_39768# a_n2312_39304# 0.02345f
C14483 a_22400_42852# a_21613_42308# 0.024416f
C14484 a_5934_30871# a_8791_42308# 0.223675f
C14485 a_8515_42308# a_8685_42308# 0.108744f
C14486 a_19864_35138# a_21589_35634# 0.150796f
C14487 EN_VIN_BSTR_P C5_P_btm 0.115337f
C14488 a_n743_46660# a_12816_46660# 4.05e-20
C14489 a_5907_46634# a_5257_43370# 0.070316f
C14490 a_4646_46812# a_8667_46634# 3.58e-21
C14491 a_3877_44458# a_8492_46660# 1.48e-21
C14492 a_12549_44172# a_13693_46688# 1.21e-19
C14493 a_768_44030# a_14543_46987# 3.15e-19
C14494 a_n881_46662# a_17339_46660# 7.38e-21
C14495 a_n1613_43370# a_765_45546# 0.205521f
C14496 a_13507_46334# a_22591_46660# 1.58e-19
C14497 a_4883_46098# a_20202_43084# 0.135688f
C14498 a_20990_47178# a_12741_44636# 5.68e-20
C14499 a_n1435_47204# a_2521_46116# 3.94e-21
C14500 a_4915_47217# a_8016_46348# 2.37e-20
C14501 a_6151_47436# a_6165_46155# 0.00218f
C14502 a_n1151_42308# a_10355_46116# 0.043227f
C14503 a_4791_45118# a_8199_44636# 0.14611f
C14504 a_2063_45854# a_10903_43370# 0.277624f
C14505 a_2779_44458# a_2813_43396# 3.22e-21
C14506 a_19615_44636# a_14021_43940# 4.32e-21
C14507 a_3600_43914# a_3499_42826# 0.125876f
C14508 a_5883_43914# a_6547_43396# 2.84e-19
C14509 a_n356_44636# a_1568_43370# 7.66e-20
C14510 a_2998_44172# a_3820_44260# 1.27e-20
C14511 a_n913_45002# a_18599_43230# 1.4e-20
C14512 en_comp a_18083_42858# 1.15e-20
C14513 a_n2017_45002# a_19164_43230# 0.048221f
C14514 a_3357_43084# a_4156_43218# 2.37e-19
C14515 a_4181_44734# VDD 0.004392f
C14516 a_n3565_39590# VCM 0.097317f
C14517 a_n4064_39616# VIN_P 0.048523f
C14518 a_n3420_38528# EN_VIN_BSTR_P 0.031973f
C14519 a_n4064_39072# C4_P_btm 1.7e-20
C14520 a_n2860_37690# a_n2956_38216# 8.73e-19
C14521 a_2711_45572# a_6194_45824# 0.013872f
C14522 a_11341_43940# a_19692_46634# 0.06f
C14523 a_8685_43396# a_5807_45002# 9.36e-20
C14524 a_n97_42460# a_4646_46812# 0.016161f
C14525 a_7287_43370# a_n2293_46634# 0.016986f
C14526 a_n2661_44458# a_n863_45724# 0.091002f
C14527 a_n2129_44697# a_n2293_45546# 3.68e-19
C14528 a_11827_44484# a_n443_42852# 1.48e-19
C14529 a_n89_44484# a_526_44458# 1.64e-20
C14530 a_17061_44734# a_15682_46116# 1.05e-20
C14531 a_3935_42891# a_584_46384# 4.23e-20
C14532 a_685_42968# a_n1151_42308# 9.34e-22
C14533 a_20556_43646# a_16327_47482# 0.014087f
C14534 a_19963_31679# a_22459_39145# 2.14e-20
C14535 a_n2946_39072# a_n4064_38528# 3.78e-20
C14536 a_n4064_39072# a_n2946_38778# 3.78e-20
C14537 a_n3565_39304# a_n2216_38778# 1e-19
C14538 a_3686_47026# VDD 4.6e-19
C14539 a_1606_42308# a_n3420_37984# 6.06e-20
C14540 a_n784_42308# a_7754_40130# 0.001644f
C14541 a_10467_46802# a_10809_44734# 4.91e-19
C14542 a_12469_46902# a_10903_43370# 1.97e-19
C14543 a_11813_46116# a_12594_46348# 1.68e-19
C14544 a_11901_46660# a_12005_46116# 1.13e-19
C14545 a_n881_46662# a_n906_45572# 3.16e-20
C14546 a_20916_46384# a_20205_31679# 2.22e-19
C14547 a_4955_46873# a_5066_45546# 0.006456f
C14548 a_22000_46634# a_22365_46825# 0.001038f
C14549 a_20841_46902# a_20820_30879# 4.77e-20
C14550 a_20273_46660# a_12741_44636# 0.540506f
C14551 a_21188_46660# a_20202_43084# 0.002416f
C14552 a_765_45546# a_n2293_46098# 0.054689f
C14553 en_comp a_22775_42308# 9.56e-20
C14554 a_n913_45002# a_22397_42558# 1.07e-20
C14555 a_17730_32519# a_22959_43396# 0.001049f
C14556 a_9313_44734# a_20922_43172# 0.011702f
C14557 a_644_44056# a_743_42282# 5.65e-22
C14558 a_10405_44172# a_10341_43396# 6.35e-20
C14559 a_11257_43940# VDD 9.66e-19
C14560 a_11322_45546# a_11787_45002# 0.035999f
C14561 a_10490_45724# a_11963_45334# 2.16e-19
C14562 a_4880_45572# a_1307_43914# 2.88e-21
C14563 a_19256_45572# a_19418_45938# 0.006453f
C14564 a_18691_45572# a_18953_45572# 0.001705f
C14565 a_2711_45572# a_6517_45366# 3.03e-19
C14566 a_14495_45572# a_6171_45002# 0.002012f
C14567 a_19177_43646# a_17339_46660# 2.77e-19
C14568 a_15682_43940# a_n357_42282# 1.36e-19
C14569 a_8791_43396# a_8199_44636# 1.65e-19
C14570 a_n4318_38216# a_n1613_43370# 1.48e-19
C14571 a_22959_46124# VDD 0.309939f
C14572 a_8746_45002# a_2063_45854# 0.058531f
C14573 a_4880_45572# a_n443_46116# 0.048165f
C14574 a_7499_43078# a_n1151_42308# 6.25e-20
C14575 a_2711_45572# a_12861_44030# 0.104124f
C14576 a_6598_45938# a_6575_47204# 1.53e-21
C14577 a_167_45260# a_n1099_45572# 2.69e-19
C14578 a_1138_42852# a_n755_45592# 0.062548f
C14579 a_1176_45822# a_997_45618# 0.140567f
C14580 a_n901_46420# a_n356_45724# 0.003091f
C14581 a_1823_45246# a_n357_42282# 0.031648f
C14582 a_n2293_46098# a_509_45822# 0.003882f
C14583 a_20708_46348# a_8049_45260# 0.006053f
C14584 a_14275_46494# a_14371_46494# 0.013793f
C14585 a_10903_43370# a_14383_46116# 2.99e-20
C14586 a_4419_46090# a_n2661_45546# 0.019708f
C14587 a_22612_30879# EN_OFFSET_CAL 0.118817f
C14588 a_n2661_46634# DATA[3] 5.46e-21
C14589 a_16547_43609# a_16664_43396# 0.161376f
C14590 a_16243_43396# a_16867_43762# 9.73e-19
C14591 a_16759_43396# a_15743_43084# 0.033478f
C14592 a_17324_43396# a_18525_43370# 0.003432f
C14593 a_20974_43370# a_20922_43172# 0.002377f
C14594 a_21381_43940# a_21195_42852# 0.238789f
C14595 a_2982_43646# a_7765_42852# 3.2e-20
C14596 a_n97_42460# a_15567_42826# 0.040819f
C14597 a_n2661_42282# a_n3674_38216# 0.051505f
C14598 a_2998_44172# a_3823_42558# 8.6e-22
C14599 a_11967_42832# a_15803_42450# 0.258862f
C14600 a_15781_43660# a_15940_43402# 0.002605f
C14601 a_10341_43396# a_20556_43646# 0.008164f
C14602 a_14543_43071# VDD 0.18866f
C14603 a_n2472_45002# a_n2433_44484# 7.88e-19
C14604 a_n2293_45010# a_n2661_44458# 0.031066f
C14605 a_n2661_45010# a_n2129_44697# 0.18531f
C14606 a_2437_43646# a_n699_43396# 0.037149f
C14607 a_6171_45002# a_17719_45144# 8.44e-20
C14608 a_18341_45572# a_18989_43940# 7.86e-20
C14609 a_13017_45260# a_14403_45348# 0.001556f
C14610 a_2903_45348# a_2809_45028# 1.26e-19
C14611 a_8696_44636# a_5891_43370# 0.084594f
C14612 a_10193_42453# a_11967_42832# 0.752992f
C14613 a_19431_45546# a_18287_44626# 6.77e-21
C14614 a_14495_45572# a_14673_44172# 5.52e-19
C14615 COMP_P a_21076_30879# 1.25e-19
C14616 a_5649_42852# a_n755_45592# 0.02386f
C14617 a_11554_42852# a_9290_44172# 0.031758f
C14618 a_2711_45572# a_14180_46812# 2.03e-20
C14619 a_10490_45724# a_11901_46660# 1.82e-20
C14620 a_11525_45546# a_11735_46660# 1.78e-20
C14621 a_11322_45546# a_11813_46116# 3.46e-20
C14622 a_2437_43646# a_22612_30879# 9.37e-20
C14623 a_2382_45260# a_n1613_43370# 2e-21
C14624 a_13348_45260# a_13507_46334# 7.06e-20
C14625 a_1307_43914# a_10227_46804# 0.081555f
C14626 a_4361_42308# a_22400_42852# 4.45e-21
C14627 a_13467_32519# a_14097_32519# 0.048755f
C14628 a_8685_43396# a_9223_42460# 2.83e-20
C14629 a_19339_43156# a_19987_42826# 0.016188f
C14630 a_3626_43646# a_11633_42308# 9.09e-19
C14631 a_19511_42282# VDD 0.244902f
C14632 a_n2109_47186# a_3315_47570# 3.55e-19
C14633 a_6151_47436# a_16023_47582# 6.16e-20
C14634 a_13381_47204# a_n1435_47204# 0.050056f
C14635 a_n971_45724# a_n89_47570# 4.31e-19
C14636 a_2063_45854# a_4883_46098# 0.116597f
C14637 a_17023_45118# a_17061_44734# 1.21e-19
C14638 a_16922_45042# a_17517_44484# 0.020096f
C14639 a_14539_43914# a_16979_44734# 0.132799f
C14640 a_626_44172# a_644_44056# 0.126386f
C14641 a_1307_43914# a_453_43940# 0.05952f
C14642 a_11823_42460# a_2982_43646# 9.47e-19
C14643 a_4223_44672# a_5205_44734# 7.73e-19
C14644 a_n2661_44458# a_9313_44734# 0.00487f
C14645 a_11691_44458# a_13857_44734# 0.049356f
C14646 a_7499_43078# a_6197_43396# 1.44e-19
C14647 a_n1059_45260# a_17973_43940# 0.004269f
C14648 a_n2017_45002# a_18079_43940# 1.02e-20
C14649 a_3065_45002# a_n2661_42282# 1.81e-19
C14650 a_5934_30871# a_n357_42282# 0.001326f
C14651 a_7963_42308# a_n755_45592# 0.003087f
C14652 a_15803_42450# a_13259_45724# 7.39e-19
C14653 a_n2302_39866# a_n2956_39304# 2.06e-19
C14654 a_8192_45572# VDD 0.004463f
C14655 a_2382_45260# a_n2293_46098# 1.97e-20
C14656 a_n23_44458# a_n2293_46634# 2.19e-20
C14657 a_n2012_44484# a_n2438_43548# 0.009651f
C14658 a_n1059_45260# a_167_45260# 1.04e-20
C14659 a_5708_44484# a_768_44030# 0.003906f
C14660 a_10193_42453# a_13259_45724# 0.284945f
C14661 a_1176_45572# a_997_45618# 0.007688f
C14662 a_1260_45572# a_n755_45592# 0.001566f
C14663 a_10210_45822# a_8049_45260# 0.01041f
C14664 a_14815_43914# a_n881_46662# 3.35e-21
C14665 a_18479_45785# a_17957_46116# 7.94e-19
C14666 a_18175_45572# a_18819_46122# 3.23e-19
C14667 a_18341_45572# a_18189_46348# 0.001747f
C14668 a_3357_43084# a_5497_46414# 0.005427f
C14669 a_453_43940# a_n443_46116# 0.004377f
C14670 a_22485_44484# a_12861_44030# 2.25e-19
C14671 a_20980_44850# a_16327_47482# 0.012339f
C14672 a_20766_44850# a_18597_46090# 0.00611f
C14673 a_22223_42860# a_21613_42308# 2.06e-21
C14674 a_n1630_35242# a_1755_42282# 6.88e-21
C14675 a_1184_42692# a_1149_42558# 1.16e-20
C14676 a_n784_42308# a_n39_42308# 4.51e-19
C14677 a_22165_42308# a_22775_42308# 5.13e-19
C14678 a_1067_42314# a_1606_42308# 0.001471f
C14679 a_4791_45118# a_765_45546# 0.052444f
C14680 a_16327_47482# a_19692_46634# 0.023298f
C14681 a_10227_46804# a_17609_46634# 1.17e-19
C14682 a_8128_46384# a_8492_46660# 0.002286f
C14683 a_n881_46662# a_10467_46802# 5.33e-19
C14684 a_33_46660# a_479_46660# 2.28e-19
C14685 a_601_46902# a_1110_47026# 2.6e-19
C14686 a_768_44030# a_5257_43370# 0.028882f
C14687 a_2107_46812# a_1983_46706# 0.212212f
C14688 a_n2438_43548# a_n2661_46098# 0.391488f
C14689 a_n133_46660# a_1799_45572# 3.14e-19
C14690 a_n1925_46634# a_3177_46902# 0.003436f
C14691 a_n743_46660# a_2443_46660# 7.25e-20
C14692 a_5807_45002# a_5907_46634# 0.00171f
C14693 a_n913_45002# a_13887_32519# 1.87e-19
C14694 a_6171_45002# a_16664_43396# 9.32e-20
C14695 a_2711_45572# a_19518_43218# 1.67e-19
C14696 a_7499_43078# a_10752_42852# 1.98e-19
C14697 a_22591_44484# a_19237_31679# 6.8e-19
C14698 a_14537_43396# a_14621_43646# 0.004541f
C14699 a_9313_44734# a_18451_43940# 4.06e-21
C14700 a_n2661_42834# a_10949_43914# 0.037251f
C14701 a_n2661_43922# a_10729_43914# 1.53e-19
C14702 a_1423_45028# a_9885_43646# 1.07e-21
C14703 a_17730_32519# a_22959_44484# 0.015145f
C14704 a_5883_43914# a_9165_43940# 0.019684f
C14705 a_19113_45348# VDD 9.31e-19
C14706 a_15051_42282# RST_Z 0.001018f
C14707 a_n2661_43922# a_n1076_46494# 1.73e-21
C14708 a_3363_44484# a_1823_45246# 0.046566f
C14709 a_19319_43548# a_19321_45002# 3.41e-19
C14710 a_18579_44172# a_17339_46660# 0.016577f
C14711 a_2889_44172# a_3090_45724# 6.33e-21
C14712 a_1423_45028# a_3503_45724# 5.37e-21
C14713 a_21101_45002# a_8049_45260# 9.79e-21
C14714 a_45_45144# a_n2293_45546# 5.47e-19
C14715 a_14309_45348# a_13259_45724# 3.49e-19
C14716 a_15004_44636# a_14840_46494# 2.04e-21
C14717 a_13720_44458# a_2324_44458# 1.95e-20
C14718 a_n1655_43396# a_n1613_43370# 0.001903f
C14719 a_4958_30871# a_n3420_39072# 0.079459f
C14720 a_n784_42308# C6_N_btm 5.52e-19
C14721 a_17609_46634# a_17339_46660# 0.010277f
C14722 a_16292_46812# a_765_45546# 2.99e-38
C14723 a_n881_46662# a_8034_45724# 0.020183f
C14724 a_3877_44458# a_5497_46414# 1.88e-19
C14725 a_4646_46812# a_5204_45822# 1.32e-19
C14726 a_4817_46660# a_4704_46090# 2.68e-19
C14727 a_4651_46660# a_5164_46348# 0.002696f
C14728 a_4955_46873# a_5068_46348# 0.081759f
C14729 a_n2661_46634# a_6945_45028# 0.03015f
C14730 a_5534_30871# VDAC_N 0.009202f
C14731 a_13507_46334# a_18147_46436# 0.001182f
C14732 a_19478_44306# a_19741_43940# 0.005795f
C14733 a_n2661_42282# a_458_43396# 7.55e-21
C14734 a_3905_42865# a_6293_42852# 2.22e-20
C14735 a_11967_42832# a_16137_43396# 0.300696f
C14736 a_10057_43914# a_10835_43094# 9.83e-19
C14737 a_2253_43940# a_2455_43940# 0.092725f
C14738 a_10555_44260# a_10555_43940# 0.001656f
C14739 a_17517_44484# a_15743_43084# 7.31e-22
C14740 a_2382_45260# a_3905_42558# 0.002037f
C14741 a_3537_45260# a_5267_42460# 3.61e-20
C14742 a_n913_45002# a_8515_42308# 0.01424f
C14743 a_3065_45002# a_3497_42558# 0.002517f
C14744 a_2711_45572# a_n913_45002# 3.09e-19
C14745 a_15037_45618# a_15903_45785# 2.5e-20
C14746 a_18083_42858# a_13661_43548# 0.009269f
C14747 a_10341_43396# a_19692_46634# 0.022785f
C14748 a_14621_43646# a_3090_45724# 1.89e-20
C14749 a_n1899_43946# a_n2661_45546# 1.44e-21
C14750 a_20512_43084# a_n357_42282# 0.005311f
C14751 a_9801_43940# a_8953_45546# 9.11e-19
C14752 a_n1329_42308# a_n1151_42308# 0.167748f
C14753 a_13003_42852# a_10227_46804# 0.012229f
C14754 a_n1853_46287# VDD 0.645231f
C14755 a_n4064_40160# a_n4209_37414# 0.055461f
C14756 a_n4315_30879# a_n3565_37414# 0.037486f
C14757 a_n4209_38502# a_n3420_37984# 0.028231f
C14758 a_1343_38525# a_3754_39466# 2.99e-19
C14759 C1_P_btm C0_N_btm 2.15e-19
C14760 C0_P_btm C0_dummy_N_btm 1.3e-19
C14761 a_8016_46348# a_10809_44734# 6.66e-20
C14762 a_8199_44636# a_6945_45028# 5.83e-20
C14763 a_13351_46090# a_2324_44458# 1.29e-20
C14764 a_14493_46090# a_14275_46494# 0.209641f
C14765 a_13759_46122# a_14840_46494# 0.102325f
C14766 a_13925_46122# a_15015_46420# 0.042415f
C14767 a_19123_46287# a_18051_46116# 8.02e-20
C14768 a_2521_46116# a_526_44458# 3.89e-20
C14769 a_2698_46116# a_2981_46116# 0.003683f
C14770 a_1176_45822# a_1337_46116# 0.026848f
C14771 a_20974_43370# a_17364_32525# 0.002207f
C14772 a_5891_43370# a_9377_42558# 0.003627f
C14773 a_8791_43396# a_8945_43396# 0.004009f
C14774 a_n2293_43922# a_6171_42473# 3.54e-20
C14775 a_11341_43940# a_5342_30871# 8.14e-20
C14776 a_11967_42832# a_n784_42308# 4.29e-21
C14777 a_15493_43396# a_18249_42858# 3.35e-20
C14778 a_17538_32519# a_22959_43396# 4.74e-19
C14779 a_3626_43646# a_17499_43370# 4.06e-20
C14780 a_8685_43396# a_13667_43396# 0.005337f
C14781 a_18451_43940# a_18599_43230# 2.19e-19
C14782 a_20990_47178# RST_Z 7.86e-20
C14783 a_19787_47423# SINGLE_ENDED 2.87e-21
C14784 a_20894_47436# START 1.67e-19
C14785 a_21259_43561# VDD 0.192954f
C14786 a_18479_45785# a_18587_45118# 0.003753f
C14787 a_18341_45572# a_18315_45260# 3.86e-19
C14788 a_18175_45572# a_18911_45144# 7.25e-20
C14789 a_13527_45546# a_13720_44458# 3.69e-21
C14790 a_11823_42460# a_14539_43914# 1.51e-19
C14791 a_10193_42453# a_18989_43940# 0.003937f
C14792 a_15861_45028# a_17801_45144# 4.92e-20
C14793 a_327_44734# a_375_42282# 0.067169f
C14794 a_2274_45254# a_1307_43914# 1.47e-19
C14795 a_6171_45002# a_11963_45334# 0.005724f
C14796 a_5111_44636# a_9482_43914# 2.65e-19
C14797 a_413_45260# a_501_45348# 1.71e-19
C14798 a_7229_43940# a_8953_45002# 7.01e-19
C14799 a_6709_45028# a_8191_45002# 9.89e-20
C14800 a_18083_42858# a_4185_45028# 4.75e-20
C14801 a_8147_43396# a_n443_42852# 0.060401f
C14802 a_16137_43396# a_13259_45724# 0.038525f
C14803 a_n3674_39304# a_n2956_39304# 0.029162f
C14804 a_8685_43396# a_n755_45592# 0.001034f
C14805 a_10991_42826# a_9290_44172# 0.045863f
C14806 a_5111_42852# a_2324_44458# 2.92e-22
C14807 a_8696_44636# a_11309_47204# 2.99e-21
C14808 a_3232_43370# a_2063_45854# 0.056568f
C14809 a_8953_45002# a_n237_47217# 9.06e-19
C14810 a_2274_45254# a_n443_46116# 0.041907f
C14811 a_2382_45260# a_4791_45118# 3.36e-20
C14812 a_413_45260# a_5815_47464# 4.35e-19
C14813 a_21350_45938# a_18479_47436# 1.16e-19
C14814 a_2437_43646# a_16588_47582# 0.00737f
C14815 a_3357_43084# a_16327_47482# 0.114502f
C14816 a_20841_45814# a_13507_46334# 3.6e-20
C14817 a_20107_45572# a_4883_46098# 5.13e-20
C14818 a_n2293_45546# a_n357_42282# 0.032623f
C14819 a_n2661_45546# a_1848_45724# 0.005986f
C14820 a_n863_45724# a_n1099_45572# 0.172847f
C14821 a_n452_45724# a_380_45546# 5.21e-19
C14822 a_7871_42858# a_7765_42852# 0.379881f
C14823 a_13678_32519# a_21671_42860# 0.014189f
C14824 a_5649_42852# a_21195_42852# 5.03e-19
C14825 a_13467_32519# a_22959_42860# 2.89e-21
C14826 a_n97_42460# a_6171_42473# 1.26e-20
C14827 a_15493_43940# a_19647_42308# 1.44e-21
C14828 a_11341_43940# a_20107_42308# 2.35e-21
C14829 a_14579_43548# a_15597_42852# 9.38e-19
C14830 a_12281_43396# a_13291_42460# 6.57e-21
C14831 a_1891_43646# a_1606_42308# 1.3e-20
C14832 a_765_45546# DATA[3] 0.004997f
C14833 a_20273_46660# RST_Z 2.21e-21
C14834 a_20107_46660# SINGLE_ENDED 2.88e-21
C14835 a_n4209_37414# a_n4064_37440# 0.265895f
C14836 a_n3565_37414# a_n3420_37440# 0.307576f
C14837 VDAC_Ni a_3726_37500# 1.5261f
C14838 a_4921_42308# VDD 0.214995f
C14839 a_n971_45724# a_1431_47204# 0.030942f
C14840 a_n237_47217# a_1209_47178# 0.206644f
C14841 a_n1741_47186# a_2952_47436# 0.010669f
C14842 a_n2109_47186# a_3160_47472# 0.054333f
C14843 a_n23_47502# a_327_47204# 0.140943f
C14844 a_n746_45260# a_1239_47204# 2.56e-19
C14845 a_n2288_47178# a_n1151_42308# 6.07e-19
C14846 a_n2661_45010# a_n2472_43914# 1.79e-21
C14847 a_1307_43914# a_14815_43914# 0.008091f
C14848 a_8696_44636# a_10807_43548# 1.09e-19
C14849 a_1423_45028# a_n2661_43922# 0.099477f
C14850 a_15765_45572# a_15682_43940# 8.25e-19
C14851 a_22775_42308# a_4185_45028# 0.023674f
C14852 a_n784_42308# a_13259_45724# 4.14e-20
C14853 a_16245_42852# a_n357_42282# 0.008838f
C14854 a_4169_42308# a_526_44458# 6.81e-19
C14855 a_5742_30871# a_n2956_39304# 5.51e-21
C14856 a_20273_45572# a_21363_46634# 2.68e-21
C14857 a_18479_45785# a_11415_45002# 0.047896f
C14858 a_5009_45028# a_4817_46660# 5.42e-22
C14859 a_20107_45572# a_21188_46660# 2.91e-21
C14860 a_11827_44484# a_n2661_46634# 3.03e-20
C14861 a_4099_45572# a_526_44458# 0.063912f
C14862 a_20841_45814# a_20623_46660# 1.29e-20
C14863 a_20528_45572# a_20107_46660# 1.27e-20
C14864 a_6171_45002# a_11901_46660# 1.49e-20
C14865 a_413_45260# a_19333_46634# 1.81e-20
C14866 a_20623_45572# a_20841_46902# 3.35e-20
C14867 a_3537_45260# a_3090_45724# 0.198803f
C14868 a_8953_45002# a_8270_45546# 0.004456f
C14869 a_13527_45546# a_13351_46090# 4.9e-19
C14870 a_13904_45546# a_12594_46348# 0.077346f
C14871 a_11525_45546# a_2324_44458# 0.005847f
C14872 a_11823_42460# a_14493_46090# 2.22e-20
C14873 a_14495_45572# a_10903_43370# 4.3e-19
C14874 a_10907_45822# a_5937_45572# 1.68e-21
C14875 a_10193_42453# a_18189_46348# 1.46e-20
C14876 a_5343_44458# a_n1613_43370# 0.03714f
C14877 a_16979_44734# a_11453_44696# 0.009676f
C14878 a_14112_44734# a_4915_47217# 4.38e-19
C14879 a_12089_42308# a_13249_42558# 2.78e-19
C14880 a_5534_30871# a_5742_30871# 0.069311f
C14881 a_12895_43230# a_13070_42354# 0.006332f
C14882 a_3080_42308# C6_N_btm 2.67e-19
C14883 a_12549_44172# a_13661_43548# 0.149087f
C14884 a_768_44030# a_5807_45002# 0.025167f
C14885 a_12891_46348# a_13747_46662# 6.08e-22
C14886 a_n1613_43370# a_n2956_39768# 3.32e-21
C14887 a_6151_47436# a_8492_46660# 0.302615f
C14888 a_6575_47204# a_7411_46660# 2.14e-19
C14889 a_7227_47204# a_7577_46660# 5.88e-19
C14890 a_4915_47217# a_10428_46928# 7.56e-19
C14891 a_18587_45118# a_14021_43940# 6.84e-23
C14892 a_7499_43078# a_10922_42852# 0.008102f
C14893 a_4223_44672# a_8333_44056# 0.122173f
C14894 a_20193_45348# a_22223_43948# 0.041425f
C14895 a_11691_44458# a_15493_43940# 4.95e-19
C14896 a_5147_45002# a_6293_42852# 8.04e-19
C14897 a_5111_44636# a_6031_43396# 0.207345f
C14898 a_3537_45260# a_6547_43396# 0.03331f
C14899 a_16751_45260# VDD 0.121848f
C14900 a_14097_32519# VCM 0.00888f
C14901 a_1606_42308# EN_VIN_BSTR_N 0.035204f
C14902 a_n784_42308# C4_P_btm 0.001073f
C14903 a_5343_44458# a_n2293_46098# 4.66e-20
C14904 a_19862_44208# a_12549_44172# 0.262561f
C14905 a_13483_43940# a_5807_45002# 1.27e-19
C14906 a_n2293_45010# a_n1099_45572# 0.002597f
C14907 a_n1059_45260# a_n863_45724# 0.162875f
C14908 a_n2956_37592# a_n2472_45546# 4.88e-19
C14909 a_n913_45002# a_n1079_45724# 2.36e-19
C14910 a_n745_45366# a_n2293_45546# 0.038459f
C14911 a_n2661_45010# a_n357_42282# 0.017732f
C14912 a_n2810_45028# a_n2956_38216# 5.73989f
C14913 en_comp a_n2661_45546# 0.001261f
C14914 a_15685_45394# a_2324_44458# 0.002859f
C14915 a_766_43646# a_584_46384# 0.006798f
C14916 a_14401_32519# a_12861_44030# 2.77e-19
C14917 a_15486_42560# a_4958_30871# 0.004787f
C14918 a_14113_42308# a_17531_42308# 8.59e-20
C14919 COMP_P a_1177_38525# 2.71e-19
C14920 a_n4318_38216# a_n4334_38304# 0.081663f
C14921 a_15764_42576# a_16269_42308# 2.28e-19
C14922 a_4915_47217# VDD 3.43172f
C14923 a_6545_47178# a_6640_46482# 9.37e-19
C14924 a_4883_46098# a_17715_44484# 0.024632f
C14925 a_13507_46334# a_17957_46116# 0.007078f
C14926 a_18597_46090# a_19900_46494# 0.039688f
C14927 a_19787_47423# a_19335_46494# 0.001054f
C14928 a_17591_47464# a_10809_44734# 0.007346f
C14929 a_18143_47464# a_6945_45028# 0.023139f
C14930 a_18479_47436# a_21137_46414# 0.002071f
C14931 a_4791_45118# a_6347_46155# 0.005265f
C14932 a_n1151_42308# a_10044_46482# 0.001342f
C14933 a_2063_45854# a_11608_46482# 0.001173f
C14934 a_4190_30871# VDAC_N 0.048476f
C14935 a_11453_44696# a_14275_46494# 6.78e-21
C14936 a_12465_44636# a_15682_46116# 4.04e-20
C14937 a_n881_46662# a_8016_46348# 0.024184f
C14938 a_6755_46942# a_14976_45028# 0.029836f
C14939 a_12549_44172# a_4185_45028# 3.66e-21
C14940 a_16979_44734# a_17324_43396# 1.03e-19
C14941 a_17767_44458# a_17499_43370# 6.82e-20
C14942 a_22959_44484# a_17538_32519# 9.27e-19
C14943 a_5495_43940# a_5745_43940# 0.014406f
C14944 a_14955_43940# a_15493_43396# 2.56e-19
C14945 a_17973_43940# a_18326_43940# 0.009992f
C14946 a_9313_44734# a_9145_43396# 0.021257f
C14947 a_375_42282# a_133_42852# 0.005083f
C14948 a_18114_32519# a_17364_32525# 0.052488f
C14949 a_11823_42460# a_11897_42308# 0.00139f
C14950 a_n2017_45002# a_17749_42852# 0.00371f
C14951 a_n1059_45260# a_17665_42852# 8.77e-19
C14952 a_20447_31679# a_22400_42852# 5.3e-20
C14953 a_2711_45572# a_15903_45785# 0.028735f
C14954 a_11962_45724# a_12791_45546# 0.124167f
C14955 a_12427_45724# a_11823_42460# 0.17307f
C14956 C1_P_btm C10_P_btm 0.31753f
C14957 C1_N_btm EN_VIN_BSTR_N 0.110046f
C14958 a_14955_43940# a_3483_46348# 0.242667f
C14959 a_12710_44260# a_12741_44636# 1.22e-20
C14960 a_14021_43940# a_11415_45002# 3.49e-20
C14961 a_4361_42308# a_13747_46662# 4.79e-20
C14962 a_n97_42460# a_19692_46634# 1.45e-19
C14963 a_n2661_42282# a_5937_45572# 0.060993f
C14964 a_n1545_43230# a_n1613_43370# 1.79e-19
C14965 a_13635_43156# a_10227_46804# 0.320228f
C14966 a_413_45260# CLK 0.033653f
C14967 a_18834_46812# VDD 0.116625f
C14968 a_5934_30871# a_n4064_37440# 0.003932f
C14969 a_1823_45246# a_3147_46376# 1.55e-20
C14970 a_167_45260# a_2698_46116# 0.019127f
C14971 a_14976_45028# a_8049_45260# 0.025611f
C14972 a_765_45546# a_6945_45028# 4.99804f
C14973 a_9313_44734# a_19273_43230# 2.85e-21
C14974 a_15493_43940# a_4190_30871# 8.96e-20
C14975 a_20512_43084# a_21356_42826# 4.04e-19
C14976 a_18184_42460# a_14113_42308# 1.64e-20
C14977 a_n97_42460# a_3457_43396# 1.01e-19
C14978 a_11341_43940# a_743_42282# 3.35e-20
C14979 a_n2833_47464# CLK_DATA 0.331592f
C14980 a_6452_43396# VDD 0.083252f
C14981 a_2711_45572# a_n2661_44458# 3.52e-21
C14982 a_n2109_45247# a_n2017_45002# 0.193269f
C14983 a_n2840_45002# a_n2810_45028# 0.161831f
C14984 a_n2293_45010# a_n1059_45260# 0.020223f
C14985 a_n2661_45010# a_n745_45366# 1.07e-20
C14986 a_21855_43396# a_4185_45028# 7.09e-21
C14987 a_21381_43940# a_n357_42282# 0.060125f
C14988 a_n2433_43396# a_n2293_45546# 9.87e-21
C14989 a_12281_43396# a_10809_44734# 4.31e-19
C14990 a_20107_42308# a_16327_47482# 4.96e-19
C14991 a_11823_42460# a_11453_44696# 0.072491f
C14992 a_13904_45546# a_12465_44636# 1.36e-20
C14993 a_14495_45572# a_4883_46098# 3.88e-20
C14994 a_14033_45822# a_12861_44030# 0.003617f
C14995 a_n1925_42282# a_n863_45724# 1.17e-19
C14996 a_9863_46634# CLK 0.001256f
C14997 a_10428_46928# DATA[5] 0.002585f
C14998 a_22591_43396# a_22959_43396# 7.52e-19
C14999 a_10341_43396# a_5342_30871# 0.001109f
C15000 a_10405_44172# a_10533_42308# 2.11e-21
C15001 a_13887_32519# a_17364_32525# 0.050078f
C15002 a_n97_42460# a_16877_43172# 0.002787f
C15003 a_n4064_37984# a_n2302_37984# 0.250408f
C15004 a_n3420_37984# a_n3607_38304# 8.36e-19
C15005 a_13291_42460# VDD 0.546706f
C15006 a_18479_45785# a_11967_42832# 0.038105f
C15007 a_626_44172# a_949_44458# 0.006992f
C15008 a_1307_43914# a_4743_44484# 0.011512f
C15009 a_9482_43914# a_10334_44484# 0.015932f
C15010 a_2711_45572# a_18451_43940# 0.010207f
C15011 a_n1059_45260# a_9313_44734# 0.089245f
C15012 a_3357_43084# a_n2293_43922# 9.05e-21
C15013 a_3537_45260# a_n356_44636# 4.16e-19
C15014 a_n2661_45010# a_3363_44484# 2.68e-20
C15015 a_7227_42308# a_4185_45028# 1.64e-19
C15016 a_18249_42858# a_n357_42282# 0.047936f
C15017 a_13113_42826# a_n443_42852# 0.001005f
C15018 a_3080_42308# C4_P_btm 5.72e-19
C15019 DATA[5] VDD 0.504354f
C15020 a_2711_45572# a_2804_46116# 1.25e-20
C15021 a_10193_42453# a_20202_43084# 0.296862f
C15022 a_4880_45572# a_n2293_46098# 0.013174f
C15023 a_14033_45822# a_14180_46812# 3.48e-22
C15024 a_14537_43396# a_n2293_46634# 0.036569f
C15025 a_16842_45938# a_3090_45724# 1.14e-19
C15026 a_2437_43646# a_10150_46912# 3.29e-20
C15027 a_3357_43084# a_8667_46634# 2.31e-20
C15028 a_7705_45326# a_2107_46812# 2.71e-20
C15029 a_413_45260# a_3055_46660# 0.002017f
C15030 a_n1655_44484# a_n2497_47436# 8.54e-19
C15031 a_5343_44458# a_4791_45118# 0.003901f
C15032 a_4743_44484# a_n443_46116# 1.56e-21
C15033 a_8975_43940# a_2063_45854# 0.149528f
C15034 a_n2661_44458# a_9313_45822# 3.78e-20
C15035 a_21005_45260# a_18597_46090# 0.034207f
C15036 a_16237_45028# a_16327_47482# 1.67e-19
C15037 a_17719_45144# a_4883_46098# 1.23e-20
C15038 a_4361_42308# a_9293_42558# 5.9e-20
C15039 a_16409_43396# a_17124_42282# 1.26e-20
C15040 a_4520_42826# a_1755_42282# 2.93e-20
C15041 a_10518_42984# a_n784_42308# 2.16e-21
C15042 a_5649_42852# a_8791_42308# 1.31e-19
C15043 a_743_42282# a_10723_42308# 0.008155f
C15044 a_10341_43396# a_20107_42308# 2.81e-20
C15045 a_18249_42858# a_18707_42852# 0.027606f
C15046 a_1847_42826# a_2725_42558# 7.35e-19
C15047 a_4190_30871# a_5742_30871# 0.029789f
C15048 a_20205_31679# a_22521_39511# 3.28e-20
C15049 a_9067_47204# a_5807_45002# 7.49e-20
C15050 a_n1435_47204# a_13675_47204# 0.012767f
C15051 a_13381_47204# a_13759_47204# 8.62e-21
C15052 a_11453_44696# a_22959_47212# 0.182671f
C15053 a_n2109_47186# a_2609_46660# 5.01e-20
C15054 a_n1151_42308# a_n2312_38680# 6.25e-20
C15055 a_1209_47178# a_1123_46634# 0.001301f
C15056 a_3160_47472# a_n1925_46634# 0.026425f
C15057 a_4700_47436# a_n2661_46634# 1.58e-20
C15058 a_584_46384# a_171_46873# 0.007683f
C15059 a_n1741_47186# a_n2661_46098# 3.12e-19
C15060 a_n746_45260# a_491_47026# 0.002692f
C15061 a_11599_46634# a_12891_46348# 0.150715f
C15062 a_14955_47212# a_12549_44172# 7.05e-20
C15063 a_14311_47204# a_768_44030# 0.033509f
C15064 a_5891_43370# a_9159_44484# 6.38e-20
C15065 a_17970_44736# a_17517_44484# 0.075165f
C15066 a_19721_31679# a_22959_44484# 4.31e-19
C15067 a_6109_44484# a_n2661_43922# 0.021636f
C15068 a_7640_43914# a_n2661_42834# 0.030156f
C15069 a_18114_32519# a_19237_31679# 8.86333f
C15070 a_16112_44458# a_16241_44484# 0.010132f
C15071 a_9482_43914# a_13565_44260# 0.003452f
C15072 a_5691_45260# a_5745_43940# 3.63e-21
C15073 a_3357_43084# a_n97_42460# 0.113127f
C15074 a_n2661_45010# a_n2433_43396# 1.83e-20
C15075 a_n2302_40160# a_n2956_38216# 0.001018f
C15076 a_n4209_39590# a_n2810_45572# 0.020489f
C15077 a_21513_45002# VDD 0.416919f
C15078 a_18494_42460# a_20107_46660# 1.14e-20
C15079 a_8701_44490# a_3090_45724# 1.21e-20
C15080 a_n2661_43922# a_4646_46812# 0.06073f
C15081 a_3422_30871# a_19321_45002# 6.52e-21
C15082 a_18479_45785# a_13259_45724# 0.004171f
C15083 a_11963_45334# a_10903_43370# 0.209081f
C15084 a_1423_45028# a_5164_46348# 8.94e-20
C15085 a_9482_43914# a_9290_44172# 0.135239f
C15086 a_1307_43914# a_8016_46348# 0.035949f
C15087 a_453_43940# a_n1613_43370# 1.01e-19
C15088 a_5205_44484# a_2324_44458# 0.523531f
C15089 a_n4318_39768# a_n2312_40392# 0.025298f
C15090 a_15682_43940# a_12861_44030# 0.016729f
C15091 a_8515_42308# a_8325_42308# 0.134955f
C15092 a_5934_30871# a_8685_42308# 0.186981f
C15093 EN_VIN_BSTR_P C6_P_btm 0.118916f
C15094 a_n2293_46634# a_3090_45724# 1.2853f
C15095 a_20843_47204# a_19692_46634# 4.52e-20
C15096 a_n743_46660# a_12991_46634# 1.55e-20
C15097 a_5167_46660# a_5257_43370# 6.3e-20
C15098 a_4646_46812# a_7927_46660# 7.75e-20
C15099 a_768_44030# a_14226_46987# 5.35e-19
C15100 a_5807_45002# a_10933_46660# 0.001833f
C15101 a_12549_44172# a_14543_46987# 3.29e-19
C15102 a_3411_47243# a_765_45546# 2.63e-19
C15103 a_13507_46334# a_11415_45002# 0.160889f
C15104 a_20894_47436# a_12741_44636# 4.32e-20
C15105 a_11453_44696# a_18280_46660# 0.005332f
C15106 a_21496_47436# a_20202_43084# 0.00124f
C15107 a_n1435_47204# a_167_45260# 1.15e-20
C15108 a_n971_45724# a_2324_44458# 0.021839f
C15109 a_n1151_42308# a_9823_46155# 0.061688f
C15110 a_2063_45854# a_11387_46155# 0.079443f
C15111 a_6298_44484# a_7112_43396# 7.71e-19
C15112 a_11967_42832# a_14021_43940# 0.030676f
C15113 a_n356_44636# a_1049_43396# 0.042597f
C15114 a_2479_44172# a_n2661_42282# 3.48e-21
C15115 a_5883_43914# a_6765_43638# 1.3e-19
C15116 a_2998_44172# a_3499_42826# 0.027036f
C15117 a_n3674_39768# a_n1644_44306# 1.74e-19
C15118 a_n2017_45002# a_19339_43156# 0.028127f
C15119 a_n913_45002# a_18817_42826# 2.27e-20
C15120 en_comp a_17701_42308# 1.94e-20
C15121 a_n1059_45260# a_18599_43230# 2.93e-19
C15122 a_3357_43084# a_3935_43218# 2.32e-19
C15123 a_n3565_39590# VREF_GND 0.041931f
C15124 a_700_44734# VDD 0.004666f
C15125 a_n3420_38528# a_n923_35174# 0.002965f
C15126 a_n4064_39072# C5_P_btm 2.13e-20
C15127 a_2711_45572# a_5907_45546# 0.01826f
C15128 a_11341_43940# a_19466_46812# 6.61e-22
C15129 a_15493_43940# a_15227_44166# 0.091653f
C15130 a_n97_42460# a_3877_44458# 3.76e-22
C15131 a_13667_43396# a_768_44030# 2.71e-19
C15132 a_21115_43940# a_19692_46634# 4.88e-20
C15133 a_6547_43396# a_n2293_46634# 0.010751f
C15134 a_14579_43548# a_12549_44172# 1.26e-21
C15135 a_10949_43914# a_13059_46348# 1.57e-20
C15136 a_n2661_44458# a_n1079_45724# 6.12e-21
C15137 a_n2433_44484# a_n2293_45546# 1.15e-19
C15138 a_n310_44484# a_526_44458# 1.02e-20
C15139 a_16241_44734# a_15682_46116# 2.24e-20
C15140 a_8387_43230# a_n971_45724# 0.001371f
C15141 a_3681_42891# a_584_46384# 0.001938f
C15142 a_743_42282# a_16327_47482# 0.026382f
C15143 a_19963_31679# a_22521_40055# 8.31e-21
C15144 a_19479_31679# a_22521_39511# 2.38e-20
C15145 a_n3420_39072# a_n4064_38528# 7.47287f
C15146 a_n2946_39072# a_n2946_38778# 0.050477f
C15147 a_1736_39043# a_2112_39137# 0.554188f
C15148 a_1343_38525# a_2684_37794# 0.224374f
C15149 a_n4064_39072# a_n3420_38528# 0.048218f
C15150 a_n1630_35242# a_2113_38308# 4.08e-20
C15151 a_n1613_43370# a_n906_45572# 2.51e-19
C15152 a_11813_46116# a_12005_46116# 0.038046f
C15153 a_11901_46660# a_10903_43370# 5.8e-19
C15154 a_11735_46660# a_12594_46348# 1.94e-19
C15155 a_10428_46928# a_10809_44734# 1.88e-19
C15156 a_4651_46660# a_5066_45546# 4.76e-19
C15157 a_768_44030# a_n755_45592# 0.202175f
C15158 a_20528_46660# a_20719_46660# 4.61e-19
C15159 a_21188_46660# a_22365_46825# 2e-20
C15160 a_20273_46660# a_20820_30879# 2.63e-19
C15161 a_20411_46873# a_12741_44636# 0.095741f
C15162 a_21363_46634# a_20202_43084# 0.048242f
C15163 a_13483_43940# a_13667_43396# 9.11e-19
C15164 a_15493_43396# a_8685_43396# 0.011009f
C15165 a_9313_44734# a_19987_42826# 0.009103f
C15166 a_20193_45348# a_20753_42852# 0.04748f
C15167 a_375_42282# a_5742_30871# 1.69e-20
C15168 a_17730_32519# a_14209_32519# 0.054558f
C15169 a_19237_31679# a_13887_32519# 0.052352f
C15170 a_20512_43084# a_20749_43396# 0.008222f
C15171 a_n2293_43922# a_5342_30871# 1.2e-20
C15172 a_22485_44484# a_17364_32525# 1e-18
C15173 en_comp a_21613_42308# 2.05e-20
C15174 a_n913_45002# a_21421_42336# 0.001645f
C15175 a_11173_43940# VDD 0.004114f
C15176 a_18479_45785# a_20273_45572# 1.17e-20
C15177 a_10490_45724# a_11787_45002# 1.44e-19
C15178 a_9049_44484# a_9482_43914# 3.58e-19
C15179 a_18691_45572# a_18787_45572# 0.013793f
C15180 a_18909_45814# a_18953_45572# 3.69e-19
C15181 a_11322_45546# a_10951_45334# 4.5e-19
C15182 a_10193_42453# a_13017_45260# 5.13e-21
C15183 a_2711_45572# a_6125_45348# 7.07e-19
C15184 a_13249_42308# a_6171_45002# 0.026329f
C15185 a_16137_43396# a_20202_43084# 5.95e-21
C15186 a_8685_43396# a_3483_46348# 6.46e-19
C15187 a_8037_42858# a_8270_45546# 9.4e-21
C15188 a_14021_43940# a_13259_45724# 0.028871f
C15189 a_14955_43940# a_n357_42282# 2.08e-21
C15190 a_n2661_42282# a_n443_42852# 0.133617f
C15191 a_8147_43396# a_8199_44636# 6.26e-20
C15192 a_10809_44734# VDD 2.67671f
C15193 a_4880_45572# a_4791_45118# 0.006889f
C15194 a_10193_42453# a_2063_45854# 0.114552f
C15195 a_8568_45546# a_n1151_42308# 4.03e-20
C15196 a_167_45260# a_380_45546# 6.63e-19
C15197 a_4185_45028# a_n2661_45546# 0.047991f
C15198 a_1208_46090# a_997_45618# 6.64e-20
C15199 a_1176_45822# a_n755_45592# 0.091892f
C15200 a_1138_42852# a_n357_42282# 0.325445f
C15201 a_n1853_46287# a_7_45899# 1.33e-19
C15202 a_2981_46116# a_526_44458# 0.077706f
C15203 a_19900_46494# a_8049_45260# 0.005334f
C15204 a_13351_46090# a_12839_46116# 7.06e-19
C15205 a_14275_46494# a_14180_46482# 0.049827f
C15206 a_14493_46090# a_14371_46494# 3.16e-19
C15207 a_14358_43442# a_4361_42308# 1.13e-20
C15208 a_16243_43396# a_16664_43396# 0.090164f
C15209 a_16977_43638# a_15743_43084# 0.042866f
C15210 a_11967_42832# a_15764_42576# 0.012941f
C15211 a_17324_43396# a_18429_43548# 1.43e-19
C15212 a_17499_43370# a_18525_43370# 1.4e-19
C15213 a_21381_43940# a_21356_42826# 0.196864f
C15214 a_3626_43646# a_5755_42852# 1.23e-20
C15215 a_2982_43646# a_7871_42858# 4.24e-20
C15216 a_n97_42460# a_5342_30871# 0.068562f
C15217 a_n2661_42282# a_n2104_42282# 4.14e-19
C15218 a_15781_43660# a_15868_43402# 0.004898f
C15219 a_10341_43396# a_743_42282# 0.017833f
C15220 a_21588_30879# EN_OFFSET_CAL 0.047538f
C15221 a_n2661_46634# DATA[2] 1.39e-19
C15222 a_13460_43230# VDD 0.276534f
C15223 en_comp a_3754_38470# 7.78e-19
C15224 a_18909_45814# a_18443_44721# 5.48e-20
C15225 a_18341_45572# a_18374_44850# 7.8e-19
C15226 a_18691_45572# a_18287_44626# 1.75e-20
C15227 a_18479_45785# a_18989_43940# 3.49e-19
C15228 a_8696_44636# a_8375_44464# 0.006586f
C15229 a_375_42282# a_n2293_42834# 0.027465f
C15230 a_13348_45260# a_13490_45394# 0.007833f
C15231 a_2809_45348# a_2809_45028# 6.96e-20
C15232 a_13017_45260# a_14309_45348# 0.002224f
C15233 a_13249_42308# a_14673_44172# 0.026424f
C15234 a_n2472_45002# a_n2661_44458# 0.002026f
C15235 a_n2661_45010# a_n2433_44484# 0.217176f
C15236 a_3357_43084# a_742_44458# 7.16e-19
C15237 a_6171_45002# a_17613_45144# 3.24e-19
C15238 a_n2216_38778# a_n2312_38680# 0.003477f
C15239 a_16823_43084# a_n443_42852# 2.55e-21
C15240 a_5649_42852# a_n357_42282# 0.011202f
C15241 a_11301_43218# a_9290_44172# 0.005694f
C15242 a_2711_45572# a_14035_46660# 1.05e-19
C15243 a_11322_45546# a_11735_46660# 5.37e-20
C15244 a_10490_45724# a_11813_46116# 1.58e-20
C15245 a_9159_45572# a_8667_46634# 1.89e-21
C15246 a_3357_43084# a_20843_47204# 0.006792f
C15247 a_2437_43646# a_21588_30879# 0.001621f
C15248 a_1667_45002# a_n881_46662# 1.43e-20
C15249 a_11963_45334# a_4883_46098# 8.43e-21
C15250 a_16019_45002# a_10227_46804# 0.001575f
C15251 a_6945_45348# a_6545_47178# 2.91e-20
C15252 a_n2661_43370# a_n1151_42308# 0.027798f
C15253 a_8560_45348# a_4791_45118# 6.07e-20
C15254 a_3626_43646# a_10149_42308# 5.71e-19
C15255 a_19339_43156# a_19164_43230# 0.233657f
C15256 a_13467_32519# a_22400_42852# 0.029855f
C15257 a_7227_42852# a_7309_42852# 0.171361f
C15258 a_743_42282# a_20356_42852# 0.001934f
C15259 a_8016_46348# DATA[4] 7.36e-22
C15260 a_n2109_47186# a_3094_47570# 6.18e-19
C15261 a_6151_47436# a_16327_47482# 3.69e-20
C15262 a_11459_47204# a_n1435_47204# 0.001005f
C15263 a_11827_44484# a_15433_44458# 0.002592f
C15264 a_626_44172# a_175_44278# 0.017096f
C15265 a_1307_43914# a_1414_42308# 0.147738f
C15266 a_11691_44458# a_13468_44734# 0.004179f
C15267 a_7499_43078# a_6293_42852# 1.55e-20
C15268 a_n2661_44458# a_9241_44734# 2.59e-19
C15269 a_n1059_45260# a_17737_43940# 6.9e-19
C15270 a_3537_45260# a_3820_44260# 0.001488f
C15271 a_21297_45572# a_19862_44208# 3.66e-20
C15272 a_2437_43646# a_15493_43940# 1.05e-21
C15273 a_6123_31319# a_n755_45592# 0.199766f
C15274 a_7963_42308# a_n357_42282# 4.75e-20
C15275 a_n2946_39866# a_n2956_38680# 3.86e-20
C15276 a_n4064_39616# a_n2956_39304# 3.3e-20
C15277 a_15764_42576# a_13259_45724# 2.69e-19
C15278 a_8120_45572# VDD 3.83e-19
C15279 a_n467_45028# a_n901_46420# 2.24e-19
C15280 a_n356_44636# a_n2293_46634# 6.35e-20
C15281 a_n913_45002# a_1823_45246# 0.041568f
C15282 a_5608_44484# a_768_44030# 0.001348f
C15283 a_11823_42460# a_14180_46482# 2.88e-20
C15284 a_12791_45546# a_12638_46436# 5.55e-20
C15285 a_1176_45572# a_n755_45592# 1.94e-19
C15286 a_9241_45822# a_8049_45260# 7.66e-19
C15287 a_11652_45724# a_11601_46155# 3.78e-19
C15288 a_18175_45572# a_17957_46116# 8.59e-20
C15289 a_18479_45785# a_18189_46348# 2.57e-19
C15290 a_18341_45572# a_17715_44484# 3.97e-20
C15291 a_1414_42308# a_n443_46116# 0.18376f
C15292 a_20512_43084# a_12861_44030# 0.005139f
C15293 a_19789_44512# a_16327_47482# 1.05e-19
C15294 a_19279_43940# a_18479_47436# 0.017993f
C15295 a_20835_44721# a_18597_46090# 0.012854f
C15296 a_11967_42832# a_13507_46334# 0.004262f
C15297 a_22165_42308# a_21613_42308# 0.027246f
C15298 a_1184_42692# a_961_42354# 0.100246f
C15299 a_564_42282# a_1755_42282# 2.36e-20
C15300 a_1067_42314# a_1221_42558# 0.008535f
C15301 a_n1630_35242# a_1606_42308# 0.032246f
C15302 a_n784_42308# a_n327_42308# 1.52e-19
C15303 a_4915_47217# a_14447_46660# 3.78e-19
C15304 a_4700_47436# a_765_45546# 0.004317f
C15305 a_4883_46098# a_11901_46660# 2.38e-19
C15306 a_18597_46090# a_3090_45724# 4.27e-20
C15307 a_16327_47482# a_19466_46812# 0.203994f
C15308 a_10227_46804# a_16292_46812# 3.76e-20
C15309 a_17591_47464# a_17609_46634# 0.014668f
C15310 a_8128_46384# a_8667_46634# 0.001141f
C15311 a_n881_46662# a_10428_46928# 0.004039f
C15312 a_5807_45002# a_5167_46660# 3.94e-19
C15313 a_n2661_46634# a_3067_47026# 0.003055f
C15314 a_33_46660# a_1110_47026# 1.46e-19
C15315 a_383_46660# a_491_47026# 0.057222f
C15316 a_948_46660# a_1983_46706# 3.51e-19
C15317 a_n2438_43548# a_1799_45572# 0.137623f
C15318 a_n1925_46634# a_2609_46660# 0.009041f
C15319 a_n743_46660# a_n2661_46098# 0.414618f
C15320 a_18989_43940# a_14021_43940# 5.23e-19
C15321 a_22591_44484# a_22959_44484# 7.52e-19
C15322 a_n2661_43922# a_10405_44172# 2.51e-20
C15323 a_n2661_42834# a_10729_43914# 0.01161f
C15324 a_9313_44734# a_18326_43940# 1.97e-20
C15325 a_n2661_43370# a_6197_43396# 5.24e-22
C15326 a_14537_43396# a_14537_43646# 0.003096f
C15327 a_22485_44484# a_19237_31679# 3.62e-20
C15328 a_5883_43914# a_8487_44056# 6.48e-19
C15329 a_1307_43914# a_12281_43396# 1.31e-19
C15330 en_comp a_4361_42308# 2.27e-19
C15331 a_n913_45002# a_22223_43396# 2.71e-20
C15332 a_22959_45036# VDD 0.30999f
C15333 a_14113_42308# RST_Z 2.01e-19
C15334 a_n2661_43922# a_n901_46420# 1.04e-20
C15335 a_2675_43914# a_3090_45724# 3.49e-22
C15336 a_1423_45028# a_3316_45546# 1.81e-19
C15337 a_21005_45260# a_8049_45260# 1.99e-20
C15338 a_15415_45028# a_n443_42852# 1.77e-21
C15339 a_13076_44458# a_2324_44458# 7.95e-21
C15340 a_5343_44458# a_6945_45028# 4.48e-20
C15341 a_n1821_43396# a_n1613_43370# 1.79e-19
C15342 a_n881_46662# VDD 2.6692f
C15343 a_7174_31319# a_n3565_39590# 5.27e-21
C15344 a_n784_42308# C5_N_btm 5.81e-19
C15345 a_16292_46812# a_17339_46660# 1.37e-19
C15346 a_3090_45724# a_19123_46287# 2.83e-19
C15347 a_22612_30879# a_10809_44734# 7.79e-20
C15348 a_3877_44458# a_5204_45822# 3.25e-19
C15349 a_4651_46660# a_5068_46348# 8.9e-19
C15350 a_4955_46873# a_4704_46090# 0.109136f
C15351 a_4646_46812# a_5164_46348# 6.79e-20
C15352 a_n743_46660# a_17957_46116# 1.41e-19
C15353 a_12465_44636# a_14537_46482# 5.66e-19
C15354 a_13507_46334# a_13259_45724# 0.023413f
C15355 a_4883_46098# a_15194_46482# 1.02e-19
C15356 a_10057_43914# a_10518_42984# 4.8e-19
C15357 a_20365_43914# a_19319_43548# 0.007317f
C15358 a_3905_42865# a_6031_43396# 4.79e-21
C15359 a_17517_44484# a_18783_43370# 9.36e-21
C15360 a_8975_43940# a_10083_42826# 5.33e-21
C15361 a_9313_44734# a_22959_43396# 0.002204f
C15362 a_n2293_43922# a_743_42282# 0.034167f
C15363 a_11341_43940# a_15037_43940# 0.00577f
C15364 a_19862_44208# a_19478_44056# 4.77e-20
C15365 a_3499_42826# a_1568_43370# 3.66e-21
C15366 a_3537_45260# a_3823_42558# 2.53e-21
C15367 a_n913_45002# a_5934_30871# 0.126791f
C15368 a_n1059_45260# a_8515_42308# 1.02e-20
C15369 a_2382_45260# a_3581_42558# 0.001326f
C15370 a_15037_45618# a_15599_45572# 6.39e-21
C15371 a_2711_45572# a_n1059_45260# 2.83e-19
C15372 a_21671_42860# a_12549_44172# 0.001174f
C15373 a_12379_42858# a_n2293_46634# 1.17e-19
C15374 a_17701_42308# a_13661_43548# 3.31e-20
C15375 a_16855_43396# a_6755_46942# 6.28e-20
C15376 a_n2472_43914# a_n2956_38216# 7.64e-21
C15377 a_9420_43940# a_8953_45546# 2.33e-19
C15378 a_15301_44260# a_2324_44458# 1.99e-19
C15379 a_14021_43940# a_18189_46348# 2.08e-20
C15380 COMP_P a_n1151_42308# 0.034f
C15381 a_13814_43218# a_10227_46804# 0.001965f
C15382 a_n2157_46122# VDD 0.42567f
C15383 a_18214_42558# CAL_N 3.01e-20
C15384 a_n4209_38502# a_n3690_38304# 2.69e-19
C15385 a_n4315_30879# a_n4334_37440# 2.61e-19
C15386 a_7174_31319# a_3726_37500# 0.002891f
C15387 C0_P_btm C0_dummy_P_btm 7.97415f
C15388 C1_P_btm C0_dummy_N_btm 1.59e-19
C15389 a_13925_46122# a_14275_46494# 0.20669f
C15390 a_13759_46122# a_15015_46420# 0.043475f
C15391 a_12594_46348# a_2324_44458# 0.001717f
C15392 a_3090_45724# a_2277_45546# 4.31e-19
C15393 a_18285_46348# a_18051_46116# 0.028958f
C15394 a_1176_45822# a_835_46155# 3.09e-19
C15395 a_1208_46090# a_1337_46116# 0.062574f
C15396 a_167_45260# a_526_44458# 0.003875f
C15397 a_11415_45002# a_10586_45546# 9.19e-19
C15398 a_22315_44484# a_22400_42852# 1.35e-22
C15399 a_18451_43940# a_18817_42826# 4.37e-22
C15400 a_8685_43396# a_10695_43548# 0.00269f
C15401 a_2982_43646# a_17324_43396# 2.59e-21
C15402 a_15493_43396# a_17333_42852# 1.04e-20
C15403 a_n97_42460# a_743_42282# 0.107736f
C15404 a_n2293_43922# a_5755_42308# 8.6e-20
C15405 a_3422_30871# a_14097_32519# 0.031284f
C15406 a_14401_32519# a_17364_32525# 7.51978f
C15407 a_17538_32519# a_14209_32519# 0.051332f
C15408 a_8791_43396# a_8873_43396# 0.005167f
C15409 a_5891_43370# a_9293_42558# 0.001253f
C15410 a_20894_47436# RST_Z 5.48e-20
C15411 SMPL_ON_N a_21589_35634# 0.399184f
C15412 a_19787_47423# START 0.220891f
C15413 a_16023_47582# CLK 0.002544f
C15414 a_19177_43646# VDD 0.004534f
C15415 a_13527_45546# a_13076_44458# 2.47e-21
C15416 a_18479_45785# a_18315_45260# 3.67e-19
C15417 a_18175_45572# a_18587_45118# 0.003125f
C15418 a_19431_45546# a_16922_45042# 2.16e-20
C15419 a_10193_42453# a_18374_44850# 1.66e-20
C15420 a_13249_42308# a_12607_44458# 3.94e-19
C15421 a_15861_45028# a_16981_45144# 9.5e-19
C15422 a_413_45260# a_375_42282# 0.112554f
C15423 a_6171_45002# a_11787_45002# 0.01986f
C15424 a_6709_45028# a_7705_45326# 0.099282f
C15425 a_7229_43940# a_8191_45002# 6.79e-19
C15426 a_17333_42852# a_3483_46348# 1.51e-19
C15427 a_17701_42308# a_4185_45028# 5.35e-20
C15428 a_7112_43396# a_n443_42852# 0.00494f
C15429 a_8685_43396# a_n357_42282# 0.319118f
C15430 a_13943_43396# a_13259_45724# 2.96e-20
C15431 a_10796_42968# a_9290_44172# 0.050429f
C15432 a_16115_45572# a_12549_44172# 1.27e-21
C15433 a_10907_45822# a_n2661_46634# 6.03e-21
C15434 a_1667_45002# a_n443_46116# 4.2e-20
C15435 a_5691_45260# a_2063_45854# 6.94e-20
C15436 a_3232_43370# a_584_46384# 0.277433f
C15437 a_413_45260# a_5129_47502# 1.79e-19
C15438 a_20731_45938# a_18597_46090# 1.8e-20
C15439 a_19479_31679# a_16327_47482# 1.04e-19
C15440 a_2437_43646# a_16763_47508# 0.014946f
C15441 a_3357_43084# a_16241_47178# 1.11e-19
C15442 a_20273_45572# a_13507_46334# 7.72e-20
C15443 a_n2661_45546# a_997_45618# 0.008847f
C15444 a_n863_45724# a_380_45546# 4.95e-19
C15445 a_n1079_45724# a_n1099_45572# 0.15766f
C15446 a_n2472_45546# a_n755_45592# 6.82e-21
C15447 a_n2293_45546# a_310_45028# 0.113595f
C15448 a_20411_46873# RST_Z 1.31e-20
C15449 a_765_45546# DATA[2] 0.006631f
C15450 a_21855_43396# a_21671_42860# 3.61e-19
C15451 a_n97_42460# a_5755_42308# 0.009194f
C15452 a_7227_42852# a_7765_42852# 0.118623f
C15453 a_13678_32519# a_21195_42852# 0.001094f
C15454 a_5649_42852# a_21356_42826# 1.42e-20
C15455 a_13467_32519# a_22223_42860# 3.77e-19
C15456 a_15493_43940# a_19511_42282# 1.21e-21
C15457 a_14579_43548# a_14853_42852# 0.002493f
C15458 a_4361_42308# a_22165_42308# 1.92e-21
C15459 a_1427_43646# a_1606_42308# 6.56e-20
C15460 a_21076_30879# a_22609_37990# 1.29e-20
C15461 a_n3565_37414# a_n3690_37440# 0.247968f
C15462 a_n4334_37440# a_n3420_37440# 0.015567f
C15463 a_n4209_37414# a_n2946_37690# 0.023544f
C15464 a_4933_42558# VDD 0.004279f
C15465 a_n2497_47436# a_n1151_42308# 0.156942f
C15466 a_n23_47502# a_n785_47204# 0.031198f
C15467 a_n237_47217# a_327_47204# 0.027301f
C15468 a_n971_45724# a_1239_47204# 0.022077f
C15469 a_n1741_47186# a_2553_47502# 0.010566f
C15470 a_n2109_47186# a_2905_45572# 0.124881f
C15471 a_n746_45260# a_1209_47178# 1.64e-19
C15472 a_15903_45785# a_15682_43940# 1.25e-19
C15473 a_1423_45028# a_n2661_42834# 1e-18
C15474 a_8696_44636# a_10949_43914# 4.65e-20
C15475 a_7499_43078# a_7499_43940# 0.003097f
C15476 a_n913_45002# a_20512_43084# 1.33e-19
C15477 a_21613_42308# a_4185_45028# 0.028903f
C15478 a_15953_42852# a_n357_42282# 0.00164f
C15479 a_15720_42674# a_2324_44458# 2.94e-22
C15480 a_20273_45572# a_20623_46660# 1.3e-20
C15481 a_18175_45572# a_11415_45002# 0.003704f
C15482 a_5093_45028# a_4651_46660# 1.49e-21
C15483 a_5009_45028# a_4955_46873# 4.28e-21
C15484 a_14537_43396# a_6755_46942# 0.120241f
C15485 a_5837_45028# a_4646_46812# 1.48e-21
C15486 a_2711_45572# a_n1925_42282# 0.019937f
C15487 a_3175_45822# a_526_44458# 0.003323f
C15488 a_8191_45002# a_8270_45546# 0.001376f
C15489 a_6171_45002# a_11813_46116# 1.01e-20
C15490 a_21188_45572# a_20107_46660# 2.1e-20
C15491 a_20623_45572# a_20273_46660# 3.64e-20
C15492 a_20841_45814# a_20841_46902# 8.24e-19
C15493 a_3357_43084# a_16721_46634# 7.55e-22
C15494 a_413_45260# a_15227_44166# 4.28e-20
C15495 a_3429_45260# a_3090_45724# 0.004791f
C15496 a_n699_43396# a_n881_46662# 6.09e-22
C15497 a_13527_45546# a_12594_46348# 0.100424f
C15498 a_11322_45546# a_2324_44458# 0.068998f
C15499 a_13249_42308# a_10903_43370# 0.211356f
C15500 a_11823_42460# a_13925_46122# 2.39e-19
C15501 a_13163_45724# a_13351_46090# 3.18e-19
C15502 a_10907_45822# a_8199_44636# 0.081841f
C15503 a_10193_42453# a_17715_44484# 0.074403f
C15504 a_10210_45822# a_5937_45572# 2.86e-19
C15505 a_9241_45822# a_8953_45546# 2.68e-20
C15506 a_14539_43914# a_11453_44696# 0.006758f
C15507 a_13113_42826# a_13070_42354# 4.26e-19
C15508 a_12545_42858# a_13575_42558# 0.001596f
C15509 a_14209_32519# a_22465_38105# 6.41e-20
C15510 a_3080_42308# C5_N_btm 3.03e-19
C15511 a_12549_44172# a_5807_45002# 0.675558f
C15512 a_12891_46348# a_13661_43548# 0.001729f
C15513 a_2747_46873# a_n2438_43548# 8.92e-19
C15514 a_6575_47204# a_5257_43370# 1.06e-19
C15515 a_4915_47217# a_10150_46912# 9.74e-20
C15516 a_6151_47436# a_8667_46634# 0.357581f
C15517 a_7227_47204# a_7715_46873# 3.86e-19
C15518 a_7903_47542# a_7411_46660# 0.001091f
C15519 a_n1741_47186# a_12251_46660# 0.011505f
C15520 a_2063_45854# a_8035_47026# 0.004006f
C15521 a_n237_47217# a_8846_46660# 7.11e-19
C15522 a_7499_43078# a_10991_42826# 0.004793f
C15523 a_626_44172# a_n97_42460# 0.005505f
C15524 a_20193_45348# a_11341_43940# 0.21261f
C15525 a_10193_42453# a_10083_42826# 0.002709f
C15526 a_2711_45572# a_19987_42826# 0.003709f
C15527 a_9313_44734# a_22959_44484# 1.37e-19
C15528 a_3537_45260# a_6765_43638# 0.025724f
C15529 a_5147_45002# a_6031_43396# 0.003581f
C15530 a_1307_43914# VDD 3.92807f
C15531 a_14097_32519# VREF_GND 0.047244f
C15532 a_1606_42308# a_11530_34132# 0.004863f
C15533 a_n784_42308# C5_P_btm 5.81e-19
C15534 a_n2661_44458# a_1823_45246# 0.036985f
C15535 a_n452_44636# a_n901_46420# 1.9e-20
C15536 a_4743_44484# a_n2293_46098# 0.002464f
C15537 a_19478_44306# a_12549_44172# 0.010691f
C15538 a_1423_45028# a_5066_45546# 3.17e-20
C15539 a_14537_43396# a_8049_45260# 3.16e-21
C15540 a_n1059_45260# a_n1079_45724# 0.003242f
C15541 a_n913_45002# a_n2293_45546# 0.043147f
C15542 a_n2017_45002# a_n863_45724# 0.111825f
C15543 a_n2956_37592# a_n2661_45546# 6.64e-20
C15544 a_n2661_45010# a_310_45028# 1.15e-19
C15545 en_comp a_n2810_45572# 2.18e-19
C15546 a_14309_45028# a_14493_46090# 1.04e-20
C15547 a_15060_45348# a_2324_44458# 0.004184f
C15548 a_21381_43940# a_12861_44030# 0.019154f
C15549 a_n443_46116# VDD 3.87014f
C15550 a_15051_42282# a_4958_30871# 0.003379f
C15551 a_14113_42308# a_17303_42282# 1.39e-19
C15552 a_n4318_38216# a_n4209_38216# 0.135236f
C15553 a_n3674_37592# a_n3565_38502# 9.8e-20
C15554 a_n1630_35242# a_n4209_38502# 3.02e-19
C15555 a_15803_42450# a_15761_42308# 2.56e-19
C15556 a_n784_42308# a_n3420_38528# 0.005039f
C15557 a_5932_42308# a_n3565_39590# 4.83e-21
C15558 a_n3674_38216# a_n4251_38528# 5.77e-20
C15559 a_11453_44696# a_14493_46090# 1.13e-21
C15560 a_12465_44636# a_2324_44458# 0.070016f
C15561 a_6491_46660# a_5066_45546# 2.85e-21
C15562 a_4883_46098# a_17583_46090# 0.012469f
C15563 a_13507_46334# a_18189_46348# 0.001569f
C15564 a_18597_46090# a_20075_46420# 0.073857f
C15565 a_18479_47436# a_20708_46348# 0.04299f
C15566 a_19386_47436# a_19335_46494# 3.45e-20
C15567 a_19787_47423# a_19553_46090# 9.41e-20
C15568 a_16588_47582# a_10809_44734# 9.65e-20
C15569 a_10227_46804# a_6945_45028# 0.220094f
C15570 a_4791_45118# a_8034_45724# 2.34e-20
C15571 a_n1151_42308# a_9823_46482# 1.61e-19
C15572 a_2063_45854# a_11387_46482# 2.86e-19
C15573 a_n881_46662# a_7920_46348# 0.025724f
C15574 a_3067_47026# a_765_45546# 0.002408f
C15575 a_8270_45546# a_8846_46660# 7.05e-19
C15576 a_6755_46942# a_3090_45724# 0.050558f
C15577 a_n743_46660# a_11415_45002# 0.038831f
C15578 a_n2661_46634# a_n2840_46090# 3.35e-19
C15579 a_768_44030# a_3483_46348# 0.281593f
C15580 a_16979_44734# a_17499_43370# 6.72e-19
C15581 a_17973_43940# a_18079_43940# 0.419086f
C15582 a_742_44458# a_743_42282# 6.63e-20
C15583 a_14539_43914# a_17324_43396# 0.008599f
C15584 a_17730_32519# a_17538_32519# 9.37324f
C15585 a_19237_31679# a_14401_32519# 0.055111f
C15586 a_19721_31679# a_14209_32519# 0.051313f
C15587 a_5013_44260# a_5745_43940# 0.007387f
C15588 a_5495_43940# a_5326_44056# 4.96e-19
C15589 a_17737_43940# a_18326_43940# 4.1e-19
C15590 a_n1059_45260# a_16877_42852# 0.058551f
C15591 a_19963_31679# a_14097_32519# 0.051059f
C15592 a_n2017_45002# a_17665_42852# 0.004242f
C15593 a_18579_44172# VDD 0.38178f
C15594 a_2711_45572# a_15599_45572# 0.045207f
C15595 a_11962_45724# a_11823_42460# 0.177935f
C15596 a_8162_45546# a_8336_45822# 9.93e-20
C15597 C0_N_btm EN_VIN_BSTR_N 0.12803f
C15598 a_13483_43940# a_3483_46348# 0.194464f
C15599 a_14021_43940# a_20202_43084# 0.020234f
C15600 a_4361_42308# a_13661_43548# 6.79e-20
C15601 a_20835_44721# a_8049_45260# 3.74e-21
C15602 a_13296_44484# a_13259_45724# 0.002753f
C15603 a_n89_44484# a_n863_45724# 8.7e-19
C15604 a_6101_44260# a_5937_45572# 9.35e-20
C15605 a_n1736_43218# a_n1613_43370# 2.47e-19
C15606 a_12895_43230# a_10227_46804# 0.152365f
C15607 a_18249_42858# a_12861_44030# 6.95e-20
C15608 a_413_45260# EN_OFFSET_CAL 0.114452f
C15609 a_17609_46634# VDD 0.501057f
C15610 a_1823_45246# a_2804_46116# 1.33e-21
C15611 a_167_45260# a_2521_46116# 0.328009f
C15612 a_3877_44458# a_3503_45724# 0.001651f
C15613 a_3090_45724# a_8049_45260# 1.23904f
C15614 a_5257_43370# a_n2661_45546# 0.003554f
C15615 a_6755_46942# a_15002_46116# 3.59e-20
C15616 a_11415_45002# a_11189_46129# 0.001065f
C15617 a_19551_46910# a_19335_46494# 6.39e-20
C15618 a_20411_46873# a_18985_46122# 1.23e-19
C15619 a_17339_46660# a_6945_45028# 6.42e-20
C15620 a_5932_42308# a_3726_37500# 0.003378f
C15621 a_9313_44734# a_18861_43218# 2.63e-19
C15622 a_15493_43940# a_21259_43561# 8.06e-20
C15623 a_20512_43084# a_20922_43172# 0.001051f
C15624 a_19862_44208# a_4361_42308# 0.006467f
C15625 a_2896_43646# a_2982_43646# 0.100706f
C15626 a_n97_42460# a_2813_43396# 0.001563f
C15627 a_14021_43940# a_16867_43762# 0.004651f
C15628 a_11341_43940# a_20301_43646# 0.001136f
C15629 a_9396_43370# VDD 0.288403f
C15630 a_11823_42460# a_13807_45067# 1.27e-21
C15631 a_13249_42308# a_14403_45348# 8.12e-19
C15632 a_n2293_45010# a_n2017_45002# 0.076023f
C15633 a_n2661_45010# a_n913_45002# 0.019536f
C15634 a_2437_43646# a_413_45260# 0.20387f
C15635 a_n2472_45002# a_n1059_45260# 7.79e-20
C15636 a_20447_31679# en_comp 2.2e-19
C15637 a_4361_42308# a_4185_45028# 0.042181f
C15638 a_3823_42558# a_n2293_46634# 8.78e-21
C15639 a_16137_43396# a_17715_44484# 1.22e-20
C15640 a_n3420_38528# SMPL_ON_P 8.16e-21
C15641 a_13258_32519# a_16327_47482# 0.019817f
C15642 a_19443_46116# VDD 0.132317f
C15643 a_13527_45546# a_12465_44636# 6.66e-22
C15644 a_12427_45724# a_11453_44696# 5.75e-21
C15645 a_15143_45578# a_13507_46334# 3.04e-21
C15646 a_13249_42308# a_4883_46098# 3.03e-20
C15647 a_8049_45260# a_15002_46116# 1.39e-19
C15648 a_14180_46482# a_14371_46494# 4.61e-19
C15649 a_526_44458# a_n863_45724# 0.801581f
C15650 a_22591_43396# a_14209_32519# 0.158752f
C15651 a_10341_43396# a_15279_43071# 0.001151f
C15652 a_22223_43396# a_17364_32525# 2.46e-19
C15653 a_n97_42460# a_16328_43172# 7.85e-19
C15654 a_17730_32519# a_22465_38105# 2.17e-19
C15655 a_n3690_38304# a_n3607_38304# 0.007692f
C15656 a_n2946_37984# a_n2302_37984# 6.68e-19
C15657 a_13003_42852# VDD 0.132655f
C15658 a_18175_45572# a_11967_42832# 4.42e-21
C15659 a_18341_45572# a_18588_44850# 5.56e-21
C15660 a_11963_45334# a_8975_43940# 4.93e-19
C15661 a_9482_43914# a_10157_44484# 0.321004f
C15662 a_626_44172# a_742_44458# 0.022141f
C15663 a_1307_43914# a_n699_43396# 0.094953f
C15664 a_2711_45572# a_18326_43940# 0.009029f
C15665 en_comp a_5891_43370# 2.34e-21
C15666 a_327_44734# a_700_44734# 0.003235f
C15667 a_n2661_45010# a_556_44484# 0.038106f
C15668 a_n2017_45002# a_9313_44734# 0.009039f
C15669 a_3357_43084# a_n2661_43922# 0.031253f
C15670 a_6761_42308# a_4185_45028# 9.41e-20
C15671 a_12545_42858# a_n443_42852# 7.04e-20
C15672 a_17333_42852# a_n357_42282# 0.05273f
C15673 a_3080_42308# C5_P_btm 3.03e-19
C15674 DATA[4] VDD 0.326957f
C15675 a_2711_45572# a_2698_46116# 6.21e-20
C15676 a_4808_45572# a_n2293_46098# 0.001218f
C15677 a_14033_45822# a_14035_46660# 0.001323f
C15678 a_13159_45002# a_n743_46660# 7.14e-21
C15679 a_3357_43084# a_7927_46660# 1.64e-20
C15680 a_2437_43646# a_9863_46634# 9.58e-21
C15681 a_4743_44484# a_4791_45118# 0.165321f
C15682 a_10057_43914# a_2063_45854# 0.06633f
C15683 a_n699_43396# a_n443_46116# 0.042248f
C15684 a_n1821_44484# a_n2497_47436# 0.001505f
C15685 a_5883_43914# a_n1151_42308# 1.46e-20
C15686 a_19929_45028# a_12861_44030# 7.5e-19
C15687 a_21101_45002# a_18479_47436# 0.001064f
C15688 a_20567_45036# a_18597_46090# 0.001626f
C15689 a_20193_45348# a_16327_47482# 0.359904f
C15690 a_11827_44484# a_10227_46804# 0.065169f
C15691 a_18315_45260# a_13507_46334# 8.76e-37
C15692 a_14309_45028# a_11453_44696# 0.004516f
C15693 a_10341_43396# a_13258_32519# 2.74e-20
C15694 a_3935_42891# a_1755_42282# 3.67e-22
C15695 a_10083_42826# a_n784_42308# 8.21e-21
C15696 a_18083_42858# a_20256_43172# 9.94e-21
C15697 a_5649_42852# a_8685_42308# 5.5e-20
C15698 a_4361_42308# a_9803_42558# 0.011987f
C15699 a_743_42282# a_10533_42308# 0.016446f
C15700 a_18599_43230# a_18861_43218# 0.001705f
C15701 a_18817_42826# a_19273_43230# 4.2e-19
C15702 a_3080_42308# a_n3420_38528# 1.75e-20
C15703 a_20692_30879# a_22459_39145# 3e-20
C15704 a_n3565_38216# VDD 0.901259f
C15705 a_14311_47204# a_12549_44172# 7.38e-20
C15706 a_13487_47204# a_768_44030# 0.371206f
C15707 a_n1435_47204# a_13569_47204# 0.011393f
C15708 a_13381_47204# a_13675_47204# 1.29e-20
C15709 a_11599_46634# a_11309_47204# 0.008095f
C15710 a_6575_47204# a_5807_45002# 1.65e-19
C15711 SMPL_ON_N a_22959_47212# 0.007483f
C15712 a_n2109_47186# a_2443_46660# 2.98e-19
C15713 a_n1741_47186# a_1799_45572# 2.42e-19
C15714 a_584_46384# a_n133_46660# 2.89e-19
C15715 a_n1151_42308# a_n2104_46634# 3.6e-20
C15716 a_n1920_47178# a_n2661_46098# 3.04e-20
C15717 a_2063_45854# a_n2438_43548# 0.033724f
C15718 a_2905_45572# a_n1925_46634# 0.029452f
C15719 a_4007_47204# a_n2661_46634# 1.08e-19
C15720 a_n746_45260# a_288_46660# 0.010226f
C15721 a_n237_47217# a_1983_46706# 8.91e-19
C15722 a_17970_44736# a_17061_44734# 1.93e-19
C15723 a_17767_44458# a_17517_44484# 0.055175f
C15724 a_18114_32519# a_22959_44484# 0.016108f
C15725 a_6109_44484# a_n2661_42834# 0.026239f
C15726 a_19721_31679# a_17730_32519# 0.051334f
C15727 a_9482_43914# a_12710_44260# 0.001272f
C15728 a_n2293_42834# a_8018_44260# 0.001899f
C15729 a_5111_44636# a_5829_43940# 1.13e-20
C15730 a_n913_45002# a_21381_43940# 5.97e-20
C15731 a_3537_45260# a_8487_44056# 2.95e-19
C15732 a_n4064_40160# a_n2956_38216# 9.27e-19
C15733 a_11967_42832# a_n743_46660# 7.36e-20
C15734 a_18184_42460# a_20107_46660# 3.9e-21
C15735 a_n2661_43922# a_3877_44458# 0.021496f
C15736 a_n2661_42834# a_4646_46812# 0.030297f
C15737 a_11827_44484# a_17339_46660# 0.031147f
C15738 a_19778_44110# a_20411_46873# 1.83e-20
C15739 a_16922_45042# a_20528_46660# 3.33e-20
C15740 a_18175_45572# a_13259_45724# 3.33e-19
C15741 a_413_45260# a_22959_46124# 0.020082f
C15742 a_n2293_45010# a_526_44458# 2.25e-19
C15743 a_20731_45938# a_8049_45260# 0.005076f
C15744 a_n967_45348# a_n967_46494# 1.79e-21
C15745 a_11787_45002# a_10903_43370# 0.003455f
C15746 a_6171_45002# a_15682_46116# 2.79e-19
C15747 a_6431_45366# a_2324_44458# 0.046214f
C15748 a_14955_43940# a_12861_44030# 0.001655f
C15749 a_4921_42308# a_5742_30871# 3.53e-20
C15750 a_5934_30871# a_8325_42308# 0.173576f
C15751 a_8515_42308# a_8337_42558# 6.01e-20
C15752 a_7963_42308# a_8685_42308# 2.62e-19
C15753 a_18194_35068# a_21589_35634# 4.88e-19
C15754 a_19120_35138# a_19864_35138# 0.081924f
C15755 EN_VIN_BSTR_P C7_P_btm 0.115875f
C15756 a_22459_39145# VIN_N 2.29e-20
C15757 a_20916_46384# a_15227_44166# 0.681561f
C15758 a_n743_46660# a_12251_46660# 3.96e-20
C15759 a_19594_46812# a_19692_46634# 0.134424f
C15760 a_5732_46660# a_5894_47026# 0.006453f
C15761 a_5167_46660# a_5429_46660# 0.001705f
C15762 a_4817_46660# a_7411_46660# 1.88e-20
C15763 a_4646_46812# a_8145_46902# 1.81e-20
C15764 a_5385_46902# a_5257_43370# 5.44e-20
C15765 a_3877_44458# a_7927_46660# 3.05e-20
C15766 a_768_44030# a_14513_46634# 8.17e-21
C15767 a_5807_45002# a_10861_46660# 0.00101f
C15768 a_12549_44172# a_14226_46987# 3.77e-19
C15769 a_3094_47243# a_765_45546# 4.26e-19
C15770 a_13507_46334# a_20202_43084# 0.205796f
C15771 a_11453_44696# a_17639_46660# 2.16e-19
C15772 a_n1435_47204# a_2202_46116# 1.01e-21
C15773 a_9067_47204# a_3483_46348# 9.45e-22
C15774 a_6151_47436# a_5204_45822# 1.22e-19
C15775 a_2063_45854# a_11133_46155# 0.026232f
C15776 a_n1151_42308# a_9569_46155# 0.05766f
C15777 a_4791_45118# a_8016_46348# 0.001293f
C15778 a_6298_44484# a_7287_43370# 0.003354f
C15779 a_20980_44850# a_20935_43940# 1.59e-19
C15780 a_5343_44458# a_8147_43396# 0.014327f
C15781 a_n356_44636# a_1209_43370# 0.025313f
C15782 a_5883_43914# a_6197_43396# 0.001031f
C15783 a_16922_45042# a_16409_43396# 4.18e-21
C15784 a_20193_45348# a_10341_43396# 0.086741f
C15785 a_742_44458# a_2813_43396# 1.77e-19
C15786 a_375_42282# a_n13_43084# 0.006217f
C15787 a_2998_44172# a_2537_44260# 3.26e-21
C15788 a_n913_45002# a_18249_42858# 4.01e-20
C15789 a_n2017_45002# a_18599_43230# 0.029677f
C15790 en_comp a_17595_43084# 2.61e-21
C15791 a_3357_43084# a_3445_43172# 5.23e-19
C15792 a_n1059_45260# a_18817_42826# 1.2e-20
C15793 a_n998_44484# VDD 1.32e-19
C15794 a_n4209_39590# VCM 0.179761f
C15795 a_n3565_39590# VREF 0.417978f
C15796 a_n3420_39616# VIN_P 0.041227f
C15797 a_n3565_38502# EN_VIN_BSTR_P 0.003421f
C15798 a_n4064_39072# C6_P_btm 2.76e-20
C15799 a_n3565_39304# C2_P_btm 1.93e-20
C15800 a_n4064_37440# a_n2956_38216# 0.001421f
C15801 a_2711_45572# a_5263_45724# 0.013854f
C15802 a_20935_43940# a_19692_46634# 6.93e-20
C15803 a_6765_43638# a_n2293_46634# 0.011639f
C15804 a_10695_43548# a_768_44030# 3.8e-21
C15805 a_n2267_44484# a_n2661_45546# 2.71e-20
C15806 a_13076_44458# a_12839_46116# 4.31e-21
C15807 a_9313_44734# a_526_44458# 4.07e-20
C15808 a_n2433_44484# a_n2956_38216# 7.79e-19
C15809 a_n2661_44458# a_n2293_45546# 0.006992f
C15810 a_n2293_43922# a_n2956_38680# 3.35e-20
C15811 a_2905_42968# a_584_46384# 3.05e-20
C15812 a_8605_42826# a_n971_45724# 0.001728f
C15813 a_5649_42852# a_12861_44030# 1.34e-19
C15814 a_20301_43646# a_16327_47482# 4.99e-19
C15815 a_17324_43396# a_11453_44696# 1.49e-21
C15816 a_n3690_39392# a_n4064_38528# 6.81e-20
C15817 a_n3420_39072# a_n2946_38778# 2.59e-20
C15818 a_n3565_39304# a_n2302_38778# 8.25e-19
C15819 a_1343_38525# a_1177_38525# 0.238422f
C15820 a_n4064_39072# a_n3690_38528# 6.81e-20
C15821 a_n2946_39072# a_n3420_38528# 2.59e-20
C15822 COMP_P VDAC_Pi 0.005217f
C15823 a_3090_45724# a_8953_45546# 0.032771f
C15824 a_10467_46802# a_6945_45028# 1.12e-19
C15825 a_11813_46116# a_10903_43370# 0.006138f
C15826 a_11735_46660# a_12005_46116# 2.1e-19
C15827 a_4955_46873# a_5210_46482# 9.61e-19
C15828 a_20916_46384# a_21071_46482# 0.006088f
C15829 a_768_44030# a_n357_42282# 0.175577f
C15830 a_4646_46812# a_5066_45546# 0.020397f
C15831 a_n743_46660# a_13259_45724# 0.025444f
C15832 a_20623_46660# a_20202_43084# 1.78e-20
C15833 a_20273_46660# a_22591_46660# 6.79e-20
C15834 a_20107_46660# a_12741_44636# 0.527863f
C15835 a_9313_44734# a_19164_43230# 0.004691f
C15836 a_n2293_42834# a_4921_42308# 2.38e-19
C15837 a_20512_43084# a_17364_32525# 1.45e-20
C15838 a_17730_32519# a_22591_43396# 7.33e-19
C15839 en_comp a_21887_42336# 2.22e-20
C15840 a_10867_43940# VDD 0.008055f
C15841 a_18175_45572# a_20273_45572# 3.92e-21
C15842 a_3775_45552# a_1423_45028# 4.78e-21
C15843 a_18479_45785# a_20107_45572# 3.61e-20
C15844 a_10490_45724# a_10951_45334# 1.32e-19
C15845 a_10193_42453# a_11963_45334# 0.007668f
C15846 a_7499_43078# a_9482_43914# 0.062333f
C15847 a_18909_45814# a_18787_45572# 3.16e-19
C15848 a_11322_45546# a_10775_45002# 6.82e-20
C15849 a_2711_45572# a_5837_45348# 3.63e-19
C15850 a_13904_45546# a_6171_45002# 3.3e-20
C15851 a_20256_43172# a_12549_44172# 5.03e-21
C15852 a_13483_43940# a_n357_42282# 1.74e-20
C15853 a_7287_43370# a_5937_45572# 8.77e-22
C15854 a_n1630_35242# a_n2312_39304# 0.002065f
C15855 a_22223_46124# VDD 0.300745f
C15856 a_8162_45546# a_n1151_42308# 0.004489f
C15857 a_5024_45822# a_n443_46116# 0.009847f
C15858 a_10180_45724# a_2063_45854# 0.002207f
C15859 a_4808_45572# a_4791_45118# 0.00122f
C15860 a_6511_45714# a_6575_47204# 2.63e-21
C15861 a_3699_46348# a_n2661_45546# 1.29e-20
C15862 a_1208_46090# a_n755_45592# 0.004994f
C15863 a_2521_46116# a_n863_45724# 9.29e-20
C15864 a_1176_45822# a_n357_42282# 0.001329f
C15865 a_n1853_46287# a_n310_45899# 9.42e-19
C15866 a_6945_45028# a_8034_45724# 4.34e-21
C15867 a_20075_46420# a_8049_45260# 0.005224f
C15868 a_12594_46348# a_12839_46116# 0.002912f
C15869 a_13925_46122# a_14371_46494# 2.28e-19
C15870 a_14579_43548# a_4361_42308# 2.32e-19
C15871 a_17499_43370# a_18429_43548# 0.012474f
C15872 a_16409_43396# a_15743_43084# 0.586918f
C15873 a_3539_42460# a_4520_42826# 0.003363f
C15874 a_3626_43646# a_5111_42852# 3.39e-20
C15875 a_n97_42460# a_15279_43071# 0.001255f
C15876 a_21381_43940# a_20922_43172# 0.00196f
C15877 a_n2661_42282# a_n4318_38216# 0.023731f
C15878 a_2998_44172# a_2903_42308# 4.71e-20
C15879 a_11967_42832# a_15486_42560# 1.23e-19
C15880 a_15681_43442# a_15868_43402# 1.84e-19
C15881 a_16137_43396# a_16664_43396# 0.002125f
C15882 a_10341_43396# a_20301_43646# 0.002799f
C15883 a_20916_46384# EN_OFFSET_CAL 8.73e-21
C15884 a_n2661_46634# DATA[1] 1.37e-19
C15885 a_n2442_46660# CLK_DATA 0.063913f
C15886 a_13635_43156# VDD 0.463701f
C15887 a_18909_45814# a_18287_44626# 8.28e-19
C15888 a_18479_45785# a_18374_44850# 3.69e-20
C15889 a_18341_45572# a_18443_44721# 3.12e-21
C15890 a_18691_45572# a_18248_44752# 2.36e-21
C15891 a_13159_45002# a_13490_45394# 2.88e-19
C15892 a_13017_45260# a_13711_45394# 2.64e-19
C15893 a_8696_44636# a_7640_43914# 9.09e-20
C15894 a_13249_42308# a_14581_44484# 1.15e-19
C15895 a_18175_45572# a_18989_43940# 6.34e-20
C15896 a_n2661_45010# a_n2661_44458# 0.090852f
C15897 a_6171_45002# a_17023_45118# 7.32e-19
C15898 a_14456_42282# a_3090_45724# 4.19e-20
C15899 a_n2860_38778# a_n2312_38680# 6.16e-19
C15900 a_13678_32519# a_n357_42282# 1.42e-19
C15901 a_11229_43218# a_9290_44172# 0.002961f
C15902 a_2711_45572# a_13885_46660# 1.07e-21
C15903 a_10490_45724# a_11735_46660# 2.75e-20
C15904 a_10193_42453# a_11901_46660# 4.59e-19
C15905 a_2437_43646# a_20916_46384# 0.010579f
C15906 a_3357_43084# a_19594_46812# 4.56e-19
C15907 a_327_44734# a_n881_46662# 3.44e-20
C15908 a_11787_45002# a_4883_46098# 1.41e-20
C15909 a_13017_45260# a_13507_46334# 2.21e-20
C15910 a_15595_45028# a_10227_46804# 0.002256f
C15911 a_3626_43646# a_9885_42308# 0.001057f
C15912 a_8685_43396# a_8685_42308# 9.74e-19
C15913 a_8387_43230# a_8483_43230# 0.013793f
C15914 a_18599_43230# a_19164_43230# 7.99e-20
C15915 a_9145_43396# a_5934_30871# 3.25e-19
C15916 a_743_42282# a_20256_42852# 1.03e-20
C15917 a_17538_32519# a_22465_38105# 2e-19
C15918 a_n1741_47186# a_2747_46873# 0.00508f
C15919 a_6151_47436# a_16241_47178# 5.05e-20
C15920 a_2063_45854# a_13507_46334# 7.95e-20
C15921 a_n815_47178# a_n89_47570# 3.25e-20
C15922 a_n452_47436# a_n310_47570# 0.007833f
C15923 a_n971_45724# a_n2312_39304# 8.21e-21
C15924 a_11459_47204# a_13381_47204# 3.65e-21
C15925 a_9313_45822# a_n1435_47204# 5.93e-19
C15926 a_16112_44458# a_14539_43914# 0.13299f
C15927 a_1307_43914# a_1467_44172# 0.228571f
C15928 a_626_44172# a_n984_44318# 7.42e-19
C15929 a_11827_44484# a_14815_43914# 0.029578f
C15930 a_7499_43078# a_6031_43396# 7.11e-20
C15931 a_11691_44458# a_13213_44734# 0.046347f
C15932 a_n2661_44458# a_8855_44734# 3.59e-19
C15933 a_3537_45260# a_3499_42826# 0.001528f
C15934 a_8191_45002# a_7845_44172# 4.75e-20
C15935 a_n1059_45260# a_15682_43940# 0.001131f
C15936 a_n2017_45002# a_17737_43940# 1.87e-21
C15937 a_2382_45260# a_n2661_42282# 2.02e-19
C15938 a_5379_42460# a_n443_42852# 9.94e-21
C15939 a_6123_31319# a_n357_42282# 0.004292f
C15940 a_7227_42308# a_n755_45592# 3.68e-19
C15941 a_n2946_39866# a_n2956_39304# 0.004782f
C15942 a_n3420_39616# a_n2956_38680# 1.52e-19
C15943 a_11682_45822# VDD 0.316586f
C15944 a_1667_45002# a_n2293_46098# 3.65e-20
C15945 a_20447_31679# a_4185_45028# 1.09e-20
C15946 a_n1059_45260# a_1823_45246# 0.021319f
C15947 a_n913_45002# a_1138_42852# 0.032304f
C15948 a_8697_45822# a_8049_45260# 0.003995f
C15949 a_1176_45572# a_n357_42282# 4.74e-21
C15950 a_n2661_43922# a_8128_46384# 4.1e-21
C15951 a_18175_45572# a_18189_46348# 0.018402f
C15952 a_18479_45785# a_17715_44484# 9.75e-21
C15953 a_3357_43084# a_5164_46348# 7.34e-20
C15954 a_2437_43646# a_6165_46155# 3.75e-20
C15955 a_1467_44172# a_n443_46116# 0.031058f
C15956 a_20766_44850# a_18479_47436# 0.007835f
C15957 a_20679_44626# a_18597_46090# 0.025074f
C15958 a_21671_42860# a_21613_42308# 9.03e-20
C15959 a_n784_42308# a_2351_42308# 0.0035f
C15960 a_22165_42308# a_21887_42336# 0.110763f
C15961 a_1067_42314# a_1149_42558# 0.004937f
C15962 a_n473_42460# a_n39_42308# 0.003935f
C15963 a_n1630_35242# a_1221_42558# 2.09e-20
C15964 a_14097_32519# a_5932_42308# 0.001859f
C15965 a_10227_46804# a_15559_46634# 7.04e-19
C15966 a_11599_46634# a_12156_46660# 2.63e-20
C15967 a_4915_47217# a_14226_46660# 1.65e-19
C15968 a_12861_44030# a_12978_47026# 6.43e-21
C15969 a_4007_47204# a_765_45546# 0.00663f
C15970 a_3080_42308# a_3754_39964# 9.9e-20
C15971 a_4883_46098# a_11813_46116# 0.019696f
C15972 a_8128_46384# a_7927_46660# 0.007223f
C15973 a_5807_45002# a_5385_46902# 2.87e-19
C15974 a_n2293_46634# a_2959_46660# 1.76e-20
C15975 a_n133_46660# a_479_46660# 3.82e-19
C15976 a_n2661_46634# a_2864_46660# 0.002851f
C15977 a_383_46660# a_288_46660# 0.049827f
C15978 a_n1021_46688# a_n2661_46098# 3.91e-20
C15979 a_601_46902# a_491_47026# 0.097745f
C15980 a_948_46660# a_2107_46812# 1.97e-20
C15981 a_n743_46660# a_1799_45572# 0.034264f
C15982 a_n1925_46634# a_2443_46660# 0.054751f
C15983 a_1123_46634# a_1983_46706# 9.93e-19
C15984 a_18374_44850# a_14021_43940# 6.68e-21
C15985 a_22591_44484# a_17730_32519# 0.156987f
C15986 a_n2661_43922# a_9672_43914# 8.49e-20
C15987 a_n2661_42834# a_10405_44172# 0.005797f
C15988 a_9313_44734# a_18079_43940# 1.98e-20
C15989 a_19721_31679# a_17538_32519# 0.051191f
C15990 a_20512_43084# a_19237_31679# 1.14e-20
C15991 a_5883_43914# a_8415_44056# 6.67e-19
C15992 a_n913_45002# a_5649_42852# 0.0586f
C15993 en_comp a_13467_32519# 1.89e-19
C15994 a_3754_39134# VDD 0.004567f
C15995 a_22223_45036# VDD 0.300162f
C15996 a_n2661_43922# a_n1641_46494# 2.64e-22
C15997 a_5891_43370# a_4185_45028# 2.79e-19
C15998 a_18533_43940# a_13661_43548# 0.046643f
C15999 a_19319_43548# a_13747_46662# 2.08e-20
C16000 a_1423_45028# a_3218_45724# 2.67e-20
C16001 a_14797_45144# a_n443_42852# 5.7e-22
C16002 a_20567_45036# a_8049_45260# 3.41e-20
C16003 a_2903_45348# a_n755_45592# 1.85e-20
C16004 a_8685_43396# a_12861_44030# 0.007455f
C16005 a_n1613_43370# VDD 4.75085f
C16006 a_n784_42308# C4_N_btm 0.001073f
C16007 a_5167_46660# a_3483_46348# 1.48e-21
C16008 a_15368_46634# a_765_45546# 5.6e-19
C16009 a_15559_46634# a_17339_46660# 1.11e-20
C16010 a_3090_45724# a_18285_46348# 1.81e-20
C16011 a_20916_46384# a_22959_46124# 7.06e-20
C16012 a_9804_47204# a_5066_45546# 1.22e-21
C16013 a_n881_46662# a_8062_46482# 0.001601f
C16014 a_21588_30879# a_10809_44734# 0.110956f
C16015 a_3877_44458# a_5164_46348# 7.65e-19
C16016 a_4646_46812# a_5068_46348# 5.4e-20
C16017 a_4651_46660# a_4704_46090# 0.013135f
C16018 a_n743_46660# a_18189_46348# 1.08e-19
C16019 a_12465_44636# a_12839_46116# 4.88e-21
C16020 a_4883_46098# a_14949_46494# 2.19e-19
C16021 a_18597_46090# a_19431_46494# 0.004523f
C16022 a_16327_47482# a_20062_46116# 1.2e-19
C16023 a_4955_46873# a_4419_46090# 7.36e-20
C16024 a_10440_44484# a_10518_42984# 1.11e-21
C16025 a_20269_44172# a_19319_43548# 0.12985f
C16026 a_8975_43940# a_8952_43230# 2.23e-20
C16027 a_10057_43914# a_10083_42826# 0.001039f
C16028 a_9313_44734# a_14209_32519# 0.068114f
C16029 a_9895_44260# a_9801_43940# 1.26e-19
C16030 a_11341_43940# a_13565_43940# 0.00518f
C16031 a_19478_44306# a_19478_44056# 0.001278f
C16032 a_19328_44172# a_19741_43940# 0.04732f
C16033 a_n1059_45260# a_5934_30871# 0.010576f
C16034 a_n2017_45002# a_8515_42308# 0.002597f
C16035 a_n913_45002# a_7963_42308# 0.044607f
C16036 a_2382_45260# a_3497_42558# 0.001486f
C16037 a_2711_45572# a_n2017_45002# 0.02728f
C16038 a_2211_45572# a_2437_43646# 5.1e-19
C16039 a_21195_42852# a_12549_44172# 2.16e-19
C16040 a_4361_42308# a_5257_43370# 7.33e-20
C16041 a_17595_43084# a_13661_43548# 2.01e-20
C16042 a_n2840_43914# a_n2956_38216# 3.88e-19
C16043 a_9801_43940# a_8199_44636# 0.048015f
C16044 a_14021_43940# a_17715_44484# 3.95e-19
C16045 a_9165_43940# a_8953_45546# 9.62e-19
C16046 a_10651_43940# a_8016_46348# 1.82e-19
C16047 a_n4318_37592# a_n1151_42308# 4.12e-21
C16048 a_n784_42308# a_584_46384# 7.55e-22
C16049 a_13569_43230# a_10227_46804# 2.95e-19
C16050 a_n2293_46098# VDD 1.7963f
C16051 C1_P_btm C0_dummy_P_btm 1.24905f
C16052 a_19332_42282# CAL_N 0.001755f
C16053 a_13759_46122# a_14275_46494# 0.105995f
C16054 a_12005_46116# a_2324_44458# 9.1e-21
C16055 a_13925_46122# a_14493_46090# 0.17072f
C16056 a_8016_46348# a_6945_45028# 4.6e-20
C16057 a_n4315_30879# a_n4209_37414# 0.039099f
C16058 a_3090_45724# a_1609_45822# 3.9e-19
C16059 a_2202_46116# a_526_44458# 2.44e-20
C16060 a_167_45260# a_2981_46116# 4.98e-19
C16061 a_1823_45246# a_n1925_42282# 0.099018f
C16062 a_21076_30879# a_8049_45260# 6.53e-20
C16063 a_18451_43940# a_18249_42858# 2.07e-20
C16064 a_8685_43396# a_9803_43646# 0.008605f
C16065 a_3626_43646# a_16977_43638# 2.8e-21
C16066 a_2982_43646# a_17499_43370# 4.15e-20
C16067 a_14401_32519# a_22959_43396# 0.016242f
C16068 a_11341_43940# a_5534_30871# 6.54e-20
C16069 a_15493_43396# a_18083_42858# 6.8e-21
C16070 a_n2661_42834# a_6171_42473# 9.02e-22
C16071 a_5891_43370# a_9803_42558# 0.002774f
C16072 a_n356_44636# a_14456_42282# 2.77e-19
C16073 a_20974_43370# a_14209_32519# 0.049701f
C16074 a_3422_30871# a_22400_42852# 0.023064f
C16075 a_19721_31679# a_22465_38105# 3.17e-19
C16076 a_19787_47423# RST_Z 5.42e-20
C16077 SMPL_ON_N a_19864_35138# 0.01194f
C16078 a_19386_47436# START 0.042951f
C16079 a_11823_42460# a_15004_44636# 2.75e-20
C16080 a_18175_45572# a_18315_45260# 0.008723f
C16081 a_10193_42453# a_18443_44721# 8.46e-19
C16082 a_8696_44636# a_16981_45144# 0.003008f
C16083 a_15861_45028# a_16886_45144# 8.28e-19
C16084 a_6171_45002# a_10951_45334# 0.00438f
C16085 a_3232_43370# a_11787_45002# 0.001844f
C16086 a_n37_45144# a_375_42282# 7.33e-19
C16087 a_3357_43084# a_5837_45028# 0.006851f
C16088 a_7229_43940# a_7705_45326# 0.203098f
C16089 a_7276_45260# a_8191_45002# 3.64e-20
C16090 a_17595_43084# a_4185_45028# 1.06e-20
C16091 a_20712_42282# a_19321_45002# 2.03e-21
C16092 a_7287_43370# a_n443_42852# 0.010578f
C16093 a_13837_43396# a_13259_45724# 0.007401f
C16094 a_3935_42891# a_2324_44458# 6.13e-22
C16095 a_10835_43094# a_9290_44172# 0.172486f
C16096 a_n3607_39392# a_n2312_39304# 5.97e-20
C16097 a_15143_45578# a_n743_46660# 7.03e-21
C16098 a_6194_45824# a_5907_46634# 8.2e-20
C16099 a_5907_45546# a_5732_46660# 1.37e-19
C16100 a_16333_45814# a_12549_44172# 3.97e-22
C16101 a_15903_45785# a_15928_47570# 6.16e-21
C16102 a_3537_45260# a_n1151_42308# 4.52e-19
C16103 a_327_44734# a_n443_46116# 4.41e-19
C16104 a_7705_45326# a_n237_47217# 5.12e-19
C16105 a_8953_45002# a_n971_45724# 1.78e-20
C16106 a_4927_45028# a_2063_45854# 5.82e-19
C16107 a_413_45260# a_4915_47217# 7.6e-19
C16108 a_22223_45572# a_16327_47482# 2.78e-19
C16109 a_20528_45572# a_18597_46090# 0.03478f
C16110 a_2437_43646# a_16023_47582# 0.00865f
C16111 a_3357_43084# a_15673_47210# 3.29e-19
C16112 a_20623_45572# a_20894_47436# 2.94e-21
C16113 a_20107_45572# a_13507_46334# 1.59e-20
C16114 a_n2661_45546# a_n755_45592# 0.14317f
C16115 a_n863_45724# a_n452_45724# 0.046903f
C16116 a_n2293_45546# a_n1099_45572# 0.004814f
C16117 a_21115_43940# a_13258_32519# 1.2e-21
C16118 a_20623_43914# a_20712_42282# 1.64e-19
C16119 a_4361_42308# a_21671_42860# 0.012186f
C16120 a_7227_42852# a_7871_42858# 2.32e-20
C16121 a_5649_42852# a_20922_43172# 8.67e-21
C16122 a_13467_32519# a_22165_42308# 0.009474f
C16123 a_3080_42308# a_2351_42308# 1.79e-19
C16124 a_10341_43396# a_15785_43172# 5.75e-19
C16125 a_20107_46660# RST_Z 1.12e-20
C16126 a_765_45546# DATA[1] 0.009245f
C16127 a_n4209_37414# a_n3420_37440# 0.245806f
C16128 a_n4334_37440# a_n3690_37440# 8.67e-19
C16129 a_3905_42558# VDD 0.176395f
C16130 a_n237_47217# a_n785_47204# 0.018044f
C16131 a_n971_45724# a_1209_47178# 0.034982f
C16132 a_n1741_47186# a_2063_45854# 0.037801f
C16133 a_n2109_47186# a_2952_47436# 0.050821f
C16134 a_n746_45260# a_327_47204# 0.022743f
C16135 a_n452_47436# a_1239_47204# 7.81e-21
C16136 a_n2833_47464# a_n1151_42308# 2.4e-19
C16137 a_15599_45572# a_15682_43940# 4.45e-19
C16138 a_15415_45028# a_15433_44458# 9.2e-19
C16139 a_626_44172# a_n2661_43922# 0.03074f
C16140 a_8696_44636# a_10729_43914# 7.58e-20
C16141 a_13249_42308# a_14485_44260# 6.05e-19
C16142 a_n2661_43370# a_n1190_44850# 1.23e-19
C16143 a_21887_42336# a_4185_45028# 8e-20
C16144 a_8515_42308# a_526_44458# 3.38e-20
C16145 a_15597_42852# a_n357_42282# 0.009386f
C16146 a_5934_30871# a_n1925_42282# 3.98e-20
C16147 a_13157_43218# a_n443_42852# 4.11e-20
C16148 a_10341_43396# CLK 4.37e-20
C16149 a_20273_45572# a_20841_46902# 5.17e-21
C16150 a_16147_45260# a_11415_45002# 0.058206f
C16151 a_5009_45028# a_4651_46660# 6.47e-22
C16152 a_n2661_43370# a_2609_46660# 7.75e-21
C16153 a_20107_45572# a_20623_46660# 1.34e-20
C16154 a_14180_45002# a_6755_46942# 2.19e-22
C16155 a_2711_45572# a_526_44458# 0.392618f
C16156 a_3065_45002# a_3090_45724# 0.475346f
C16157 a_3357_43084# a_16388_46812# 5.22e-20
C16158 a_6171_45002# a_11735_46660# 1.67e-20
C16159 a_3232_43370# a_11813_46116# 6.78e-22
C16160 a_20623_45572# a_20411_46873# 6.29e-19
C16161 a_4223_44672# a_n881_46662# 1.75e-20
C16162 a_13904_45546# a_10903_43370# 0.081466f
C16163 a_13163_45724# a_12594_46348# 0.053634f
C16164 a_10490_45724# a_2324_44458# 0.015189f
C16165 a_11823_42460# a_13759_46122# 1.12e-19
C16166 a_9241_45822# a_5937_45572# 0.010703f
C16167 a_8697_45822# a_8953_45546# 0.006215f
C16168 a_10210_45822# a_8199_44636# 0.012124f
C16169 a_n699_43396# a_n1613_43370# 0.008801f
C16170 a_16112_44458# a_11453_44696# 8.57e-20
C16171 a_18287_44626# a_4883_46098# 1.92e-21
C16172 a_12545_42858# a_13070_42354# 5.71e-19
C16173 a_3080_42308# C4_N_btm 5.72e-19
C16174 a_12891_46348# a_5807_45002# 0.044188f
C16175 a_2747_46873# a_n743_46660# 1.24e-19
C16176 a_4915_47217# a_9863_46634# 8.01e-20
C16177 a_6151_47436# a_7927_46660# 0.182356f
C16178 a_n1435_47204# a_6540_46812# 2.44e-21
C16179 a_7227_47204# a_7411_46660# 0.011806f
C16180 a_6491_46660# a_7577_46660# 4.53e-20
C16181 a_n1741_47186# a_12469_46902# 4.21e-19
C16182 a_n1151_42308# a_6969_46634# 2.33e-19
C16183 a_2063_45854# a_7832_46660# 0.011867f
C16184 a_n237_47217# a_8601_46660# 1.58e-19
C16185 a_11691_44458# a_11341_43940# 4.94e-19
C16186 a_7499_43078# a_10796_42968# 0.030705f
C16187 a_20193_45348# a_21115_43940# 0.01963f
C16188 a_375_42282# a_104_43370# 0.001385f
C16189 a_2711_45572# a_19164_43230# 0.006484f
C16190 a_n356_44636# a_895_43940# 0.026898f
C16191 a_9313_44734# a_17730_32519# 3.13e-20
C16192 a_3537_45260# a_6197_43396# 0.337459f
C16193 a_n913_45002# a_8685_43396# 0.03156f
C16194 a_16019_45002# VDD 0.174085f
C16195 COMP_P RST_Z 0.034203f
C16196 a_14097_32519# VREF 2.43e-19
C16197 a_n784_42308# C6_P_btm 5.52e-19
C16198 a_22469_40625# a_21076_30879# 6.02e-20
C16199 a_n1177_44458# a_n1076_46494# 3.46e-22
C16200 a_n699_43396# a_n2293_46098# 0.001069f
C16201 a_n2661_44458# a_1138_42852# 0.026505f
C16202 a_15433_44458# a_15368_46634# 1.7e-19
C16203 a_15493_43396# a_12549_44172# 0.079226f
C16204 a_3499_42826# a_n2293_46634# 0.022726f
C16205 a_n2661_42282# a_n2956_39768# 6.98e-20
C16206 a_4185_45348# a_n1925_42282# 1.16e-20
C16207 a_n2661_45010# a_n1099_45572# 7.2e-21
C16208 a_n1059_45260# a_n2293_45546# 0.076047f
C16209 a_n2956_37592# a_n2810_45572# 0.048284f
C16210 a_15493_43940# a_n881_46662# 4.43e-21
C16211 a_14976_45348# a_2324_44458# 0.002969f
C16212 a_3080_42308# a_584_46384# 0.010326f
C16213 a_3626_43646# a_n971_45724# 4.16e-20
C16214 a_19741_43940# a_12861_44030# 2.77e-20
C16215 a_4791_45118# VDD 3.05095f
C16216 a_14113_42308# a_4958_30871# 0.058048f
C16217 a_15764_42576# a_15761_42308# 2.36e-20
C16218 a_n3674_37592# a_n4334_38528# 6.44e-20
C16219 a_5934_30871# a_n4315_30879# 8.24e-21
C16220 a_11453_44696# a_13925_46122# 3.96e-21
C16221 a_12465_44636# a_14840_46494# 2.12e-20
C16222 a_6545_47178# a_5066_45546# 0.021464f
C16223 a_4883_46098# a_15682_46116# 0.06363f
C16224 a_13507_46334# a_17715_44484# 0.003011f
C16225 a_18479_47436# a_19900_46494# 0.001423f
C16226 a_18597_46090# a_19335_46494# 0.036056f
C16227 a_10227_46804# a_21137_46414# 1.29e-19
C16228 a_19787_47423# a_18985_46122# 5.06e-20
C16229 a_19386_47436# a_19553_46090# 2.56e-20
C16230 a_16763_47508# a_10809_44734# 2.22e-19
C16231 a_17591_47464# a_6945_45028# 0.025004f
C16232 a_2063_45854# a_10586_45546# 0.056181f
C16233 a_n1151_42308# a_9241_46436# 5.09e-19
C16234 a_n881_46662# a_6419_46155# 0.019005f
C16235 a_2864_46660# a_765_45546# 8.25e-19
C16236 a_8270_45546# a_8601_46660# 8.69e-20
C16237 a_6755_46942# a_15009_46634# 0.012747f
C16238 a_n2956_39768# a_n2840_46090# 6.87e-19
C16239 a_12549_44172# a_3483_46348# 0.185475f
C16240 a_17737_43940# a_18079_43940# 0.001885f
C16241 a_14539_43914# a_17499_43370# 0.005043f
C16242 a_18114_32519# a_14209_32519# 0.054602f
C16243 a_5013_44260# a_5326_44056# 7.61e-19
C16244 a_17730_32519# a_20974_43370# 0.016457f
C16245 a_n1059_45260# a_16245_42852# 0.130348f
C16246 a_n913_45002# a_15953_42852# 1.61e-20
C16247 a_n2017_45002# a_16877_42852# 5.23e-19
C16248 a_19963_31679# a_22400_42852# 3.97e-20
C16249 a_11652_45724# a_11823_42460# 0.035142f
C16250 a_11962_45724# a_12427_45724# 0.064229f
C16251 a_10193_42453# a_13249_42308# 0.001874f
C16252 a_8162_45546# a_6977_45572# 1.1e-19
C16253 a_2711_45572# a_15297_45822# 1.6e-19
C16254 C0_dummy_N_btm EN_VIN_BSTR_N 0.026355f
C16255 a_12429_44172# a_3483_46348# 9.13e-22
C16256 a_20556_43646# a_19321_45002# 4.6e-19
C16257 a_4361_42308# a_5807_45002# 2.93e-22
C16258 a_n23_44458# a_n443_42852# 0.002324f
C16259 a_n310_44484# a_n863_45724# 1.13e-19
C16260 a_6453_43914# a_2324_44458# 0.010794f
C16261 a_5841_44260# a_5937_45572# 1.15e-20
C16262 a_n4318_38680# a_n1613_43370# 1.09e-19
C16263 a_9127_43156# a_4883_46098# 0.011077f
C16264 a_13113_42826# a_10227_46804# 0.159547f
C16265 a_8649_43218# a_n971_45724# 3.91e-20
C16266 a_413_45260# DATA[5] 0.0381f
C16267 a_16292_46812# VDD 0.123916f
C16268 a_1823_45246# a_2698_46116# 2.13e-21
C16269 a_15009_46634# a_8049_45260# 2.77e-21
C16270 a_11813_46116# a_11608_46482# 9.21e-19
C16271 a_3877_44458# a_3316_45546# 9.66e-20
C16272 a_11415_45002# a_9290_44172# 0.031886f
C16273 a_20411_46873# a_18819_46122# 2.15e-20
C16274 a_19551_46910# a_19553_46090# 2.94e-19
C16275 a_19123_46287# a_19335_46494# 3.12e-19
C16276 a_6123_31319# a_n4064_37440# 2.49e-19
C16277 a_5934_30871# a_n3420_37440# 7.32e-19
C16278 a_19862_44208# a_13467_32519# 2.46e-19
C16279 a_9313_44734# a_17749_42852# 6.88e-20
C16280 a_3422_30871# a_22223_42860# 0.002205f
C16281 a_20623_43914# a_20556_43646# 3.65e-19
C16282 a_11341_43940# a_4190_30871# 0.00376f
C16283 a_7845_44172# a_7765_42852# 1.24e-19
C16284 a_20512_43084# a_19987_42826# 0.11919f
C16285 a_14021_43940# a_16664_43396# 0.003073f
C16286 a_n97_42460# a_2437_43396# 1.3e-19
C16287 a_8791_43396# VDD 0.191045f
C16288 a_n2293_45010# a_n2109_45247# 0.068458f
C16289 a_n2661_45010# a_n1059_45260# 0.021417f
C16290 a_21513_45002# a_413_45260# 2.28e-21
C16291 a_n2472_45002# a_n2017_45002# 4.25e-20
C16292 a_10193_42453# a_17613_45144# 2.06e-20
C16293 a_8696_44636# a_1423_45028# 0.095059f
C16294 a_11823_42460# a_13490_45067# 6.19e-21
C16295 a_13467_32519# a_4185_45028# 0.033397f
C16296 a_3318_42354# a_n2293_46634# 2.67e-19
C16297 a_n4318_39304# a_n2956_38216# 0.023138f
C16298 a_19647_42308# a_16327_47482# 1.59e-19
C16299 a_13904_45546# a_4883_46098# 1.69e-20
C16300 a_10907_45822# a_10227_46804# 2.47e-19
C16301 a_14955_43396# a_5342_30871# 0.002466f
C16302 a_10341_43396# a_5534_30871# 2.97e-19
C16303 a_15095_43370# a_15567_42826# 0.167909f
C16304 a_13887_32519# a_14209_32519# 0.086073f
C16305 a_5649_42852# a_17364_32525# 6.86e-20
C16306 a_3457_43396# a_n2293_42282# 3.86e-19
C16307 a_3626_43646# a_3863_42891# 5.26e-19
C16308 a_n97_42460# a_15785_43172# 3.4e-19
C16309 a_n2946_37984# a_n4064_37984# 0.053263f
C16310 a_n3420_37984# a_n2302_37984# 2.4e-19
C16311 a_11787_45002# a_8975_43940# 4.91e-20
C16312 a_16147_45260# a_11967_42832# 6.48e-20
C16313 a_9482_43914# a_9838_44484# 0.175591f
C16314 a_1307_43914# a_4223_44672# 0.747516f
C16315 a_2711_45572# a_18079_43940# 0.006173f
C16316 a_3065_45002# a_n356_44636# 2.39e-19
C16317 a_n2661_45010# a_484_44484# 0.002755f
C16318 a_3357_43084# a_n2661_42834# 0.081135f
C16319 a_413_45260# a_700_44734# 3.75e-19
C16320 a_18214_42558# a_17339_46660# 8.1e-20
C16321 a_18083_42858# a_n357_42282# 0.026806f
C16322 a_3080_42308# C6_P_btm 2.67e-19
C16323 DATA[3] VDD 0.309692f
C16324 a_3175_45822# a_167_45260# 2.8e-19
C16325 a_5263_45724# a_1823_45246# 2e-20
C16326 a_5024_45822# a_n2293_46098# 0.001497f
C16327 a_13017_45260# a_n743_46660# 6.48e-21
C16328 a_13777_45326# a_n2293_46634# 1.56e-21
C16329 a_17478_45572# a_19466_46812# 2.38e-21
C16330 a_3357_43084# a_8145_46902# 2.87e-21
C16331 a_3429_45260# a_2959_46660# 5.07e-19
C16332 a_7229_43940# a_2107_46812# 4.89e-21
C16333 a_3065_45002# a_3699_46634# 8.84e-21
C16334 a_n2293_42834# a_n881_46662# 4.05e-20
C16335 a_n699_43396# a_4791_45118# 0.024838f
C16336 a_n1190_44850# a_n2497_47436# 1.37e-19
C16337 a_18545_45144# a_12861_44030# 1.5e-19
C16338 a_21005_45260# a_18479_47436# 0.015257f
C16339 a_18494_42460# a_18597_46090# 3.29e-19
C16340 a_11691_44458# a_16327_47482# 0.536141f
C16341 a_17719_45144# a_13507_46334# 8.16e-21
C16342 a_13807_45067# a_11453_44696# 2e-19
C16343 a_16547_43609# a_16522_42674# 4.2e-20
C16344 a_16243_43396# a_17124_42282# 1.48e-20
C16345 a_3681_42891# a_1755_42282# 1.9e-20
C16346 a_8952_43230# a_n784_42308# 1.44e-22
C16347 a_15743_43084# a_15890_42674# 0.001174f
C16348 a_18083_42858# a_18707_42852# 9.73e-19
C16349 a_5649_42852# a_8325_42308# 7.52e-20
C16350 a_4361_42308# a_9223_42460# 0.009506f
C16351 a_10341_43396# a_19647_42308# 2.22e-20
C16352 a_18817_42826# a_18861_43218# 3.69e-19
C16353 a_18249_42858# a_19273_43230# 2.36e-20
C16354 a_743_42282# a_10545_42558# 7.22e-19
C16355 a_20205_31679# a_22459_39145# 2.38e-20
C16356 a_20692_30879# a_22521_40055# 1.07e-20
C16357 a_n4334_38304# VDD 0.385989f
C16358 a_12861_44030# a_768_44030# 0.260776f
C16359 a_7903_47542# a_5807_45002# 1.29e-20
C16360 a_13487_47204# a_12549_44172# 0.036506f
C16361 a_13381_47204# a_13569_47204# 3.03e-20
C16362 SMPL_ON_N a_11453_44696# 0.147722f
C16363 a_22731_47423# a_22959_47212# 0.08444f
C16364 a_n1151_42308# a_n2293_46634# 0.02925f
C16365 a_n237_47217# a_2107_46812# 0.086093f
C16366 a_n2109_47186# a_n2661_46098# 3.71e-19
C16367 a_327_47204# a_383_46660# 0.001388f
C16368 a_584_46384# a_n2438_43548# 0.099362f
C16369 a_2063_45854# a_n743_46660# 1.58762f
C16370 a_3815_47204# a_n2661_46634# 9.75e-20
C16371 a_n971_45724# a_288_46660# 9.88e-20
C16372 a_5111_44636# a_5745_43940# 5.27e-19
C16373 a_5147_45002# a_5829_43940# 6.15e-19
C16374 a_3537_45260# a_8415_44056# 3.72e-19
C16375 a_17970_44736# a_16241_44734# 1.65e-20
C16376 a_16979_44734# a_17517_44484# 0.109784f
C16377 a_5891_43370# a_5708_44484# 4.97e-20
C16378 a_10193_42453# a_19700_43370# 7.43e-21
C16379 a_18114_32519# a_17730_32519# 9.1497f
C16380 a_1307_43914# a_15493_43940# 0.057588f
C16381 a_7640_43914# a_9159_44484# 8.4e-20
C16382 a_9482_43914# a_12603_44260# 0.002516f
C16383 a_n2293_42834# a_7911_44260# 0.00163f
C16384 a_5289_44734# a_n2661_43922# 1.98e-35
C16385 a_n4334_40480# a_n2956_38216# 6.67e-19
C16386 a_n2661_42834# a_3877_44458# 2.79e-19
C16387 a_6298_44484# a_3090_45724# 0.013998f
C16388 a_3422_30871# a_13747_46662# 1.93e-19
C16389 a_5891_43370# a_5257_43370# 0.001693f
C16390 a_20980_44850# a_19321_45002# 6.29e-21
C16391 a_16147_45260# a_13259_45724# 0.033344f
C16392 a_3357_43084# a_5066_45546# 0.033559f
C16393 a_20528_45572# a_8049_45260# 0.004485f
C16394 a_10951_45334# a_10903_43370# 0.005295f
C16395 a_11787_45002# a_11387_46155# 3.57e-19
C16396 a_6171_45002# a_2324_44458# 2.73828f
C16397 a_413_45260# a_10809_44734# 0.333257f
C16398 a_13483_43940# a_12861_44030# 1.39e-19
C16399 a_7963_42308# a_8325_42308# 0.002341f
C16400 a_6123_31319# a_8685_42308# 1.64e-19
C16401 EN_VIN_BSTR_N a_21589_35634# 2.66e-19
C16402 a_18194_35068# a_19864_35138# 0.045378f
C16403 EN_VIN_BSTR_P C8_P_btm 0.090252f
C16404 a_4646_46812# a_7577_46660# 0.002516f
C16405 a_2107_46812# a_8270_45546# 0.047835f
C16406 a_12549_44172# a_14513_46634# 0.008065f
C16407 a_768_44030# a_14180_46812# 0.009222f
C16408 a_19321_45002# a_19692_46634# 0.040279f
C16409 a_19594_46812# a_19466_46812# 0.100902f
C16410 a_4817_46660# a_5257_43370# 4.13e-19
C16411 a_5167_46660# a_5263_46660# 0.013793f
C16412 a_5385_46902# a_5429_46660# 3.69e-19
C16413 a_3877_44458# a_8145_46902# 1.22e-20
C16414 a_13507_46334# a_22365_46825# 0.033904f
C16415 a_n1435_47204# a_1823_45246# 1.9e-20
C16416 a_4915_47217# a_6165_46155# 3.17e-20
C16417 a_6151_47436# a_5164_46348# 5.71e-20
C16418 a_n1151_42308# a_9625_46129# 0.046431f
C16419 a_4791_45118# a_7920_46348# 1.09e-19
C16420 a_2063_45854# a_11189_46129# 0.294233f
C16421 a_6298_44484# a_6547_43396# 0.002809f
C16422 a_n23_44458# a_n229_43646# 8.22e-20
C16423 a_18579_44172# a_15493_43940# 0.377126f
C16424 a_n356_44636# a_458_43396# 0.001988f
C16425 a_5883_43914# a_6293_42852# 4.78e-19
C16426 a_5343_44458# a_7112_43396# 1.78e-21
C16427 a_375_42282# a_n1076_43230# 1.84e-20
C16428 a_n4318_39768# a_n3674_39768# 3.06574f
C16429 a_2675_43914# a_3499_42826# 0.010775f
C16430 a_2998_44172# a_2253_44260# 2.04e-20
C16431 a_n2661_44458# a_8685_43396# 3.35e-20
C16432 a_11691_44458# a_10341_43396# 1.54e-19
C16433 a_13249_42308# a_n784_42308# 1.26e-20
C16434 a_3232_43370# a_9127_43156# 4.38e-21
C16435 a_3357_43084# a_n2293_42282# 0.146926f
C16436 a_n1059_45260# a_18249_42858# 0.002769f
C16437 a_n913_45002# a_17333_42852# 2.15e-20
C16438 a_n2017_45002# a_18817_42826# 0.018518f
C16439 a_n1243_44484# VDD 7.26e-20
C16440 a_n4209_39590# VREF_GND 0.083908f
C16441 a_n3420_39072# C5_P_btm 0.001006f
C16442 a_n4064_39072# C7_P_btm 0.072179f
C16443 a_n3565_39304# C3_P_btm 3.19e-20
C16444 a_2711_45572# a_4099_45572# 0.176427f
C16445 a_n2946_37690# a_n2956_38216# 0.004064f
C16446 a_22315_44484# a_4185_45028# 0.002812f
C16447 a_11341_43940# a_15227_44166# 0.04747f
C16448 a_10555_44260# a_3090_45724# 0.041801f
C16449 a_20623_43914# a_19692_46634# 0.007357f
C16450 a_6197_43396# a_n2293_46634# 0.05355f
C16451 a_9803_43646# a_768_44030# 5.37e-20
C16452 a_n2433_44484# a_n2472_45546# 3.17e-20
C16453 a_n2661_44458# a_n2956_38216# 0.009784f
C16454 a_n2293_43922# a_n2956_39304# 4.52e-20
C16455 a_14673_44172# a_2324_44458# 0.015622f
C16456 a_11967_42832# a_9290_44172# 0.0995f
C16457 a_8037_42858# a_n971_45724# 7.81e-19
C16458 a_13678_32519# a_12861_44030# 6.9e-20
C16459 a_4190_30871# a_16327_47482# 0.335014f
C16460 a_17499_43370# a_11453_44696# 8.56e-21
C16461 a_19479_31679# a_22459_39145# 1.76e-20
C16462 a_n3565_39304# a_n4064_38528# 0.029566f
C16463 a_n3420_39072# a_n3420_38528# 0.127439f
C16464 a_n4064_39072# a_n3565_38502# 0.030685f
C16465 a_3090_45724# a_5937_45572# 0.002157f
C16466 a_10428_46928# a_6945_45028# 8.06e-21
C16467 a_11735_46660# a_10903_43370# 0.002577f
C16468 a_11813_46116# a_11387_46155# 0.080527f
C16469 a_n881_46662# a_n310_45899# 5.94e-19
C16470 a_20916_46384# a_20850_46482# 4.71e-19
C16471 a_4955_46873# a_4365_46436# 7.84e-21
C16472 a_n743_46660# a_14383_46116# 0.00314f
C16473 a_12549_44172# a_n357_42282# 1.1e-19
C16474 a_3877_44458# a_5066_45546# 6.79e-20
C16475 a_20841_46902# a_20202_43084# 3.14e-20
C16476 a_19551_46910# a_12741_44636# 2.24e-19
C16477 a_20273_46660# a_11415_45002# 2.53e-20
C16478 a_20107_46660# a_20820_30879# 2.92e-20
C16479 en_comp a_21335_42336# 2.22e-20
C16480 a_22591_44484# a_22591_43396# 2.73e-20
C16481 a_22485_44484# a_14209_32519# 4.86e-19
C16482 a_14955_43940# a_9145_43396# 1.77e-19
C16483 a_13857_44734# a_13635_43156# 2.1e-21
C16484 a_9313_44734# a_19339_43156# 0.01152f
C16485 a_13565_43940# a_n97_42460# 1.86e-21
C16486 a_17730_32519# a_13887_32519# 0.053953f
C16487 a_n2293_43922# a_5534_30871# 0.271171f
C16488 a_20974_43370# a_17538_32519# 0.001842f
C16489 a_1307_43914# a_5742_30871# 2.36e-20
C16490 a_10651_43940# VDD 0.003431f
C16491 a_10193_42453# a_11787_45002# 0.0195f
C16492 a_7227_45028# a_1423_45028# 0.009712f
C16493 a_18175_45572# a_20107_45572# 4.32e-19
C16494 a_10490_45724# a_10775_45002# 1.62e-19
C16495 a_8746_45002# a_10951_45334# 7.44e-20
C16496 a_18909_45814# a_19418_45938# 2.6e-19
C16497 a_18341_45572# a_18787_45572# 2.28e-19
C16498 a_18479_45785# a_18953_45572# 0.002424f
C16499 a_2711_45572# a_5365_45348# 3.34e-19
C16500 a_13527_45546# a_6171_45002# 3.83e-20
C16501 a_7871_42858# a_8270_45546# 8.9e-21
C16502 a_16823_43084# a_17339_46660# 7.42e-19
C16503 a_18695_43230# a_13661_43548# 2.15e-19
C16504 a_12429_44172# a_n357_42282# 5.79e-21
C16505 a_6547_43396# a_5937_45572# 6.63e-19
C16506 a_n1630_35242# a_n2312_40392# 0.033733f
C16507 a_6945_45028# VDD 1.30257f
C16508 a_10053_45546# a_2063_45854# 1.55e-19
C16509 a_5024_45822# a_4791_45118# 1.87e-20
C16510 a_6472_45840# a_6575_47204# 6.84e-21
C16511 a_6598_45938# a_6851_47204# 1.17e-21
C16512 a_3483_46348# a_n2661_45546# 0.163728f
C16513 a_472_46348# a_997_45618# 6.4e-19
C16514 a_167_45260# a_n863_45724# 0.424358f
C16515 a_n1853_46287# a_n23_45546# 7.5e-20
C16516 a_1138_42852# a_n1099_45572# 3.41e-20
C16517 a_n2293_46098# a_7_45899# 3.19e-19
C16518 a_19335_46494# a_8049_45260# 0.001373f
C16519 a_13925_46122# a_14180_46482# 0.056391f
C16520 a_9290_44172# a_13259_45724# 0.272297f
C16521 a_12005_46116# a_12839_46116# 6e-19
C16522 a_13759_46122# a_14371_46494# 3.82e-19
C16523 a_n4064_37984# C1_P_btm 8.65e-20
C16524 a_14955_43396# a_743_42282# 3.11e-20
C16525 a_17499_43370# a_17324_43396# 0.234322f
C16526 a_16547_43609# a_15743_43084# 0.028834f
C16527 a_10341_43396# a_4190_30871# 0.090771f
C16528 a_3539_42460# a_3935_42891# 2.26e-20
C16529 a_3626_43646# a_4520_42826# 4.31e-20
C16530 a_2982_43646# a_5755_42852# 1.01e-20
C16531 a_n97_42460# a_5534_30871# 0.109695f
C16532 a_21381_43940# a_19987_42826# 1.97e-19
C16533 a_9313_44734# a_22465_38105# 0.002447f
C16534 a_n2661_42282# a_n2472_42282# 0.028691f
C16535 a_2889_44172# a_2903_42308# 3.69e-22
C16536 a_11967_42832# a_15051_42282# 1.9e-19
C16537 a_11341_43940# a_14635_42282# 4.84e-20
C16538 a_n2661_46634# DATA[0] 0.012107f
C16539 a_12895_43230# VDD 0.212352f
C16540 a_413_45260# a_22959_45036# 0.024709f
C16541 a_6171_45002# a_16922_45042# 0.00895f
C16542 a_2437_43646# a_949_44458# 0.038046f
C16543 a_n2840_45002# a_n2661_44458# 0.003602f
C16544 a_n2661_45010# a_n4318_40392# 8.18e-22
C16545 a_18909_45814# a_18248_44752# 1.74e-19
C16546 a_18479_45785# a_18443_44721# 7.52e-19
C16547 a_18175_45572# a_18374_44850# 3.73e-19
C16548 a_18341_45572# a_18287_44626# 3.7e-20
C16549 a_9482_43914# a_n2661_43370# 2.58e-19
C16550 a_1307_43914# a_n2293_42834# 0.089964f
C16551 a_2304_45348# a_2448_45028# 6.84e-19
C16552 a_13017_45260# a_13490_45394# 2.62e-19
C16553 a_10193_42453# a_17325_44484# 1.97e-19
C16554 COMP_P a_20820_30879# 8.52e-20
C16555 a_n2302_38778# a_n2312_38680# 0.161815f
C16556 a_4361_42308# a_n755_45592# 0.035265f
C16557 a_10193_42453# a_11813_46116# 0.02832f
C16558 a_10907_45822# a_10467_46802# 4.68e-20
C16559 a_10210_45822# a_10623_46897# 3.91e-20
C16560 a_5437_45600# a_3090_45724# 5.24e-20
C16561 a_3357_43084# a_19321_45002# 0.030763f
C16562 a_n913_45002# a_768_44030# 2.6e-19
C16563 a_21513_45002# a_20916_46384# 1.63e-20
C16564 a_413_45260# a_n881_46662# 0.026808f
C16565 a_327_44734# a_n1613_43370# 3.68e-20
C16566 a_10951_45334# a_4883_46098# 2.01e-20
C16567 a_15415_45028# a_10227_46804# 0.001754f
C16568 a_n2293_42834# a_n443_46116# 9.36e-19
C16569 a_5755_42852# a_5837_42852# 0.171361f
C16570 a_8387_43230# a_8292_43218# 0.049827f
C16571 a_8605_42826# a_8483_43230# 3.16e-19
C16572 a_18817_42826# a_19164_43230# 0.051162f
C16573 a_8685_43396# a_8325_42308# 3.75e-20
C16574 a_n97_42460# a_19647_42308# 6.61e-19
C16575 a_n1741_47186# a_2487_47570# 2.13e-19
C16576 a_n815_47178# a_n310_47570# 9.52e-19
C16577 a_11031_47542# a_n1435_47204# 2.39e-19
C16578 a_6151_47436# a_15673_47210# 0.002744f
C16579 a_15004_44636# a_14539_43914# 0.001002f
C16580 a_375_42282# a_175_44278# 0.017991f
C16581 a_626_44172# a_n809_44244# 1.91e-19
C16582 a_1307_43914# a_1115_44172# 0.115939f
C16583 a_11691_44458# a_n2293_43922# 0.02314f
C16584 a_n2661_44458# a_8783_44734# 1.49e-19
C16585 a_n913_45002# a_13483_43940# 9.64e-21
C16586 a_n1059_45260# a_14955_43940# 8.05e-22
C16587 a_n2017_45002# a_15682_43940# 2.7e-20
C16588 a_5267_42460# a_n443_42852# 7.84e-22
C16589 a_6761_42308# a_n755_45592# 2.19e-19
C16590 a_7227_42308# a_n357_42282# 7.15e-20
C16591 a_n3420_39616# a_n2956_39304# 9.34e-19
C16592 a_11280_45822# VDD 0.004437f
C16593 a_327_44734# a_n2293_46098# 1.74e-19
C16594 a_22959_45572# a_4185_45028# 3.35e-19
C16595 a_556_44484# a_768_44030# 0.001175f
C16596 a_n1059_45260# a_1138_42852# 0.004009f
C16597 a_n2017_45002# a_1823_45246# 0.024027f
C16598 a_n967_45348# a_n1076_46494# 4.41e-20
C16599 a_9159_45572# a_5066_45546# 0.040307f
C16600 a_11823_42460# a_12379_46436# 4.72e-19
C16601 a_1260_45572# a_n1099_45572# 5.75e-20
C16602 a_8336_45822# a_8049_45260# 4e-19
C16603 a_16147_45260# a_18189_46348# 0.129202f
C16604 a_12561_45572# a_10809_44734# 1.38e-19
C16605 a_1115_44172# a_n443_46116# 6.13e-20
C16606 a_5013_44260# a_584_46384# 1.69e-19
C16607 a_18753_44484# a_16327_47482# 7.32e-19
C16608 a_20835_44721# a_18479_47436# 0.007754f
C16609 a_20640_44752# a_18597_46090# 0.027095f
C16610 a_18204_44850# a_11453_44696# 1.39e-19
C16611 a_21195_42852# a_21613_42308# 7.21e-19
C16612 a_21671_42860# a_21887_42336# 1.89e-21
C16613 a_1576_42282# a_1184_42692# 0.033078f
C16614 a_1067_42314# a_961_42354# 0.13675f
C16615 a_n784_42308# a_2123_42473# 0.216332f
C16616 a_n4318_38680# a_n4334_38304# 3.4e-19
C16617 a_n473_42460# a_n327_42308# 0.013377f
C16618 a_n1630_35242# a_1149_42558# 2.88e-20
C16619 a_4883_46098# a_11735_46660# 2.67e-19
C16620 a_16327_47482# a_15227_44166# 0.239667f
C16621 a_10227_46804# a_15368_46634# 0.003141f
C16622 a_18479_47436# a_3090_45724# 1.24e-20
C16623 a_3815_47204# a_765_45546# 0.003873f
C16624 a_n881_46662# a_9863_46634# 0.001329f
C16625 a_8128_46384# a_8145_46902# 0.012246f
C16626 a_n2293_46634# a_3177_46902# 1.62e-20
C16627 a_n743_46660# a_645_46660# 0.002128f
C16628 a_33_46660# a_491_47026# 0.027606f
C16629 a_n1925_46634# a_n2661_46098# 0.059432f
C16630 a_1123_46634# a_2107_46812# 0.002783f
C16631 a_n2661_46634# a_3524_46660# 0.0105f
C16632 a_5807_45002# a_4817_46660# 2.58e-19
C16633 a_n1059_45260# a_5649_42852# 0.030637f
C16634 a_n913_45002# a_13678_32519# 0.023168f
C16635 a_6171_45002# a_15743_43084# 1.19e-20
C16636 a_n2661_43922# a_9028_43914# 3.15e-20
C16637 a_22485_44484# a_17730_32519# 0.091577f
C16638 a_n2661_42834# a_9672_43914# 0.009389f
C16639 a_n2661_43370# a_6031_43396# 4.62e-21
C16640 a_18114_32519# a_17538_32519# 0.052981f
C16641 a_5883_43914# a_7499_43940# 0.04798f
C16642 a_11691_44458# a_n97_42460# 1.21e-19
C16643 a_1307_43914# a_10849_43646# 9.39e-19
C16644 a_7754_39300# VDD 0.048307f
C16645 a_11827_44484# VDD 0.615802f
C16646 a_13258_32519# a_22459_39145# 2.2e-19
C16647 a_19319_43548# a_13661_43548# 0.189089f
C16648 a_1423_45028# a_2957_45546# 1.39e-20
C16649 a_18494_42460# a_8049_45260# 1.4e-19
C16650 a_14537_43396# a_n443_42852# 0.03432f
C16651 a_2809_45348# a_n755_45592# 7.33e-20
C16652 a_13105_45348# a_13259_45724# 1.66e-19
C16653 a_12607_44458# a_2324_44458# 4.05e-20
C16654 a_n1809_43762# a_n1613_43370# 0.012235f
C16655 a_n1557_42282# a_n2312_39304# 1.92e-20
C16656 a_3411_47243# VDD 2.18e-20
C16657 a_7174_31319# a_n4209_39590# 8.87e-22
C16658 a_n784_42308# C3_N_btm 0.001962f
C16659 a_3633_46660# a_1823_45246# 6.58e-20
C16660 a_3090_45724# a_17829_46910# 1.43e-19
C16661 a_14976_45028# a_765_45546# 3.1e-19
C16662 a_8128_46384# a_5066_45546# 0.032968f
C16663 a_21588_30879# a_22223_46124# 1.77e-19
C16664 a_20916_46384# a_10809_44734# 0.038071f
C16665 a_3877_44458# a_5068_46348# 1.58e-19
C16666 a_4646_46812# a_4704_46090# 0.01107f
C16667 a_n743_46660# a_17715_44484# 0.01357f
C16668 a_13507_46334# a_15194_46482# 2.67e-19
C16669 a_4883_46098# a_14537_46482# 1.2e-19
C16670 a_18597_46090# a_19240_46482# 0.025784f
C16671 a_n1435_47204# a_n2293_45546# 1.57e-19
C16672 a_n1151_42308# a_2277_45546# 1.18e-22
C16673 a_2905_45572# a_2307_45899# 9.36e-20
C16674 a_584_46384# a_603_45572# 3.31e-19
C16675 a_10440_44484# a_10083_42826# 9.38e-21
C16676 a_10334_44484# a_10518_42984# 1.38e-22
C16677 a_19862_44208# a_19319_43548# 0.049274f
C16678 a_19478_44306# a_18533_43940# 3.55e-20
C16679 a_9313_44734# a_22591_43396# 0.001502f
C16680 a_8975_43940# a_9127_43156# 8.61e-21
C16681 a_n2661_42834# a_743_42282# 1.34e-20
C16682 a_9801_44260# a_9801_43940# 6.96e-20
C16683 a_11341_43940# a_11257_43940# 2.31e-19
C16684 a_15493_43396# a_19478_44056# 3.41e-19
C16685 a_3232_43370# a_1755_42282# 1.63e-20
C16686 a_3065_45002# a_3823_42558# 0.198186f
C16687 a_n913_45002# a_6123_31319# 0.21316f
C16688 a_n1059_45260# a_7963_42308# 5.71e-20
C16689 a_n2017_45002# a_5934_30871# 0.007182f
C16690 a_15037_45618# a_15225_45822# 7.47e-21
C16691 a_10341_43396# a_15227_44166# 0.068268f
C16692 a_21356_42826# a_12549_44172# 2.29e-20
C16693 a_10555_43940# a_8016_46348# 3.45e-19
C16694 a_9165_43940# a_5937_45572# 1.38e-20
C16695 a_n1736_42282# a_n1151_42308# 1.63e-20
C16696 a_15597_42852# a_12861_44030# 5.41e-19
C16697 a_11136_42852# a_10227_46804# 0.012196f
C16698 a_n2472_46090# VDD 0.224658f
C16699 C1_P_btm C0_P_btm 11.2332f
C16700 a_18907_42674# CAL_N 7.78e-19
C16701 a_13759_46122# a_14493_46090# 0.053479f
C16702 a_10903_43370# a_2324_44458# 0.038342f
C16703 a_1343_38525# VDAC_Pi 0.035744f
C16704 a_765_45546# a_18051_46116# 0.006713f
C16705 a_3090_45724# a_n443_42852# 0.269331f
C16706 a_19123_46287# a_19240_46482# 0.157972f
C16707 a_22959_46660# a_8049_45260# 2.87e-20
C16708 a_1138_42852# a_n1925_42282# 1.19e-20
C16709 a_472_46348# a_1337_46116# 2.04e-19
C16710 a_1823_45246# a_526_44458# 1.93329f
C16711 a_19386_47436# RST_Z 6.35e-20
C16712 a_18597_46090# START 0.020125f
C16713 a_7542_44172# a_7309_42852# 6.74e-21
C16714 a_18326_43940# a_18249_42858# 8.19e-22
C16715 a_8685_43396# a_9145_43396# 0.201058f
C16716 a_3626_43646# a_16409_43396# 3.02e-21
C16717 a_2982_43646# a_16759_43396# 7.55e-21
C16718 a_20974_43370# a_22591_43396# 0.046632f
C16719 a_11341_43940# a_14543_43071# 8.65e-21
C16720 a_15493_43396# a_17701_42308# 4.48e-20
C16721 a_18451_43940# a_17333_42852# 4.67e-20
C16722 a_3737_43940# a_3681_42891# 2.18e-20
C16723 a_n97_42460# a_4190_30871# 0.140814f
C16724 a_n2661_42834# a_5755_42308# 1.09e-20
C16725 a_5891_43370# a_9223_42460# 0.13879f
C16726 a_n356_44636# a_13575_42558# 1.46e-19
C16727 a_14401_32519# a_14209_32519# 10.7535f
C16728 a_17538_32519# a_13887_32519# 0.051087f
C16729 a_3422_30871# a_20836_43172# 2.5e-20
C16730 a_18114_32519# a_22465_38105# 2.37e-19
C16731 a_13527_45546# a_12607_44458# 8.08e-22
C16732 a_11823_42460# a_13720_44458# 7.98e-20
C16733 a_18909_45814# a_16922_45042# 3.62e-20
C16734 a_10193_42453# a_18287_44626# 5.37e-19
C16735 a_8696_44636# a_16886_45144# 0.00316f
C16736 a_15861_45028# a_16237_45028# 0.062212f
C16737 a_16147_45260# a_18315_45260# 4.61e-19
C16738 a_6171_45002# a_10775_45002# 0.008718f
C16739 a_3232_43370# a_10951_45334# 5.7e-20
C16740 a_413_45260# a_1307_43914# 0.080885f
C16741 a_7229_43940# a_6709_45028# 0.136786f
C16742 a_5205_44484# a_8191_45002# 2.44e-20
C16743 a_16795_42852# a_4185_45028# 4.48e-21
C16744 a_6547_43396# a_n443_42852# 0.006641f
C16745 a_13749_43396# a_13259_45724# 0.002234f
C16746 a_5649_42852# a_n1925_42282# 0.001675f
C16747 a_3681_42891# a_2324_44458# 9.45e-22
C16748 a_10518_42984# a_9290_44172# 0.04331f
C16749 a_10341_42308# a_8953_45546# 0.006033f
C16750 a_413_45260# a_n443_46116# 0.369976f
C16751 a_3537_45260# a_3160_47472# 1.25e-21
C16752 a_5111_44636# a_2063_45854# 0.004291f
C16753 a_8191_45002# a_n971_45724# 0.015833f
C16754 a_14495_45572# a_n743_46660# 6.59e-20
C16755 a_7227_45028# a_4646_46812# 0.305597f
C16756 a_3775_45552# a_3877_44458# 0.002726f
C16757 a_15765_45572# a_12549_44172# 3.88e-21
C16758 a_21188_45572# a_18597_46090# 0.00956f
C16759 a_20731_45938# a_18479_47436# 0.007339f
C16760 a_2437_43646# a_16327_47482# 0.046662f
C16761 a_3357_43084# a_15811_47375# 2.81e-19
C16762 a_20841_45814# a_20894_47436# 3.24e-21
C16763 a_n2661_45546# a_n357_42282# 0.044767f
C16764 a_n2293_45546# a_380_45546# 4.68e-20
C16765 a_n1079_45724# a_n452_45724# 6.61e-19
C16766 a_n2956_38216# a_n1099_45572# 3.28e-19
C16767 a_20269_44172# a_7174_31319# 7.85e-21
C16768 a_4905_42826# a_1755_42282# 1.01e-19
C16769 a_4361_42308# a_21195_42852# 0.020952f
C16770 a_5649_42852# a_19987_42826# 3.08e-20
C16771 a_13467_32519# a_21671_42860# 0.015185f
C16772 a_743_42282# a_n2293_42282# 0.058933f
C16773 a_11341_43940# a_19511_42282# 3.14e-21
C16774 a_3080_42308# a_2123_42473# 3.08e-20
C16775 a_10341_43396# a_14635_42282# 1.31e-19
C16776 a_19862_44208# a_21335_42336# 6.38e-20
C16777 a_21076_30879# a_22609_38406# 5.77e-21
C16778 a_19123_46287# START 0.003458f
C16779 a_765_45546# DATA[0] 6.38e-19
C16780 a_n4334_37440# a_n3565_37414# 0.001292f
C16781 a_n4209_37414# a_n3690_37440# 0.046103f
C16782 a_3581_42558# VDD 0.006789f
C16783 a_n237_47217# a_n23_47502# 0.056864f
C16784 a_n746_45260# a_n785_47204# 0.198992f
C16785 a_n971_45724# a_327_47204# 0.075444f
C16786 a_n1741_47186# a_584_46384# 0.021978f
C16787 a_n2109_47186# a_2553_47502# 0.04572f
C16788 a_n2017_45002# a_20512_43084# 4.16e-19
C16789 en_comp a_3422_30871# 0.357746f
C16790 a_1423_45028# a_9159_44484# 0.037664f
C16791 a_13249_42308# a_14021_43940# 0.07296f
C16792 a_626_44172# a_n2661_42834# 0.032386f
C16793 a_8696_44636# a_10405_44172# 2.24e-20
C16794 a_375_42282# a_n2293_43922# 3e-19
C16795 a_18114_32519# a_19721_31679# 0.051894f
C16796 a_14537_43396# a_15146_44811# 8.25e-19
C16797 a_n2661_43370# a_n1809_44850# 0.002228f
C16798 a_21335_42336# a_4185_45028# 8e-20
C16799 a_5934_30871# a_526_44458# 3.53e-19
C16800 a_14097_32519# a_20692_30879# 0.051423f
C16801 a_12991_43230# a_n443_42852# 1.9e-19
C16802 a_14853_42852# a_n357_42282# 5.87e-19
C16803 a_20273_45572# a_20273_46660# 4.74e-19
C16804 a_11136_45572# a_3483_46348# 0.020129f
C16805 a_n2661_44458# a_768_44030# 0.028401f
C16806 a_n2661_43370# a_2443_46660# 1.76e-21
C16807 a_13777_45326# a_6755_46942# 1.05e-21
C16808 a_2680_45002# a_3090_45724# 0.003269f
C16809 a_20623_45572# a_20107_46660# 2.63e-20
C16810 a_3357_43084# a_13059_46348# 1.83e-20
C16811 a_2779_44458# a_n881_46662# 3.56e-21
C16812 a_13527_45546# a_10903_43370# 0.035694f
C16813 a_12791_45546# a_12594_46348# 0.026771f
C16814 a_8746_45002# a_2324_44458# 0.34917f
C16815 a_10193_42453# a_15682_46116# 7.91e-19
C16816 a_11823_42460# a_13351_46090# 1.2e-19
C16817 a_8697_45822# a_5937_45572# 0.019555f
C16818 a_9241_45822# a_8199_44636# 1.53e-20
C16819 a_10907_45822# a_8016_46348# 1.99e-20
C16820 a_4223_44672# a_n1613_43370# 0.022154f
C16821 a_15004_44636# a_11453_44696# 3.53e-21
C16822 a_18248_44752# a_4883_46098# 1.47e-21
C16823 a_12379_42858# a_13575_42558# 1.06e-19
C16824 a_12545_42858# a_12563_42308# 1.83e-19
C16825 a_12089_42308# a_13070_42354# 9.69e-20
C16826 a_4190_30871# a_n3420_39616# 1.16e-20
C16827 a_13887_32519# a_22465_38105# 0.005089f
C16828 a_3080_42308# C3_N_btm 0.027071f
C16829 a_11309_47204# a_5807_45002# 0.032739f
C16830 a_6491_46660# a_7715_46873# 1.43e-20
C16831 a_6151_47436# a_8145_46902# 0.178565f
C16832 a_n1435_47204# a_5732_46660# 1.28e-20
C16833 a_6545_47178# a_7577_46660# 3.97e-20
C16834 a_n1741_47186# a_11901_46660# 0.034005f
C16835 a_n1151_42308# a_6755_46942# 0.142929f
C16836 a_n971_45724# a_8846_46660# 5.95e-19
C16837 a_17613_45144# a_14021_43940# 4.87e-21
C16838 a_7499_43078# a_10835_43094# 0.028158f
C16839 a_20193_45348# a_20935_43940# 0.016238f
C16840 a_n356_44636# a_2479_44172# 8.76e-21
C16841 a_18479_45785# a_19700_43370# 0.004581f
C16842 a_375_42282# a_n97_42460# 0.039466f
C16843 a_2711_45572# a_19339_43156# 0.020184f
C16844 a_16241_44734# a_16335_44484# 1.26e-19
C16845 a_3537_45260# a_6293_42852# 0.01772f
C16846 a_n1059_45260# a_8685_43396# 0.036086f
C16847 a_15595_45028# VDD 0.156299f
C16848 a_14097_32519# VIN_N 0.053964f
C16849 a_1606_42308# EN_VIN_BSTR_P 0.035204f
C16850 a_n784_42308# C7_P_btm 0.002308f
C16851 a_n1630_35242# a_21589_35634# 0.015148f
C16852 a_22521_40599# a_21076_30879# 7.82e-20
C16853 a_n2661_44458# a_1176_45822# 8.11e-22
C16854 a_n1352_44484# a_n1641_46494# 2.48e-20
C16855 a_4223_44672# a_n2293_46098# 0.422068f
C16856 a_19328_44172# a_12549_44172# 0.012953f
C16857 a_15146_44811# a_3090_45724# 1.56e-19
C16858 a_13777_45326# a_8049_45260# 4.46e-20
C16859 a_n2661_45010# a_380_45546# 3.48e-21
C16860 a_n745_45366# a_n2661_45546# 0.00237f
C16861 a_n2017_45002# a_n2293_45546# 1.75e-19
C16862 a_n2293_45010# a_n863_45724# 0.090522f
C16863 a_n2810_45028# a_n2810_45572# 0.063288f
C16864 a_4699_43561# a_584_46384# 7.44e-19
C16865 a_21205_44306# a_12861_44030# 3.21e-19
C16866 a_14403_45348# a_2324_44458# 0.0023f
C16867 a_14309_45028# a_13759_46122# 1.57e-20
C16868 a_4700_47436# VDD 0.086132f
C16869 a_15890_42674# a_16104_42674# 0.097745f
C16870 a_15803_42450# a_17124_42282# 0.00132f
C16871 a_n3674_37592# a_n4209_38502# 7.92e-20
C16872 a_15486_42560# a_15761_42308# 0.007416f
C16873 a_15959_42545# a_16522_42674# 0.049827f
C16874 a_14113_42308# a_16269_42308# 0.004499f
C16875 a_5932_42308# a_n4209_39590# 8.09e-22
C16876 a_11453_44696# a_13759_46122# 9.57e-21
C16877 a_12465_44636# a_15015_46420# 8.41e-21
C16878 a_6151_47436# a_5066_45546# 0.019067f
C16879 a_4883_46098# a_2324_44458# 0.074521f
C16880 a_13507_46334# a_17583_46090# 0.004113f
C16881 a_18597_46090# a_19553_46090# 0.021441f
C16882 a_18479_47436# a_20075_46420# 0.061108f
C16883 a_10227_46804# a_20708_46348# 0.001063f
C16884 a_19787_47423# a_18819_46122# 1.83e-20
C16885 a_16588_47582# a_6945_45028# 0.011591f
C16886 a_19386_47436# a_18985_46122# 6.11e-19
C16887 a_16023_47582# a_10809_44734# 5.41e-20
C16888 a_n1151_42308# a_8049_45260# 0.075767f
C16889 a_n881_46662# a_6165_46155# 2.6e-19
C16890 a_n1613_43370# a_6419_46155# 0.013016f
C16891 a_3524_46660# a_765_45546# 0.002975f
C16892 a_6755_46942# a_14084_46812# 0.052304f
C16893 a_n2293_46634# a_12741_44636# 3.52e-21
C16894 a_n2840_46634# a_n2840_46090# 0.026152f
C16895 a_768_44030# a_2804_46116# 0.001471f
C16896 a_12891_46348# a_3483_46348# 0.053153f
C16897 a_n1059_45260# a_15953_42852# 0.005616f
C16898 a_n913_45002# a_15597_42852# 6.49e-20
C16899 a_n2017_45002# a_16245_42852# 0.003157f
C16900 a_22591_44484# a_20974_43370# 6.26e-19
C16901 a_18287_44626# a_16137_43396# 8.65e-23
C16902 a_17737_43940# a_17973_43940# 0.22264f
C16903 a_626_44172# a_n2293_42282# 7.4e-21
C16904 a_14539_43914# a_16759_43396# 0.012597f
C16905 a_10193_42453# a_17124_42282# 3.1e-19
C16906 a_17730_32519# a_14401_32519# 0.086728f
C16907 a_19721_31679# a_13887_32519# 0.051264f
C16908 a_5013_44260# a_5025_43940# 0.011829f
C16909 a_5244_44056# a_5326_44056# 0.004767f
C16910 a_22485_44484# a_17538_32519# 0.002174f
C16911 a_18114_32519# a_22591_43396# 6.25e-19
C16912 a_11525_45546# a_11823_42460# 0.001062f
C16913 a_7230_45938# a_6977_45572# 4.61e-19
C16914 a_8162_45546# a_6905_45572# 4.64e-20
C16915 a_11322_45546# a_12791_45546# 5.08e-20
C16916 a_2711_45572# a_15225_45822# 7.31e-20
C16917 a_11750_44172# a_3483_46348# 2.37e-21
C16918 a_n97_42460# a_15227_44166# 0.044664f
C16919 a_21487_43396# a_13747_46662# 0.009398f
C16920 a_19095_43396# a_13661_43548# 0.048302f
C16921 a_20749_43396# a_12549_44172# 0.018798f
C16922 a_5837_43396# a_5257_43370# 1.77e-21
C16923 a_743_42282# a_19321_45002# 1.16e-19
C16924 a_n356_44636# a_n443_42852# 0.262144f
C16925 a_20640_44752# a_8049_45260# 2.15e-21
C16926 a_5891_43370# a_n755_45592# 0.062112f
C16927 a_5663_43940# a_2324_44458# 0.010841f
C16928 a_n3674_39304# a_n1613_43370# 2.21e-20
C16929 a_12545_42858# a_10227_46804# 0.03565f
C16930 a_18083_42858# a_12861_44030# 2.04e-22
C16931 a_413_45260# DATA[4] 0.037695f
C16932 a_15559_46634# VDD 0.301657f
C16933 a_1823_45246# a_2521_46116# 5.42e-19
C16934 a_2202_46116# a_167_45260# 0.159883f
C16935 a_11813_46116# a_11387_46482# 1.25e-20
C16936 a_18285_46348# a_19335_46494# 1.12e-20
C16937 a_19123_46287# a_19553_46090# 1.56e-20
C16938 a_16751_46987# a_10809_44734# 4.31e-19
C16939 a_9313_44734# a_17665_42852# 5.16e-20
C16940 a_21115_43940# a_4190_30871# 0.01145f
C16941 a_20623_43914# a_743_42282# 1.51e-19
C16942 a_14021_43940# a_19700_43370# 0.007203f
C16943 a_11341_43940# a_21259_43561# 0.00271f
C16944 a_7845_44172# a_7871_42858# 5.57e-21
C16945 a_20512_43084# a_19164_43230# 1.84e-20
C16946 a_3422_30871# a_22165_42308# 0.00669f
C16947 a_15493_43396# a_4361_42308# 3.03e-20
C16948 a_8147_43396# VDD 0.393534f
C16949 a_n2472_45002# a_n2109_45247# 0.001038f
C16950 a_n2661_45010# a_n2017_45002# 0.087596f
C16951 a_n2840_45002# a_n1059_45260# 2.05e-21
C16952 a_19963_31679# en_comp 1.68e-19
C16953 a_10193_42453# a_17023_45118# 0.027968f
C16954 a_6469_45572# a_n2661_43370# 3.64e-21
C16955 a_5342_30871# a_13059_46348# 1.53e-19
C16956 a_n3565_38502# SMPL_ON_P 8.06e-19
C16957 a_19511_42282# a_16327_47482# 0.089559f
C16958 a_n2661_43922# CLK 1.98e-19
C16959 a_5907_45546# a_768_44030# 1.57e-21
C16960 a_11652_45724# a_11453_44696# 0.01055f
C16961 a_12791_45546# a_12465_44636# 5.57e-21
C16962 a_13527_45546# a_4883_46098# 9.93e-20
C16963 a_13249_42308# a_13507_46334# 2.05e-20
C16964 a_10210_45822# a_10227_46804# 0.006028f
C16965 a_n1925_42282# a_n2956_38216# 3.5e-20
C16966 a_526_44458# a_n2293_45546# 1.47e-19
C16967 a_14955_43396# a_15279_43071# 4.47e-19
C16968 a_13887_32519# a_22591_43396# 0.006001f
C16969 a_10341_43396# a_14543_43071# 6.95e-20
C16970 a_15095_43370# a_5342_30871# 0.238762f
C16971 a_n97_42460# a_14635_42282# 0.077798f
C16972 a_13678_32519# a_17364_32525# 0.050075f
C16973 a_22223_43396# a_14209_32519# 0.001768f
C16974 a_14579_43548# a_16795_42852# 4.68e-21
C16975 a_n3420_37984# a_n4064_37984# 8.18485f
C16976 a_18175_45572# a_18588_44850# 1.76e-20
C16977 a_10951_45334# a_8975_43940# 2.96e-20
C16978 a_1307_43914# a_2779_44458# 0.332183f
C16979 a_2711_45572# a_17973_43940# 0.011171f
C16980 a_375_42282# a_742_44458# 1.19e-20
C16981 a_9482_43914# a_5883_43914# 0.003705f
C16982 a_n2661_45010# a_n89_44484# 1.47e-19
C16983 a_4169_42308# a_1823_45246# 0.002692f
C16984 a_12379_42858# a_n443_42852# 2.06e-19
C16985 a_17701_42308# a_n357_42282# 0.026888f
C16986 a_1606_42308# a_10903_43370# 1.35e-20
C16987 a_3080_42308# C7_P_btm 0.002948f
C16988 DATA[2] VDD 0.3216f
C16989 a_4099_45572# a_1823_45246# 0.047087f
C16990 a_2711_45572# a_167_45260# 0.003442f
C16991 a_7499_43078# a_11415_45002# 4.24e-20
C16992 a_13556_45296# a_n2293_46634# 0.00155f
C16993 a_14537_43396# a_n2661_46634# 7.41e-21
C16994 a_3357_43084# a_7577_46660# 1.08e-20
C16995 a_2437_43646# a_8667_46634# 1.27e-20
C16996 a_3537_45260# a_2609_46660# 4.52e-20
C16997 a_3065_45002# a_2959_46660# 2.84e-20
C16998 a_3429_45260# a_3177_46902# 3.58e-20
C16999 a_8103_44636# a_n1151_42308# 2.41e-19
C17000 a_4223_44672# a_4791_45118# 0.399086f
C17001 a_2779_44458# a_n443_46116# 0.00406f
C17002 a_10334_44484# a_2063_45854# 4.46e-36
C17003 a_n1809_44850# a_n2497_47436# 0.00201f
C17004 a_19113_45348# a_16327_47482# 1.22e-19
C17005 a_20567_45036# a_18479_47436# 2.48e-20
C17006 a_18184_42460# a_18597_46090# 0.020766f
C17007 a_16922_45042# a_4883_46098# 4.62e-20
C17008 a_13490_45067# a_11453_44696# 4.23e-19
C17009 a_n2293_42834# a_n1613_43370# 0.123758f
C17010 a_2905_42968# a_1755_42282# 2.89e-20
C17011 a_9127_43156# a_n784_42308# 1.7e-20
C17012 a_15743_43084# a_15959_42545# 0.00371f
C17013 a_1847_42826# a_2351_42308# 0.120686f
C17014 a_4361_42308# a_8791_42308# 0.009181f
C17015 a_16137_43396# a_17124_42282# 6.71e-20
C17016 a_10341_43396# a_19511_42282# 1.05e-21
C17017 a_5342_30871# a_14097_32519# 0.028503f
C17018 a_14209_32519# a_5934_30871# 0.004208f
C17019 a_743_42282# a_9885_42558# 0.006242f
C17020 a_8049_45260# START 1.99e-20
C17021 a_20205_31679# a_22521_40055# 9e-21
C17022 a_n4209_38216# VDD 0.833976f
C17023 a_7227_47204# a_5807_45002# 1.09e-19
C17024 a_12861_44030# a_12549_44172# 1.20253f
C17025 a_13717_47436# a_768_44030# 0.029731f
C17026 a_13487_47204# a_12891_46348# 1.6e-19
C17027 a_16023_47582# a_n881_46662# 1.58e-20
C17028 a_22731_47423# a_11453_44696# 0.048111f
C17029 a_584_46384# a_n743_46660# 0.42078f
C17030 a_n2109_47186# a_1799_45572# 1.89e-19
C17031 a_n237_47217# a_948_46660# 6.91e-20
C17032 a_n1151_42308# a_n2442_46660# 6.91e-20
C17033 a_n2288_47178# a_n2661_46098# 2.56e-20
C17034 a_n785_47204# a_383_46660# 0.001568f
C17035 a_327_47204# a_601_46902# 0.003002f
C17036 a_2124_47436# a_n2438_43548# 3.55e-19
C17037 a_2553_47502# a_n1925_46634# 4.04e-20
C17038 a_n971_45724# a_1983_46706# 0.004287f
C17039 a_3785_47178# a_n2661_46634# 7.96e-20
C17040 a_18114_32519# a_22591_44484# 0.018563f
C17041 a_15004_44636# a_15146_44484# 0.007833f
C17042 a_16979_44734# a_17061_44734# 0.171361f
C17043 a_14539_43914# a_17517_44484# 6.45e-19
C17044 a_9482_43914# a_12495_44260# 0.002157f
C17045 a_16019_45002# a_15493_43940# 3.46e-19
C17046 a_5147_45002# a_5745_43940# 0.007407f
C17047 a_3232_43370# a_3737_43940# 6.52e-19
C17048 a_n2017_45002# a_21381_43940# 3.18e-20
C17049 a_2437_43646# a_n97_42460# 0.201806f
C17050 a_5111_44636# a_5326_44056# 2.81e-20
C17051 a_21613_42308# a_n357_42282# 3.71e-20
C17052 a_n4315_30879# a_n2956_38216# 0.025091f
C17053 a_n2302_40160# a_n2810_45572# 7.76e-19
C17054 a_21350_45938# VDD 7.19e-19
C17055 a_5518_44484# a_3090_45724# 9.17e-21
C17056 a_21398_44850# a_13747_46662# 0.011329f
C17057 a_17786_45822# a_13259_45724# 0.001706f
C17058 a_21188_45572# a_8049_45260# 0.015577f
C17059 a_n2661_45010# a_526_44458# 0.703081f
C17060 a_10775_45002# a_10903_43370# 3.83e-19
C17061 a_3232_43370# a_2324_44458# 0.410727f
C17062 a_11341_43940# a_4915_47217# 3.68e-20
C17063 a_12429_44172# a_12861_44030# 0.108591f
C17064 a_1423_45028# a_4419_46090# 3.66e-20
C17065 a_6761_42308# a_8791_42308# 6.62e-21
C17066 a_6123_31319# a_8325_42308# 6.08e-19
C17067 a_7227_42308# a_8685_42308# 7.46e-20
C17068 COMP_P a_4958_30871# 0.02709f
C17069 a_18194_35068# a_19120_35138# 0.558402f
C17070 EN_VIN_BSTR_N a_19864_35138# 0.573134f
C17071 EN_VIN_BSTR_P C9_P_btm 0.226529f
C17072 a_n2661_46634# a_3090_45724# 6.05e-20
C17073 a_768_44030# a_14035_46660# 0.270355f
C17074 a_19321_45002# a_19466_46812# 0.130025f
C17075 a_19594_46812# a_19333_46634# 0.060858f
C17076 a_12549_44172# a_14180_46812# 0.023435f
C17077 a_n743_46660# a_11901_46660# 9.04e-20
C17078 a_4646_46812# a_7715_46873# 0.058457f
C17079 a_4651_46660# a_7411_46660# 1.59e-21
C17080 a_5385_46902# a_5263_46660# 3.16e-19
C17081 a_5807_45002# a_12156_46660# 0.002125f
C17082 a_3877_44458# a_7577_46660# 2.44e-19
C17083 a_4955_46873# a_5257_43370# 2.43e-21
C17084 a_10227_46804# a_21542_46660# 0.002879f
C17085 a_18597_46090# a_12741_44636# 0.267775f
C17086 a_13507_46334# a_20885_46660# 4.28e-19
C17087 a_n1435_47204# a_1138_42852# 1.06e-20
C17088 a_5129_47502# a_5204_45822# 2.88e-19
C17089 a_n1151_42308# a_8953_45546# 0.120628f
C17090 a_2063_45854# a_9290_44172# 0.655982f
C17091 a_4791_45118# a_6419_46155# 0.371259f
C17092 a_6298_44484# a_6765_43638# 0.001141f
C17093 a_1414_42308# a_n2661_42282# 1.17e-20
C17094 a_5883_43914# a_6031_43396# 0.001063f
C17095 a_5343_44458# a_7287_43370# 2.75e-19
C17096 a_16922_45042# a_16243_43396# 6.03e-22
C17097 a_9313_44734# a_20974_43370# 1.96e-19
C17098 a_3422_30871# a_19862_44208# 0.030442f
C17099 a_2998_44172# a_1525_44260# 4.65e-22
C17100 a_5111_44636# a_10083_42826# 0.005394f
C17101 a_3232_43370# a_8387_43230# 1.01e-22
C17102 a_n913_45002# a_18083_42858# 6.19e-20
C17103 a_n2017_45002# a_18249_42858# 0.545311f
C17104 a_n1059_45260# a_17333_42852# 0.270324f
C17105 a_7_44811# VDD 0.001865f
C17106 a_n4209_39590# VREF 0.860047f
C17107 a_n3565_39590# VIN_P 0.068367f
C17108 a_n4209_38502# EN_VIN_BSTR_P 0.002888f
C17109 a_n3565_38502# a_n1532_35090# 1.48e-19
C17110 a_n4064_39072# C8_P_btm 7.96e-19
C17111 a_n3420_39072# C6_P_btm 0.054459f
C17112 a_n3565_39304# C4_P_btm 5.85e-20
C17113 a_2711_45572# a_3175_45822# 7.71e-19
C17114 a_n3420_37440# a_n2956_38216# 0.001161f
C17115 a_n2302_37690# a_n2810_45572# 5.35e-19
C17116 a_3422_30871# a_4185_45028# 0.176529f
C17117 a_9145_43396# a_768_44030# 0.004455f
C17118 a_20365_43914# a_19692_46634# 0.001873f
C17119 a_6293_42852# a_n2293_46634# 0.014742f
C17120 a_n2433_44484# a_n2661_45546# 3.06e-20
C17121 a_n2661_43922# a_n2956_39304# 1.05e-20
C17122 a_n4318_40392# a_n2956_38216# 0.027558f
C17123 a_1847_42826# a_584_46384# 4.79e-19
C17124 a_n722_43218# a_n1151_42308# 3.54e-19
C17125 a_21855_43396# a_12861_44030# 9.83e-19
C17126 a_21259_43561# a_16327_47482# 4.28e-20
C17127 a_19700_43370# a_13507_46334# 4.92e-21
C17128 a_14581_44484# a_2324_44458# 1.05e-20
C17129 a_13213_44734# a_10809_44734# 1.94e-20
C17130 a_14673_44172# a_14840_46494# 2.17e-21
C17131 a_3067_47026# VDD 0.132018f
C17132 a_n4334_39392# a_n4064_38528# 7.84e-19
C17133 a_n3690_39392# a_n3420_38528# 7.84e-19
C17134 a_n2946_39072# a_n3565_38502# 9.15e-19
C17135 a_n2302_39072# a_n4209_38502# 9.15e-19
C17136 a_n3420_39072# a_n3690_38528# 0.017537f
C17137 a_n4209_39304# a_n2302_38778# 0.001019f
C17138 a_1736_39587# a_2684_37794# 0.565517f
C17139 a_n4064_39072# a_n4334_38528# 0.00115f
C17140 a_n3565_39304# a_n2946_38778# 9.15e-19
C17141 a_n4064_39616# a_n3565_38216# 0.028071f
C17142 a_1736_39043# comp_n 0.005064f
C17143 a_n1630_35242# a_n2302_37984# 5.02e-20
C17144 a_10150_46912# a_6945_45028# 5.48e-20
C17145 a_11735_46660# a_11387_46155# 1.2e-19
C17146 a_3090_45724# a_8199_44636# 0.030057f
C17147 a_n881_46662# a_n23_45546# 3.9e-19
C17148 a_20623_46660# a_20885_46660# 0.001705f
C17149 a_21188_46660# a_21350_47026# 0.006453f
C17150 a_20411_46873# a_11415_45002# 4.84e-20
C17151 a_19123_46287# a_12741_44636# 3.1e-21
C17152 a_20273_46660# a_20202_43084# 8.55e-20
C17153 a_20107_46660# a_22591_46660# 3.89e-21
C17154 a_13483_43940# a_9145_43396# 0.002944f
C17155 a_22485_44484# a_22591_43396# 0.025074f
C17156 a_9313_44734# a_18599_43230# 0.008115f
C17157 a_14401_32519# a_17538_32519# 0.052152f
C17158 a_19237_31679# a_13678_32519# 0.052466f
C17159 a_20512_43084# a_14209_32519# 0.006512f
C17160 en_comp a_7174_31319# 5.65154f
C17161 a_n913_45002# a_22775_42308# 7.44e-19
C17162 a_10555_43940# VDD 0.002652f
C17163 a_6598_45938# a_1423_45028# 2.06e-21
C17164 a_10193_42453# a_10951_45334# 1.8e-20
C17165 a_8746_45002# a_10775_45002# 2.04e-20
C17166 a_18341_45572# a_19418_45938# 1.46e-19
C17167 a_18479_45785# a_18787_45572# 0.004823f
C17168 a_2711_45572# a_5105_45348# 1.42e-19
C17169 a_10490_45724# a_8953_45002# 4.57e-19
C17170 a_13163_45724# a_6171_45002# 1.51e-20
C17171 a_743_42282# a_13059_46348# 2.35e-20
C17172 a_11750_44172# a_n357_42282# 2.28e-21
C17173 a_6765_43638# a_5937_45572# 9.53e-19
C17174 a_n3674_37592# a_n2312_39304# 0.026622f
C17175 a_5742_30871# a_4791_45118# 3.2e-20
C17176 a_21137_46414# VDD 0.219745f
C17177 a_2211_45572# a_n443_46116# 1.46e-19
C17178 a_9049_44484# a_2063_45854# 3.38e-20
C17179 a_6598_45938# a_6491_46660# 1.3e-21
C17180 a_2711_45572# a_11459_47204# 3.52e-21
C17181 a_6511_45714# a_7227_47204# 7.86e-21
C17182 a_n1853_46287# a_n356_45724# 0.011459f
C17183 a_472_46348# a_n755_45592# 3.56e-20
C17184 a_3147_46376# a_n2661_45546# 6.59e-20
C17185 a_805_46414# a_n357_42282# 6.63e-19
C17186 a_1176_45822# a_n1099_45572# 5.28e-20
C17187 a_n2293_46098# a_n310_45899# 7.73e-19
C17188 a_19553_46090# a_8049_45260# 0.002856f
C17189 a_13759_46122# a_14180_46482# 0.086708f
C17190 a_10903_43370# a_12839_46116# 0.115226f
C17191 a_15095_43370# a_743_42282# 2.85e-19
C17192 a_16243_43396# a_15743_43084# 0.600668f
C17193 a_10341_43396# a_21259_43561# 0.00679f
C17194 a_648_43396# a_685_42968# 5.58e-19
C17195 a_3539_42460# a_3681_42891# 4.58e-21
C17196 a_3626_43646# a_3935_42891# 0.002569f
C17197 a_2982_43646# a_5111_42852# 2.74e-20
C17198 a_n97_42460# a_14543_43071# 7.94e-21
C17199 a_n2661_42282# a_n3674_38680# 0.00768f
C17200 a_11967_42832# a_14113_42308# 0.003103f
C17201 a_16759_43396# a_17324_43396# 7.99e-20
C17202 a_16409_43396# a_18525_43370# 1.15e-20
C17203 a_n2661_46634# CLK_DATA 3.38e-19
C17204 a_13113_42826# VDD 0.217254f
C17205 a_18175_45572# a_18443_44721# 9.32e-21
C17206 a_18341_45572# a_18248_44752# 3.18e-20
C17207 a_18479_45785# a_18287_44626# 0.024431f
C17208 a_13017_45260# a_13105_45348# 2.63e-19
C17209 a_1423_45028# a_2809_45028# 8.35e-21
C17210 a_7499_43078# a_11967_42832# 5.46e-21
C17211 a_n2840_45002# a_n4318_40392# 4.48e-19
C17212 a_n2661_45010# a_n2840_44458# 3.06e-19
C17213 a_2437_43646# a_742_44458# 0.081793f
C17214 a_6171_45002# a_16501_45348# 2.67e-19
C17215 a_413_45260# a_22223_45036# 2.66e-19
C17216 a_n4064_38528# a_n2312_38680# 0.22404f
C17217 a_4361_42308# a_n357_42282# 0.069224f
C17218 a_n2293_42282# a_n2956_38680# 3.4e-20
C17219 a_10793_43218# a_9290_44172# 0.001055f
C17220 a_10193_42453# a_11735_46660# 0.001441f
C17221 a_10907_45822# a_10428_46928# 4.91e-20
C17222 a_10210_45822# a_10467_46802# 4.57e-20
C17223 a_n1059_45260# a_768_44030# 2.61e-19
C17224 a_n913_45002# a_12549_44172# 7.26e-19
C17225 a_2437_43646# a_20843_47204# 0.004179f
C17226 a_3357_43084# a_19452_47524# 1.74e-19
C17227 a_n37_45144# a_n881_46662# 3.17e-19
C17228 a_413_45260# a_n1613_43370# 0.046335f
C17229 a_10775_45002# a_4883_46098# 1.52e-21
C17230 a_16751_45260# a_16327_47482# 1.87e-19
C17231 a_14797_45144# a_10227_46804# 0.003451f
C17232 a_n2293_42834# a_4791_45118# 0.046352f
C17233 a_18249_42858# a_19164_43230# 0.118759f
C17234 a_3626_43646# a_15890_42674# 0.003304f
C17235 a_n97_42460# a_19511_42282# 7.78e-21
C17236 a_8037_42858# a_8483_43230# 2.28e-19
C17237 a_14401_32519# a_22465_38105# 8.57e-20
C17238 a_6419_46155# DATA[3] 9.23e-21
C17239 a_18214_42558# VDD 0.295211f
C17240 a_n356_44636# CAL_N 5.72e-19
C17241 a_n815_47178# a_n2312_39304# 8.4e-20
C17242 a_9313_45822# a_11459_47204# 0.210847f
C17243 a_9863_47436# a_n1435_47204# 2.39e-19
C17244 a_6151_47436# a_15811_47375# 1.9e-19
C17245 a_n1741_47186# a_2266_47570# 2.25e-19
C17246 a_n2109_47186# a_2747_46873# 0.087441f
C17247 a_11691_44458# a_n2661_43922# 0.038882f
C17248 a_375_42282# a_n984_44318# 1.76e-20
C17249 a_1307_43914# a_644_44056# 1.94e-20
C17250 a_18114_32519# a_9313_44734# 1.28e-20
C17251 a_n2661_44458# a_8333_44734# 9.44e-20
C17252 a_n913_45002# a_12429_44172# 1.57e-21
C17253 a_n1059_45260# a_13483_43940# 1.59e-20
C17254 a_3065_45002# a_3499_42826# 3.27e-19
C17255 a_3823_42558# a_n443_42852# 9.86e-21
C17256 a_6761_42308# a_n357_42282# 5.14e-21
C17257 a_14113_42308# a_13259_45724# 0.00391f
C17258 a_n3565_39590# a_n2956_38680# 0.021577f
C17259 a_10907_45822# VDD 0.352181f
C17260 a_413_45260# a_n2293_46098# 0.034414f
C17261 a_n2017_45002# a_1138_42852# 1.31e-19
C17262 a_19963_31679# a_4185_45028# 9.16e-19
C17263 a_6194_45824# a_n2661_45546# 4.12e-20
C17264 a_1176_45572# a_n1099_45572# 5.07e-20
C17265 a_1525_44260# a_n2497_47436# 4.47e-19
C17266 a_895_43940# a_n1151_42308# 6.25e-21
C17267 a_18681_44484# a_16327_47482# 0.001931f
C17268 a_20679_44626# a_18479_47436# 0.018117f
C17269 a_20362_44736# a_18597_46090# 3.05e-20
C17270 a_17517_44484# a_11453_44696# 0.014468f
C17271 a_2437_43646# a_5204_45822# 3.52e-20
C17272 a_16147_45260# a_17715_44484# 0.020415f
C17273 a_1067_42314# a_1184_42692# 0.147283f
C17274 a_n784_42308# a_1755_42282# 0.073102f
C17275 a_n1630_35242# a_961_42354# 3.02e-19
C17276 a_13507_46334# a_11813_46116# 1.34e-19
C17277 a_10227_46804# a_14976_45028# 0.536884f
C17278 a_16327_47482# a_18834_46812# 3.5e-20
C17279 a_6151_47436# a_13059_46348# 1.9e-19
C17280 a_3785_47178# a_765_45546# 0.004672f
C17281 a_8128_46384# a_7577_46660# 0.023306f
C17282 a_5807_45002# a_4955_46873# 4.29e-20
C17283 a_n2438_43548# a_1110_47026# 2.49e-19
C17284 a_n743_46660# a_479_46660# 0.004337f
C17285 a_1123_46634# a_948_46660# 0.234322f
C17286 a_33_46660# a_288_46660# 0.056391f
C17287 a_n1925_46634# a_1799_45572# 0.035794f
C17288 a_n2293_46634# a_2609_46660# 1.11e-20
C17289 a_n2661_46634# a_3699_46634# 0.009256f
C17290 a_n2312_38680# a_n2661_46098# 0.003978f
C17291 a_18287_44626# a_14021_43940# 2.78e-20
C17292 a_22485_44484# a_22591_44484# 0.15878f
C17293 a_n2661_43922# a_8333_44056# 7.64e-20
C17294 a_n2661_42834# a_9028_43914# 0.009687f
C17295 a_9313_44734# a_17737_43940# 1.96e-20
C17296 a_19721_31679# a_14401_32519# 0.053967f
C17297 a_5883_43914# a_6671_43940# 0.051304f
C17298 a_7499_43078# a_9114_42852# 2.49e-19
C17299 a_1307_43914# a_10765_43646# 8.56e-19
C17300 a_n913_45002# a_21855_43396# 3.57e-20
C17301 a_n2017_45002# a_5649_42852# 0.03149f
C17302 a_21359_45002# VDD 0.319372f
C17303 a_5891_43370# a_3483_46348# 0.005051f
C17304 a_19319_43548# a_5807_45002# 1.9e-20
C17305 a_1423_45028# a_1848_45724# 8.69e-22
C17306 a_18184_42460# a_8049_45260# 6.28e-23
C17307 a_2304_45348# a_n755_45592# 2.24e-19
C17308 a_8975_43940# a_2324_44458# 0.005091f
C17309 a_n356_44636# a_8199_44636# 2.05e-19
C17310 a_4223_44672# a_6945_45028# 1.31e-20
C17311 a_n2012_43396# a_n1613_43370# 2.53e-19
C17312 a_n1557_42282# a_n2312_40392# 2.63e-20
C17313 a_10341_43396# a_4915_47217# 2.29e-20
C17314 a_3094_47243# VDD 6.34e-20
C17315 a_n784_42308# C2_N_btm 0.005178f
C17316 a_6755_46942# a_12741_44636# 0.131965f
C17317 a_4955_46873# a_3699_46348# 1.24e-20
C17318 a_3090_45724# a_765_45546# 0.001007f
C17319 a_15368_46634# a_15312_46660# 1.11e-19
C17320 a_768_44030# a_n1925_42282# 0.145535f
C17321 a_n881_46662# a_5210_46155# 1.33e-19
C17322 a_3877_44458# a_4704_46090# 3.8e-19
C17323 a_20916_46384# a_22223_46124# 5.13e-19
C17324 a_n743_46660# a_17583_46090# 4.13e-19
C17325 a_21588_30879# a_6945_45028# 1.26e-19
C17326 a_4883_46098# a_12839_46116# 1.63e-19
C17327 a_13507_46334# a_14949_46494# 2.9e-19
C17328 a_18597_46090# a_16375_45002# 0.105669f
C17329 a_11599_46634# a_20850_46155# 7e-21
C17330 a_16327_47482# a_20850_46482# 2.1e-19
C17331 a_n443_46116# a_n23_45546# 0.118272f
C17332 a_2905_45572# a_1990_45899# 1.24e-19
C17333 a_584_46384# a_509_45572# 3.56e-19
C17334 a_4646_46812# a_4419_46090# 1.97e-19
C17335 a_10334_44484# a_10083_42826# 5.56e-20
C17336 a_19478_44306# a_19319_43548# 0.005956f
C17337 a_11967_42832# a_15781_43660# 0.026392f
C17338 a_17517_44484# a_17324_43396# 7.13e-22
C17339 a_9313_44734# a_13887_32519# 0.191376f
C17340 a_1241_43940# a_1443_43940# 0.092725f
C17341 a_19328_44172# a_19478_44056# 0.003538f
C17342 a_11341_43940# a_11173_43940# 1.36e-19
C17343 a_n1059_45260# a_6123_31319# 0.001842f
C17344 a_n913_45002# a_7227_42308# 0.052824f
C17345 a_3065_45002# a_3318_42354# 0.146272f
C17346 a_n2017_45002# a_7963_42308# 0.003883f
C17347 en_comp a_5932_42308# 0.233106f
C17348 a_n2661_42282# VDD 0.406474f
C17349 a_20922_43172# a_12549_44172# 6.03e-19
C17350 a_10991_42826# a_n2293_46634# 4.93e-20
C17351 a_16414_43172# a_13661_43548# 2.69e-21
C17352 a_n3674_38216# a_n1151_42308# 6.62e-20
C17353 a_13157_43218# a_10227_46804# 0.001903f
C17354 a_n914_42852# a_n1613_43370# 1.3e-19
C17355 a_9801_43940# a_8016_46348# 4.95e-19
C17356 a_11341_43940# a_10809_44734# 1.55e-19
C17357 a_n2840_46090# VDD 0.295278f
C17358 a_18727_42674# CAL_N 0.001564f
C17359 a_13759_46122# a_13925_46122# 0.576786f
C17360 a_6419_46155# a_6945_45028# 1.24e-19
C17361 a_10903_43370# a_14840_46494# 8.02e-21
C17362 a_18285_46348# a_19240_46482# 2.07e-21
C17363 a_17339_46660# a_18051_46116# 0.040259f
C17364 a_19123_46287# a_16375_45002# 1.65e-19
C17365 a_12741_44636# a_8049_45260# 0.037594f
C17366 a_1138_42852# a_526_44458# 0.039045f
C17367 a_472_46348# a_835_46155# 0.005265f
C17368 a_18079_43940# a_18249_42858# 7.49e-20
C17369 a_18326_43940# a_17333_42852# 7.02e-19
C17370 a_18451_43940# a_18083_42858# 2.66e-22
C17371 a_2982_43646# a_16977_43638# 3.11e-21
C17372 a_3626_43646# a_16547_43609# 3.44e-21
C17373 a_14401_32519# a_22591_43396# 0.01561f
C17374 a_11341_43940# a_13460_43230# 2.23e-21
C17375 a_15493_43396# a_17595_43084# 1.05e-20
C17376 a_n2293_43922# a_4921_42308# 1.79e-19
C17377 a_5891_43370# a_8791_42308# 7.71e-19
C17378 a_n356_44636# a_13070_42354# 1.4e-19
C17379 a_20974_43370# a_13887_32519# 0.033282f
C17380 a_8685_43396# a_8423_43396# 2.34e-19
C17381 a_18597_46090# RST_Z 1.14e-19
C17382 a_18479_47436# SINGLE_ENDED 0.040779f
C17383 SMPL_ON_N a_18194_35068# 3.71e-19
C17384 a_15673_47210# CLK 3.17e-19
C17385 a_18780_47178# START 0.01578f
C17386 a_16823_43084# VDD 0.159922f
C17387 a_18341_45572# a_16922_45042# 3.38e-20
C17388 a_16147_45260# a_17719_45144# 0.049848f
C17389 a_8696_44636# a_16237_45028# 3.7e-19
C17390 a_11823_42460# a_13076_44458# 1.17e-19
C17391 a_10193_42453# a_18248_44752# 0.004992f
C17392 a_2711_45572# a_9313_44734# 0.036278f
C17393 a_6598_45938# a_6109_44484# 6.27e-20
C17394 a_6469_45572# a_5883_43914# 3.18e-21
C17395 a_3232_43370# a_10775_45002# 1.54e-20
C17396 a_3537_45260# a_9482_43914# 3.66e-21
C17397 a_7276_45260# a_6709_45028# 0.215102f
C17398 a_6171_45002# a_8953_45002# 0.034987f
C17399 a_6431_45366# a_8191_45002# 8.63e-21
C17400 a_7174_31319# a_13661_43548# 1.16e-20
C17401 a_5649_42852# a_526_44458# 0.058712f
C17402 a_6765_43638# a_n443_42852# 0.00334f
C17403 a_2905_42968# a_2324_44458# 8.09e-22
C17404 a_10083_42826# a_9290_44172# 0.136441f
C17405 a_n2302_39072# a_n2312_39304# 0.130454f
C17406 a_n37_45144# a_n443_46116# 3.75e-19
C17407 a_413_45260# a_4791_45118# 2.6e-19
C17408 a_3429_45260# a_3160_47472# 3.37e-21
C17409 a_5147_45002# a_2063_45854# 1.79e-19
C17410 a_7229_43940# a_n237_47217# 4.29e-19
C17411 a_7705_45326# a_n971_45724# 5.33e-21
C17412 a_13249_42308# a_n743_46660# 4.93e-20
C17413 a_6598_45938# a_4646_46812# 6.19e-19
C17414 a_15903_45785# a_12549_44172# 3.38e-20
C17415 a_16223_45938# a_n881_46662# 8.49e-19
C17416 a_21363_45546# a_18597_46090# 0.001567f
C17417 a_21513_45002# a_16327_47482# 0.013118f
C17418 a_2437_43646# a_16241_47178# 0.004738f
C17419 a_3357_43084# a_15507_47210# 4.74e-19
C17420 a_20273_45572# a_20894_47436# 1.81e-21
C17421 a_n2661_45546# a_310_45028# 0.035423f
C17422 a_n2293_45546# a_n452_45724# 2.19e-20
C17423 a_n1079_45724# a_n863_45724# 0.091159f
C17424 a_n2472_45546# a_n1099_45572# 9.27e-20
C17425 a_20623_43914# a_13258_32519# 1.97e-21
C17426 a_3080_42308# a_1755_42282# 0.047244f
C17427 a_4361_42308# a_21356_42826# 0.017293f
C17428 a_13467_32519# a_21195_42852# 0.034759f
C17429 a_5649_42852# a_19164_43230# 5.64e-21
C17430 a_14021_43940# a_17124_42282# 4.98e-21
C17431 a_n97_42460# a_4921_42308# 3.35e-20
C17432 a_10341_43396# a_13291_42460# 7.32e-20
C17433 a_20820_30879# a_22609_37990# 1.17e-20
C17434 a_18285_46348# START 0.001916f
C17435 a_19123_46287# RST_Z 4.05e-21
C17436 a_n4209_37414# a_n3565_37414# 6.90997f
C17437 a_3497_42558# VDD 0.007751f
C17438 a_n971_45724# a_n785_47204# 0.385455f
C17439 a_n746_45260# a_n23_47502# 0.148631f
C17440 a_n1741_47186# a_2124_47436# 0.009997f
C17441 a_n2109_47186# a_2063_45854# 0.045645f
C17442 a_14537_43396# a_15433_44458# 0.018743f
C17443 a_8696_44636# a_9672_43914# 4.19e-20
C17444 a_14797_45144# a_14815_43914# 3.57e-20
C17445 a_13249_42308# a_13829_44260# 7.14e-19
C17446 a_375_42282# a_n2661_43922# 0.024229f
C17447 a_13904_45546# a_14021_43940# 1.09e-21
C17448 a_n2661_43370# a_n2012_44484# 8.13e-19
C17449 a_7174_31319# a_4185_45028# 0.027406f
C17450 a_13622_42852# a_n357_42282# 1.14e-19
C17451 a_7963_42308# a_526_44458# 5.22e-20
C17452 a_22400_42852# a_20692_30879# 8.51e-20
C17453 a_14097_32519# a_20205_31679# 0.051224f
C17454 a_6123_31319# a_n1925_42282# 3.21e-20
C17455 a_20273_45572# a_20411_46873# 6.47e-19
C17456 a_11064_45572# a_3483_46348# 0.002687f
C17457 a_16377_45572# a_11415_45002# 4.28e-19
C17458 a_20107_45572# a_20273_46660# 8.09e-19
C17459 a_13556_45296# a_6755_46942# 0.103107f
C17460 a_20193_45348# a_19321_45002# 0.489018f
C17461 a_16981_45144# a_13661_43548# 2.68e-21
C17462 a_n2661_43370# a_n2661_46098# 1.87e-20
C17463 a_11691_44458# a_19594_46812# 1.96e-19
C17464 a_n2661_44458# a_12549_44172# 4.11e-20
C17465 a_2382_45260# a_3090_45724# 0.002468f
C17466 a_2437_43646# a_16721_46634# 1.5e-22
C17467 a_413_45260# a_16292_46812# 1.24e-20
C17468 a_20841_45814# a_20107_46660# 1.73e-21
C17469 a_7229_43940# a_8270_45546# 1.4e-36
C17470 a_949_44458# a_n881_46662# 1.39e-19
C17471 a_10193_42453# a_2324_44458# 0.041338f
C17472 a_13163_45724# a_10903_43370# 0.06577f
C17473 a_11823_42460# a_12594_46348# 0.081079f
C17474 a_8697_45822# a_8199_44636# 0.067739f
C17475 a_10210_45822# a_8016_46348# 0.003734f
C17476 a_13720_44458# a_11453_44696# 1.26e-20
C17477 a_9313_44734# a_9313_45822# 1.19e-20
C17478 a_12089_42308# a_12563_42308# 0.03299f
C17479 a_12379_42858# a_13070_42354# 6.78e-21
C17480 a_5649_42852# a_21973_42336# 0.001208f
C17481 a_13887_32519# a_22397_42558# 0.002537f
C17482 a_3080_42308# C2_N_btm 0.108823f
C17483 a_2747_46873# a_n1925_46634# 0.007371f
C17484 a_6491_46660# a_7411_46660# 2.68e-21
C17485 a_6151_47436# a_7577_46660# 0.578207f
C17486 a_4915_47217# a_8667_46634# 4.1e-20
C17487 a_6545_47178# a_7715_46873# 0.003195f
C17488 a_n1435_47204# a_5907_46634# 3.08e-20
C17489 a_n1741_47186# a_11813_46116# 0.004098f
C17490 a_n1151_42308# a_10249_46116# 0.060327f
C17491 a_n237_47217# a_8270_45546# 0.552109f
C17492 a_n971_45724# a_8601_46660# 5.7e-19
C17493 a_22223_45036# a_22223_43948# 6.3e-19
C17494 a_20193_45348# a_20623_43914# 0.048456f
C17495 a_7499_43078# a_10518_42984# 0.03265f
C17496 a_9313_44734# a_22485_44484# 2.92e-21
C17497 a_1307_43914# a_104_43370# 7.32e-21
C17498 a_n699_43396# a_n2661_42282# 4.19e-21
C17499 a_18479_45785# a_19268_43646# 0.12682f
C17500 a_2711_45572# a_18599_43230# 4e-19
C17501 a_16241_44734# a_16241_44484# 6.96e-20
C17502 a_14673_44172# a_16335_44484# 6.01e-19
C17503 a_11827_44484# a_15493_43940# 0.010315f
C17504 a_3537_45260# a_6031_43396# 0.034593f
C17505 a_n2017_45002# a_8685_43396# 2.66e-19
C17506 a_3232_43370# a_3539_42460# 1.57e-22
C17507 a_15415_45028# VDD 0.191729f
C17508 a_1606_42308# a_n923_35174# 0.002555f
C17509 a_n1630_35242# a_19864_35138# 0.020191f
C17510 a_n784_42308# C8_P_btm 6.79e-20
C17511 a_4235_43370# a_584_46384# 0.016368f
C17512 a_2982_43646# a_n971_45724# 3.56e-20
C17513 a_1512_43396# a_n2497_47436# 9.13e-21
C17514 a_n1177_44458# a_n1641_46494# 4.88e-19
C17515 a_2779_44458# a_n2293_46098# 2.44e-20
C17516 a_15433_44458# a_3090_45724# 0.001223f
C17517 a_18451_43940# a_12549_44172# 0.013387f
C17518 a_11787_45002# a_10586_45546# 3.84e-19
C17519 a_13556_45296# a_8049_45260# 8.2e-22
C17520 a_3602_45348# a_526_44458# 7.3e-19
C17521 a_n2661_45010# a_n452_45724# 4.16e-21
C17522 a_n2810_45028# a_n2840_45546# 5.19e-19
C17523 a_n913_45002# a_n2661_45546# 9.6e-19
C17524 a_14309_45348# a_2324_44458# 0.001898f
C17525 a_11341_43940# a_n881_46662# 6.61e-21
C17526 a_4007_47204# VDD 0.41212f
C17527 a_15803_42450# a_16522_42674# 0.089677f
C17528 a_9803_42558# a_7174_31319# 4.88e-21
C17529 a_15959_42545# a_16104_42674# 0.057222f
C17530 a_14113_42308# a_16197_42308# 0.002157f
C17531 a_15764_42576# a_17124_42282# 1e-19
C17532 a_6123_31319# a_n4315_30879# 7.4e-21
C17533 a_11453_44696# a_13351_46090# 8.02e-21
C17534 a_12465_44636# a_14275_46494# 0.00587f
C17535 a_4883_46098# a_14840_46494# 0.004918f
C17536 a_13507_46334# a_15682_46116# 0.022078f
C17537 a_19386_47436# a_18819_46122# 1.81e-21
C17538 a_18479_47436# a_19335_46494# 1.52e-20
C17539 a_18597_46090# a_18985_46122# 0.027318f
C17540 a_16327_47482# a_10809_44734# 0.036039f
C17541 a_16763_47508# a_6945_45028# 0.01658f
C17542 a_4791_45118# a_5527_46155# 2.63e-19
C17543 a_n881_46662# a_5497_46414# 0.001017f
C17544 a_n1613_43370# a_6165_46155# 3.04e-19
C17545 a_3699_46634# a_765_45546# 0.002795f
C17546 a_6755_46942# a_13607_46688# 0.129798f
C17547 a_11309_47204# a_3483_46348# 1.47e-20
C17548 a_768_44030# a_2698_46116# 0.001262f
C17549 a_16979_44734# a_16409_43396# 6.95e-19
C17550 a_22485_44484# a_20974_43370# 0.101193f
C17551 a_14673_44172# a_3626_43646# 4.56e-21
C17552 a_14539_43914# a_16977_43638# 0.013865f
C17553 a_18114_32519# a_13887_32519# 0.054996f
C17554 a_5244_44056# a_5025_43940# 6.46e-21
C17555 a_20512_43084# a_17538_32519# 5.55e-20
C17556 a_22591_44484# a_14401_32519# 0.001482f
C17557 a_n2017_45002# a_15953_42852# 9.63e-19
C17558 a_19479_31679# a_14097_32519# 0.05096f
C17559 a_n1059_45260# a_15597_42852# 0.056846f
C17560 a_n913_45002# a_14853_42852# 7.37e-19
C17561 a_19279_43940# VDD 0.302681f
C17562 a_2711_45572# a_15037_45618# 0.005856f
C17563 a_11322_45546# a_11823_42460# 0.133185f
C17564 a_11652_45724# a_11962_45724# 0.002072f
C17565 a_10490_45724# a_12791_45546# 8.97e-21
C17566 a_10807_43548# a_3483_46348# 1.08e-20
C17567 a_5565_43396# a_5257_43370# 2.14e-19
C17568 a_15037_43940# a_13059_46348# 4.6e-20
C17569 a_5891_43370# a_n357_42282# 0.304889f
C17570 a_20362_44736# a_8049_45260# 1.72e-21
C17571 a_5495_43940# a_2324_44458# 8.3e-21
C17572 a_n13_43084# a_n1613_43370# 4.63e-20
C17573 a_12089_42308# a_10227_46804# 5.68e-19
C17574 a_413_45260# DATA[3] 0.037695f
C17575 a_15368_46634# VDD 0.324877f
C17576 a_6123_31319# a_n3420_37440# 0.00105f
C17577 a_1823_45246# a_167_45260# 0.155648f
C17578 a_11813_46116# a_10586_45546# 7.37e-19
C17579 a_6755_46942# a_16375_45002# 8.39e-21
C17580 a_19123_46287# a_18985_46122# 0.215692f
C17581 a_18285_46348# a_19553_46090# 7.38e-22
C17582 a_16434_46987# a_10809_44734# 9.15e-19
C17583 a_20365_43914# a_743_42282# 0.001315f
C17584 a_20935_43940# a_4190_30871# 6.17e-21
C17585 a_21115_43940# a_21259_43561# 1.55e-19
C17586 a_20623_43914# a_20301_43646# 0.002259f
C17587 a_15037_43940# a_15095_43370# 1.6e-19
C17588 a_14021_43940# a_19268_43646# 0.007741f
C17589 a_19862_44208# a_21487_43396# 0.00184f
C17590 a_7542_44172# a_7871_42858# 6.14e-20
C17591 a_3422_30871# a_21671_42860# 0.199876f
C17592 a_1568_43370# a_1512_43396# 5.16e-20
C17593 a_4905_42826# a_3539_42460# 4.19e-20
C17594 a_n97_42460# a_6452_43396# 5.26e-20
C17595 a_n2293_43922# a_13291_42460# 5.94e-19
C17596 w_11334_34010# RST_Z 0.00509f
C17597 a_7112_43396# VDD 0.273193f
C17598 a_16223_45938# a_1307_43914# 2.89e-19
C17599 a_10193_42453# a_16922_45042# 0.035103f
C17600 a_6229_45572# a_n2661_43370# 4.04e-19
C17601 a_n2472_45002# a_n2293_45010# 0.177252f
C17602 a_n2661_45010# a_n2109_45247# 0.025907f
C17603 a_n2840_45002# a_n2017_45002# 1.31e-20
C17604 a_21487_43396# a_4185_45028# 2.21e-21
C17605 a_8685_43396# a_526_44458# 0.04962f
C17606 a_17303_42282# a_18597_46090# 4.04e-19
C17607 a_10341_43396# a_10809_44734# 4.7e-21
C17608 a_n2661_42834# CLK 3.56e-20
C17609 a_11823_42460# a_12465_44636# 0.127538f
C17610 a_11525_45546# a_11453_44696# 5.01e-19
C17611 a_13904_45546# a_13507_46334# 2.05e-20
C17612 a_8049_45260# a_16375_45002# 0.026933f
C17613 a_14205_43396# a_5342_30871# 1.54e-19
C17614 a_22223_43396# a_22591_43396# 7.52e-19
C17615 a_10341_43396# a_13460_43230# 3.71e-20
C17616 a_15095_43370# a_15279_43071# 0.105784f
C17617 a_12281_43396# a_12545_42858# 0.029151f
C17618 a_n97_42460# a_13291_42460# 0.419357f
C17619 a_21855_43396# a_17364_32525# 7.4e-20
C17620 a_4361_42308# a_20749_43396# 3.4e-19
C17621 a_14579_43548# a_16414_43172# 1.1e-20
C17622 a_2982_43646# a_3863_42891# 5.25e-19
C17623 a_5649_42852# a_14209_32519# 4.85e-19
C17624 a_n3420_37984# a_n2946_37984# 0.238664f
C17625 a_n3690_38304# a_n4064_37984# 0.085872f
C17626 a_6755_46942# RST_Z 1.33e-19
C17627 a_11136_42852# VDD 0.132515f
C17628 a_10775_45002# a_8975_43940# 4.88e-21
C17629 a_1307_43914# a_949_44458# 0.028157f
C17630 a_2711_45572# a_17737_43940# 0.005447f
C17631 a_2382_45260# a_n356_44636# 2.62e-19
C17632 a_327_44734# a_7_44811# 9.51e-20
C17633 a_2437_43646# a_n2661_43922# 0.033401f
C17634 a_5932_42308# a_4185_45028# 0.118319f
C17635 a_3905_42308# a_1823_45246# 0.003168f
C17636 a_17595_43084# a_n357_42282# 0.007854f
C17637 a_10341_42308# a_n443_42852# 2.65e-20
C17638 a_3080_42308# C8_P_btm 0.006767f
C17639 a_949_44458# a_n443_46116# 0.045448f
C17640 a_6298_44484# a_n1151_42308# 0.009717f
C17641 DATA[1] VDD 0.321585f
C17642 a_3175_45822# a_1823_45246# 2.41e-19
C17643 a_1609_45572# a_167_45260# 2.26e-19
C17644 a_17478_45572# a_15227_44166# 0.009301f
C17645 a_9482_43914# a_n2293_46634# 6.32e-20
C17646 a_3357_43084# a_7715_46873# 6.39e-20
C17647 a_3429_45260# a_2609_46660# 6.06e-22
C17648 a_3537_45260# a_2443_46660# 3.5e-19
C17649 a_5205_44484# a_2107_46812# 1.38e-20
C17650 a_3065_45002# a_3177_46902# 8.4e-21
C17651 a_18494_42460# a_18479_47436# 2.53e-21
C17652 a_19778_44110# a_18597_46090# 0.006796f
C17653 a_8387_43230# a_n784_42308# 2.3e-21
C17654 a_16137_43396# a_16522_42674# 0.001223f
C17655 a_4361_42308# a_8685_42308# 0.014949f
C17656 a_15743_43084# a_15803_42450# 1.96e-19
C17657 a_18083_42858# a_19273_43230# 2.56e-19
C17658 a_1847_42826# a_2123_42473# 0.004599f
C17659 a_18249_42858# a_17749_42852# 4.27e-20
C17660 a_743_42282# a_9377_42558# 0.00119f
C17661 a_8049_45260# RST_Z 0.002763f
C17662 a_12861_44030# a_12891_46348# 0.053595f
C17663 a_6851_47204# a_5807_45002# 7.21e-20
C17664 a_13717_47436# a_12549_44172# 0.002227f
C17665 a_n1435_47204# a_768_44030# 6.95e-20
C17666 a_16327_47482# a_n881_46662# 0.195459f
C17667 a_22223_47212# a_11453_44696# 0.057984f
C17668 a_12465_44636# a_22959_47212# 3.19e-20
C17669 a_22731_47423# SMPL_ON_N 0.194951f
C17670 a_n237_47217# a_1123_46634# 0.003027f
C17671 a_n1151_42308# a_n2472_46634# 1.07e-20
C17672 a_n2497_47436# a_n2661_46098# 0.026032f
C17673 a_327_47204# a_33_46660# 0.001418f
C17674 a_1431_47204# a_n2438_43548# 5.68e-21
C17675 a_n971_45724# a_2107_46812# 0.06261f
C17676 a_2063_45854# a_n1925_46634# 0.064288f
C17677 a_3381_47502# a_n2661_46634# 2.12e-20
C17678 a_n746_45260# a_948_46660# 0.001665f
C17679 a_2905_45572# a_n2293_46634# 8.29e-19
C17680 a_n3607_38528# VDD 2.79e-20
C17681 a_14539_43914# a_17061_44734# 0.020462f
C17682 a_18114_32519# a_22485_44484# 0.020813f
C17683 a_10193_42453# a_15743_43084# 0.027326f
C17684 a_9241_44734# a_9313_44734# 5.24e-19
C17685 a_1307_43914# a_11341_43940# 2.31482f
C17686 a_9482_43914# a_11816_44260# 0.003029f
C17687 a_16112_44458# a_17517_44484# 1.99e-21
C17688 a_13249_42308# a_13837_43396# 8.11e-20
C17689 a_3537_45260# a_6671_43940# 0.00223f
C17690 a_21887_42336# a_n357_42282# 3.8e-20
C17691 a_n4064_40160# a_n2810_45572# 7.36e-19
C17692 a_1423_45028# a_4185_45028# 0.016283f
C17693 a_n2661_43370# a_11415_45002# 0.092334f
C17694 a_5343_44458# a_3090_45724# 0.023693f
C17695 a_20980_44850# a_13747_46662# 0.001171f
C17696 a_16377_45572# a_13259_45724# 0.002102f
C17697 a_21363_45546# a_8049_45260# 0.013686f
C17698 a_11963_45334# a_9290_44172# 1.31e-19
C17699 a_9482_43914# a_9625_46129# 2.09e-19
C17700 a_644_44056# a_n1613_43370# 1.52e-20
C17701 a_6171_45002# a_15015_46420# 2.21e-20
C17702 a_5691_45260# a_2324_44458# 0.013607f
C17703 a_413_45260# a_6945_45028# 1.33e-19
C17704 a_1443_43940# a_n746_45260# 3.72e-20
C17705 a_6761_42308# a_8685_42308# 3.39e-20
C17706 a_7227_42308# a_8325_42308# 4.47e-20
C17707 a_14097_32519# a_13258_32519# 0.051815f
C17708 EN_VIN_BSTR_P C10_P_btm 0.320569f
C17709 EN_VIN_BSTR_N a_19120_35138# 0.652984f
C17710 a_11530_34132# a_19864_35138# 0.201937f
C17711 a_12549_44172# a_14035_46660# 0.026143f
C17712 a_13747_46662# a_19692_46634# 0.001071f
C17713 a_19594_46812# a_15227_44166# 0.073663f
C17714 a_n743_46660# a_11813_46116# 0.003585f
C17715 a_4646_46812# a_7411_46660# 0.266058f
C17716 a_4651_46660# a_5257_43370# 2.06e-19
C17717 a_5385_46902# a_5894_47026# 2.6e-19
C17718 a_4817_46660# a_5263_46660# 2.28e-19
C17719 a_19321_45002# a_19333_46634# 0.001085f
C17720 a_3877_44458# a_7715_46873# 2.82e-20
C17721 a_768_44030# a_13885_46660# 0.029614f
C17722 a_19452_47524# a_19466_46812# 4e-19
C17723 a_5807_45002# a_10425_46660# 2.9e-19
C17724 a_2583_47243# a_765_45546# 2e-19
C17725 a_11453_44696# a_20731_47026# 0.026307f
C17726 a_10227_46804# a_21297_46660# 6.03e-19
C17727 a_13507_46334# a_20719_46660# 7.51e-19
C17728 a_n1435_47204# a_1176_45822# 2.97e-20
C17729 a_4915_47217# a_5204_45822# 4.09e-20
C17730 a_4791_45118# a_6165_46155# 0.291653f
C17731 a_n1151_42308# a_5937_45572# 0.11638f
C17732 a_2063_45854# a_10355_46116# 9.15e-21
C17733 a_6298_44484# a_6197_43396# 0.002222f
C17734 a_11691_44458# a_14955_43396# 6.92e-19
C17735 a_4223_44672# a_8147_43396# 0.001199f
C17736 a_18579_44172# a_11341_43940# 0.030765f
C17737 a_5343_44458# a_6547_43396# 3.36e-21
C17738 a_10193_42453# a_1606_42308# 1.31e-19
C17739 a_2479_44172# a_3499_42826# 0.004494f
C17740 a_895_43940# a_2537_44260# 7.13e-20
C17741 a_21398_44850# a_19862_44208# 9.39e-19
C17742 a_9313_44734# a_14401_32519# 0.00363f
C17743 a_5111_44636# a_8952_43230# 1.01e-19
C17744 a_n1059_45260# a_18083_42858# 0.021784f
C17745 a_n913_45002# a_17701_42308# 1.16e-19
C17746 a_n2017_45002# a_17333_42852# 0.314084f
C17747 a_n310_44811# VDD 0.001779f
C17748 a_n3565_38502# a_n1386_35608# 1.73e-19
C17749 a_n4064_39072# C9_P_btm 7.29e-20
C17750 a_n3420_39072# C7_P_btm 9.48e-19
C17751 a_n3565_39304# C5_P_btm 3.17e-19
C17752 a_n4064_37440# a_n2810_45572# 1.13e-20
C17753 a_791_42968# a_584_46384# 4.57e-19
C17754 a_7871_42858# a_n971_45724# 2.7e-19
C17755 a_20365_43914# a_19466_46812# 5.98e-19
C17756 a_6031_43396# a_n2293_46634# 0.037881f
C17757 a_9145_43396# a_12549_44172# 6.67e-19
C17758 a_n2661_42834# a_n2956_39304# 5.57e-20
C17759 a_n2661_44458# a_n2661_45546# 0.032856f
C17760 a_n2840_44458# a_n2956_38216# 0.004419f
C17761 a_4361_42308# a_12861_44030# 0.005354f
C17762 a_19177_43646# a_16327_47482# 7.13e-19
C17763 a_19268_43646# a_13507_46334# 2.35e-21
C17764 a_n2293_43922# a_10809_44734# 2.24e-19
C17765 a_14673_44172# a_15015_46420# 2.63e-21
C17766 a_n3690_39392# a_n3690_38528# 0.050585f
C17767 a_1239_39043# comp_n 0.38743f
C17768 a_n3420_39072# a_n3565_38502# 0.034254f
C17769 a_1736_39587# a_1177_38525# 0.001279f
C17770 a_n4064_39072# a_n4209_38502# 0.030674f
C17771 a_n4209_39304# a_n4064_38528# 0.029379f
C17772 a_n3565_39304# a_n3420_38528# 0.028052f
C17773 a_n4064_39616# a_n4334_38304# 8e-19
C17774 a_2864_46660# VDD 0.076834f
C17775 COMP_P a_7754_40130# 1.45e-19
C17776 a_n881_46662# a_n356_45724# 0.002904f
C17777 a_10768_47026# a_10903_43370# 7.21e-21
C17778 a_11813_46116# a_11189_46129# 0.009001f
C17779 a_9863_46634# a_6945_45028# 1.05e-19
C17780 a_5807_45002# a_21167_46155# 1.15e-20
C17781 a_20273_46660# a_22365_46825# 7.72e-20
C17782 a_20841_46902# a_20885_46660# 3.69e-19
C17783 a_20623_46660# a_20719_46660# 0.013793f
C17784 a_18285_46348# a_12741_44636# 8.73e-21
C17785 a_20411_46873# a_20202_43084# 1.99e-21
C17786 a_20107_46660# a_11415_45002# 2.81e-22
C17787 a_12429_44172# a_9145_43396# 1.63e-19
C17788 a_22485_44484# a_13887_32519# 5.15e-23
C17789 a_10807_43548# a_10695_43548# 0.159782f
C17790 a_9313_44734# a_18817_42826# 0.003505f
C17791 a_14401_32519# a_20974_43370# 0.118041f
C17792 a_20193_45348# a_14097_32519# 4.63e-20
C17793 a_20512_43084# a_22591_43396# 5.83e-19
C17794 en_comp a_20712_42282# 4.59e-20
C17795 a_n913_45002# a_21613_42308# 0.259761f
C17796 a_9801_43940# VDD 0.19512f
C17797 a_6667_45809# a_1423_45028# 8.66e-22
C17798 a_10193_42453# a_10775_45002# 1.13e-21
C17799 a_18175_45572# a_18787_45572# 3.82e-19
C17800 a_16147_45260# a_18953_45572# 2.59e-20
C17801 a_10180_45724# a_10951_45334# 6.34e-19
C17802 a_17478_45572# a_2437_43646# 1.42e-21
C17803 a_12791_45546# a_6171_45002# 9.74e-21
C17804 a_8746_45002# a_8953_45002# 0.257529f
C17805 a_10807_43548# a_n357_42282# 0.031251f
C17806 a_3499_42826# a_n443_42852# 0.023367f
C17807 a_6197_43396# a_5937_45572# 2.15e-19
C17808 a_3080_42308# a_2324_44458# 1.53e-21
C17809 a_3626_43646# a_10903_43370# 0.001928f
C17810 a_n3674_37592# a_n2312_40392# 0.035844f
C17811 a_22469_40625# RST_Z 8.08e-20
C17812 a_20708_46348# VDD 0.093079f
C17813 a_7499_43078# a_2063_45854# 0.478913f
C17814 a_1990_45572# a_n443_46116# 3.19e-20
C17815 a_7227_45028# a_6151_47436# 0.006424f
C17816 a_2711_45572# a_9313_45822# 0.016843f
C17817 a_6667_45809# a_6491_46660# 1.51e-21
C17818 a_6598_45938# a_6545_47178# 9.57e-19
C17819 a_6511_45714# a_6851_47204# 1.94e-21
C17820 a_6472_45840# a_7227_47204# 4.49e-20
C17821 a_167_45260# a_n2293_45546# 0.681309f
C17822 a_n2293_46098# a_n23_45546# 0.00525f
C17823 a_472_46348# a_n357_42282# 0.001836f
C17824 a_2804_46116# a_n2661_45546# 1.07e-20
C17825 a_1823_45246# a_n863_45724# 0.207189f
C17826 a_376_46348# a_n755_45592# 1.77e-21
C17827 a_1176_45822# a_380_45546# 2.97e-19
C17828 a_18985_46122# a_8049_45260# 0.006692f
C17829 a_13759_46122# a_12638_46436# 1.15e-20
C17830 a_10903_43370# a_11601_46155# 2.78e-19
C17831 a_2675_43914# a_2713_42308# 8.11e-22
C17832 a_14205_43396# a_743_42282# 2.22e-20
C17833 a_16243_43396# a_18783_43370# 2.36e-21
C17834 a_3626_43646# a_3681_42891# 0.001623f
C17835 a_16137_43396# a_15743_43084# 0.029757f
C17836 a_2982_43646# a_4520_42826# 3.49e-20
C17837 a_n2661_42282# a_n2840_42282# 0.173771f
C17838 a_n97_42460# a_13460_43230# 1.61e-19
C17839 a_16977_43638# a_17324_43396# 0.051162f
C17840 a_16409_43396# a_18429_43548# 1.76e-19
C17841 a_n3674_39768# a_n1630_35242# 1.64e-19
C17842 a_10341_43396# a_19177_43646# 2.93e-19
C17843 a_n3420_37984# C1_P_btm 1.26e-19
C17844 a_n2956_39768# CLK_DATA 0.015401f
C17845 a_12545_42858# VDD 0.285703f
C17846 a_18479_45785# a_18248_44752# 0.002693f
C17847 a_18175_45572# a_18287_44626# 2.34e-19
C17848 a_1423_45028# a_2448_45028# 6.07e-21
C17849 a_n2840_45002# a_n2840_44458# 0.025171f
C17850 a_6171_45002# a_16405_45348# 2.48e-19
C17851 a_12563_42308# a_3090_45724# 4.38e-21
C17852 a_n2946_38778# a_n2312_38680# 0.024631f
C17853 a_n2293_42282# a_n2956_39304# 4.17e-20
C17854 a_13467_32519# a_n357_42282# 0.002449f
C17855 a_15940_43402# a_n443_42852# 0.005303f
C17856 a_10553_43218# a_9290_44172# 0.002152f
C17857 VDAC_Pi w_1575_34946# 5.84e-19
C17858 a_10210_45822# a_10428_46928# 2.06e-20
C17859 a_4880_45572# a_3090_45724# 0.002202f
C17860 a_2437_43646# a_19594_46812# 0.003991f
C17861 a_3357_43084# a_13747_46662# 7.23e-19
C17862 a_n2017_45002# a_768_44030# 1.14e-19
C17863 a_n1059_45260# a_12549_44172# 2.03e-19
C17864 a_n143_45144# a_n881_46662# 7.46e-19
C17865 a_14537_43396# a_10227_46804# 0.094463f
C17866 a_8953_45002# a_4883_46098# 0.013985f
C17867 a_1307_43914# a_16327_47482# 3.53e-20
C17868 a_8037_42858# a_8292_43218# 0.064178f
C17869 a_18817_42826# a_18599_43230# 0.209641f
C17870 a_18083_42858# a_19987_42826# 6.28e-21
C17871 a_18249_42858# a_19339_43156# 0.042415f
C17872 a_3626_43646# a_15959_42545# 0.005102f
C17873 a_5111_42852# a_5193_42852# 0.171361f
C17874 a_17333_42852# a_19164_43230# 3.85e-20
C17875 a_4190_30871# a_19326_42852# 1.16e-19
C17876 a_19332_42282# VDD 0.227361f
C17877 a_n1741_47186# a_n89_47570# 3.69e-19
C17878 a_n1605_47204# a_n2312_39304# 0.001342f
C17879 a_11031_47542# a_11459_47204# 0.001175f
C17880 a_9067_47204# a_n1435_47204# 0.001005f
C17881 a_6151_47436# a_15507_47210# 0.003878f
C17882 a_11691_44458# a_n2661_42834# 0.018854f
C17883 a_1307_43914# a_175_44278# 8.72e-21
C17884 a_5343_44458# a_n356_44636# 5.46e-20
C17885 a_n2661_44458# a_8238_44734# 5.96e-19
C17886 a_7229_43940# a_7845_44172# 1.1e-20
C17887 a_n2017_45002# a_13483_43940# 1.15e-21
C17888 a_n913_45002# a_11750_44172# 9.36e-22
C17889 a_2382_45260# a_3820_44260# 0.001415f
C17890 a_13657_42558# a_13259_45724# 0.023664f
C17891 a_5934_30871# a_n863_45724# 2.07e-20
C17892 a_3318_42354# a_n443_42852# 1.12e-21
C17893 a_n3565_39590# a_n2956_39304# 0.072956f
C17894 a_10210_45822# VDD 0.323342f
C17895 a_3905_42865# a_584_46384# 4.97e-20
C17896 a_1241_44260# a_n2497_47436# 0.001773f
C17897 a_n3674_39768# a_n971_45724# 2.61e-20
C17898 a_n37_45144# a_n2293_46098# 4.54e-20
C17899 a_n2661_45010# a_167_45260# 6.95e-20
C17900 a_n467_45028# a_n1853_46287# 1.67e-19
C17901 a_10193_42453# a_12839_46116# 2.22e-20
C17902 a_1609_45572# a_n863_45724# 1.88e-19
C17903 a_5907_45546# a_n2661_45546# 3.27e-19
C17904 a_20640_44752# a_18479_47436# 0.018112f
C17905 a_20159_44458# a_18597_46090# 1.48e-20
C17906 a_18579_44172# a_16327_47482# 0.043297f
C17907 a_17061_44734# a_11453_44696# 0.005756f
C17908 a_2437_43646# a_5164_46348# 3.03e-20
C17909 a_17786_45822# a_17715_44484# 0.001664f
C17910 a_16147_45260# a_17583_46090# 1.41e-20
C17911 a_22959_42860# a_13258_32519# 7.81e-21
C17912 a_1067_42314# a_1576_42282# 0.017282f
C17913 a_n1630_35242# a_1184_42692# 0.003096f
C17914 a_n784_42308# a_1606_42308# 15.027599f
C17915 a_564_42282# a_961_42354# 0.003943f
C17916 a_21195_42852# a_21335_42336# 8.75e-20
C17917 COMP_P a_n39_42308# 5.96e-21
C17918 a_3080_42308# a_2113_38308# 1.02e-19
C17919 a_11599_46634# a_19692_46634# 0.069066f
C17920 a_16327_47482# a_17609_46634# 0.001241f
C17921 a_10227_46804# a_3090_45724# 0.320681f
C17922 a_16023_47582# a_16292_46812# 7.28e-19
C17923 a_3381_47502# a_765_45546# 0.002383f
C17924 a_8128_46384# a_7715_46873# 0.006283f
C17925 a_n881_46662# a_8667_46634# 5.47e-20
C17926 a_n1925_46634# a_645_46660# 4.33e-19
C17927 a_n2438_43548# a_n935_46688# 6.37e-19
C17928 a_383_46660# a_948_46660# 7.99e-20
C17929 a_n2104_46634# a_n2661_46098# 1.32e-19
C17930 a_171_46873# a_288_46660# 0.159893f
C17931 a_n133_46660# a_491_47026# 9.73e-19
C17932 a_n2293_46634# a_2443_46660# 1.47e-20
C17933 a_n2661_46634# a_2959_46660# 0.006729f
C17934 a_5807_45002# a_4651_46660# 8.13e-19
C17935 a_18248_44752# a_14021_43940# 1.74e-20
C17936 a_5883_43914# a_5829_43940# 0.009634f
C17937 a_n2661_42834# a_8333_44056# 0.007771f
C17938 a_9313_44734# a_15682_43940# 1.54e-19
C17939 a_18114_32519# a_14401_32519# 0.087478f
C17940 a_n2293_42834# a_8147_43396# 7.84e-19
C17941 a_20512_43084# a_22591_44484# 2.48e-20
C17942 a_14539_43914# a_15301_44260# 6.38e-21
C17943 a_7499_43078# a_10793_43218# 3.95e-19
C17944 a_1307_43914# a_10341_43396# 2.19e-19
C17945 a_n913_45002# a_4361_42308# 0.250497f
C17946 a_21101_45002# VDD 0.2903f
C17947 a_8375_44464# a_3483_46348# 0.003197f
C17948 a_15463_44811# a_12741_44636# 2.47e-19
C17949 a_18797_44260# a_13661_43548# 0.002056f
C17950 a_7845_44172# a_8270_45546# 1.29e-19
C17951 a_13777_45326# a_n443_42852# 1.94e-21
C17952 a_19778_44110# a_8049_45260# 2.13e-20
C17953 a_2232_45348# a_n755_45592# 1.57e-19
C17954 a_13720_44458# a_13925_46122# 1.08e-20
C17955 a_10057_43914# a_2324_44458# 1.41e-19
C17956 a_104_43370# a_n1613_43370# 1.95e-19
C17957 a_3626_43646# a_4883_46098# 4.8e-20
C17958 a_5742_30871# a_n4209_38216# 4.02e-21
C17959 a_n784_42308# C1_N_btm 0.027772f
C17960 a_4955_46873# a_3483_46348# 1.84e-20
C17961 a_4646_46812# a_4185_45028# 1.6e-20
C17962 a_3090_45724# a_17339_46660# 0.019979f
C17963 a_15227_44166# a_16388_46812# 0.02839f
C17964 a_15009_46634# a_765_45546# 6.36e-21
C17965 a_14976_45028# a_15312_46660# 0.01024f
C17966 a_16292_46812# a_16751_46987# 6.64e-19
C17967 a_768_44030# a_526_44458# 0.341438f
C17968 a_n881_46662# a_6640_46482# 6.85e-19
C17969 a_20916_46384# a_6945_45028# 0.036695f
C17970 a_n743_46660# a_15682_46116# 0.051046f
C17971 a_n2438_43548# a_2324_44458# 0.00362f
C17972 a_20843_47204# a_10809_44734# 9.21e-19
C17973 a_13507_46334# a_14537_46482# 7.17e-19
C17974 a_16327_47482# a_19443_46116# 0.012553f
C17975 a_18597_46090# a_18243_46436# 6.59e-20
C17976 a_10227_46804# a_15002_46116# 4.37e-19
C17977 a_n443_46116# a_n356_45724# 0.113738f
C17978 a_n1151_42308# a_n443_42852# 0.001061f
C17979 a_2905_45572# a_2277_45546# 5.92e-19
C17980 a_3877_44458# a_4419_46090# 6.31e-19
C17981 a_10157_44484# a_10083_42826# 1.72e-19
C17982 a_15493_43396# a_19319_43548# 0.120111f
C17983 a_17517_44484# a_17499_43370# 1.98e-19
C17984 a_11967_42832# a_15681_43442# 1.86e-19
C17985 a_18579_44172# a_10341_43396# 0.023217f
C17986 a_9313_44734# a_22223_43396# 1.02e-20
C17987 a_11341_43940# a_10867_43940# 3.41e-19
C17988 a_2382_45260# a_3823_42558# 0.058499f
C17989 a_n913_45002# a_6761_42308# 0.350952f
C17990 a_n1059_45260# a_7227_42308# 1.26e-19
C17991 a_n2017_45002# a_6123_31319# 0.007053f
C17992 a_3065_45002# a_2903_42308# 2.87e-19
C17993 a_10907_45822# a_12649_45572# 4.44e-21
C17994 a_8791_45572# a_8696_44636# 1.87e-19
C17995 a_1184_42692# a_n971_45724# 2.87e-20
C17996 a_14955_43396# a_15227_44166# 0.001876f
C17997 a_10796_42968# a_n2293_46634# 6.09e-20
C17998 a_15567_42826# a_13661_43548# 1.39e-23
C17999 a_19987_42826# a_12549_44172# 6.54e-20
C18000 a_12991_43230# a_10227_46804# 1.79e-19
C18001 a_14021_43940# a_2324_44458# 8.72e-19
C18002 a_18057_42282# CAL_N 3.79e-19
C18003 a_17303_42282# a_22469_40625# 4.4e-19
C18004 a_18285_46348# a_16375_45002# 0.003864f
C18005 a_376_46348# a_835_46155# 6.64e-19
C18006 a_472_46348# a_518_46155# 0.006879f
C18007 a_20820_30879# a_8049_45260# 1.76e-19
C18008 a_18079_43940# a_17333_42852# 1.33e-20
C18009 a_18326_43940# a_18083_42858# 1e-20
C18010 a_3626_43646# a_16243_43396# 5.34e-20
C18011 a_2982_43646# a_16409_43396# 5.61e-21
C18012 a_20974_43370# a_22223_43396# 0.04256f
C18013 a_11341_43940# a_13635_43156# 3.77e-20
C18014 a_5891_43370# a_8685_42308# 0.048111f
C18015 a_n356_44636# a_12563_42308# 2.77e-19
C18016 a_14401_32519# a_13887_32519# 0.07508f
C18017 a_9396_43370# a_10341_43396# 5.02e-19
C18018 a_21845_43940# a_13678_32519# 1.2e-19
C18019 a_8685_43396# a_8317_43396# 2.29e-19
C18020 a_18780_47178# RST_Z 1.31e-19
C18021 SMPL_ON_N EN_VIN_BSTR_N 1.61e-19
C18022 a_15811_47375# CLK 4.17e-19
C18023 a_18479_47436# START 0.313639f
C18024 a_18479_45785# a_16922_45042# 0.02321f
C18025 a_16147_45260# a_17613_45144# 0.028566f
C18026 a_15861_45028# a_11691_44458# 2.17e-19
C18027 a_11823_42460# a_12883_44458# 0.026633f
C18028 a_10193_42453# a_17970_44736# 9.16e-19
C18029 a_6511_45714# a_7640_43914# 3.14e-19
C18030 a_7276_45260# a_7229_43940# 0.322065f
C18031 a_5205_44484# a_6709_45028# 0.095031f
C18032 a_6171_45002# a_8191_45002# 0.024424f
C18033 a_3232_43370# a_8953_45002# 0.012103f
C18034 a_15567_42826# a_4185_45028# 9.4e-21
C18035 a_5932_42308# a_5257_43370# 3.61e-20
C18036 a_6197_43396# a_n443_42852# 0.007993f
C18037 a_2075_43172# a_2324_44458# 1.36e-20
C18038 a_8952_43230# a_9290_44172# 2.21e-19
C18039 a_10341_42308# a_8199_44636# 1.19e-19
C18040 a_n4064_39072# a_n2312_39304# 0.094407f
C18041 a_n143_45144# a_n443_46116# 0.001224f
C18042 a_413_45260# a_4700_47436# 8.97e-20
C18043 a_3429_45260# a_2905_45572# 4.46e-19
C18044 a_4558_45348# a_2063_45854# 8.06e-22
C18045 a_3065_45002# a_3160_47472# 1.34e-21
C18046 a_13904_45546# a_n743_46660# 1.24e-20
C18047 a_5263_45724# a_5167_46660# 4.57e-21
C18048 a_6667_45809# a_4646_46812# 3.86e-19
C18049 a_6598_45938# a_3877_44458# 4.85e-19
C18050 a_15599_45572# a_12549_44172# 5.18e-22
C18051 a_21188_45572# a_18479_47436# 0.005114f
C18052 a_20731_45938# a_10227_46804# 8.16e-20
C18053 a_20885_45572# a_16327_47482# 0.002535f
C18054 a_20623_45572# a_18597_46090# 0.046479f
C18055 a_2437_43646# a_15673_47210# 0.007104f
C18056 a_3357_43084# a_11599_46634# 9.81e-19
C18057 a_20107_45572# a_20894_47436# 1.49e-21
C18058 a_19431_45546# a_11453_44696# 3.07e-21
C18059 a_16020_45572# a_n881_46662# 0.013745f
C18060 a_n2661_45546# a_n1099_45572# 0.068604f
C18061 a_n2293_45546# a_n863_45724# 0.17075f
C18062 a_20269_44172# a_20107_42308# 3.94e-19
C18063 a_20365_43914# a_13258_32519# 6.32e-21
C18064 a_4699_43561# a_1755_42282# 2.85e-21
C18065 a_21487_43396# a_21671_42860# 3.61e-19
C18066 a_5649_42852# a_19339_43156# 2.62e-21
C18067 a_4361_42308# a_20922_43172# 0.00325f
C18068 a_13467_32519# a_21356_42826# 0.001409f
C18069 a_n1557_42282# a_961_42354# 1.02e-20
C18070 a_3539_42460# a_n784_42308# 2.97e-20
C18071 a_19862_44208# a_20712_42282# 3.07e-21
C18072 a_3080_42308# a_1606_42308# 4.87174f
C18073 a_15095_43370# a_15785_43172# 0.002407f
C18074 a_n4209_37414# a_n4334_37440# 0.253282f
C18075 a_13059_46348# CLK 2.07e-20
C18076 a_18285_46348# RST_Z 1.19e-20
C18077 a_5379_42460# VDD 0.213136f
C18078 a_18494_42460# CAL_N 0.001361f
C18079 a_n746_45260# a_n237_47217# 0.285294f
C18080 a_n971_45724# a_n23_47502# 0.225828f
C18081 a_n452_47436# a_n785_47204# 0.03755f
C18082 a_n1741_47186# a_1431_47204# 0.014137f
C18083 a_n2109_47186# a_584_46384# 0.352889f
C18084 a_n815_47178# a_327_47204# 1.12e-19
C18085 a_8696_44636# a_9028_43914# 4.56e-21
C18086 a_14537_43396# a_14815_43914# 0.015948f
C18087 a_1307_43914# a_n2293_43922# 0.022859f
C18088 a_13249_42308# a_13565_44260# 0.002149f
C18089 a_375_42282# a_n2661_42834# 0.035547f
C18090 a_20712_42282# a_4185_45028# 1.64e-19
C18091 a_6123_31319# a_526_44458# 1.83e-19
C18092 a_22400_42852# a_20205_31679# 4.56e-20
C18093 a_20273_45572# a_20107_46660# 0.001469f
C18094 a_16211_45572# a_11415_45002# 8.47e-19
C18095 a_1423_45028# a_5257_43370# 0.020778f
C18096 a_n2661_43370# a_1799_45572# 9.48e-20
C18097 a_20107_45572# a_20411_46873# 0.001307f
C18098 a_9482_43914# a_6755_46942# 0.01168f
C18099 a_11691_44458# a_19321_45002# 0.064467f
C18100 a_16886_45144# a_13661_43548# 2.62e-21
C18101 a_17023_45118# a_n743_46660# 5.2e-19
C18102 a_413_45260# a_15559_46634# 2.31e-21
C18103 a_2437_43646# a_16388_46812# 1.36e-19
C18104 a_10180_45724# a_2324_44458# 0.064932f
C18105 a_12791_45546# a_10903_43370# 0.042213f
C18106 a_12427_45724# a_12594_46348# 0.040872f
C18107 a_11823_42460# a_12005_46116# 0.010777f
C18108 a_13249_42308# a_9290_44172# 0.033421f
C18109 a_8336_45822# a_8199_44636# 2.62e-19
C18110 a_6977_45572# a_5937_45572# 4.29e-19
C18111 a_949_44458# a_n1613_43370# 6.55e-22
C18112 a_13076_44458# a_11453_44696# 9.33e-21
C18113 a_14539_43914# a_12465_44636# 0.054102f
C18114 a_18248_44752# a_13507_46334# 1.76e-21
C18115 a_n356_44636# a_10227_46804# 4.54e-19
C18116 a_13678_32519# a_21973_42336# 3.77e-19
C18117 a_12379_42858# a_12563_42308# 2.54e-20
C18118 a_22959_43396# a_22775_42308# 2.94e-20
C18119 a_12089_42308# a_11633_42558# 0.003531f
C18120 a_5649_42852# a_22465_38105# 7.91e-21
C18121 a_3080_42308# C1_N_btm 0.011373f
C18122 a_768_44030# a_13759_47204# 5.98e-19
C18123 a_6491_46660# a_5257_43370# 0.1719f
C18124 a_6151_47436# a_7715_46873# 0.025823f
C18125 a_n1435_47204# a_5167_46660# 2.1e-20
C18126 a_n1151_42308# a_10554_47026# 2.53e-20
C18127 a_n1741_47186# a_11735_46660# 0.029236f
C18128 a_2063_45854# a_6999_46987# 4.27e-21
C18129 a_16922_45042# a_14021_43940# 0.11663f
C18130 a_11827_44484# a_22223_43948# 0.003019f
C18131 a_21359_45002# a_15493_43940# 8.21e-21
C18132 a_1307_43914# a_n97_42460# 0.23336f
C18133 a_20193_45348# a_20365_43914# 0.025746f
C18134 a_22223_45036# a_11341_43940# 7.11e-20
C18135 a_375_42282# a_n1352_43396# 9.86e-21
C18136 a_18479_45785# a_15743_43084# 0.001697f
C18137 a_7499_43078# a_10083_42826# 0.375624f
C18138 a_9313_44734# a_20512_43084# 0.028182f
C18139 a_14673_44172# a_16241_44484# 9.76e-19
C18140 a_4223_44672# a_n2661_42282# 0.064384f
C18141 a_17517_44484# a_18204_44850# 6.24e-19
C18142 a_n356_44636# a_453_43940# 0.02089f
C18143 a_2711_45572# a_18817_42826# 0.001093f
C18144 a_3232_43370# a_3626_43646# 0.204337f
C18145 a_14797_45144# VDD 0.124624f
C18146 a_n1630_35242# a_19120_35138# 7.97e-19
C18147 a_n784_42308# C9_P_btm 9.31e-20
C18148 a_22469_40625# a_20820_30879# 2.62e-20
C18149 a_n229_43646# a_n1151_42308# 4.13e-20
C18150 a_n97_42460# a_n443_46116# 0.131756f
C18151 a_4093_43548# a_584_46384# 0.00472f
C18152 a_n1177_44458# a_n1423_46090# 9.12e-21
C18153 a_949_44458# a_n2293_46098# 4.44e-20
C18154 a_14815_43914# a_3090_45724# 9.92e-21
C18155 a_18326_43940# a_12549_44172# 0.013334f
C18156 a_10951_45334# a_10586_45546# 2.24e-20
C18157 a_9482_43914# a_8049_45260# 2.04e-21
C18158 a_3495_45348# a_526_44458# 0.002123f
C18159 a_18533_43940# a_12861_44030# 1.12e-19
C18160 a_13711_45394# a_2324_44458# 6.14e-19
C18161 en_comp a_20692_30879# 2.56e-19
C18162 a_2437_43646# a_3316_45546# 7.08e-22
C18163 a_n1059_45260# a_n2661_45546# 0.003807f
C18164 a_n2293_45010# a_n2293_45546# 0.257189f
C18165 a_n2661_45010# a_n863_45724# 0.345234f
C18166 a_3815_47204# VDD 0.260661f
C18167 a_15803_42450# a_16104_42674# 9.73e-19
C18168 a_15764_42576# a_16522_42674# 0.05936f
C18169 a_9223_42460# a_7174_31319# 4.88e-21
C18170 a_n4318_37592# a_n4064_38528# 0.020352f
C18171 a_15051_42282# a_15521_42308# 0.007399f
C18172 a_14113_42308# a_15761_42308# 9.35e-19
C18173 a_n1613_43370# a_5497_46414# 0.003931f
C18174 a_11453_44696# a_12594_46348# 2.02e-20
C18175 a_12465_44636# a_14493_46090# 0.008365f
C18176 a_4883_46098# a_15015_46420# 0.010147f
C18177 a_13507_46334# a_2324_44458# 0.033576f
C18178 a_10227_46804# a_20075_46420# 1.19e-20
C18179 a_18479_47436# a_19553_46090# 1.71e-19
C18180 a_18597_46090# a_18819_46122# 0.230891f
C18181 a_16241_47178# a_10809_44734# 7.12e-21
C18182 a_16023_47582# a_6945_45028# 0.00884f
C18183 a_4791_45118# a_5210_46155# 6.75e-22
C18184 a_n881_46662# a_5204_45822# 0.089827f
C18185 a_2959_46660# a_765_45546# 0.002438f
C18186 a_6755_46942# a_12816_46660# 0.061031f
C18187 a_768_44030# a_2521_46116# 0.008186f
C18188 a_15682_43940# a_17737_43940# 1.13e-19
C18189 a_22485_44484# a_14401_32519# 0.01705f
C18190 a_5891_43370# a_9803_43646# 0.011447f
C18191 a_14539_43914# a_16409_43396# 0.031761f
C18192 a_18579_44172# a_n97_42460# 0.005302f
C18193 a_20512_43084# a_20974_43370# 0.020132f
C18194 a_375_42282# a_n2293_42282# 5.08e-19
C18195 a_13249_42308# a_15051_42282# 4.99e-21
C18196 a_11823_42460# a_15890_42674# 1.45e-19
C18197 a_3905_42865# a_5025_43940# 4.14e-19
C18198 a_18114_32519# a_22223_43396# 4.85e-19
C18199 a_n2017_45002# a_15597_42852# 0.004498f
C18200 a_5111_44636# a_8495_42852# 2.05e-20
C18201 a_n1059_45260# a_14853_42852# 0.003368f
C18202 a_n913_45002# a_13622_42852# 4.2e-19
C18203 a_19479_31679# a_22400_42852# 3.1e-20
C18204 a_20766_44850# VDD 0.197657f
C18205 a_11525_45546# a_11962_45724# 0.095856f
C18206 a_10490_45724# a_11823_42460# 0.022778f
C18207 a_11322_45546# a_12427_45724# 0.010517f
C18208 a_2711_45572# a_14033_45822# 7.91e-19
C18209 a_10949_43914# a_3483_46348# 1.95e-20
C18210 a_4190_30871# a_19321_45002# 6.81e-20
C18211 a_13565_43940# a_13059_46348# 0.011241f
C18212 a_20556_43646# a_13661_43548# 8.75e-19
C18213 a_20159_44458# a_8049_45260# 6.75e-22
C18214 a_5013_44260# a_2324_44458# 1.86e-20
C18215 a_n1076_43230# a_n1613_43370# 0.224215f
C18216 a_12379_42858# a_10227_46804# 0.298444f
C18217 a_413_45260# DATA[2] 0.048779f
C18218 a_14976_45028# VDD 0.484864f
C18219 a_1138_42852# a_167_45260# 0.250282f
C18220 a_1823_45246# a_2202_46116# 0.25354f
C18221 a_11735_46660# a_10586_45546# 0.001215f
C18222 a_1799_45572# a_2307_45899# 1.33e-19
C18223 a_19123_46287# a_18819_46122# 0.172712f
C18224 a_16721_46634# a_10809_44734# 0.004449f
C18225 a_18285_46348# a_18985_46122# 5.57e-21
C18226 a_7542_44172# a_7227_42852# 2.27e-20
C18227 a_20365_43914# a_20301_43646# 0.001115f
C18228 a_20269_44172# a_743_42282# 7.1e-21
C18229 a_20623_43914# a_4190_30871# 6.24e-20
C18230 a_4905_42826# a_3626_43646# 1.99e-19
C18231 a_n97_42460# a_9396_43370# 1.44e-20
C18232 a_14021_43940# a_15743_43084# 0.045789f
C18233 a_3422_30871# a_21195_42852# 0.289298f
C18234 a_3080_42308# a_3539_42460# 0.037567f
C18235 a_15493_43396# a_19095_43396# 1.29e-19
C18236 a_19862_44208# a_20556_43646# 0.009839f
C18237 a_9313_44734# a_16245_42852# 2.19e-19
C18238 a_1568_43370# a_648_43396# 4.6e-20
C18239 a_15493_43940# a_16823_43084# 6.79e-20
C18240 w_1575_34946# RST_Z 0.001495f
C18241 a_7287_43370# VDD 0.457521f
C18242 a_10193_42453# a_16501_45348# 0.009694f
C18243 a_n2661_45010# a_n2293_45010# 0.400159f
C18244 a_n4209_38502# SMPL_ON_P 0.001002f
C18245 a_5534_30871# a_13059_46348# 1.92e-19
C18246 a_21887_42336# a_12861_44030# 2.1e-21
C18247 a_8415_44056# a_n443_42852# 1.8e-19
C18248 a_n4318_39304# a_n2810_45572# 0.023142f
C18249 a_19319_43548# a_n357_42282# 1.18e-21
C18250 a_18051_46116# VDD 0.189782f
C18251 a_4099_45572# a_768_44030# 4.61e-22
C18252 a_11322_45546# a_11453_44696# 0.004775f
C18253 a_12427_45724# a_12465_44636# 1.45e-19
C18254 a_12791_45546# a_4883_46098# 8.52e-20
C18255 a_13527_45546# a_13507_46334# 0.001293f
C18256 a_n1925_42282# a_n2661_45546# 0.181908f
C18257 a_12379_46436# a_12638_46436# 0.093752f
C18258 a_14358_43442# a_5342_30871# 2.31e-19
C18259 a_5649_42852# a_22591_43396# 2.81e-19
C18260 a_22223_43396# a_13887_32519# 0.154411f
C18261 a_12281_43396# a_12089_42308# 0.210903f
C18262 a_10341_43396# a_13635_43156# 2.32e-19
C18263 a_15095_43370# a_5534_30871# 1.69e-19
C18264 a_13678_32519# a_14209_32519# 0.048492f
C18265 a_4361_42308# a_17364_32525# 4.28e-20
C18266 a_14579_43548# a_15567_42826# 4.33e-19
C18267 a_n2661_42282# a_5742_30871# 3.56e-20
C18268 a_8667_46634# DATA[4] 3.49e-19
C18269 a_10775_45002# a_10057_43914# 0.010331f
C18270 a_2711_45572# a_15682_43940# 0.038198f
C18271 a_1307_43914# a_742_44458# 0.355379f
C18272 a_8953_45002# a_8975_43940# 0.001233f
C18273 a_n913_45002# a_5891_43370# 0.255618f
C18274 a_327_44734# a_n310_44811# 1.25e-19
C18275 a_2437_43646# a_n2661_42834# 0.033942f
C18276 a_6171_42473# a_4185_45028# 6.87e-20
C18277 a_18727_42674# a_17339_46660# 8.21e-21
C18278 a_16795_42852# a_n357_42282# 0.180926f
C18279 a_3080_42308# C9_P_btm 9.33e-20
C18280 a_742_44458# a_n443_46116# 0.018829f
C18281 DATA[0] VDD 1.05526f
C18282 a_2711_45572# a_1823_45246# 0.262616f
C18283 a_10951_45334# a_n743_46660# 3.01e-20
C18284 a_1423_45028# a_5807_45002# 2.15e-19
C18285 a_15861_45028# a_15227_44166# 0.208121f
C18286 a_18911_45144# a_18597_46090# 4.8e-20
C18287 a_16922_45042# a_13507_46334# 4.88e-20
C18288 a_14309_45028# a_12465_44636# 0.001972f
C18289 a_413_45260# a_3067_47026# 0.005586f
C18290 a_3065_45002# a_2609_46660# 4.49e-20
C18291 a_3429_45260# a_2443_46660# 2.96e-21
C18292 a_3357_43084# a_7411_46660# 2.31e-20
C18293 a_2437_43646# a_8145_46902# 8.67e-21
C18294 a_1847_42826# a_1755_42282# 2.18e-19
C18295 a_8605_42826# a_n784_42308# 4.32e-21
C18296 a_15743_43084# a_15764_42576# 0.006278f
C18297 a_2075_43172# a_1606_42308# 4.06e-19
C18298 a_4361_42308# a_8325_42308# 0.020707f
C18299 a_16664_43396# a_14113_42308# 2.4e-20
C18300 a_13887_32519# a_5934_30871# 2.14e-19
C18301 a_5534_30871# a_14097_32519# 0.041746f
C18302 a_17333_42852# a_17749_42852# 0.002387f
C18303 a_18249_42858# a_17665_42852# 3.34e-20
C18304 a_743_42282# a_9293_42558# 9.79e-19
C18305 a_n4251_38528# VDD 3.95e-19
C18306 a_6151_47436# a_13747_46662# 1.38e-19
C18307 a_n1435_47204# a_12549_44172# 0.072753f
C18308 a_6491_46660# a_5807_45002# 0.01567f
C18309 a_13717_47436# a_12891_46348# 3.83e-20
C18310 a_13381_47204# a_768_44030# 5.3e-20
C18311 a_16241_47178# a_n881_46662# 1.39e-21
C18312 a_12465_44636# a_11453_44696# 0.084038f
C18313 a_22223_47212# SMPL_ON_N 0.00103f
C18314 a_n971_45724# a_948_46660# 6.67e-20
C18315 a_n237_47217# a_383_46660# 3.31e-20
C18316 a_n2833_47464# a_n2661_46098# 1.96e-20
C18317 a_n785_47204# a_33_46660# 0.008206f
C18318 a_1239_47204# a_n2438_43548# 1.77e-19
C18319 a_1431_47204# a_n743_46660# 0.00119f
C18320 a_584_46384# a_n1925_46634# 0.047378f
C18321 a_n1151_42308# a_n2661_46634# 0.832521f
C18322 a_n746_45260# a_1123_46634# 4.1e-19
C18323 a_n2497_47436# a_1799_45572# 1.83e-20
C18324 a_15415_45028# a_15493_43940# 1.94e-21
C18325 a_10193_42453# a_18783_43370# 0.007846f
C18326 a_6109_44484# a_5708_44484# 0.002689f
C18327 a_14539_43914# a_16241_44734# 0.006538f
C18328 a_9482_43914# a_11173_44260# 0.043729f
C18329 a_n2293_42834# a_n2661_42282# 0.026231f
C18330 a_13249_42308# a_13749_43396# 3.84e-19
C18331 a_18114_32519# a_20512_43084# 5.22e-19
C18332 a_3537_45260# a_5829_43940# 3.27e-20
C18333 a_n4334_40480# a_n2810_45572# 5.22e-19
C18334 a_21335_42336# a_n357_42282# 2.03e-19
C18335 a_7174_31319# a_n755_45592# 2.56e-20
C18336 a_11691_44458# a_13059_46348# 0.015799f
C18337 a_4743_44484# a_3090_45724# 0.05313f
C18338 a_18911_45144# a_19123_46287# 7.75e-20
C18339 a_6109_44484# a_5257_43370# 0.001517f
C18340 a_16211_45572# a_13259_45724# 0.004313f
C18341 a_20623_45572# a_8049_45260# 0.01128f
C18342 a_n984_44318# a_n881_46662# 8.92e-19
C18343 a_10951_45334# a_11189_46129# 4.23e-21
C18344 a_11787_45002# a_9290_44172# 4.62e-19
C18345 a_9482_43914# a_8953_45546# 1.61e-19
C18346 a_175_44278# a_n1613_43370# 2.35e-19
C18347 a_413_45260# a_21137_46414# 4e-22
C18348 a_6171_45002# a_14275_46494# 1.21e-20
C18349 a_4927_45028# a_2324_44458# 3.2e-20
C18350 a_1241_43940# a_n746_45260# 4.29e-20
C18351 a_6761_42308# a_8325_42308# 5.55e-19
C18352 a_5934_30871# a_8515_42308# 0.222946f
C18353 a_22400_42852# a_13258_32519# 0.039664f
C18354 a_11530_34132# a_19120_35138# 0.480251f
C18355 EN_VIN_BSTR_N a_18194_35068# 0.340036f
C18356 a_6151_47436# a_4419_46090# 4.28e-20
C18357 a_12891_46348# a_14035_46660# 1.12e-20
C18358 a_4646_46812# a_5257_43370# 0.024804f
C18359 a_13661_43548# a_19692_46634# 0.093373f
C18360 a_13747_46662# a_19466_46812# 0.869986f
C18361 a_12549_44172# a_13885_46660# 0.036345f
C18362 a_n743_46660# a_11735_46660# 1.24e-19
C18363 a_3877_44458# a_7411_46660# 4.74e-19
C18364 a_19321_45002# a_15227_44166# 0.145462f
C18365 a_4817_46660# a_5894_47026# 1.46e-19
C18366 a_5807_45002# a_10185_46660# 6.99e-19
C18367 a_2266_47243# a_765_45546# 3.3e-19
C18368 a_11453_44696# a_20528_46660# 0.016145f
C18369 a_18479_47436# a_12741_44636# 0.020666f
C18370 a_13507_46334# a_21350_47026# 3.44e-19
C18371 a_4915_47217# a_5164_46348# 2.37e-20
C18372 a_n443_46116# a_5204_45822# 0.020803f
C18373 a_2063_45854# a_9823_46155# 3.28e-19
C18374 a_4791_45118# a_5497_46414# 0.056648f
C18375 a_n1151_42308# a_8199_44636# 0.161616f
C18376 a_19279_43940# a_15493_43940# 0.019758f
C18377 a_5343_44458# a_6765_43638# 9.35e-22
C18378 a_4223_44672# a_7112_43396# 3.59e-20
C18379 a_6298_44484# a_6293_42852# 2.36e-20
C18380 a_9313_44734# a_21381_43940# 0.028978f
C18381 a_11691_44458# a_15095_43370# 1.02e-20
C18382 a_20980_44850# a_19862_44208# 1.48e-19
C18383 a_22223_45036# a_10341_43396# 2.09e-19
C18384 a_5111_44636# a_9127_43156# 4.76e-19
C18385 a_3232_43370# a_8037_42858# 2.1e-22
C18386 a_n913_45002# a_17595_43084# 1.88e-20
C18387 a_n1059_45260# a_17701_42308# 0.073596f
C18388 a_n2017_45002# a_18083_42858# 0.03192f
C18389 en_comp a_5342_30871# 0.032532f
C18390 a_n23_44458# VDD 0.169093f
C18391 a_n4064_40160# VCM 0.121302f
C18392 a_n4209_39590# VIN_P 0.105382f
C18393 a_n4209_38502# a_n1532_35090# 9.11e-20
C18394 a_n3565_38502# a_n1838_35608# 1.42e-19
C18395 a_n3420_39072# C8_P_btm 8.3e-20
C18396 a_n3565_39304# C6_P_btm 0.080378f
C18397 a_n4064_39072# C10_P_btm 1.08e-19
C18398 a_n3565_37414# a_n2956_38216# 0.001835f
C18399 a_685_42968# a_584_46384# 0.00804f
C18400 a_20269_44172# a_19466_46812# 2.46e-20
C18401 a_9145_43396# a_12891_46348# 0.001541f
C18402 a_19862_44208# a_19692_46634# 0.027038f
C18403 a_13467_32519# a_12861_44030# 9.12e-21
C18404 a_17678_43396# a_16327_47482# 0.001965f
C18405 a_15743_43084# a_13507_46334# 0.158635f
C18406 a_16409_43396# a_11453_44696# 8.34e-21
C18407 a_n2661_43922# a_10809_44734# 0.073946f
C18408 a_14673_44172# a_14275_46494# 3.31e-21
C18409 a_8696_44636# CLK 0.006002f
C18410 a_1239_39043# a_1736_39043# 0.08488f
C18411 a_n3565_39304# a_n3690_38528# 6.38e-20
C18412 a_n3420_39072# a_n4334_38528# 0.008604f
C18413 a_1239_39587# a_1177_38525# 3.88e-21
C18414 a_n3690_39392# a_n3565_38502# 6.38e-20
C18415 a_n4064_39616# a_n4209_38216# 0.027937f
C18416 a_n3420_39616# a_n3565_38216# 0.028042f
C18417 a_n2302_39072# a_n2216_39072# 0.011479f
C18418 a_3524_46660# VDD 0.278519f
C18419 a_n881_46662# a_3503_45724# 0.001143f
C18420 a_11186_47026# a_11133_46155# 1.37e-19
C18421 a_3090_45724# a_8016_46348# 0.0122f
C18422 a_11813_46116# a_9290_44172# 4.46e-19
C18423 a_n1613_43370# a_n356_45724# 4.43e-20
C18424 a_5807_45002# a_20850_46155# 6.12e-21
C18425 a_3877_44458# a_4365_46436# 9.48e-20
C18426 a_20841_46902# a_20719_46660# 3.16e-19
C18427 a_19692_46634# a_4185_45028# 4.25e-20
C18428 a_20107_46660# a_20202_43084# 4.38e-20
C18429 a_10949_43914# a_10695_43548# 2.27e-19
C18430 a_9313_44734# a_18249_42858# 0.007699f
C18431 a_21381_43940# a_20974_43370# 0.02221f
C18432 a_1307_43914# a_10533_42308# 1.27e-21
C18433 a_20193_45348# a_22400_42852# 0.05078f
C18434 a_17730_32519# a_13678_32519# 0.054146f
C18435 a_10807_43548# a_9803_43646# 3.09e-19
C18436 a_20512_43084# a_13887_32519# 8.15e-19
C18437 a_n356_44636# a_945_42968# 2.2e-19
C18438 a_5883_43914# a_9114_42852# 8.7e-21
C18439 a_n913_45002# a_21887_42336# 0.060677f
C18440 en_comp a_20107_42308# 4.59e-20
C18441 a_9420_43940# VDD 0.0046f
C18442 a_6511_45714# a_1423_45028# 4.54e-21
C18443 a_10180_45724# a_10775_45002# 0.073185f
C18444 a_16147_45260# a_18787_45572# 4.04e-20
C18445 a_18479_45785# a_17668_45572# 1.16e-19
C18446 a_11823_42460# a_6171_45002# 0.123118f
C18447 a_10193_42453# a_8953_45002# 0.001294f
C18448 a_8746_45002# a_8191_45002# 7.28e-19
C18449 a_4699_43561# a_2324_44458# 1.33e-20
C18450 a_6293_42852# a_5937_45572# 1.17e-19
C18451 a_n1630_35242# SMPL_ON_N 0.076872f
C18452 a_4958_30871# w_11334_34010# 0.003841f
C18453 a_n4064_37440# VCM 0.020152f
C18454 a_22521_40599# RST_Z 2.23e-19
C18455 a_19900_46494# VDD 0.279179f
C18456 a_6598_45938# a_6151_47436# 0.173467f
C18457 a_6667_45809# a_6545_47178# 1.61e-19
C18458 a_6472_45840# a_6851_47204# 5.75e-21
C18459 a_6511_45714# a_6491_46660# 5.95e-22
C18460 a_n2293_46098# a_n356_45724# 0.022803f
C18461 a_376_46348# a_n357_42282# 2.8e-19
C18462 a_2698_46116# a_n2661_45546# 9.6e-20
C18463 a_n1076_46494# a_n755_45592# 6.77e-20
C18464 a_472_46348# a_310_45028# 3.57e-19
C18465 a_4185_45028# a_20692_30879# 1.35e-19
C18466 a_1138_42852# a_n863_45724# 0.135594f
C18467 a_12741_44636# a_n443_42852# 7.1e-20
C18468 a_2324_44458# a_10586_45546# 0.436403f
C18469 a_18819_46122# a_8049_45260# 0.003213f
C18470 a_13351_46090# a_12638_46436# 0.001216f
C18471 a_11387_46155# a_11601_46155# 0.005572f
C18472 a_9313_44734# a_21125_42558# 2.22e-19
C18473 a_15682_43940# a_16877_42852# 2.72e-20
C18474 a_2479_44172# a_2903_42308# 2.23e-20
C18475 a_14358_43442# a_743_42282# 1.97e-20
C18476 a_16409_43396# a_17324_43396# 0.118759f
C18477 a_16243_43396# a_18525_43370# 4.59e-21
C18478 a_n97_42460# a_13635_43156# 0.001861f
C18479 a_n4318_39768# a_n1630_35242# 1.81e-19
C18480 a_9145_43396# a_4361_42308# 1.15e-19
C18481 a_10341_43396# a_17678_43396# 2.66e-19
C18482 a_n2840_46634# CLK_DATA 9e-19
C18483 a_12089_42308# VDD 0.807892f
C18484 a_11823_42460# a_14673_44172# 7.39e-20
C18485 a_18175_45572# a_18248_44752# 8.43e-19
C18486 a_2711_45572# a_20512_43084# 7.39e-20
C18487 a_6171_45002# a_16321_45348# 3.7e-19
C18488 a_n3420_38528# a_n2312_38680# 0.009774f
C18489 a_15868_43402# a_n443_42852# 3.07e-19
C18490 a_4808_45572# a_3090_45724# 2.21e-19
C18491 a_3357_43084# a_13661_43548# 2.72e-20
C18492 a_2437_43646# a_19321_45002# 0.009654f
C18493 a_n2017_45002# a_12549_44172# 5.58e-20
C18494 a_19479_31679# a_13747_46662# 8.06e-20
C18495 a_n467_45028# a_n881_46662# 0.008624f
C18496 a_n143_45144# a_n1613_43370# 4.99e-21
C18497 a_413_45260# a_3094_47243# 5.44e-19
C18498 a_14180_45002# a_10227_46804# 0.002579f
C18499 a_n2661_43370# a_2063_45854# 0.039988f
C18500 a_18249_42858# a_18599_43230# 0.210876f
C18501 a_7765_42852# a_8292_43218# 0.157652f
C18502 a_18083_42858# a_19164_43230# 0.101963f
C18503 a_3626_43646# a_15803_42450# 0.006237f
C18504 a_2982_43646# a_15890_42674# 9.89e-20
C18505 a_4190_30871# a_14097_32519# 0.031855f
C18506 a_5111_42852# a_4649_42852# 1.58e-19
C18507 a_17333_42852# a_19339_43156# 4.42e-21
C18508 a_18907_42674# VDD 0.148872f
C18509 a_n1741_47186# a_n310_47570# 5.79e-19
C18510 a_n1605_47204# a_n2312_40392# 2.12e-19
C18511 SMPL_ON_P a_n2312_39304# 0.040801f
C18512 a_11031_47542# a_9313_45822# 0.063846f
C18513 a_6575_47204# a_n1435_47204# 5.93e-19
C18514 a_6151_47436# a_11599_46634# 0.008629f
C18515 a_n699_43396# a_n23_44458# 2.43e-20
C18516 a_n2661_44458# a_5891_43370# 0.013115f
C18517 a_10193_42453# a_3626_43646# 0.13905f
C18518 a_11691_44458# a_11649_44734# 4.78e-19
C18519 a_626_44172# a_n1899_43946# 2.19e-20
C18520 a_7229_43940# a_7542_44172# 0.086946f
C18521 a_n2017_45002# a_12429_44172# 3.24e-21
C18522 a_n913_45002# a_10807_43548# 0.023237f
C18523 a_n1059_45260# a_11750_44172# 1.48e-21
C18524 a_2382_45260# a_3499_42826# 0.040227f
C18525 a_3357_43084# a_19862_44208# 9.13e-21
C18526 a_5932_42308# a_n755_45592# 0.040158f
C18527 a_n4209_39590# a_n2956_38680# 0.020934f
C18528 a_13333_42558# a_13259_45724# 8.98e-20
C18529 a_9241_45822# VDD 0.003665f
C18530 a_3600_43914# a_584_46384# 3.17e-19
C18531 a_n143_45144# a_n2293_46098# 2.2e-21
C18532 a_n2293_45010# a_1138_42852# 9.98e-19
C18533 a_3357_43084# a_4185_45028# 0.027077f
C18534 a_n2012_44484# a_n2293_46634# 8.23e-19
C18535 a_6109_44484# a_5807_45002# 3.89e-20
C18536 a_18245_44484# a_16327_47482# 3.03e-19
C18537 a_20362_44736# a_18479_47436# 1.52e-20
C18538 a_2437_43646# a_5068_46348# 1.07e-20
C18539 a_n2293_43922# a_n1613_43370# 2.76e-19
C18540 a_16147_45260# a_15682_46116# 2.64e-19
C18541 a_17478_45572# a_10809_44734# 1.1e-21
C18542 a_n2661_43922# a_n881_46662# 4.12e-19
C18543 a_5263_45724# a_n2661_45546# 6.45e-19
C18544 a_8192_45572# a_5066_45546# 0.001238f
C18545 a_10193_42453# a_11601_46155# 0.002905f
C18546 a_21356_42826# a_21335_42336# 0.00235f
C18547 a_22223_42860# a_13258_32519# 1.75e-20
C18548 a_564_42282# a_1184_42692# 0.00104f
C18549 a_n3674_37592# a_961_42354# 1.74e-21
C18550 a_12800_43218# a_12563_42308# 5.38e-19
C18551 a_n1630_35242# a_1576_42282# 1.99e-20
C18552 COMP_P a_n327_42308# 3.18e-21
C18553 a_11136_42852# a_5742_30871# 6.68e-19
C18554 a_11599_46634# a_19466_46812# 0.453656f
C18555 a_10227_46804# a_15009_46634# 0.02057f
C18556 a_16327_47482# a_16292_46812# 0.027563f
C18557 a_17591_47464# a_3090_45724# 5.31e-19
C18558 a_n1151_42308# a_765_45546# 1.7705f
C18559 a_8128_46384# a_7411_46660# 0.019875f
C18560 a_n881_46662# a_7927_46660# 0.017621f
C18561 a_n1925_46634# a_479_46660# 8.56e-19
C18562 a_n2438_43548# a_491_47026# 8.49e-19
C18563 a_601_46902# a_948_46660# 0.051162f
C18564 a_n743_46660# a_n935_46688# 0.001334f
C18565 a_n2293_46634# a_n2661_46098# 0.022053f
C18566 a_n133_46660# a_288_46660# 0.086708f
C18567 a_n2661_46634# a_3177_46902# 0.00699f
C18568 a_5807_45002# a_4646_46812# 0.032485f
C18569 a_6298_44484# a_7499_43940# 3.16e-19
C18570 a_17970_44736# a_14021_43940# 2.51e-21
C18571 a_5883_43914# a_5745_43940# 0.007922f
C18572 a_4223_44672# a_9801_43940# 3.24e-20
C18573 a_9313_44734# a_14955_43940# 1.56e-20
C18574 a_n2293_42834# a_7112_43396# 6.84e-20
C18575 a_20512_43084# a_22485_44484# 0.004999f
C18576 a_14539_43914# a_15037_44260# 8.96e-19
C18577 a_7499_43078# a_10553_43218# 1.15e-19
C18578 a_n2661_42834# a_8018_44260# 2.37e-19
C18579 a_n1059_45260# a_4361_42308# 0.033614f
C18580 a_n913_45002# a_13467_32519# 0.024166f
C18581 a_20447_31679# a_17364_32525# 0.054026f
C18582 en_comp a_743_42282# 1.86e-20
C18583 a_3754_39466# VDD 0.009313f
C18584 a_21005_45260# VDD 0.184261f
C18585 a_7640_43914# a_3483_46348# 0.003497f
C18586 a_n2293_43922# a_n2293_46098# 7.21e-22
C18587 a_15146_44811# a_12741_44636# 1.05e-19
C18588 a_1414_42308# a_3090_45724# 8.03e-21
C18589 a_21845_43940# a_12549_44172# 0.003853f
C18590 a_7542_44172# a_8270_45546# 4.69e-19
C18591 a_18533_44260# a_13661_43548# 7.69e-20
C18592 a_1307_43914# a_3503_45724# 1.08e-21
C18593 a_1423_45028# a_n755_45592# 0.032517f
C18594 a_18911_45144# a_8049_45260# 1.78e-20
C18595 a_13556_45296# a_n443_42852# 2.5e-20
C18596 a_13720_44458# a_13759_46122# 1.69e-22
C18597 a_n97_42460# a_n1613_43370# 0.011527f
C18598 a_3080_42308# a_n2312_39304# 4.02e-21
C18599 a_n784_42308# C0_N_btm 0.281635f
C18600 a_3877_44458# a_4185_45028# 0.338483f
C18601 a_14084_46812# a_765_45546# 7.01e-21
C18602 a_15227_44166# a_13059_46348# 5.76e-19
C18603 a_16292_46812# a_16434_46987# 0.005572f
C18604 a_3090_45724# a_15312_46660# 9.66e-19
C18605 a_n881_46662# a_6419_46482# 3.32e-21
C18606 a_20916_46384# a_21137_46414# 0.118131f
C18607 a_n743_46660# a_2324_44458# 0.036195f
C18608 a_19594_46812# a_10809_44734# 0.042242f
C18609 a_16750_47204# a_6945_45028# 7.64e-20
C18610 a_n1613_43370# a_6640_46482# 7.81e-19
C18611 a_18479_47436# a_16375_45002# 2.07e-21
C18612 a_16327_47482# a_20254_46482# 0.001965f
C18613 a_18597_46090# a_18147_46436# 5.21e-20
C18614 a_n443_46116# a_3503_45724# 1.86e-19
C18615 a_2063_45854# a_2307_45899# 4.37e-19
C18616 a_19328_44172# a_19319_43548# 0.033025f
C18617 a_9313_44734# a_5649_42852# 0.028023f
C18618 a_20193_45348# a_22223_42860# 0.017179f
C18619 a_8975_43940# a_8037_42858# 2.54e-20
C18620 a_18451_43940# a_18533_43940# 0.171361f
C18621 a_11341_43940# a_10651_43940# 7.77e-20
C18622 a_5111_44636# a_1755_42282# 2.47e-19
C18623 a_3065_45002# a_2713_42308# 3.6e-19
C18624 a_2382_45260# a_3318_42354# 0.028613f
C18625 a_n2017_45002# a_7227_42308# 0.005025f
C18626 a_n1059_45260# a_6761_42308# 6.76e-21
C18627 a_n913_45002# a_6773_42558# 0.003807f
C18628 a_10907_45822# a_12561_45572# 4.22e-21
C18629 a_n4318_38216# a_n1151_42308# 9.61e-21
C18630 a_n97_42460# a_n2293_46098# 0.333817f
C18631 a_15095_43370# a_15227_44166# 0.022423f
C18632 a_10835_43094# a_n2293_46634# 8.49e-20
C18633 a_19164_43230# a_12549_44172# 1.3e-20
C18634 a_12281_43396# a_3090_45724# 0.027472f
C18635 a_12800_43218# a_10227_46804# 2.53e-19
C18636 a_3422_30871# a_n357_42282# 0.122733f
C18637 a_1736_39587# VDAC_Pi 0.009393f
C18638 a_17531_42308# CAL_N 7.31e-19
C18639 a_13351_46090# a_13759_46122# 0.043782f
C18640 a_11189_46129# a_2324_44458# 2.84e-19
C18641 a_10903_43370# a_14275_46494# 3.08e-20
C18642 a_17829_46910# a_16375_45002# 1.99e-19
C18643 a_18285_46348# a_18243_46436# 0.002179f
C18644 a_1138_42852# a_1431_46436# 6.23e-19
C18645 a_376_46348# a_518_46155# 0.005572f
C18646 a_18079_43940# a_18083_42858# 7.22e-20
C18647 a_2982_43646# a_16547_43609# 9.82e-21
C18648 a_14401_32519# a_22223_43396# 0.006786f
C18649 a_20974_43370# a_5649_42852# 0.186094f
C18650 a_5891_43370# a_8325_42308# 0.053347f
C18651 a_14539_43914# a_15890_42674# 3.49e-22
C18652 a_3626_43646# a_16137_43396# 0.003078f
C18653 a_17538_32519# a_13678_32519# 0.051187f
C18654 a_8791_43396# a_10341_43396# 1.01e-19
C18655 a_8685_43396# a_8229_43396# 1.2e-19
C18656 a_n97_42460# a_17678_43396# 2.62e-19
C18657 a_18479_47436# RST_Z 1.77e-19
C18658 a_10227_46804# SINGLE_ENDED 1.93e-19
C18659 a_15507_47210# CLK 6.68e-19
C18660 a_18143_47464# START 0.006044f
C18661 SMPL_ON_N a_11530_34132# 2.32e-19
C18662 a_6511_45714# a_6109_44484# 1.17e-19
C18663 a_8696_44636# a_11691_44458# 0.141053f
C18664 a_18175_45572# a_16922_45042# 5.86e-20
C18665 a_16147_45260# a_17023_45118# 0.040001f
C18666 a_11823_42460# a_12607_44458# 0.01822f
C18667 a_11962_45724# a_13076_44458# 1.5e-19
C18668 a_6431_45366# a_6709_45028# 0.112564f
C18669 a_6171_45002# a_7705_45326# 0.009164f
C18670 a_5205_44484# a_7229_43940# 0.006973f
C18671 a_3232_43370# a_8191_45002# 0.045343f
C18672 a_5342_30871# a_4185_45028# 0.067871f
C18673 a_20107_42308# a_13661_43548# 3.89e-19
C18674 a_6293_42852# a_n443_42852# 0.033407f
C18675 a_4361_42308# a_n1925_42282# 0.08654f
C18676 a_1847_42826# a_2324_44458# 3.13e-21
C18677 a_9127_43156# a_9290_44172# 0.003077f
C18678 a_10796_42968# a_8953_45546# 2.18e-20
C18679 a_n2946_39072# a_n2312_39304# 0.020842f
C18680 a_n467_45028# a_n443_46116# 1.81e-19
C18681 a_413_45260# a_4007_47204# 4.35e-19
C18682 a_3065_45002# a_2905_45572# 0.004116f
C18683 a_4574_45260# a_2063_45854# 6.45e-20
C18684 a_5205_44484# a_n237_47217# 1.8e-20
C18685 a_7229_43940# a_n971_45724# 7.24e-21
C18686 a_4558_45348# a_584_46384# 2.74e-19
C18687 a_13527_45546# a_n743_46660# 8.32e-20
C18688 a_6511_45714# a_4646_46812# 0.421269f
C18689 a_6667_45809# a_3877_44458# 7.89e-19
C18690 a_2711_45572# a_5732_46660# 2.43e-20
C18691 a_3357_43084# a_14955_47212# 2.77e-19
C18692 a_2437_43646# a_15811_47375# 0.006582f
C18693 a_20841_45814# a_18597_46090# 0.024341f
C18694 a_20719_45572# a_16327_47482# 0.001951f
C18695 a_21363_45546# a_18479_47436# 0.001869f
C18696 a_17478_45572# a_n881_46662# 0.11503f
C18697 a_n2661_45546# a_380_45546# 0.012814f
C18698 a_n2293_45546# a_n1079_45724# 5.25e-19
C18699 a_n2810_45572# a_n1099_45572# 0.001228f
C18700 a_n2956_38216# a_n863_45724# 0.001226f
C18701 a_13467_32519# a_20922_43172# 5.27e-19
C18702 a_20269_44172# a_13258_32519# 1.75e-21
C18703 a_20623_43914# a_19511_42282# 1.33e-21
C18704 a_4235_43370# a_1755_42282# 6.88e-21
C18705 a_21487_43396# a_21195_42852# 0.01192f
C18706 a_5111_42852# a_5755_42852# 1.15e-19
C18707 a_5649_42852# a_18599_43230# 9.69e-21
C18708 a_4361_42308# a_19987_42826# 1.33e-19
C18709 a_n1557_42282# a_1184_42692# 1.23e-19
C18710 a_15493_43940# a_19332_42282# 2.75e-21
C18711 a_19862_44208# a_20107_42308# 2.1e-21
C18712 a_15095_43370# a_14635_42282# 0.001265f
C18713 a_9145_43396# a_13622_42852# 5.7e-20
C18714 a_20820_30879# a_22609_38406# 5.26e-21
C18715 a_7754_39300# a_5700_37509# 2.64e-19
C18716 a_5267_42460# VDD 0.170631f
C18717 a_18184_42460# CAL_N 7.63e-19
C18718 a_n2497_47436# a_2063_45854# 4e-20
C18719 a_n815_47178# a_n785_47204# 0.123817f
C18720 a_n971_45724# a_n237_47217# 0.134971f
C18721 a_n1741_47186# a_1239_47204# 0.022889f
C18722 a_n2109_47186# a_2124_47436# 0.037038f
C18723 a_15037_45618# a_14955_43940# 3.52e-21
C18724 a_1307_43914# a_n2661_43922# 0.023892f
C18725 a_9482_43914# a_15463_44811# 0.005265f
C18726 a_14976_45348# a_14539_43914# 4.77e-20
C18727 a_2711_45572# a_21381_43940# 4.03e-21
C18728 a_413_45260# a_19279_43940# 1.83e-21
C18729 a_20447_31679# a_19237_31679# 0.051563f
C18730 a_20107_42308# a_4185_45028# 1.64e-19
C18731 a_15486_42560# a_2324_44458# 5.07e-20
C18732 a_18504_43218# a_n357_42282# 0.003243f
C18733 a_7227_42308# a_526_44458# 5.53e-20
C18734 a_20107_45572# a_20107_46660# 0.001171f
C18735 a_19113_45348# a_19321_45002# 0.147788f
C18736 a_16237_45028# a_13661_43548# 5.58e-19
C18737 a_20193_45348# a_13747_46662# 0.049365f
C18738 a_16922_45042# a_n743_46660# 2.99e-19
C18739 a_n2661_44458# a_11309_47204# 1.64e-20
C18740 a_413_45260# a_15368_46634# 4.42e-20
C18741 a_2437_43646# a_13059_46348# 7.82e-20
C18742 a_10053_45546# a_2324_44458# 0.008381f
C18743 a_11962_45724# a_12594_46348# 0.177228f
C18744 a_12427_45724# a_12005_46116# 0.01091f
C18745 a_11823_42460# a_10903_43370# 1.16382f
C18746 a_6905_45572# a_5937_45572# 9.25e-20
C18747 a_12883_44458# a_11453_44696# 1.4e-20
C18748 a_n2661_43922# a_n443_46116# 0.044169f
C18749 a_n2293_43922# a_4791_45118# 3.57e-19
C18750 a_n2293_42282# a_4921_42308# 2.29e-20
C18751 a_12089_42308# a_11551_42558# 0.109508f
C18752 a_14209_32519# a_22775_42308# 1.21e-19
C18753 a_13678_32519# a_22465_38105# 0.034429f
C18754 a_3080_42308# C0_N_btm 0.018211f
C18755 a_768_44030# a_13675_47204# 5.16e-20
C18756 a_12549_44172# a_13759_47204# 3.89e-19
C18757 a_9804_47204# a_5807_45002# 0.039093f
C18758 a_n2312_39304# a_n2438_43548# 0.052323f
C18759 a_6151_47436# a_7411_46660# 0.330209f
C18760 a_4915_47217# a_8145_46902# 5.23e-20
C18761 a_n1435_47204# a_5385_46902# 3.12e-20
C18762 a_6545_47178# a_5257_43370# 8.38e-19
C18763 a_n971_45724# a_8270_45546# 0.251101f
C18764 a_n1151_42308# a_10623_46897# 1.42e-19
C18765 a_n237_47217# a_8023_46660# 1.98e-19
C18766 a_2063_45854# a_6682_46987# 8.35e-21
C18767 a_11827_44484# a_11341_43940# 0.231114f
C18768 a_n2661_44458# a_10807_43548# 1.72e-19
C18769 a_20193_45348# a_20269_44172# 0.002705f
C18770 a_n356_44636# a_1414_42308# 0.179164f
C18771 a_9049_44484# a_9127_43156# 1.35e-22
C18772 a_2711_45572# a_18249_42858# 0.001642f
C18773 a_7499_43078# a_8952_43230# 0.054554f
C18774 a_18479_45785# a_18783_43370# 2.61e-19
C18775 a_3232_43370# a_3540_43646# 0.00217f
C18776 a_14537_43396# VDD 0.779752f
C18777 a_n1630_35242# a_18194_35068# 0.465356f
C18778 a_n784_42308# C10_P_btm 1.34e-19
C18779 a_22521_40599# a_20820_30879# 3.31e-20
C18780 a_n97_42460# a_4791_45118# 0.02536f
C18781 a_1756_43548# a_584_46384# 0.00975f
C18782 a_n2129_44697# a_n1076_46494# 2.07e-21
C18783 a_n1177_44458# a_n1991_46122# 9.68e-22
C18784 a_19319_43548# a_12861_44030# 0.024237f
C18785 a_13490_45394# a_2324_44458# 6.46e-19
C18786 en_comp a_20205_31679# 1.91e-19
C18787 a_n2017_45002# a_n2661_45546# 0.001101f
C18788 a_n2472_45002# a_n2293_45546# 3.35e-19
C18789 a_n2661_45010# a_n1079_45724# 5.36e-21
C18790 a_13348_45260# a_8049_45260# 7.18e-21
C18791 a_10775_45002# a_10586_45546# 1.57e-19
C18792 a_18079_43940# a_12549_44172# 0.008672f
C18793 a_3785_47178# VDD 0.387755f
C18794 a_8791_42308# a_7174_31319# 9.76e-21
C18795 a_15764_42576# a_16104_42674# 0.029366f
C18796 a_14113_42308# a_15521_42308# 0.002088f
C18797 a_1606_42308# a_n3420_39072# 0.001872f
C18798 a_n881_46662# a_5164_46348# 0.03104f
C18799 a_n1613_43370# a_5204_45822# 0.002482f
C18800 a_11453_44696# a_12005_46116# 4.21e-21
C18801 a_12465_44636# a_13925_46122# 0.018086f
C18802 a_n1435_47204# a_n1533_46116# 3.18e-20
C18803 a_4883_46098# a_14275_46494# 0.006919f
C18804 a_13507_46334# a_14840_46494# 0.005149f
C18805 a_10227_46804# a_19335_46494# 8.56e-21
C18806 a_18597_46090# a_17957_46116# 0.018356f
C18807 a_18479_47436# a_18985_46122# 2.08e-19
C18808 a_16327_47482# a_6945_45028# 0.111399f
C18809 a_15673_47210# a_10809_44734# 4.01e-20
C18810 a_18780_47178# a_18819_46122# 1.69e-19
C18811 a_n1741_47186# a_12839_46116# 0.113988f
C18812 a_4791_45118# a_6640_46482# 0.001342f
C18813 a_2063_45854# a_9823_46482# 1.18e-21
C18814 a_10249_46116# a_12816_46660# 4.52e-20
C18815 a_3177_46902# a_765_45546# 0.001508f
C18816 a_6755_46942# a_12991_46634# 0.077634f
C18817 a_n2293_46634# a_11415_45002# 0.001066f
C18818 a_n2661_46634# a_12741_44636# 2.1e-19
C18819 a_768_44030# a_167_45260# 0.014856f
C18820 a_5891_43370# a_9145_43396# 0.049186f
C18821 a_n2661_43922# a_9396_43370# 9.06e-21
C18822 a_9313_44734# a_8685_43396# 0.124273f
C18823 a_14539_43914# a_16547_43609# 0.01221f
C18824 a_16979_44734# a_16243_43396# 3.15e-20
C18825 a_n356_44636# a_12281_43396# 2.72e-19
C18826 a_19721_31679# a_13678_32519# 0.051384f
C18827 a_10193_42453# a_13921_42308# 0.002387f
C18828 a_20512_43084# a_14401_32519# 5.21e-19
C18829 a_13249_42308# a_14113_42308# 2.26e-19
C18830 a_11823_42460# a_15959_42545# 9.34e-20
C18831 a_1307_43914# a_3445_43172# 1.01e-21
C18832 a_2998_44172# a_5326_44056# 9.84e-20
C18833 a_n1059_45260# a_13622_42852# 1.72e-19
C18834 a_20835_44721# VDD 0.198384f
C18835 a_10490_45724# a_12427_45724# 0.108721f
C18836 a_11322_45546# a_11962_45724# 0.270736f
C18837 a_11525_45546# a_11652_45724# 0.138143f
C18838 a_8746_45002# a_11823_42460# 2.13e-21
C18839 a_7499_43078# a_13249_42308# 1.99e-20
C18840 a_2711_45572# a_12016_45572# 2.58e-19
C18841 C0_dummy_P_btm EN_VIN_BSTR_P 0.026355f
C18842 a_10729_43914# a_3483_46348# 1.6e-21
C18843 a_743_42282# a_13661_43548# 0.132115f
C18844 a_7640_43914# a_n357_42282# 8.82e-19
C18845 a_5244_44056# a_2324_44458# 1.7e-20
C18846 a_n901_43156# a_n1613_43370# 0.281398f
C18847 a_10341_42308# a_10227_46804# 0.004877f
C18848 a_413_45260# DATA[1] 0.004906f
C18849 a_3090_45724# VDD 2.05725f
C18850 a_1176_45822# a_167_45260# 0.091673f
C18851 a_n2661_46098# a_2277_45546# 5.6e-20
C18852 a_12991_46634# a_8049_45260# 1.12e-20
C18853 a_4646_46812# a_n755_45592# 8.29e-20
C18854 a_1799_45572# a_1990_45899# 8.94e-19
C18855 a_n2293_46098# a_5204_45822# 0.008417f
C18856 a_19123_46287# a_17957_46116# 2.21e-20
C18857 a_18285_46348# a_18819_46122# 1.08e-19
C18858 a_16388_46812# a_10809_44734# 0.013923f
C18859 a_19862_44208# a_743_42282# 4.04e-19
C18860 a_20269_44172# a_20301_43646# 4.32e-19
C18861 a_20365_43914# a_4190_30871# 1.62e-20
C18862 a_4699_43561# a_3539_42460# 0.109444f
C18863 a_14021_43940# a_18783_43370# 0.006778f
C18864 a_3080_42308# a_3626_43646# 0.092602f
C18865 a_n97_42460# a_8791_43396# 6.57e-22
C18866 a_n2661_42282# a_n13_43084# 5.65e-21
C18867 a_3422_30871# a_21356_42826# 0.024863f
C18868 a_1049_43396# a_648_43396# 5.57e-19
C18869 a_1209_43370# a_1512_43396# 0.001377f
C18870 a_1568_43370# a_548_43396# 1.89e-20
C18871 a_6547_43396# VDD 0.219105f
C18872 a_16020_45572# a_16019_45002# 6.19e-19
C18873 a_15861_45028# a_16751_45260# 0.044248f
C18874 a_10193_42453# a_16405_45348# 0.001843f
C18875 a_n2661_45010# a_n2472_45002# 0.065751f
C18876 a_n2840_45002# a_n2293_45010# 2.81e-19
C18877 a_19479_31679# en_comp 1.32e-19
C18878 a_743_42282# a_4185_45028# 0.031243f
C18879 a_21671_42860# a_19692_46634# 1.06e-19
C18880 a_14543_43071# a_13059_46348# 4.18e-19
C18881 a_15002_46116# VDD 4.6e-19
C18882 a_10490_45724# a_11453_44696# 6.39e-21
C18883 a_11962_45724# a_12465_44636# 1.34e-21
C18884 a_11823_42460# a_4883_46098# 1.64e-19
C18885 a_13163_45724# a_13507_46334# 4.48e-19
C18886 a_526_44458# a_n2661_45546# 0.071855f
C18887 a_n1925_42282# a_n2810_45572# 3.89e-20
C18888 a_14579_43548# a_5342_30871# 0.041574f
C18889 a_5649_42852# a_13887_32519# 0.004879f
C18890 a_12281_43396# a_12379_42858# 0.036584f
C18891 a_14205_43396# a_5534_30871# 1.04e-19
C18892 a_13467_32519# a_17364_32525# 0.050014f
C18893 a_4361_42308# a_22959_43396# 1.39e-19
C18894 a_15095_43370# a_14543_43071# 1.43e-19
C18895 a_21855_43396# a_14209_32519# 2.74e-19
C18896 a_n3690_38304# a_n3420_37984# 0.414894f
C18897 a_8953_45002# a_10057_43914# 0.001204f
C18898 a_6171_45002# a_14539_43914# 3.43e-19
C18899 a_n1059_45260# a_5891_43370# 0.186322f
C18900 a_327_44734# a_n23_44458# 0.141544f
C18901 a_3357_43084# a_5708_44484# 0.005179f
C18902 a_5934_30871# a_1823_45246# 3.73e-20
C18903 a_5755_42308# a_4185_45028# 1.64e-19
C18904 a_18057_42282# a_17339_46660# 1.93e-19
C18905 a_10991_42826# a_n443_42852# 1.25e-19
C18906 a_16414_43172# a_n357_42282# 0.005649f
C18907 a_3080_42308# C10_P_btm 1.34e-19
C18908 a_n452_44636# a_n443_46116# 1.47e-20
C18909 a_5343_44458# a_n1151_42308# 1.19e-19
C18910 a_1176_45572# a_167_45260# 0.00195f
C18911 a_3733_45822# a_n2293_46098# 5.15e-19
C18912 a_19778_44110# a_18479_47436# 0.038618f
C18913 a_11827_44484# a_16327_47482# 0.107078f
C18914 a_18587_45118# a_18597_46090# 6.25e-19
C18915 a_6945_45348# a_n1613_43370# 1.51e-19
C18916 a_413_45260# a_2864_46660# 9.11e-21
C18917 a_6171_45002# a_2107_46812# 0.023061f
C18918 a_2680_45002# a_2609_46660# 1.09e-20
C18919 a_3065_45002# a_2443_46660# 2.64e-21
C18920 a_2437_43646# a_7577_46660# 1.39e-20
C18921 a_3357_43084# a_5257_43370# 0.894879f
C18922 a_10775_45002# a_n743_46660# 1.84e-21
C18923 a_8696_44636# a_15227_44166# 0.203885f
C18924 a_17478_45572# a_17609_46634# 8.56e-20
C18925 CLK_DATA VDD 0.422202f
C18926 a_1847_42826# a_1606_42308# 0.025123f
C18927 a_8037_42858# a_n784_42308# 6.19e-21
C18928 a_15743_43084# a_15486_42560# 6.65e-19
C18929 a_5649_42852# a_8515_42308# 5.44e-20
C18930 a_743_42282# a_9803_42558# 0.010183f
C18931 a_18083_42858# a_17749_42852# 3.87e-19
C18932 a_17333_42852# a_17665_42852# 0.001922f
C18933 a_3422_30871# a_n4064_37440# 0.032121f
C18934 a_2684_37794# VDD 0.286898f
C18935 a_n1435_47204# a_12891_46348# 0.001028f
C18936 a_6545_47178# a_5807_45002# 0.030195f
C18937 a_13381_47204# a_12549_44172# 0.135267f
C18938 a_15673_47210# a_n881_46662# 7.77e-20
C18939 a_12465_44636# SMPL_ON_N 0.006167f
C18940 a_22223_47212# a_22731_47423# 0.011229f
C18941 a_n971_45724# a_1123_46634# 1.3e-19
C18942 a_n785_47204# a_171_46873# 1.04e-19
C18943 a_n23_47502# a_33_46660# 0.001405f
C18944 a_327_47204# a_n133_46660# 0.006131f
C18945 a_1209_47178# a_n2438_43548# 4.34e-19
C18946 a_1239_47204# a_n743_46660# 8.16e-20
C18947 a_3160_47472# a_n2661_46634# 0.026361f
C18948 a_n746_45260# a_383_46660# 0.011439f
C18949 a_21811_47423# a_11453_44696# 0.005338f
C18950 a_4883_46098# a_22959_47212# 8.05e-21
C18951 a_14539_43914# a_14673_44172# 0.205935f
C18952 a_10193_42453# a_18525_43370# 2.7e-19
C18953 a_2711_45572# a_5649_42852# 1.3e-19
C18954 a_5826_44734# a_5708_44484# 1.98e-20
C18955 a_16112_44458# a_16241_44734# 0.062574f
C18956 a_9482_43914# a_10555_44260# 0.088693f
C18957 a_6109_44484# a_5608_44484# 4.33e-19
C18958 a_18479_45785# a_3626_43646# 4.26e-20
C18959 a_n998_44484# a_n2661_43922# 3.71e-19
C18960 a_n1059_45260# a_18533_43940# 5.26e-21
C18961 a_3537_45260# a_5745_43940# 1.23e-19
C18962 a_n4315_30879# a_n2810_45572# 0.024132f
C18963 a_7174_31319# a_n357_42282# 4.25e-19
C18964 a_20731_45938# VDD 0.142103f
C18965 a_1423_45028# a_3483_46348# 0.110369f
C18966 a_n699_43396# a_3090_45724# 0.058797f
C18967 a_19279_43940# a_20916_46384# 1.62e-21
C18968 a_11967_42832# a_n2293_46634# 6.03e-20
C18969 a_5826_44734# a_5257_43370# 0.003375f
C18970 a_18494_42460# a_17339_46660# 8.02e-20
C18971 a_20841_45814# a_8049_45260# 0.008238f
C18972 en_comp a_n2956_38680# 3.44e-19
C18973 a_n809_44244# a_n881_46662# 3.25e-20
C18974 a_10951_45334# a_9290_44172# 0.136064f
C18975 a_n984_44318# a_n1613_43370# 0.245331f
C18976 a_6171_45002# a_14493_46090# 6.27e-21
C18977 a_413_45260# a_20708_46348# 2.68e-21
C18978 a_5111_44636# a_2324_44458# 0.090721f
C18979 a_10949_43914# a_12861_44030# 8.34e-19
C18980 a_5379_42460# a_5742_30871# 7.37e-20
C18981 a_7963_42308# a_8515_42308# 8.26e-20
C18982 a_11530_34132# a_18194_35068# 0.4004f
C18983 CAL_P RST_Z 0.551895f
C18984 a_3877_44458# a_5257_43370# 0.142219f
C18985 a_13661_43548# a_19466_46812# 0.011727f
C18986 a_5807_45002# a_19692_46634# 6.61e-19
C18987 a_13747_46662# a_19333_46634# 0.011849f
C18988 a_5732_46660# a_6540_46812# 2.56e-19
C18989 a_5167_46660# a_5275_47026# 0.057222f
C18990 a_12549_44172# a_13170_46660# 2.28e-19
C18991 a_11453_44696# a_22000_46634# 0.008499f
C18992 a_18597_46090# a_11415_45002# 0.061694f
C18993 a_13507_46334# a_19636_46660# 4.68e-19
C18994 a_4915_47217# a_5068_46348# 6.9e-20
C18995 a_4791_45118# a_5204_45822# 0.053732f
C18996 a_n1151_42308# a_8349_46414# 0.095055f
C18997 a_2063_45854# a_9569_46155# 5.78e-20
C18998 a_n443_46116# a_5164_46348# 1.86e-20
C18999 a_6298_44484# a_6031_43396# 0.001377f
C19000 a_7542_44172# a_7845_44172# 0.137004f
C19001 a_5343_44458# a_6197_43396# 1.12e-20
C19002 a_4223_44672# a_7287_43370# 2.11e-19
C19003 a_2127_44172# a_2537_44260# 0.007617f
C19004 a_10057_43914# a_3626_43646# 2.08e-20
C19005 a_11827_44484# a_10341_43396# 3.05e-19
C19006 a_5111_44636# a_8387_43230# 0.001241f
C19007 a_n913_45002# a_16795_42852# 7.33e-21
C19008 a_n1059_45260# a_17595_43084# 0.049f
C19009 a_n2017_45002# a_17701_42308# 0.132871f
C19010 a_n356_44636# VDD 1.17667f
C19011 a_n4064_40160# VREF_GND 0.493568f
C19012 a_n4209_38502# a_n1386_35608# 1.52e-19
C19013 a_n4209_39304# C5_P_btm 1.83e-19
C19014 a_n3420_39072# C9_P_btm 5.77e-20
C19015 a_n3565_39304# C7_P_btm 0.001136f
C19016 a_15940_43402# a_10227_46804# 1.75e-19
C19017 a_17433_43396# a_16327_47482# 2.95e-19
C19018 a_18783_43370# a_13507_46334# 6.51e-20
C19019 a_16547_43609# a_11453_44696# 2.27e-20
C19020 a_14673_44172# a_14493_46090# 4.72e-21
C19021 a_n2661_42834# a_10809_44734# 0.14417f
C19022 a_n2661_44458# a_n2840_45546# 2.89e-19
C19023 a_n2840_44458# a_n2661_45546# 3.06e-19
C19024 a_n4318_40392# a_n2810_45572# 0.02461f
C19025 a_19862_44208# a_19466_46812# 4.57e-20
C19026 a_n3565_39304# a_n3565_38502# 0.041674f
C19027 a_n3420_39072# a_n4209_38502# 0.032647f
C19028 a_n4209_39304# a_n3420_38528# 0.029412f
C19029 a_n3420_39616# a_n4334_38304# 4.87e-19
C19030 a_n4064_39072# a_n2216_39072# 0.005565f
C19031 a_3699_46634# VDD 0.347281f
C19032 a_n3674_37592# a_n4064_37984# 0.020548f
C19033 a_19594_46812# a_19443_46116# 1.96e-19
C19034 a_n2293_46634# a_13259_45724# 0.032341f
C19035 a_768_44030# a_n863_45724# 0.020071f
C19036 a_n743_46660# a_12839_46116# 0.011568f
C19037 a_4955_46873# a_3873_46454# 1.98e-20
C19038 a_n881_46662# a_3316_45546# 6.79e-20
C19039 a_11186_47026# a_11189_46129# 3.64e-19
C19040 a_8667_46634# a_6945_45028# 5.95e-20
C19041 a_20273_46660# a_20719_46660# 2.28e-19
C19042 a_20841_46902# a_21350_47026# 2.6e-19
C19043 a_20107_46660# a_22365_46825# 4.87e-21
C19044 a_19123_46287# a_11415_45002# 5.55e-20
C19045 a_10729_43914# a_10695_43548# 0.00999f
C19046 a_10807_43548# a_9145_43396# 0.290878f
C19047 a_9313_44734# a_17333_42852# 0.010555f
C19048 a_n2293_42834# a_5379_42460# 1.97e-21
C19049 a_14021_43940# a_3626_43646# 1.24e-20
C19050 a_19237_31679# a_13467_32519# 0.052472f
C19051 a_n1761_44111# a_743_42282# 1.3e-19
C19052 a_n356_44636# a_873_42968# 2.03e-19
C19053 a_n2293_43922# a_12895_43230# 0.001356f
C19054 a_20193_45348# a_20836_43172# 9.63e-20
C19055 a_3422_30871# a_20749_43396# 1.42e-19
C19056 a_21381_43940# a_14401_32519# 4.91e-20
C19057 a_20512_43084# a_22223_43396# 0.001484f
C19058 a_n913_45002# a_21335_42336# 0.062808f
C19059 en_comp a_13258_32519# 0.007613f
C19060 a_9165_43940# VDD 0.192035f
C19061 a_6472_45840# a_1423_45028# 3.3e-21
C19062 a_18175_45572# a_17668_45572# 1.93e-20
C19063 a_7499_43078# a_11787_45002# 4.1e-20
C19064 a_18691_45572# a_18799_45938# 0.057222f
C19065 a_18479_45785# a_17568_45572# 5.46e-20
C19066 a_12427_45724# a_6171_45002# 8.61e-21
C19067 a_10180_45724# a_8953_45002# 0.107499f
C19068 a_11823_42460# a_3232_43370# 0.002063f
C19069 a_n4064_37440# VREF_GND 0.048151f
C19070 a_16328_43172# a_13661_43548# 1.62e-19
C19071 a_10729_43914# a_n357_42282# 4.51e-22
C19072 a_6031_43396# a_5937_45572# 0.010894f
C19073 a_2982_43646# a_10903_43370# 3.15e-19
C19074 a_n784_42308# a_n2312_40392# 7.39e-19
C19075 a_4958_30871# w_1575_34946# 0.00296f
C19076 CAL_N RST_Z 0.058301f
C19077 a_20075_46420# VDD 0.347847f
C19078 a_8162_45546# a_2063_45854# 2.61e-19
C19079 a_6667_45809# a_6151_47436# 0.1609f
C19080 a_6472_45840# a_6491_46660# 7.23e-22
C19081 a_6511_45714# a_6545_47178# 4.48e-20
C19082 a_n2293_46098# a_3503_45724# 0.01404f
C19083 a_1823_45246# a_n2293_45546# 0.234971f
C19084 a_472_46348# a_n1099_45572# 0.005608f
C19085 a_805_46414# a_380_45546# 5.77e-19
C19086 a_376_46348# a_310_45028# 5.66e-19
C19087 a_n901_46420# a_n755_45592# 0.002034f
C19088 a_1176_45822# a_n863_45724# 2.47e-19
C19089 a_4185_45028# a_20205_31679# 8.52e-20
C19090 a_17957_46116# a_8049_45260# 4.87e-20
C19091 a_12594_46348# a_12638_46436# 0.049443f
C19092 a_11189_46129# a_12839_46116# 8.15e-20
C19093 a_13351_46090# a_12379_46436# 2.98e-20
C19094 a_11387_46155# a_11315_46155# 6.64e-19
C19095 a_15682_43940# a_16245_42852# 6.93e-20
C19096 a_14579_43548# a_743_42282# 3.98e-19
C19097 a_16409_43396# a_17499_43370# 0.042737f
C19098 a_16977_43638# a_16759_43396# 0.209641f
C19099 a_16243_43396# a_18429_43548# 6.92e-21
C19100 a_16137_43396# a_18525_43370# 2.8e-19
C19101 a_2982_43646# a_3681_42891# 0.006879f
C19102 a_3905_42865# a_1755_42282# 5.4e-20
C19103 a_n97_42460# a_12895_43230# 1.91e-20
C19104 a_n3674_39768# a_n3674_37592# 0.024722f
C19105 a_16547_43609# a_17324_43396# 5.47e-21
C19106 a_3539_42460# a_1847_42826# 1.09e-20
C19107 a_10341_43396# a_17433_43396# 1.6e-19
C19108 a_13747_46662# CLK 3.82e-20
C19109 a_12379_42858# VDD 0.484153f
C19110 a_18175_45572# a_17970_44736# 2.35e-20
C19111 a_11787_45002# a_11915_45394# 0.004764f
C19112 a_11963_45334# a_n2661_43370# 2.8e-19
C19113 a_1307_43914# a_5837_45028# 1.79e-20
C19114 en_comp a_20193_45348# 6.75e-20
C19115 a_6171_45002# a_14309_45028# 0.00276f
C19116 a_21542_45572# a_19721_31679# 3.76e-20
C19117 a_9306_43218# a_9290_44172# 1.97e-21
C19118 a_15231_43396# a_n443_42852# 4.71e-19
C19119 a_n3690_38528# a_n2312_38680# 5.77e-19
C19120 a_11551_42558# a_3090_45724# 6.89e-20
C19121 a_10210_45822# a_9863_46634# 2.83e-20
C19122 a_3357_43084# a_5807_45002# 0.071743f
C19123 a_n2293_45010# a_768_44030# 0.03517f
C19124 a_21513_45002# a_19321_45002# 0.002479f
C19125 a_2437_43646# a_19452_47524# 0.001463f
C19126 a_n467_45028# a_n1613_43370# 0.004184f
C19127 a_6171_45002# a_11453_44696# 1.39146f
C19128 a_7705_45326# a_4883_46098# 4.33e-20
C19129 a_13777_45326# a_10227_46804# 9.51e-19
C19130 a_n2661_43370# a_584_46384# 0.034714f
C19131 a_11361_45348# a_2063_45854# 6.44e-22
C19132 a_18249_42858# a_18817_42826# 0.16939f
C19133 a_18083_42858# a_19339_43156# 0.042271f
C19134 a_7871_42858# a_8292_43218# 0.086377f
C19135 a_8685_43396# a_8515_42308# 5.84e-21
C19136 a_3626_43646# a_15764_42576# 0.002707f
C19137 a_2982_43646# a_15959_42545# 2.23e-19
C19138 a_4520_42826# a_4649_42852# 0.062574f
C19139 a_7765_42852# a_7573_43172# 1.97e-19
C19140 a_17333_42852# a_18599_43230# 3.68e-19
C19141 a_21381_43940# a_21421_42336# 1.07e-19
C19142 a_18727_42674# VDD 0.181095f
C19143 a_n1151_42308# a_10227_46804# 0.458569f
C19144 a_n2109_47186# a_n89_47570# 2.32e-19
C19145 SMPL_ON_P a_n2312_40392# 4.89949f
C19146 a_n1741_47186# a_n2312_39304# 0.005742f
C19147 a_9863_47436# a_9313_45822# 0.049145f
C19148 a_7903_47542# a_n1435_47204# 2.39e-19
C19149 a_6151_47436# a_14955_47212# 0.192081f
C19150 a_n699_43396# a_n356_44636# 0.044884f
C19151 a_n2661_44458# a_8375_44464# 0.003111f
C19152 a_626_44172# a_n1761_44111# 3.66e-23
C19153 a_11827_44484# a_n2293_43922# 0.028646f
C19154 a_1307_43914# a_n809_44244# 5.87e-21
C19155 a_7229_43940# a_7281_43914# 0.164835f
C19156 a_n1059_45260# a_10807_43548# 0.031771f
C19157 a_n2017_45002# a_11750_44172# 1.48e-22
C19158 a_n913_45002# a_10949_43914# 0.001202f
C19159 a_5932_42308# a_n357_42282# 6.58e-19
C19160 a_6123_31319# a_n863_45724# 8.96e-21
C19161 a_6171_42473# a_n755_45592# 1.56e-19
C19162 a_n4209_39590# a_n2956_39304# 0.022939f
C19163 a_13249_42558# a_13259_45724# 8.98e-20
C19164 a_8697_45822# VDD 0.189893f
C19165 a_17364_32525# VCM 0.035838f
C19166 a_2998_44172# a_584_46384# 0.181241f
C19167 a_7845_44172# a_n971_45724# 1.69e-20
C19168 a_261_44278# a_n2497_47436# 0.002478f
C19169 a_20159_44458# a_18479_47436# 3.97e-21
C19170 a_18005_44484# a_16327_47482# 0.001967f
C19171 a_11967_42832# a_18597_46090# 0.021692f
C19172 a_3422_30871# a_12861_44030# 0.018986f
C19173 a_14673_44172# a_11453_44696# 0.001076f
C19174 a_n2661_43922# a_n1613_43370# 0.113996f
C19175 a_16147_45260# a_2324_44458# 1.7e-19
C19176 a_15861_45028# a_10809_44734# 8.82e-22
C19177 a_n2661_42834# a_n881_46662# 6.26e-20
C19178 a_8336_45822# a_8034_45724# 8.44e-21
C19179 a_10193_42453# a_11315_46155# 7.86e-19
C19180 a_4099_45572# a_n2661_45546# 0.008087f
C19181 a_n967_45348# a_n1991_46122# 1.72e-20
C19182 a_n2661_45010# a_1823_45246# 1.68e-19
C19183 a_9313_44734# a_768_44030# 0.044729f
C19184 a_n467_45028# a_n2293_46098# 2.4e-21
C19185 a_19479_31679# a_4185_45028# 0.03554f
C19186 a_n745_45366# a_n1076_46494# 5.48e-20
C19187 a_22165_42308# a_13258_32519# 0.004531f
C19188 a_n3674_37592# a_1184_42692# 1.16e-19
C19189 a_11136_42852# a_11323_42473# 8.95e-19
C19190 a_n1630_35242# a_1067_42314# 4.97e-19
C19191 a_11599_46634# a_19333_46634# 0.001374f
C19192 a_16241_47178# a_16292_46812# 3.13e-19
C19193 a_10227_46804# a_14084_46812# 1.42e-19
C19194 a_16327_47482# a_15559_46634# 0.001169f
C19195 a_4915_47217# a_13059_46348# 0.021189f
C19196 a_3160_47472# a_765_45546# 0.027219f
C19197 a_n881_46662# a_8145_46902# 0.003327f
C19198 a_n2438_43548# a_288_46660# 0.013776f
C19199 a_n1021_46688# a_n935_46688# 0.006584f
C19200 a_33_46660# a_948_46660# 0.117156f
C19201 a_n133_46660# a_1983_46706# 6.11e-21
C19202 a_n2293_46634# a_1799_45572# 0.001265f
C19203 a_n2661_46634# a_2609_46660# 0.045654f
C19204 a_5807_45002# a_3877_44458# 0.034811f
C19205 a_n2442_46660# a_n2661_46098# 6.94e-20
C19206 a_n743_46660# a_491_47026# 6.49e-20
C19207 a_6298_44484# a_6671_43940# 4.34e-19
C19208 a_9313_44734# a_13483_43940# 1.18e-20
C19209 a_n2293_42834# a_7287_43370# 7.97e-19
C19210 a_1307_43914# a_14955_43396# 5.43e-20
C19211 a_14539_43914# a_14761_44260# 3.61e-19
C19212 a_22315_44484# a_19237_31679# 4.46e-20
C19213 a_11827_44484# a_n97_42460# 4.56e-20
C19214 a_n2661_42834# a_7911_44260# 4.06e-19
C19215 a_n2017_45002# a_4361_42308# 0.004087f
C19216 a_7754_39632# VDD 0.205733f
C19217 a_20567_45036# VDD 0.237324f
C19218 a_15433_44458# a_12741_44636# 0.004093f
C19219 a_6109_44484# a_3483_46348# 0.003232f
C19220 a_n2661_43922# a_n2293_46098# 0.026124f
C19221 a_15037_43940# a_13661_43548# 2.04e-19
C19222 a_7281_43914# a_8270_45546# 1.81e-20
C19223 a_17538_32519# a_12549_44172# 1.42e-19
C19224 a_1307_43914# a_3316_45546# 1.38e-19
C19225 a_9482_43914# a_n443_42852# 1.75e-19
C19226 a_18587_45118# a_8049_45260# 2.06e-21
C19227 a_1423_45028# a_n357_42282# 2.14e-20
C19228 a_1145_45348# a_n755_45592# 7.7e-19
C19229 a_626_44172# a_997_45618# 1.07e-19
C19230 a_14539_43914# a_10903_43370# 3.63e-21
C19231 a_n447_43370# a_n1613_43370# 7.94e-19
C19232 a_3080_42308# a_n2312_40392# 5.51e-21
C19233 a_3626_43646# a_13507_46334# 0.04477f
C19234 a_22775_42308# a_22465_38105# 0.330766f
C19235 a_21613_42308# a_21973_42336# 0.001645f
C19236 a_2583_47243# VDD 2.18e-20
C19237 a_n784_42308# C0_dummy_N_btm 2.62e-20
C19238 a_3877_44458# a_3699_46348# 0.084544f
C19239 a_4646_46812# a_3483_46348# 0.048267f
C19240 a_6755_46942# a_11415_45002# 0.02226f
C19241 a_17609_46634# a_16388_46812# 2.5e-19
C19242 a_13607_46688# a_765_45546# 2.05e-20
C19243 a_15009_46634# a_15312_46660# 0.001377f
C19244 a_n881_46662# a_5066_45546# 0.801045f
C19245 a_20916_46384# a_20708_46348# 0.189941f
C19246 a_n743_46660# a_14840_46494# 0.010488f
C19247 a_19321_45002# a_10809_44734# 0.035502f
C19248 a_20843_47204# a_6945_45028# 0.003967f
C19249 a_2107_46812# a_10903_43370# 9.6e-21
C19250 a_4883_46098# a_14371_46494# 2.3e-19
C19251 a_18597_46090# a_13259_45724# 1.02e-19
C19252 a_11599_46634# a_20062_46116# 6.27e-19
C19253 a_16327_47482# a_20009_46494# 2.95e-19
C19254 a_n1151_42308# a_n906_45572# 0.002303f
C19255 a_n443_46116# a_3316_45546# 3.74e-19
C19256 a_n2661_42282# a_104_43370# 5.48e-21
C19257 a_20193_45348# a_22165_42308# 0.252856f
C19258 a_9313_44734# a_13678_32519# 0.097255f
C19259 a_18326_43940# a_18533_43940# 0.001502f
C19260 a_19328_44172# a_19808_44306# 0.001696f
C19261 a_18451_43940# a_19319_43548# 1.99e-20
C19262 a_5111_44636# a_1606_42308# 1.35e-20
C19263 a_n2017_45002# a_6761_42308# 0.006728f
C19264 a_n913_45002# a_6481_42558# 0.005099f
C19265 a_2382_45260# a_2903_42308# 1.98e-20
C19266 a_6511_45714# a_3357_43084# 1.21e-20
C19267 a_n4064_37984# EN_VIN_BSTR_P 0.031746f
C19268 a_10752_42852# a_10227_46804# 1.7e-19
C19269 a_6671_43940# a_5937_45572# 0.06027f
C19270 a_14205_43396# a_15227_44166# 1.11e-19
C19271 a_19339_43156# a_12549_44172# 1.24e-20
C19272 a_10518_42984# a_n2293_46634# 4.29e-20
C19273 a_743_42282# a_5257_43370# 1.37e-19
C19274 a_5342_30871# a_5807_45002# 1.35e-22
C19275 a_21076_30879# VDD 1.17389f
C19276 a_12594_46348# a_13759_46122# 9.6e-19
C19277 a_9290_44172# a_2324_44458# 0.026216f
C19278 a_10903_43370# a_14493_46090# 1.62e-20
C19279 a_7174_31319# a_n4064_37440# 1.84e-19
C19280 a_17303_42282# CAL_N 0.003472f
C19281 a_19123_46287# a_13259_45724# 6.59e-21
C19282 a_765_45546# a_16375_45002# 0.008153f
C19283 a_18285_46348# a_18147_46436# 0.001014f
C19284 a_1138_42852# a_1337_46436# 1.4e-19
C19285 a_11415_45002# a_8049_45260# 0.426371f
C19286 a_17973_43940# a_18083_42858# 5.46e-19
C19287 a_2982_43646# a_16243_43396# 7.65e-20
C19288 a_14401_32519# a_5649_42852# 3.64e-19
C19289 a_15493_43396# a_15567_42826# 4.1e-20
C19290 a_10555_44260# a_10796_42968# 6.32e-21
C19291 a_14539_43914# a_15959_42545# 3.47e-21
C19292 a_n356_44636# a_11551_42558# 1.46e-19
C19293 a_19721_31679# a_22775_42308# 3.9e-21
C19294 a_20974_43370# a_13678_32519# 0.020999f
C19295 a_5891_43370# a_8337_42558# 4.22e-21
C19296 a_8685_43396# a_7466_43396# 3.33e-20
C19297 a_n97_42460# a_17433_43396# 1.55e-19
C19298 a_18143_47464# RST_Z 2.7e-19
C19299 a_11599_46634# CLK 6.41e-19
C19300 a_10227_46804# START 0.088203f
C19301 a_17486_43762# VDD 4.6e-19
C19302 a_16115_45572# a_16237_45028# 4.93e-20
C19303 a_11823_42460# a_8975_43940# 7.95e-20
C19304 a_16147_45260# a_16922_45042# 0.016249f
C19305 a_12427_45724# a_12607_44458# 3.74e-21
C19306 a_10193_42453# a_16979_44734# 0.016398f
C19307 a_6472_45840# a_6109_44484# 7.09e-20
C19308 a_n967_45348# a_375_42282# 0.001506f
C19309 a_6431_45366# a_7229_43940# 1.72e-19
C19310 a_6171_45002# a_6709_45028# 0.021915f
C19311 a_3232_43370# a_7705_45326# 0.02181f
C19312 a_15567_42826# a_3483_46348# 8.48e-21
C19313 a_13291_42460# a_13059_46348# 0.007788f
C19314 a_13258_32519# a_13661_43548# 6.71e-21
C19315 a_20256_43172# a_19692_46634# 4.35e-19
C19316 a_5755_42308# a_5257_43370# 3.66e-19
C19317 a_6031_43396# a_n443_42852# 0.020526f
C19318 a_4361_42308# a_526_44458# 0.072573f
C19319 a_10835_43094# a_8953_45546# 5.45e-21
C19320 a_8387_43230# a_9290_44172# 1.54e-20
C19321 a_n3420_39072# a_n2312_39304# 6.52e-19
C19322 a_19237_31679# VCM 0.03748f
C19323 a_413_45260# a_3815_47204# 5.94e-19
C19324 a_3537_45260# a_2063_45854# 1.21e-20
C19325 a_4574_45260# a_584_46384# 0.001263f
C19326 a_7276_45260# a_n971_45724# 2.9e-22
C19327 a_21188_45572# a_10227_46804# 1.59e-21
C19328 a_3357_43084# a_14311_47204# 1.17e-19
C19329 a_2437_43646# a_15507_47210# 0.027848f
C19330 a_20623_45572# a_18479_47436# 0.007543f
C19331 a_20273_45572# a_18597_46090# 0.048762f
C19332 a_15861_45028# a_n881_46662# 0.153795f
C19333 a_8746_45002# a_2107_46812# 0.020783f
C19334 a_5263_45724# a_4817_46660# 2.13e-19
C19335 a_6472_45840# a_4646_46812# 0.129446f
C19336 a_13163_45724# a_n743_46660# 1.17e-20
C19337 a_15037_45618# a_768_44030# 1.6e-21
C19338 a_n2661_45546# a_n452_45724# 0.007419f
C19339 a_n2840_45546# a_n1099_45572# 3.93e-20
C19340 a_n2956_38216# a_n1079_45724# 5.55e-20
C19341 a_n2472_45546# a_n863_45724# 1.45e-19
C19342 a_13467_32519# a_19987_42826# 5.32e-19
C19343 a_19862_44208# a_13258_32519# 3.59e-19
C19344 a_1568_43370# a_2351_42308# 3.07e-21
C19345 a_4093_43548# a_1755_42282# 1.31e-21
C19346 a_5649_42852# a_18817_42826# 1.52e-20
C19347 a_4361_42308# a_19164_43230# 1.97e-20
C19348 a_12281_43396# a_12800_43218# 9.09e-21
C19349 a_15095_43370# a_13291_42460# 6.1e-21
C19350 a_14205_43396# a_14635_42282# 6.79e-20
C19351 a_21076_30879# a_22469_39537# 8.69e-20
C19352 a_17339_46660# START 0.00197f
C19353 a_765_45546# RST_Z 0.002113f
C19354 a_7754_39300# a_5088_37509# 1.3e-19
C19355 a_n971_45724# a_n746_45260# 0.393354f
C19356 a_n1605_47204# a_n785_47204# 2e-19
C19357 a_n452_47436# a_n237_47217# 0.061523f
C19358 a_n1741_47186# a_1209_47178# 0.046323f
C19359 a_n2109_47186# a_1431_47204# 0.050586f
C19360 a_n2497_47436# a_584_46384# 0.06459f
C19361 a_n815_47178# a_n23_47502# 9.5e-20
C19362 a_3823_42558# VDD 0.170296f
C19363 a_n2293_42834# a_n23_44458# 8.19e-21
C19364 a_1423_45028# a_3363_44484# 8.49e-19
C19365 a_13556_45296# a_15433_44458# 0.1084f
C19366 a_1307_43914# a_n2661_42834# 3.43601f
C19367 a_9482_43914# a_15146_44811# 0.006879f
C19368 a_2711_45572# a_19741_43940# 0.005487f
C19369 a_n913_45002# a_3422_30871# 0.145467f
C19370 a_13258_32519# a_4185_45028# 0.068774f
C19371 a_15051_42282# a_2324_44458# 2.79e-19
C19372 a_17141_43172# a_n357_42282# 7.19e-19
C19373 a_11691_44458# a_13747_46662# 3.75e-19
C19374 a_13159_45002# a_6755_46942# 1.18e-21
C19375 a_20193_45348# a_13661_43548# 1.38e-20
C19376 a_16501_45348# a_n743_46660# 8.3e-19
C19377 a_413_45260# a_14976_45028# 3.29e-20
C19378 a_9049_44484# a_2324_44458# 0.102942f
C19379 a_12427_45724# a_10903_43370# 0.083943f
C19380 a_11962_45724# a_12005_46116# 1.83e-19
C19381 a_11652_45724# a_12594_46348# 5.18e-20
C19382 a_6469_45572# a_5937_45572# 1.2e-19
C19383 a_n452_44636# a_n1613_43370# 0.001807f
C19384 a_12607_44458# a_11453_44696# 7.57e-20
C19385 a_n2661_42834# a_n443_46116# 0.075503f
C19386 a_n2661_43922# a_4791_45118# 0.034957f
C19387 a_22591_43396# a_22775_42308# 1.54e-19
C19388 a_10341_42308# a_11633_42558# 2.57e-19
C19389 a_12089_42308# a_5742_30871# 1.26e-19
C19390 a_14209_32519# a_21613_42308# 9.39e-21
C19391 a_13678_32519# a_22397_42558# 0.001628f
C19392 a_3080_42308# C0_dummy_N_btm 1.48e-19
C19393 a_15928_47570# a_16119_47582# 4.61e-19
C19394 a_12891_46348# a_13759_47204# 1.25e-20
C19395 a_768_44030# a_13569_47204# 8.63e-20
C19396 a_12549_44172# a_13675_47204# 5.51e-19
C19397 a_8128_46384# a_5807_45002# 0.023925f
C19398 a_n2312_40392# a_n2438_43548# 6.39e-22
C19399 a_4883_46098# a_2107_46812# 2.95673f
C19400 a_4915_47217# a_7577_46660# 1.88e-19
C19401 a_n1435_47204# a_4817_46660# 1.96e-20
C19402 a_6151_47436# a_5257_43370# 0.009542f
C19403 a_2063_45854# a_6969_46634# 0.00119f
C19404 a_n1151_42308# a_10467_46802# 0.031981f
C19405 a_21359_45002# a_11341_43940# 1.28e-20
C19406 a_n2661_44458# a_10949_43914# 1.28e-19
C19407 a_11827_44484# a_21115_43940# 0.005833f
C19408 a_2711_45572# a_17333_42852# 2.07e-20
C19409 a_7499_43078# a_9127_43156# 0.08498f
C19410 a_17061_44734# a_17517_44484# 0.004238f
C19411 a_20193_45348# a_19862_44208# 0.041264f
C19412 a_n356_44636# a_1467_44172# 0.061333f
C19413 a_3232_43370# a_2982_43646# 0.416054f
C19414 a_5111_44636# a_3539_42460# 2.98e-20
C19415 a_14180_45002# VDD 0.151315f
C19416 a_n1630_35242# EN_VIN_BSTR_N 0.009773f
C19417 a_1568_43370# a_584_46384# 0.057089f
C19418 a_13105_45348# a_2324_44458# 2.03e-19
C19419 a_6945_45348# a_6945_45028# 0.009798f
C19420 a_n2661_45010# a_n2293_45546# 0.014846f
C19421 a_3357_43084# a_n755_45592# 0.00172f
C19422 a_n2109_45247# a_n2661_45546# 0.003324f
C19423 a_n2293_45010# a_n2472_45546# 3.35e-19
C19424 a_n2472_45002# a_n2956_38216# 0.00378f
C19425 a_2809_45348# a_526_44458# 0.001579f
C19426 a_13159_45002# a_8049_45260# 4.59e-21
C19427 a_18989_43940# a_19123_46287# 2.88e-20
C19428 a_17973_43940# a_12549_44172# 0.015874f
C19429 a_11967_42832# a_6755_46942# 0.030705f
C19430 a_20193_45348# a_4185_45028# 0.015456f
C19431 a_n1177_44458# a_n1853_46287# 5.46e-23
C19432 a_n2267_44484# a_n1641_46494# 4.94e-19
C19433 a_n2661_44458# a_376_46348# 9.54e-22
C19434 a_3381_47502# VDD 0.197761f
C19435 a_14113_42308# a_17124_42282# 4.43e-19
C19436 a_8685_42308# a_7174_31319# 4.88e-21
C19437 a_n4318_37592# a_n3420_38528# 0.024768f
C19438 a_n3674_38216# a_n4064_38528# 0.020875f
C19439 a_n881_46662# a_5068_46348# 0.078135f
C19440 a_n1613_43370# a_5164_46348# 3.39e-19
C19441 a_11453_44696# a_10903_43370# 0.040346f
C19442 a_12465_44636# a_13759_46122# 0.018063f
C19443 a_4883_46098# a_14493_46090# 0.00233f
C19444 a_13507_46334# a_15015_46420# 0.005128f
C19445 a_16327_47482# a_21137_46414# 1.42e-20
C19446 a_10227_46804# a_19553_46090# 4.1e-21
C19447 a_18479_47436# a_18819_46122# 6.05e-20
C19448 a_15811_47375# a_10809_44734# 0.049971f
C19449 a_16241_47178# a_6945_45028# 0.011279f
C19450 a_18597_46090# a_18189_46348# 4.44e-19
C19451 a_n443_46116# a_5066_45546# 0.130975f
C19452 a_n1151_42308# a_8034_45724# 0.040415f
C19453 a_4791_45118# a_6419_46482# 9.06e-19
C19454 a_9804_47204# a_3483_46348# 6.33e-21
C19455 a_6755_46942# a_12251_46660# 0.033714f
C19456 a_2609_46660# a_765_45546# 0.009946f
C19457 a_22612_30879# a_21076_30879# 0.056101f
C19458 a_16979_44734# a_16137_43396# 8.54e-22
C19459 a_1307_43914# a_n2293_42282# 0.004191f
C19460 a_n2661_43922# a_8791_43396# 3e-20
C19461 a_n2661_42834# a_9396_43370# 8.6e-21
C19462 a_14539_43914# a_16243_43396# 0.029808f
C19463 a_20512_43084# a_21381_43940# 0.019564f
C19464 a_11823_42460# a_15803_42450# 8.2e-20
C19465 a_18114_32519# a_13678_32519# 0.055126f
C19466 a_3600_43914# a_3992_43940# 0.016359f
C19467 a_5891_43370# a_8423_43396# 7.18e-21
C19468 a_13249_42308# a_13657_42558# 0.002219f
C19469 a_10193_42453# a_13657_42308# 5.7e-19
C19470 a_16112_44458# a_16547_43609# 1.97e-19
C19471 a_2998_44172# a_5025_43940# 5.5e-20
C19472 a_20679_44626# VDD 0.439119f
C19473 a_10490_45724# a_11962_45724# 0.114064f
C19474 a_10193_42453# a_11823_42460# 0.235429f
C19475 a_11322_45546# a_11652_45724# 0.26844f
C19476 a_7227_45028# a_8192_45572# 7.21e-20
C19477 a_2711_45572# a_11778_45572# 8.22e-19
C19478 C0_P_btm EN_VIN_BSTR_P 0.12803f
C19479 a_4190_30871# a_13747_46662# 4.43e-21
C19480 a_743_42282# a_5807_45002# 2.41e-20
C19481 a_20301_43646# a_13661_43548# 0.072262f
C19482 a_6109_44484# a_n357_42282# 1.45e-19
C19483 a_3905_42865# a_2324_44458# 1.55e-19
C19484 a_n1641_43230# a_n1613_43370# 0.152896f
C19485 a_10922_42852# a_10227_46804# 0.159426f
C19486 a_n2293_42282# a_n443_46116# 2.82e-20
C19487 a_15009_46634# VDD 0.205396f
C19488 a_1138_42852# a_1823_45246# 7.31e-20
C19489 a_1208_46090# a_167_45260# 0.001892f
C19490 a_3877_44458# a_n755_45592# 0.001347f
C19491 a_6755_46942# a_13259_45724# 0.021651f
C19492 a_4646_46812# a_n357_42282# 0.030404f
C19493 a_1799_45572# a_2277_45546# 2.46e-19
C19494 a_8270_45546# a_10037_46155# 4.27e-20
C19495 a_n2293_46098# a_5164_46348# 2.77e-19
C19496 a_19123_46287# a_18189_46348# 1.43e-20
C19497 a_18285_46348# a_17957_46116# 0.12677f
C19498 a_13059_46348# a_10809_44734# 0.003202f
C19499 a_16721_46634# a_6945_45028# 6e-20
C19500 a_5932_42308# a_n4064_37440# 1.17e-19
C19501 a_19478_44306# a_743_42282# 1.05e-20
C19502 a_20269_44172# a_4190_30871# 4.64e-20
C19503 a_4235_43370# a_3539_42460# 0.005553f
C19504 a_4699_43561# a_3626_43646# 5.64e-20
C19505 a_4905_42826# a_2982_43646# 1.34e-19
C19506 a_n97_42460# a_8147_43396# 8.39e-22
C19507 a_14021_43940# a_18525_43370# 0.007346f
C19508 a_21398_44850# a_21356_42826# 1.64e-20
C19509 a_n2661_42282# a_n1076_43230# 2.25e-20
C19510 a_3422_30871# a_20922_43172# 0.045027f
C19511 a_9313_44734# a_15597_42852# 4.48e-19
C19512 a_15493_43396# a_20556_43646# 1.31e-20
C19513 a_11341_43940# a_16823_43084# 2.12e-19
C19514 a_6765_43638# VDD 0.218204f
C19515 a_8696_44636# a_16751_45260# 0.265287f
C19516 a_15861_45028# a_1307_43914# 0.067929f
C19517 a_10193_42453# a_16321_45348# 9.06e-20
C19518 a_n2840_45002# a_n2472_45002# 7.52e-19
C19519 a_n4064_38528# w_1575_34946# 7.84e-19
C19520 a_21195_42852# a_19692_46634# 6.29e-21
C19521 a_13460_43230# a_13059_46348# 5.21e-21
C19522 a_10617_44484# CLK 6.69e-19
C19523 a_2711_45572# a_768_44030# 0.529995f
C19524 a_3775_45552# a_n881_46662# 0.002767f
C19525 a_8746_45002# a_11453_44696# 0.002934f
C19526 a_8696_44636# a_4915_47217# 0.02426f
C19527 a_8049_45260# a_13259_45724# 0.895805f
C19528 a_14358_43442# a_5534_30871# 0.002889f
C19529 a_5649_42852# a_22223_43396# 0.165664f
C19530 a_14205_43396# a_14543_43071# 9.94e-20
C19531 a_12281_43396# a_10341_42308# 2.53e-20
C19532 a_15095_43370# a_13460_43230# 5.97e-21
C19533 a_14579_43548# a_15279_43071# 0.108607f
C19534 a_13678_32519# a_13887_32519# 10.751599f
C19535 a_4361_42308# a_14209_32519# 8.23e-20
C19536 a_12800_43218# VDD 0.078978f
C19537 a_19431_45546# a_17517_44484# 1.08e-20
C19538 a_2711_45572# a_13483_43940# 1.84e-21
C19539 a_14403_45348# a_14309_45028# 1.26e-19
C19540 a_327_44734# a_n356_44636# 0.085841f
C19541 a_6171_45002# a_16112_44458# 5.94e-20
C19542 a_8953_45002# a_10440_44484# 1.69e-19
C19543 a_n2017_45002# a_5891_43370# 0.065487f
C19544 a_10796_42968# a_n443_42852# 1.54e-19
C19545 a_15567_42826# a_n357_42282# 0.008527f
C19546 a_1606_42308# a_9290_44172# 9.18e-20
C19547 a_5883_43914# a_584_46384# 2.91e-20
C19548 a_11691_44458# a_11599_46634# 7.06e-20
C19549 a_18315_45260# a_18597_46090# 1.77e-20
C19550 a_21359_45002# a_16327_47482# 2.1e-19
C19551 SINGLE_ENDED VDD 0.210835f
C19552 a_5093_45028# a_n881_46662# 8.78e-20
C19553 a_3232_43370# a_2107_46812# 0.026265f
C19554 a_413_45260# a_3524_46660# 4.83e-21
C19555 a_2680_45002# a_2443_46660# 3.28e-21
C19556 a_2437_43646# a_7715_46873# 2.14e-19
C19557 a_8953_45002# a_n743_46660# 0.001504f
C19558 a_16223_45938# a_15368_46634# 6.08e-20
C19559 a_9482_43914# a_n2661_46634# 9.45e-19
C19560 a_15861_45028# a_17609_46634# 2.54e-19
C19561 a_3638_45822# a_n2293_46098# 4.88e-19
C19562 a_15743_43084# a_15051_42282# 5.67e-19
C19563 a_17333_42852# a_16877_42852# 0.003649f
C19564 a_5649_42852# a_5934_30871# 0.058776f
C19565 a_743_42282# a_9223_42460# 0.010592f
C19566 a_13887_32519# a_6123_31319# 1.56e-19
C19567 a_17701_42308# a_17749_42852# 0.004244f
C19568 a_18083_42858# a_17665_42852# 2.63e-19
C19569 a_4361_42308# a_4169_42308# 7.22e-19
C19570 a_1177_38525# VDD 0.373535f
C19571 a_6151_47436# a_5807_45002# 0.099462f
C19572 a_13381_47204# a_12891_46348# 0.002658f
C19573 a_11459_47204# a_12549_44172# 1.19e-20
C19574 a_9313_45822# a_768_44030# 2.99e-20
C19575 a_n1435_47204# a_11309_47204# 1.78e-20
C19576 a_15811_47375# a_n881_46662# 1.05e-19
C19577 a_12465_44636# a_22731_47423# 0.002949f
C19578 a_2063_45854# a_n2293_46634# 0.004931f
C19579 a_n971_45724# a_383_46660# 1.21e-19
C19580 a_n237_47217# a_33_46660# 7.19e-21
C19581 a_n23_47502# a_171_46873# 0.001553f
C19582 a_n785_47204# a_n133_46660# 0.001087f
C19583 a_327_47204# a_n2438_43548# 2.1e-19
C19584 a_1209_47178# a_n743_46660# 9.52e-20
C19585 a_1431_47204# a_n1925_46634# 1.02e-20
C19586 a_2905_45572# a_n2661_46634# 0.029475f
C19587 a_n746_45260# a_601_46902# 0.004287f
C19588 a_4883_46098# a_11453_44696# 0.071224f
C19589 a_15415_45028# a_11341_43940# 7.47e-21
C19590 a_16112_44458# a_14673_44172# 0.077293f
C19591 a_10193_42453# a_18429_43548# 0.002926f
C19592 a_14537_43396# a_15493_43940# 8.79e-19
C19593 a_9482_43914# a_9895_44260# 0.005015f
C19594 a_11823_42460# a_16137_43396# 6.91e-20
C19595 a_n1243_44484# a_n2661_43922# 2.55e-19
C19596 a_n998_44484# a_n2661_42834# 2.81e-19
C19597 a_5147_45002# a_3737_43940# 2.51e-20
C19598 a_20712_42282# a_n357_42282# 0.173926f
C19599 a_20528_45572# VDD 0.08228f
C19600 a_1423_45028# a_3147_46376# 8.68e-21
C19601 a_3602_45348# a_1823_45246# 0.001718f
C19602 a_20273_45572# a_8049_45260# 0.040989f
C19603 a_18579_44172# a_19321_45002# 0.00855f
C19604 a_4223_44672# a_3090_45724# 0.269823f
C19605 a_18184_42460# a_17339_46660# 3.97e-20
C19606 a_14127_45572# a_13259_45724# 2.92e-19
C19607 a_n2956_37592# a_n2956_38680# 0.047258f
C19608 en_comp a_n2956_39304# 8.4e-19
C19609 a_10775_45002# a_9290_44172# 0.215292f
C19610 a_9482_43914# a_8199_44636# 0.276776f
C19611 a_n809_44244# a_n1613_43370# 0.291484f
C19612 a_6171_45002# a_13925_46122# 2.53e-20
C19613 a_5147_45002# a_2324_44458# 0.056065f
C19614 a_10729_43914# a_12861_44030# 3.15e-20
C19615 a_5267_42460# a_5742_30871# 1.46e-20
C19616 a_7963_42308# a_5934_30871# 0.002785f
C19617 a_1606_42308# a_15051_42282# 1.09e-19
C19618 a_20256_43172# a_20107_42308# 1.36e-19
C19619 a_6123_31319# a_8515_42308# 8.12e-20
C19620 a_22400_42852# a_19511_42282# 2.86e-21
C19621 a_11530_34132# EN_VIN_BSTR_N 1.02927f
C19622 a_5807_45002# a_19466_46812# 0.178376f
C19623 a_13661_43548# a_19333_46634# 0.011985f
C19624 a_13747_46662# a_15227_44166# 0.05203f
C19625 a_5385_46902# a_5275_47026# 0.097745f
C19626 a_5907_46634# a_6540_46812# 0.017547f
C19627 a_5167_46660# a_5072_46660# 0.049827f
C19628 a_3877_44458# a_5429_46660# 0.00211f
C19629 a_12891_46348# a_13170_46660# 2.99e-19
C19630 a_12549_44172# a_12925_46660# 3.4e-20
C19631 a_n2661_46634# a_12816_46660# 5.55e-19
C19632 a_n881_46662# a_13059_46348# 0.642888f
C19633 a_11453_44696# a_21188_46660# 0.047802f
C19634 a_10227_46804# a_12741_44636# 0.188309f
C19635 a_18597_46090# a_20202_43084# 0.04177f
C19636 a_13507_46334# a_18900_46660# 9.83e-19
C19637 a_6545_47178# a_3483_46348# 2.08e-20
C19638 a_4915_47217# a_4704_46090# 5.74e-20
C19639 a_n2109_47186# a_2324_44458# 0.004259f
C19640 a_2063_45854# a_9625_46129# 0.001267f
C19641 a_n443_46116# a_5068_46348# 9.9e-19
C19642 a_4791_45118# a_5164_46348# 0.42219f
C19643 a_n1151_42308# a_8016_46348# 0.580516f
C19644 a_21359_45002# a_10341_43396# 7.35e-21
C19645 a_20835_44721# a_15493_43940# 7.97e-20
C19646 a_19279_43940# a_11341_43940# 0.003029f
C19647 a_1414_42308# a_3499_42826# 0.023314f
C19648 a_5343_44458# a_6293_42852# 1.91e-20
C19649 a_4223_44672# a_6547_43396# 3.73e-19
C19650 a_11823_42460# a_n784_42308# 5.93e-20
C19651 a_2127_44172# a_2253_44260# 0.013015f
C19652 a_375_42282# a_n1853_43023# 2.99e-20
C19653 a_18579_44172# a_20623_43914# 1.89e-20
C19654 a_n2661_42834# a_10867_43940# 6.15e-20
C19655 a_n1059_45260# a_16795_42852# 0.182174f
C19656 a_n2017_45002# a_17595_43084# 0.016123f
C19657 en_comp a_5534_30871# 0.021896f
C19658 a_n1655_44484# VDD 1.27e-19
C19659 a_n4315_30879# VCM 0.473529f
C19660 a_n4064_40160# VREF 1.12e-19
C19661 a_n4209_38502# a_n1838_35608# 1.6e-19
C19662 a_n4209_39304# C6_P_btm 0.001067f
C19663 a_n3565_39304# C8_P_btm 1.15e-19
C19664 a_n3420_39072# C10_P_btm 3.37e-20
C19665 a_22469_40625# a_13259_45724# 1.39e-19
C19666 a_n4209_37414# a_n2956_38216# 4.59e-21
C19667 a_15868_43402# a_10227_46804# 2.96e-20
C19668 a_16823_43084# a_16327_47482# 0.535969f
C19669 a_21487_43396# a_12861_44030# 7.46e-20
C19670 a_16243_43396# a_11453_44696# 1.19e-21
C19671 a_14673_44172# a_13925_46122# 2.92e-21
C19672 a_11649_44734# a_10809_44734# 2.53e-19
C19673 a_n2661_43922# a_6945_45028# 1.07e-19
C19674 a_18989_43940# a_8049_45260# 6.26e-20
C19675 a_5891_43370# a_526_44458# 1.12739f
C19676 a_15493_43396# a_19692_46634# 0.001909f
C19677 a_15493_43940# a_3090_45724# 0.255251f
C19678 a_n809_44244# a_n2293_46098# 1.32e-20
C19679 a_n3565_39590# a_n3565_38216# 0.031123f
C19680 a_n3420_39616# a_n4209_38216# 0.027924f
C19681 a_n4064_39072# a_n2860_39072# 0.003765f
C19682 a_2959_46660# VDD 0.19762f
C19683 a_20273_46660# a_21350_47026# 1.46e-19
C19684 a_20411_46873# a_20719_46660# 2.12e-19
C19685 a_4817_46660# a_526_44458# 4.05e-20
C19686 a_19321_45002# a_19443_46116# 0.003684f
C19687 a_4955_46873# a_n1925_42282# 6.24e-20
C19688 a_n743_46660# a_11601_46155# 6.77e-19
C19689 a_18285_46348# a_11415_45002# 1.48e-20
C19690 a_17339_46660# a_12741_44636# 0.032832f
C19691 a_22485_44484# a_13678_32519# 3.76e-22
C19692 a_10405_44172# a_10695_43548# 1.89e-19
C19693 a_20512_43084# a_5649_42852# 0.141324f
C19694 a_9313_44734# a_18083_42858# 0.05022f
C19695 a_n2293_42834# a_5267_42460# 5.73e-21
C19696 a_3422_30871# a_17364_32525# 0.007014f
C19697 a_20193_45348# a_20573_43172# 1.16e-20
C19698 en_comp a_19647_42308# 4.59e-20
C19699 a_n913_45002# a_7174_31319# 0.02792f
C19700 a_19431_45546# a_19256_45572# 0.233657f
C19701 a_18909_45814# a_18799_45938# 0.097745f
C19702 a_7499_43078# a_10951_45334# 0.008335f
C19703 a_16147_45260# a_17668_45572# 5.57e-19
C19704 a_18691_45572# a_18596_45572# 0.049827f
C19705 a_11962_45724# a_6171_45002# 8.2e-19
C19706 a_10053_45546# a_8953_45002# 0.009534f
C19707 a_11206_38545# RST_Z 0.382319f
C19708 a_n3420_37440# VCM 0.033198f
C19709 a_10405_44172# a_n357_42282# 2.3e-20
C19710 a_4093_43548# a_2324_44458# 1.63e-20
C19711 a_n4064_37440# VREF 1.56e-19
C19712 a_19335_46494# VDD 0.198512f
C19713 a_12791_45546# a_n1741_47186# 1.89e-19
C19714 a_3775_45552# a_n443_46116# 9.26e-22
C19715 a_7230_45938# a_2063_45854# 0.016263f
C19716 a_6511_45714# a_6151_47436# 0.3215f
C19717 a_6472_45840# a_6545_47178# 6.79e-20
C19718 a_2711_45572# a_9067_47204# 1.64e-21
C19719 a_7227_45028# a_4915_47217# 4.56e-21
C19720 a_n2293_46098# a_3316_45546# 0.008121f
C19721 a_167_45260# a_n2661_45546# 0.084316f
C19722 a_472_46348# a_380_45546# 3.1e-21
C19723 a_376_46348# a_n1099_45572# 6.04e-21
C19724 a_1138_42852# a_n2293_45546# 0.021487f
C19725 a_10903_43370# a_14180_46482# 0.001228f
C19726 a_18189_46348# a_8049_45260# 0.030061f
C19727 a_12594_46348# a_12379_46436# 0.04209f
C19728 a_11189_46129# a_11601_46155# 0.007009f
C19729 a_1414_42308# a_3318_42354# 0.001376f
C19730 a_16243_43396# a_17324_43396# 0.102355f
C19731 a_16409_43396# a_16759_43396# 0.20669f
C19732 a_2982_43646# a_2905_42968# 3.17e-20
C19733 a_10341_43396# a_16823_43084# 0.044262f
C19734 a_19319_43548# a_19987_42826# 8.72e-20
C19735 a_n97_42460# a_13113_42826# 4.45e-21
C19736 a_9313_44734# a_22775_42308# 0.011571f
C19737 a_11967_42832# a_14456_42282# 4.2e-20
C19738 a_n4318_39768# a_n3674_37592# 0.024842f
C19739 a_16547_43609# a_17499_43370# 1.26e-20
C19740 a_3626_43646# a_1847_42826# 3.62e-21
C19741 a_n1441_43940# COMP_P 2.51e-20
C19742 a_16137_43396# a_18429_43548# 9.56e-19
C19743 a_10341_42308# VDD 0.931019f
C19744 a_16147_45260# a_17970_44736# 2.03e-19
C19745 a_18175_45572# a_17767_44458# 6.65e-20
C19746 a_11787_45002# a_n2661_43370# 0.00108f
C19747 a_6171_45002# a_13807_45067# 1.73e-19
C19748 a_9114_42852# a_8953_45546# 1.98e-19
C19749 a_9061_43230# a_9290_44172# 2.91e-21
C19750 a_20556_43646# a_n357_42282# 4.02e-19
C19751 a_743_42282# a_n755_45592# 0.160592f
C19752 a_n3565_38502# a_n2312_38680# 0.134976f
C19753 a_5742_30871# a_3090_45724# 7.9e-19
C19754 a_n2302_37984# SMPL_ON_P 5.6e-20
C19755 a_15143_45578# a_6755_46942# 2.33e-21
C19756 a_8746_45002# a_10384_47026# 5.86e-21
C19757 a_3260_45572# a_3090_45724# 6.23e-19
C19758 a_2437_43646# a_13747_46662# 0.008951f
C19759 a_n659_45366# a_n881_46662# 8.3e-19
C19760 a_3232_43370# a_11453_44696# 0.132496f
C19761 a_13556_45296# a_10227_46804# 0.013693f
C19762 a_1307_43914# a_15811_47375# 1.46e-19
C19763 a_5837_45028# a_4791_45118# 5.56e-20
C19764 a_18083_42858# a_18599_43230# 0.113784f
C19765 a_3626_43646# a_15486_42560# 0.005343f
C19766 a_2982_43646# a_15803_42450# 4.86e-19
C19767 a_743_42282# a_20256_43172# 0.00713f
C19768 a_17333_42852# a_18817_42826# 1.28e-19
C19769 a_8685_43396# a_5934_30871# 4.81e-19
C19770 a_7466_43396# a_6123_31319# 4.05e-20
C19771 a_18057_42282# VDD 0.130308f
C19772 a_n2109_47186# a_n310_47570# 9.67e-19
C19773 a_n1741_47186# a_n2312_40392# 4.79e-19
C19774 a_n1920_47178# a_n2312_39304# 0.157528f
C19775 a_9067_47204# a_9313_45822# 0.013659f
C19776 a_7227_47204# a_n1435_47204# 0.001005f
C19777 a_6151_47436# a_14311_47204# 0.136645f
C19778 a_10193_42453# a_2982_43646# 0.231527f
C19779 a_n2661_44458# a_7640_43914# 0.005176f
C19780 a_11827_44484# a_n2661_43922# 0.32722f
C19781 a_11691_44458# a_10617_44484# 1.65e-20
C19782 a_626_44172# a_n2065_43946# 1.31e-21
C19783 a_375_42282# a_n1899_43946# 8.99e-21
C19784 a_n2017_45002# a_10807_43548# 0.0319f
C19785 a_7229_43940# a_6453_43914# 0.001044f
C19786 a_5205_44484# a_7542_44172# 3.34e-20
C19787 a_6171_42473# a_n357_42282# 0.010166f
C19788 a_5755_42308# a_n755_45592# 3.68e-19
C19789 a_14456_42282# a_13259_45724# 5.4e-19
C19790 a_8336_45822# VDD 0.004437f
C19791 a_17364_32525# VREF_GND 0.048253f
C19792 a_2889_44172# a_584_46384# 4.84e-20
C19793 a_7542_44172# a_n971_45724# 4.49e-21
C19794 a_n1441_43940# a_n2497_47436# 0.004491f
C19795 a_2437_43646# a_4419_46090# 3.77e-20
C19796 a_19279_43940# a_16327_47482# 0.446333f
C19797 a_19006_44850# a_18597_46090# 3.17e-20
C19798 a_21398_44850# a_12861_44030# 2.74e-20
C19799 a_n2661_42834# a_n1613_43370# 0.112184f
C19800 a_16842_45938# a_17715_44484# 4.81e-20
C19801 a_8696_44636# a_10809_44734# 0.117876f
C19802 a_17478_45572# a_6945_45028# 2.17e-21
C19803 a_12791_45546# a_10586_45546# 9.22e-21
C19804 a_3175_45822# a_n2661_45546# 2.16e-19
C19805 a_15143_45578# a_8049_45260# 0.001756f
C19806 a_n967_45348# a_n1853_46287# 3.76e-21
C19807 a_8975_43940# a_2107_46812# 0.075583f
C19808 a_n2661_45010# a_1138_42852# 0.017849f
C19809 a_9313_44734# a_12549_44172# 3.97e-19
C19810 a_n2293_42834# a_3090_45724# 0.023056f
C19811 a_3357_43084# a_3483_46348# 0.030022f
C19812 a_1307_43914# a_13059_46348# 0.04241f
C19813 a_n913_45002# a_n1076_46494# 8.43e-20
C19814 a_n745_45366# a_n901_46420# 7.11e-19
C19815 a_21671_42860# a_13258_32519# 6.52e-20
C19816 a_564_42282# a_1067_42314# 1.81e-19
C19817 a_n327_42558# a_1184_42692# 1.76e-19
C19818 a_n784_42308# a_961_42354# 0.038477f
C19819 a_10227_46804# a_13607_46688# 0.027032f
C19820 a_11599_46634# a_15227_44166# 0.101252f
C19821 a_15673_47210# a_16292_46812# 1.35e-19
C19822 a_15811_47375# a_17609_46634# 4.73e-20
C19823 a_16327_47482# a_15368_46634# 2.32e-20
C19824 a_2905_45572# a_765_45546# 0.039575f
C19825 a_n2661_46634# a_2443_46660# 0.021792f
C19826 a_n133_46660# a_2107_46812# 2.94e-21
C19827 a_601_46902# a_383_46660# 0.209641f
C19828 a_n2438_43548# a_1983_46706# 0.057412f
C19829 a_33_46660# a_1123_46634# 0.041798f
C19830 a_n2472_46634# a_n2661_46098# 2.78e-21
C19831 a_n743_46660# a_288_46660# 0.024827f
C19832 a_171_46873# a_948_46660# 5.47e-21
C19833 a_n1925_46634# a_n935_46688# 6.05e-19
C19834 a_n881_46662# a_7577_46660# 0.028487f
C19835 a_15415_45028# a_10341_43396# 3.51e-21
C19836 a_1423_45028# a_9803_43646# 3.46e-20
C19837 a_16979_44734# a_14021_43940# 3.43e-21
C19838 a_9313_44734# a_12429_44172# 9.29e-21
C19839 a_4223_44672# a_9165_43940# 1.39e-19
C19840 a_n2293_42834# a_6547_43396# 3.28e-20
C19841 a_1307_43914# a_15095_43370# 1.5e-20
C19842 a_3422_30871# a_19237_31679# 1.04e-19
C19843 a_n2293_43922# a_n2661_42282# 0.133253f
C19844 a_n356_44636# a_15493_43940# 9.87e-21
C19845 a_n2661_42834# a_7584_44260# 1.21e-19
C19846 a_n913_45002# a_21487_43396# 7.6e-21
C19847 a_19963_31679# a_17364_32525# 0.053794f
C19848 a_20447_31679# a_14209_32519# 0.051502f
C19849 a_n2017_45002# a_13467_32519# 2.68e-20
C19850 en_comp a_4190_30871# 0.086973f
C19851 a_18494_42460# VDD 0.73193f
C19852 a_4958_30871# CAL_P 0.007236f
C19853 a_14815_43914# a_12741_44636# 0.003697f
C19854 a_n2661_42834# a_n2293_46098# 0.029385f
C19855 a_n2661_43922# a_n2472_46090# 5.03e-21
C19856 a_5826_44734# a_3483_46348# 8.07e-19
C19857 a_20974_43370# a_12549_44172# 0.061866f
C19858 a_13565_43940# a_13661_43548# 0.017205f
C19859 a_1307_43914# a_3218_45724# 6.18e-21
C19860 a_626_44172# a_n755_45592# 0.100613f
C19861 a_18315_45260# a_8049_45260# 1.23e-20
C19862 a_2903_45348# a_n863_45724# 1.21e-20
C19863 a_1145_45348# a_n357_42282# 1.17e-20
C19864 a_13076_44458# a_13351_46090# 3.69e-21
C19865 a_10157_44484# a_2324_44458# 2.29e-21
C19866 a_n1352_43396# a_n1613_43370# 0.244933f
C19867 a_14205_43396# a_4915_47217# 8.72e-21
C19868 a_21887_42336# a_21973_42336# 0.006584f
C19869 a_21613_42308# a_22465_38105# 0.026117f
C19870 a_2266_47243# VDD 6.34e-20
C19871 a_n784_42308# C0_dummy_P_btm 2.62e-20
C19872 a_3877_44458# a_3483_46348# 0.083955f
C19873 a_10249_46116# a_11415_45002# 1.8e-20
C19874 a_16292_46812# a_16388_46812# 0.318472f
C19875 a_12816_46660# a_765_45546# 3.23e-20
C19876 a_n881_46662# a_5431_46482# 9.41e-19
C19877 a_n743_46660# a_15015_46420# 0.007103f
C19878 a_19594_46812# a_6945_45028# 0.014072f
C19879 a_n1925_46634# a_2324_44458# 8.77e-20
C19880 a_n1613_43370# a_5066_45546# 0.015391f
C19881 a_4883_46098# a_14180_46482# 0.001483f
C19882 a_16327_47482# a_19597_46482# 0.001903f
C19883 a_10227_46804# a_16375_45002# 7.63e-19
C19884 a_584_46384# a_1990_45899# 4.9e-19
C19885 a_n1151_42308# a_n1013_45572# 0.002324f
C19886 a_n443_46116# a_3218_45724# 9.08e-19
C19887 a_2063_45854# a_2277_45546# 0.057116f
C19888 a_n23_44458# a_n13_43084# 7.92e-19
C19889 a_19279_43940# a_10341_43396# 9.98e-20
C19890 a_n2661_42282# a_n97_42460# 0.025699f
C19891 a_9313_44734# a_21855_43396# 2.95e-19
C19892 a_9838_44484# a_9127_43156# 8.54e-21
C19893 a_3905_42865# a_3539_42460# 0.022817f
C19894 a_5883_43914# a_8952_43230# 3.2e-19
C19895 a_2382_45260# a_2713_42308# 1.18e-20
C19896 a_n913_45002# a_5932_42308# 0.220872f
C19897 a_n2017_45002# a_6773_42558# 0.001353f
C19898 a_3499_42826# VDD 0.333472f
C19899 a_n1630_35242# a_n971_45724# 0.028303f
C19900 a_n4064_37984# a_n923_35174# 0.005035f
C19901 a_11554_42852# a_10227_46804# 2.46e-19
C19902 a_n2293_42282# a_n1613_43370# 6.65e-20
C19903 a_5829_43940# a_5937_45572# 0.006959f
C19904 a_16867_43762# a_6755_46942# 2.42e-19
C19905 a_18599_43230# a_12549_44172# 3.17e-20
C19906 a_10083_42826# a_n2293_46634# 6.79e-20
C19907 a_5534_30871# a_13661_43548# 4.79e-20
C19908 a_22959_46660# VDD 0.299681f
C19909 a_10903_43370# a_13925_46122# 0.001937f
C19910 a_12594_46348# a_13351_46090# 2.97e-19
C19911 a_10355_46116# a_2324_44458# 3.32e-21
C19912 a_1343_38525# a_3754_39964# 3.37e-19
C19913 a_n4064_39072# a_n4064_37984# 0.044699f
C19914 a_n2293_46098# a_5066_45546# 0.140248f
C19915 a_472_46348# a_526_44458# 3.38e-21
C19916 a_1208_46090# a_1431_46436# 0.011458f
C19917 a_1176_45822# a_1337_46436# 9.42e-19
C19918 a_20202_43084# a_8049_45260# 0.042894f
C19919 a_17339_46660# a_16375_45002# 0.0296f
C19920 a_19692_46634# a_n357_42282# 1.03e-19
C19921 a_18285_46348# a_13259_45724# 3.76e-21
C19922 a_4958_30871# CAL_N 0.039702f
C19923 a_20974_43370# a_21855_43396# 0.029556f
C19924 a_n97_42460# a_16823_43084# 0.205258f
C19925 a_11341_43940# a_12545_42858# 1.16e-20
C19926 a_21381_43940# a_5649_42852# 1.8e-20
C19927 a_n356_44636# a_5742_30871# 0.120133f
C19928 a_14539_43914# a_15803_42450# 1.18e-22
C19929 a_2982_43646# a_16137_43396# 5.37e-19
C19930 a_14401_32519# a_13678_32519# 0.050672f
C19931 a_8685_43396# a_7221_43396# 7.37e-21
C19932 a_10227_46804# RST_Z 7.13e-19
C19933 a_14955_47212# CLK 3.68e-19
C19934 a_17591_47464# START 5.79e-19
C19935 a_16333_45814# a_16237_45028# 5.69e-20
C19936 a_16855_45546# a_11691_44458# 5.15e-22
C19937 a_10193_42453# a_14539_43914# 0.278963f
C19938 a_11962_45724# a_12607_44458# 5.74e-21
C19939 a_16147_45260# a_16501_45348# 9.04e-19
C19940 a_6194_45824# a_6109_44484# 1.36e-19
C19941 a_n913_45002# a_1423_45028# 1.35e-22
C19942 a_6171_45002# a_7229_43940# 0.010208f
C19943 a_3232_43370# a_6709_45028# 0.086072f
C19944 a_5111_44636# a_8953_45002# 3.17e-19
C19945 a_5342_30871# a_3483_46348# 8.76e-19
C19946 a_5534_30871# a_4185_45028# 0.05188f
C19947 a_19647_42308# a_13661_43548# 5.53e-21
C19948 a_2813_43396# a_n755_45592# 6.23e-21
C19949 a_1512_43396# a_n443_42852# 3.67e-19
C19950 a_10518_42984# a_8953_45546# 9.33e-20
C19951 a_8605_42826# a_9290_44172# 9.78e-21
C19952 a_10796_42968# a_8199_44636# 1.77e-20
C19953 a_n3690_39392# a_n2312_39304# 4.25e-19
C19954 a_19237_31679# VREF_GND 0.0061f
C19955 a_3357_43084# a_13487_47204# 5.65e-19
C19956 a_6171_45002# a_n237_47217# 1.47e-19
C19957 a_413_45260# a_3785_47178# 7.03e-19
C19958 a_3429_45260# a_2063_45854# 6.96e-22
C19959 a_5205_44484# a_n971_45724# 9.71e-22
C19960 a_3537_45260# a_584_46384# 0.108506f
C19961 a_20107_45572# a_18597_46090# 0.069963f
C19962 a_2437_43646# a_11599_46634# 0.006609f
C19963 a_20841_45814# a_18479_47436# 0.011134f
C19964 a_21363_45546# a_10227_46804# 3.24e-21
C19965 a_19610_45572# a_16327_47482# 0.00341f
C19966 a_18341_45572# a_11453_44696# 0.026938f
C19967 a_8696_44636# a_n881_46662# 0.178516f
C19968 a_14033_45822# a_768_44030# 0.005149f
C19969 a_2711_45572# a_5167_46660# 1.79e-20
C19970 a_6472_45840# a_3877_44458# 2.74e-20
C19971 a_6194_45824# a_4646_46812# 9.75e-21
C19972 a_12791_45546# a_n743_46660# 6.76e-20
C19973 a_14495_45572# a_n2293_46634# 5.19e-21
C19974 a_15037_45618# a_12549_44172# 7.69e-21
C19975 a_n2661_45546# a_n863_45724# 0.045552f
C19976 a_n2956_38216# a_n2293_45546# 0.005455f
C19977 a_2982_43646# a_n784_42308# 0.026817f
C19978 a_19862_44208# a_19647_42308# 1.12e-20
C19979 a_1756_43548# a_1755_42282# 1.07e-19
C19980 a_14358_43442# a_14635_42282# 9.06e-19
C19981 a_5649_42852# a_18249_42858# 2.71e-20
C19982 a_4361_42308# a_19339_43156# 3.07e-21
C19983 a_15493_43940# a_18727_42674# 1.18e-21
C19984 a_11341_43940# a_19332_42282# 5.32e-21
C19985 a_4520_42826# a_5111_42852# 0.047152f
C19986 a_n3674_39768# a_n4064_39072# 2.52e-21
C19987 a_14205_43396# a_13291_42460# 6.79e-20
C19988 a_21076_30879# a_22821_38993# 1.66e-19
C19989 VDAC_Pi VDAC_P 2.7e-19
C19990 a_3318_42354# VDD 0.203036f
C19991 a_n452_47436# a_n746_45260# 0.187792f
C19992 a_n1741_47186# a_327_47204# 0.013765f
C19993 a_n2109_47186# a_1239_47204# 0.080115f
C19994 a_n815_47178# a_n237_47217# 0.005891f
C19995 SMPL_ON_P a_n785_47204# 1.53e-19
C19996 a_9482_43914# a_15433_44458# 0.20244f
C19997 a_13556_45296# a_14815_43914# 0.378519f
C19998 a_11823_42460# a_14021_43940# 0.034191f
C19999 a_n2293_42834# a_n356_44636# 0.027771f
C20000 a_n1059_45260# a_3422_30871# 7.02e-20
C20001 a_19963_31679# a_19237_31679# 0.05162f
C20002 a_20447_31679# a_17730_32519# 0.051365f
C20003 a_19647_42308# a_4185_45028# 1.64e-19
C20004 a_9159_45572# a_3483_46348# 0.006021f
C20005 a_11691_44458# a_13661_43548# 0.263889f
C20006 a_18479_45785# a_18280_46660# 5.88e-20
C20007 a_22223_45036# a_19321_45002# 5.03e-20
C20008 a_20193_45348# a_5807_45002# 1.07e-19
C20009 a_18114_32519# a_12549_44172# 0.001232f
C20010 a_16405_45348# a_n743_46660# 7.86e-19
C20011 a_19113_45348# a_13747_46662# 2.83e-19
C20012 a_6171_45002# a_8270_45546# 0.027058f
C20013 a_3357_43084# a_14513_46634# 2.21e-20
C20014 a_413_45260# a_3090_45724# 0.135828f
C20015 en_comp a_15227_44166# 4.89e-21
C20016 a_7499_43078# a_2324_44458# 0.018394f
C20017 a_11962_45724# a_10903_43370# 0.357882f
C20018 a_11525_45546# a_12594_46348# 2.4e-19
C20019 a_6229_45572# a_5937_45572# 5.31e-19
C20020 a_n1352_44484# a_n1613_43370# 0.232498f
C20021 a_8975_43940# a_11453_44696# 0.027482f
C20022 a_13720_44458# a_12465_44636# 0.019702f
C20023 a_n2661_42834# a_4791_45118# 0.024946f
C20024 a_22591_43396# a_21613_42308# 2.05e-21
C20025 a_10341_42308# a_11551_42558# 1.68e-19
C20026 a_20749_43396# a_20712_42282# 1.09e-20
C20027 a_13887_32519# a_22775_42308# 0.006279f
C20028 a_12089_42308# a_11323_42473# 2.1e-19
C20029 a_13467_32519# a_21973_42336# 0.00115f
C20030 a_3080_42308# C0_dummy_P_btm 1.48e-19
C20031 a_12549_44172# a_13569_47204# 0.005506f
C20032 a_12891_46348# a_13675_47204# 2.93e-20
C20033 a_4915_47217# a_7715_46873# 3.51e-19
C20034 a_n1435_47204# a_4955_46873# 4.48e-20
C20035 a_5815_47464# a_5257_43370# 8.52e-20
C20036 a_2063_45854# a_6755_46942# 0.131005f
C20037 a_n1151_42308# a_10428_46928# 0.011222f
C20038 a_n356_44636# a_1115_44172# 0.006316f
C20039 a_n2661_44458# a_10729_43914# 1.94e-19
C20040 a_11827_44484# a_20935_43940# 0.003973f
C20041 a_742_44458# a_n2661_42282# 8.96e-21
C20042 a_7499_43078# a_8387_43230# 0.008868f
C20043 a_2711_45572# a_18083_42858# 4.96e-19
C20044 a_n699_43396# a_3499_42826# 1.7e-19
C20045 a_5111_44636# a_3626_43646# 1.57e-19
C20046 a_3232_43370# a_2896_43646# 1.75e-19
C20047 C10_N_btm VDD 2.40001f
C20048 a_13777_45326# VDD 0.145151f
C20049 a_n1630_35242# a_11530_34132# 0.029967f
C20050 VDAC_N a_21076_30879# 0.003547f
C20051 a_1049_43396# a_584_46384# 0.148494f
C20052 a_11915_45394# a_2324_44458# 8.14e-19
C20053 a_3357_43084# a_n357_42282# 0.010127f
C20054 a_n2293_45010# a_n2661_45546# 0.003149f
C20055 a_n2661_45010# a_n2956_38216# 0.005195f
C20056 a_2437_43646# a_1848_45724# 0.007112f
C20057 a_n2472_45002# a_n2472_45546# 0.026152f
C20058 a_13017_45260# a_8049_45260# 4.13e-20
C20059 a_n1644_44306# a_n2438_43548# 1.68e-20
C20060 a_17737_43940# a_12549_44172# 0.007227f
C20061 a_n2267_44484# a_n1423_46090# 5.61e-21
C20062 a_n2129_44697# a_n1641_46494# 1.53e-21
C20063 a_n2661_44458# a_n1076_46494# 3.36e-21
C20064 a_n1151_42308# VDD 2.57238f
C20065 a_14113_42308# a_16522_42674# 0.183181f
C20066 a_8325_42308# a_7174_31319# 4.88e-21
C20067 a_n881_46662# a_4704_46090# 0.049125f
C20068 a_n1613_43370# a_5068_46348# 1.7e-19
C20069 a_11453_44696# a_11387_46155# 3.7e-21
C20070 a_4883_46098# a_13925_46122# 0.006732f
C20071 a_13507_46334# a_14275_46494# 0.004384f
C20072 a_16327_47482# a_20708_46348# 0.001227f
C20073 a_18597_46090# a_17715_44484# 2.16e-20
C20074 a_10227_46804# a_18985_46122# 1.14e-20
C20075 a_15673_47210# a_6945_45028# 0.056077f
C20076 a_15507_47210# a_10809_44734# 6.3e-20
C20077 a_4791_45118# a_5066_45546# 0.238282f
C20078 a_2063_45854# a_8049_45260# 0.037406f
C20079 a_n1151_42308# a_8283_46482# 0.003687f
C20080 a_768_44030# a_1823_45246# 0.287407f
C20081 a_22612_30879# a_22959_46660# 6.06e-19
C20082 a_21588_30879# a_21076_30879# 8.21286f
C20083 a_6755_46942# a_12469_46902# 0.042969f
C20084 a_2443_46660# a_765_45546# 0.004286f
C20085 a_10249_46116# a_12251_46660# 1.57e-19
C20086 a_8128_46384# a_3483_46348# 1.2e-20
C20087 a_n2661_42834# a_8791_43396# 4.78e-20
C20088 a_n2661_43922# a_8147_43396# 2.31e-21
C20089 a_14539_43914# a_16137_43396# 0.004691f
C20090 a_3600_43914# a_3737_43940# 0.126609f
C20091 a_10193_42453# a_11897_42308# 0.00383f
C20092 a_13249_42308# a_13333_42558# 0.004402f
C20093 a_5891_43370# a_8317_43396# 5.61e-21
C20094 a_11823_42460# a_15764_42576# 4.46e-19
C20095 a_19279_43940# a_n97_42460# 1.72e-21
C20096 a_2998_44172# a_3992_43940# 5.62e-19
C20097 en_comp a_14635_42282# 4.34e-21
C20098 a_n1059_45260# a_18504_43218# 2.15e-20
C20099 a_20640_44752# VDD 0.246486f
C20100 a_10490_45724# a_11652_45724# 0.044431f
C20101 a_11322_45546# a_11525_45546# 0.055031f
C20102 a_7227_45028# a_8120_45572# 1.01e-19
C20103 a_8746_45002# a_11962_45724# 1.72e-21
C20104 a_10180_45724# a_11823_42460# 1.16e-20
C20105 a_2711_45572# a_11688_45572# 7.53e-19
C20106 C1_P_btm EN_VIN_BSTR_P 0.110046f
C20107 a_9672_43914# a_3483_46348# 0.125466f
C20108 a_15493_43940# a_21076_30879# 1.4e-20
C20109 a_4190_30871# a_13661_43548# 0.147163f
C20110 a_n23_44458# a_n23_45546# 6.98e-19
C20111 a_n1423_42826# a_n1613_43370# 0.15981f
C20112 a_10991_42826# a_10227_46804# 0.152133f
C20113 a_15567_42826# a_12861_44030# 0.004897f
C20114 a_14084_46812# VDD 0.087769f
C20115 a_n4064_39072# C0_P_btm 8.17e-21
C20116 a_1176_45822# a_1823_45246# 1.52e-20
C20117 a_472_46348# a_2521_46116# 5.15e-21
C20118 a_1208_46090# a_2202_46116# 0.001619f
C20119 a_n2661_46098# a_n443_42852# 9.75e-20
C20120 a_1799_45572# a_1609_45822# 0.079527f
C20121 a_3877_44458# a_n357_42282# 1.85e-23
C20122 a_8270_45546# a_9751_46155# 3.2e-20
C20123 a_18285_46348# a_18189_46348# 0.118603f
C20124 a_16388_46812# a_6945_45028# 3.6e-19
C20125 a_15227_46910# a_10809_44734# 0.006323f
C20126 a_9313_44734# a_14853_42852# 4.55e-21
C20127 a_15493_43396# a_743_42282# 1.59e-19
C20128 a_19862_44208# a_4190_30871# 0.023868f
C20129 a_458_43396# a_648_43396# 0.045837f
C20130 a_4235_43370# a_3626_43646# 1.4e-19
C20131 a_14021_43940# a_18429_43548# 0.00816f
C20132 a_4093_43548# a_3539_42460# 0.001457f
C20133 a_3080_42308# a_2982_43646# 0.095684f
C20134 a_n2661_42282# a_n901_43156# 5.27e-20
C20135 a_n97_42460# a_7112_43396# 0.002373f
C20136 a_3422_30871# a_19987_42826# 0.006447f
C20137 a_4223_44672# a_3823_42558# 7.52e-22
C20138 a_6197_43396# VDD 0.408793f
C20139 a_16680_45572# a_16751_45260# 9.83e-19
C20140 a_15861_45028# a_16019_45002# 0.04712f
C20141 a_8696_44636# a_1307_43914# 0.030679f
C20142 a_n2840_45002# a_n2661_45010# 0.189331f
C20143 a_19332_42282# a_16327_47482# 6.14e-19
C20144 a_17303_42282# a_10227_46804# 8.27e-21
C20145 a_20712_42282# a_12861_44030# 7.11e-22
C20146 a_15781_43660# a_2324_44458# 4.8e-19
C20147 a_5934_30871# a_768_44030# 3.24e-23
C20148 a_21356_42826# a_19692_46634# 5.5e-20
C20149 a_13635_43156# a_13059_46348# 3.86e-20
C20150 a_4190_30871# a_4185_45028# 0.16524f
C20151 a_743_42282# a_3483_46348# 2.47e-22
C20152 a_19240_46482# VDD 0.077608f
C20153 a_2711_45572# a_12549_44172# 2.05236f
C20154 a_7227_45028# a_n881_46662# 5.19e-19
C20155 a_3775_45552# a_n1613_43370# 1.56e-20
C20156 a_10193_42453# a_11453_44696# 0.071253f
C20157 a_11962_45724# a_4883_46098# 9.92e-21
C20158 a_11823_42460# a_13507_46334# 1.48e-19
C20159 a_8049_45260# a_14383_46116# 0.002486f
C20160 a_4905_42826# a_5193_42852# 0.016389f
C20161 a_14579_43548# a_5534_30871# 0.030066f
C20162 a_14358_43442# a_14543_43071# 0.001166f
C20163 a_10341_43396# a_12545_42858# 8.88e-20
C20164 a_9028_43914# a_9223_42460# 3.81e-21
C20165 a_13467_32519# a_14209_32519# 0.048306f
C20166 a_20556_43646# a_20749_43396# 0.018955f
C20167 a_13678_32519# a_22223_43396# 0.004894f
C20168 a_4361_42308# a_22591_43396# 2.7e-19
C20169 a_21855_43396# a_13887_32519# 3.59e-19
C20170 a_10752_42852# VDD 4.6e-19
C20171 a_1423_45028# a_n2661_44458# 0.164701f
C20172 a_2711_45572# a_12429_44172# 3.56e-22
C20173 a_14309_45348# a_14309_45028# 6.96e-20
C20174 a_9482_43914# a_5343_44458# 2.61e-20
C20175 a_n37_45144# a_n23_44458# 4.88e-19
C20176 a_413_45260# a_n356_44636# 5.61e-19
C20177 a_6171_45002# a_15004_44636# 4.14e-20
C20178 a_n1059_45260# a_7640_43914# 6.31e-21
C20179 a_6123_31319# a_1823_45246# 3.21e-20
C20180 a_5337_42558# a_4185_45028# 3.05e-19
C20181 a_17303_42282# a_17339_46660# 9.87e-21
C20182 a_10835_43094# a_n443_42852# 1.88e-19
C20183 a_5342_30871# a_n357_42282# 0.039779f
C20184 a_22612_30879# C10_N_btm 1.5848f
C20185 START VDD 0.114358f
C20186 a_n699_43396# a_n1151_42308# 0.022019f
C20187 a_21101_45002# a_16327_47482# 1.72e-19
C20188 a_n913_45002# a_4646_46812# 7.74e-20
C20189 a_8191_45002# a_n743_46660# 6.12e-22
C20190 a_5691_45260# a_2107_46812# 1.52e-20
C20191 a_413_45260# a_3699_46634# 3.59e-20
C20192 a_2437_43646# a_7411_46660# 7.33e-20
C20193 a_2382_45260# a_2443_46660# 8.11e-22
C20194 a_16020_45572# a_15368_46634# 5.92e-20
C20195 a_16855_45546# a_15227_44166# 8.57e-19
C20196 a_1260_45572# a_1138_42852# 0.001766f
C20197 a_3775_45552# a_n2293_46098# 0.003338f
C20198 a_7871_42858# a_n784_42308# 4.17e-21
C20199 a_15743_43084# a_14113_42308# 5.99e-20
C20200 a_5649_42852# a_7963_42308# 5.44e-20
C20201 a_743_42282# a_8791_42308# 0.008346f
C20202 a_10341_43396# a_19332_42282# 2.01e-21
C20203 a_13678_32519# a_5934_30871# 2.14e-19
C20204 a_17701_42308# a_17665_42852# 0.002723f
C20205 a_17595_43084# a_17749_42852# 0.010303f
C20206 a_17333_42852# a_16245_42852# 1.21e-20
C20207 a_4361_42308# a_3905_42308# 3.53e-19
C20208 a_5066_45546# DATA[3] 7.36e-22
C20209 a_3422_30871# a_n3420_37440# 0.0344f
C20210 a_n2216_38778# VDD 0.004173f
C20211 a_4915_47217# a_13747_46662# 0.710704f
C20212 a_11459_47204# a_12891_46348# 1.33e-19
C20213 a_15507_47210# a_n881_46662# 2.15e-19
C20214 a_12465_44636# a_22223_47212# 0.175138f
C20215 a_n1741_47186# a_1983_46706# 1.98e-20
C20216 a_n971_45724# a_601_46902# 1.1e-19
C20217 a_n746_45260# a_33_46660# 0.035747f
C20218 a_n237_47217# a_171_46873# 9.39e-20
C20219 a_n23_47502# a_n133_46660# 0.001147f
C20220 a_n785_47204# a_n2438_43548# 3.7e-19
C20221 a_327_47204# a_n743_46660# 9.48e-19
C20222 a_1239_47204# a_n1925_46634# 4.34e-20
C20223 a_584_46384# a_n2293_46634# 0.374996f
C20224 a_21496_47436# a_11453_44696# 4.71e-20
C20225 a_14797_45144# a_11341_43940# 1.37e-20
C20226 a_15004_44636# a_14673_44172# 0.039287f
C20227 a_10193_42453# a_17324_43396# 9.84e-20
C20228 a_11823_42460# a_13943_43396# 0.006456f
C20229 a_9482_43914# a_9801_44260# 0.003952f
C20230 a_18479_45785# a_2982_43646# 2.74e-20
C20231 a_n1243_44484# a_n2661_42834# 1.91e-19
C20232 a_20447_31679# a_17538_32519# 0.051306f
C20233 a_20107_42308# a_n357_42282# 5.18e-19
C20234 a_21188_45572# VDD 0.288663f
C20235 a_1423_45028# a_2804_46116# 1.3e-21
C20236 a_3495_45348# a_1823_45246# 2.54e-19
C20237 a_5093_45028# a_n2293_46098# 0.00251f
C20238 a_2779_44458# a_3090_45724# 5.81e-20
C20239 a_18315_45260# a_18285_46348# 5.03e-22
C20240 a_22485_44484# a_12549_44172# 2.07e-20
C20241 a_18753_44484# a_13661_43548# 0.00166f
C20242 a_16922_45042# a_20411_46873# 1.1e-20
C20243 a_20107_45572# a_8049_45260# 0.024509f
C20244 a_14033_45572# a_13259_45724# 2.45e-19
C20245 a_n2956_37592# a_n2956_39304# 0.044994f
C20246 a_n2810_45028# a_n2956_38680# 0.043221f
C20247 a_n1549_44318# a_n1613_43370# 0.16289f
C20248 a_6171_45002# a_13759_46122# 4.55e-20
C20249 a_413_45260# a_20075_46420# 4.37e-21
C20250 a_4558_45348# a_2324_44458# 9.57e-20
C20251 a_8953_45002# a_9290_44172# 0.002181f
C20252 a_11173_44260# a_2063_45854# 0.00917f
C20253 a_3823_42558# a_5742_30871# 1.54e-20
C20254 a_6123_31319# a_5934_30871# 15.8951f
C20255 a_13661_43548# a_15227_44166# 0.805606f
C20256 a_5907_46634# a_5732_46660# 0.233657f
C20257 a_5807_45002# a_19333_46634# 5.26e-20
C20258 a_4817_46660# a_5275_47026# 0.031068f
C20259 a_13747_46662# a_18834_46812# 0.00381f
C20260 a_3877_44458# a_5263_46660# 0.004328f
C20261 a_4646_46812# a_5894_47026# 2.49e-19
C20262 a_12891_46348# a_12925_46660# 4.23e-19
C20263 a_n2661_46634# a_12991_46634# 2.4e-19
C20264 a_7_47243# a_765_45546# 1.52e-21
C20265 a_11453_44696# a_21363_46634# 0.027075f
C20266 a_18479_47436# a_11415_45002# 0.033153f
C20267 a_10227_46804# a_20820_30879# 3.25e-20
C20268 a_13507_46334# a_18280_46660# 0.004063f
C20269 a_6151_47436# a_3483_46348# 2.14e-20
C20270 a_4791_45118# a_5068_46348# 0.003762f
C20271 a_n443_46116# a_4704_46090# 0.017894f
C20272 a_2063_45854# a_8953_45546# 5.65e-19
C20273 a_n1151_42308# a_7920_46348# 0.085186f
C20274 a_20679_44626# a_15493_43940# 1.03e-19
C20275 a_19279_43940# a_21115_43940# 1.52e-19
C20276 a_7281_43914# a_7542_44172# 0.060549f
C20277 a_18579_44172# a_20365_43914# 1.9e-19
C20278 a_n23_44458# a_104_43370# 1.77e-20
C20279 a_5343_44458# a_6031_43396# 9.7e-21
C20280 a_11827_44484# a_14955_43396# 5.17e-21
C20281 a_375_42282# a_n2157_42858# 2.28e-21
C20282 a_7499_43078# a_1606_42308# 5.24e-20
C20283 a_1414_42308# a_2537_44260# 4.33e-19
C20284 a_n2661_42834# a_10651_43940# 5.65e-20
C20285 a_5111_44636# a_8037_42858# 2.31e-19
C20286 a_3537_45260# a_8952_43230# 3.58e-20
C20287 a_n913_45002# a_15567_42826# 6.93e-20
C20288 a_n1059_45260# a_16414_43172# 0.094309f
C20289 a_n2017_45002# a_16795_42852# 6.5e-19
C20290 a_n1821_44484# VDD 4.61e-20
C20291 a_n4315_30879# VREF_GND 0.168163f
C20292 a_n4209_39304# C7_P_btm 0.184297f
C20293 a_n3565_39304# C9_P_btm 1.64e-19
C20294 a_22521_40599# a_13259_45724# 3.75e-19
C20295 a_n3565_37414# a_n2810_45572# 1.88e-20
C20296 a_16137_43396# a_11453_44696# 2.08e-20
C20297 a_15231_43396# a_10227_46804# 9.49e-20
C20298 a_17021_43396# a_16327_47482# 0.001903f
C20299 a_n2661_42834# a_6945_45028# 4.26e-20
C20300 a_14673_44172# a_13759_46122# 1.65e-20
C20301 a_8375_44464# a_526_44458# 5.01e-22
C20302 a_11341_43940# a_14976_45028# 2.74e-20
C20303 a_15493_43396# a_19466_46812# 2.36e-21
C20304 a_n4334_39392# a_n4334_38528# 0.050585f
C20305 a_n3565_39304# a_n4209_38502# 5.79402f
C20306 a_n2946_39072# a_n2860_39072# 0.011479f
C20307 a_n4209_39304# a_n3565_38502# 0.029672f
C20308 a_n3420_39072# a_n2216_39072# 7.08e-20
C20309 a_3177_46902# VDD 0.200982f
C20310 a_n3674_37592# a_n3420_37984# 0.172946f
C20311 a_n784_42308# a_n4064_37984# 0.00652f
C20312 a_n881_46662# a_2957_45546# 2.67e-20
C20313 a_10768_47026# a_9290_44172# 3.45e-19
C20314 a_8145_46902# a_6945_45028# 3.44e-20
C20315 a_6755_46942# a_17715_44484# 2.63e-19
C20316 a_15227_44166# a_4185_45028# 3.86e-20
C20317 a_20107_46660# a_20719_46660# 3.82e-19
C20318 a_768_44030# a_n2293_45546# 3.42e-20
C20319 a_n743_46660# a_11315_46155# 1.84e-19
C20320 a_5807_45002# a_20062_46116# 1.96e-20
C20321 a_10729_43914# a_9145_43396# 2.31e-20
C20322 a_14955_43940# a_8685_43396# 2.16e-19
C20323 a_14021_43940# a_2982_43646# 0.00345f
C20324 a_9313_44734# a_17701_42308# 0.008094f
C20325 a_n2293_42834# a_3823_42558# 2.98e-20
C20326 a_17730_32519# a_13467_32519# 0.054292f
C20327 a_20512_43084# a_13678_32519# 0.059475f
C20328 a_n2293_43922# a_12545_42858# 0.022686f
C20329 a_n1059_45260# a_7174_31319# 5.53e-20
C20330 en_comp a_19511_42282# 2.68e-20
C20331 a_n913_45002# a_20712_42282# 0.003267f
C20332 a_20447_31679# a_22465_38105# 4.46e-19
C20333 a_5907_45546# a_1423_45028# 3.15e-20
C20334 a_7499_43078# a_10775_45002# 0.00194f
C20335 a_17786_45822# a_17668_45572# 1.98e-20
C20336 a_18341_45572# a_18799_45938# 0.027606f
C20337 a_18691_45572# a_19256_45572# 7.99e-20
C20338 a_11652_45724# a_6171_45002# 0.072138f
C20339 a_9049_44484# a_8953_45002# 0.031391f
C20340 VDAC_P RST_Z 0.158793f
C20341 a_n3420_37440# VREF_GND 0.033872f
C20342 a_20749_43396# a_19692_46634# 3.6e-20
C20343 a_3626_43646# a_9290_44172# 0.014922f
C20344 a_19553_46090# VDD 0.204238f
C20345 a_6598_45938# a_4915_47217# 1.39e-21
C20346 a_6472_45840# a_6151_47436# 0.045851f
C20347 a_11823_42460# a_n1741_47186# 9.63e-19
C20348 a_6812_45938# a_2063_45854# 0.026385f
C20349 a_n2293_46098# a_3218_45724# 0.007233f
C20350 a_2202_46116# a_n2661_45546# 6.86e-21
C20351 a_1176_45822# a_n2293_45546# 2.19e-20
C20352 a_n1076_46494# a_n1099_45572# 3.72e-20
C20353 a_376_46348# a_380_45546# 0.011689f
C20354 a_805_46414# a_n863_45724# 8.12e-20
C20355 a_11415_45002# a_n443_42852# 1.47e-20
C20356 a_17715_44484# a_8049_45260# 0.03139f
C20357 a_12005_46116# a_12379_46436# 0.038694f
C20358 a_11189_46129# a_11315_46155# 0.005516f
C20359 a_10903_43370# a_12638_46436# 0.006548f
C20360 a_6945_45028# a_5066_45546# 0.018752f
C20361 a_9290_44172# a_11601_46155# 8.23e-19
C20362 a_9313_44734# a_21613_42308# 0.001498f
C20363 a_1414_42308# a_2903_42308# 1.7e-19
C20364 a_18326_43940# a_18504_43218# 2.4e-20
C20365 a_15781_43660# a_15743_43084# 0.050751f
C20366 a_16409_43396# a_16977_43638# 0.17072f
C20367 a_16243_43396# a_17499_43370# 0.043633f
C20368 a_16137_43396# a_17324_43396# 1.29e-20
C20369 a_19319_43548# a_19164_43230# 7.09e-19
C20370 a_n97_42460# a_12545_42858# 3.58e-19
C20371 a_16547_43609# a_16759_43396# 9.49e-19
C20372 a_8685_43396# a_5649_42852# 2.05e-20
C20373 a_10341_43396# a_17021_43396# 4.33e-19
C20374 a_21588_30879# SINGLE_ENDED 0.001491f
C20375 a_5807_45002# CLK 0.033646f
C20376 a_10922_42852# VDD 0.216186f
C20377 a_10951_45334# a_n2661_43370# 0.004229f
C20378 a_10907_45822# a_n2661_43922# 2.58e-19
C20379 a_16147_45260# a_17767_44458# 1.74e-19
C20380 a_1307_43914# a_5009_45028# 2.65e-20
C20381 a_20447_31679# a_19721_31679# 0.070259f
C20382 a_6171_45002# a_13490_45067# 3.54e-19
C20383 a_743_42282# a_n357_42282# 0.067793f
C20384 a_n4334_38528# a_n2312_38680# 6.16e-20
C20385 a_11323_42473# a_3090_45724# 4.17e-20
C20386 a_14635_42282# a_4185_45028# 9.41e-20
C20387 a_n4064_37984# SMPL_ON_P 7.33e-21
C20388 a_14495_45572# a_6755_46942# 2.1e-21
C20389 a_8746_45002# a_8270_45546# 0.017581f
C20390 a_17034_45572# a_n743_46660# 2.11e-19
C20391 a_2211_45572# a_3090_45724# 1.16e-19
C20392 a_20731_45938# a_20916_46384# 8.76e-21
C20393 a_2437_43646# a_13661_43548# 0.003998f
C20394 a_21513_45002# a_13747_46662# 0.02166f
C20395 a_n2661_45010# a_768_44030# 0.015059f
C20396 a_20719_45572# a_19321_45002# 1.72e-19
C20397 a_n967_45348# a_n881_46662# 6.86e-19
C20398 a_n659_45366# a_n1613_43370# 0.001198f
C20399 a_9482_43914# a_10227_46804# 0.032461f
C20400 a_7229_43940# a_4883_46098# 6.78e-21
C20401 a_5009_45028# a_n443_46116# 4.3e-20
C20402 a_5093_45028# a_4791_45118# 0.007375f
C20403 a_8137_45348# a_n1151_42308# 5.47e-21
C20404 a_17333_42852# a_18249_42858# 0.311255f
C20405 a_18083_42858# a_18817_42826# 0.0532f
C20406 a_3626_43646# a_15051_42282# 0.009723f
C20407 a_2982_43646# a_15764_42576# 3.1e-19
C20408 a_n97_42460# a_19332_42282# 2.35e-20
C20409 a_14401_32519# a_22775_42308# 3.78e-20
C20410 a_3935_42891# a_4149_42891# 0.005572f
C20411 a_7227_42852# a_7573_43172# 0.013377f
C20412 a_4185_45028# EN_OFFSET_CAL 4.56e-21
C20413 a_17531_42308# VDD 0.262303f
C20414 a_n237_47217# a_4883_46098# 0.181672f
C20415 a_n1920_47178# a_n2312_40392# 7.09e-19
C20416 a_n2109_47186# a_n2312_39304# 0.06316f
C20417 a_6575_47204# a_9313_45822# 0.017088f
C20418 a_6151_47436# a_13487_47204# 0.038134f
C20419 a_9067_47204# a_11031_47542# 6.46e-21
C20420 a_6851_47204# a_n1435_47204# 2.24e-19
C20421 a_4915_47217# a_11599_46634# 0.015066f
C20422 a_949_44458# a_n23_44458# 3.38e-20
C20423 a_n2661_44458# a_6109_44484# 0.004386f
C20424 a_375_42282# a_n1761_44111# 1.36e-19
C20425 a_n1352_44484# a_n1243_44484# 0.007416f
C20426 a_n1177_44458# a_n998_44484# 0.007399f
C20427 a_n452_44636# a_7_44811# 6.64e-19
C20428 a_11827_44484# a_n2661_42834# 0.046936f
C20429 a_12607_44458# a_15004_44636# 1.81e-20
C20430 a_5205_44484# a_7281_43914# 0.008497f
C20431 a_n913_45002# a_10405_44172# 2.38e-20
C20432 a_n1059_45260# a_10729_43914# 5.14e-23
C20433 a_13575_42558# a_13259_45724# 0.097619f
C20434 a_5755_42308# a_n357_42282# 4.82e-20
C20435 a_n2302_40160# a_n2956_38680# 6.16e-19
C20436 a_7174_31319# a_n1925_42282# 2.64e-20
C20437 a_14209_32519# VCM 0.007464f
C20438 a_20980_44850# a_12861_44030# 7.8e-21
C20439 a_2675_43914# a_584_46384# 7.8e-20
C20440 a_n3674_39768# SMPL_ON_P 0.03705f
C20441 a_n630_44306# a_n2497_47436# 3.9e-19
C20442 a_20766_44850# a_16327_47482# 0.17113f
C20443 a_11967_42832# a_18479_47436# 0.017885f
C20444 a_15861_45028# a_6945_45028# 5.7e-21
C20445 a_2711_45572# a_n2661_45546# 0.359276f
C20446 a_14495_45572# a_8049_45260# 0.004043f
C20447 a_11823_42460# a_10586_45546# 0.005505f
C20448 a_n967_45348# a_n2157_46122# 1.95e-20
C20449 a_10057_43914# a_2107_46812# 7.24e-20
C20450 a_16019_45002# a_13059_46348# 4.51e-21
C20451 a_9313_44734# a_12891_46348# 2.52e-21
C20452 a_413_45260# a_21076_30879# 0.141502f
C20453 a_n913_45002# a_n901_46420# 6.07e-19
C20454 a_n1059_45260# a_n1076_46494# 3.89e-20
C20455 a_n2661_44458# a_4646_46812# 0.05901f
C20456 a_19987_42826# a_7174_31319# 6.85e-20
C20457 a_21195_42852# a_13258_32519# 1.05e-19
C20458 a_n784_42308# a_1184_42692# 0.026118f
C20459 a_564_42282# a_n1630_35242# 0.156633f
C20460 a_196_42282# a_961_42354# 1.2e-21
C20461 a_22165_42308# a_19511_42282# 1.52e-19
C20462 a_n881_46662# a_7715_46873# 0.02091f
C20463 a_n1613_43370# a_7577_46660# 3.27e-20
C20464 a_4883_46098# a_8270_45546# 0.278829f
C20465 a_11599_46634# a_18834_46812# 0.012948f
C20466 a_15811_47375# a_16292_46812# 0.080078f
C20467 a_10227_46804# a_12816_46660# 0.253017f
C20468 a_16327_47482# a_14976_45028# 1.2e-20
C20469 a_6151_47436# a_14513_46634# 3.62e-20
C20470 a_12861_44030# a_19692_46634# 0.097215f
C20471 a_2952_47436# a_765_45546# 0.004287f
C20472 a_n1151_42308# a_14447_46660# 0.003689f
C20473 a_n2438_43548# a_2107_46812# 0.111283f
C20474 a_33_46660# a_383_46660# 0.20669f
C20475 a_n133_46660# a_948_46660# 0.102355f
C20476 a_n2661_46634# a_n2661_46098# 0.066513f
C20477 a_171_46873# a_1123_46634# 1.13e-20
C20478 a_n2312_38680# a_n935_46688# 7.7e-20
C20479 a_n743_46660# a_1983_46706# 0.001758f
C20480 a_1423_45028# a_9145_43396# 3.76e-21
C20481 a_5518_44484# a_5829_43940# 1.88e-20
C20482 a_14539_43914# a_14021_43940# 0.043922f
C20483 a_9313_44734# a_11750_44172# 2.81e-21
C20484 a_1307_43914# a_14205_43396# 1.03e-20
C20485 a_8696_44636# a_13635_43156# 2.2e-22
C20486 a_3422_30871# a_22959_44484# 2.88e-19
C20487 a_n2661_42834# a_6756_44260# 1.06e-19
C20488 a_22315_44484# a_17730_32519# 0.001043f
C20489 VDAC_Pi VDD 0.591846f
C20490 a_18184_42460# VDD 2.05053f
C20491 a_4181_44734# a_4185_45028# 5.69e-19
C20492 a_14112_44734# a_12741_44636# 7.78e-19
C20493 a_5289_44734# a_3483_46348# 5.06e-20
C20494 a_14401_32519# a_12549_44172# 0.004427f
C20495 a_1307_43914# a_2957_45546# 1.73e-20
C20496 a_17719_45144# a_8049_45260# 3.83e-20
C20497 a_626_44172# a_n357_42282# 0.551369f
C20498 a_501_45348# a_n755_45592# 5.21e-19
C20499 a_2809_45348# a_n863_45724# 1.93e-19
C20500 a_4640_45348# a_n2661_45546# 0.003021f
C20501 a_13159_45002# a_n443_42852# 1.23e-20
C20502 a_9838_44484# a_2324_44458# 4.19e-20
C20503 a_13076_44458# a_12594_46348# 4.02e-22
C20504 a_n1177_43370# a_n1613_43370# 0.325171f
C20505 a_2982_43646# a_13507_46334# 0.063751f
C20506 a_14358_43442# a_4915_47217# 3.86e-20
C20507 a_5742_30871# a_1177_38525# 1.05e-19
C20508 a_21613_42308# a_22397_42558# 0.001996f
C20509 a_21887_42336# a_22465_38105# 7.29e-21
C20510 a_7174_31319# a_n4315_30879# 6.67e-21
C20511 a_n784_42308# C0_P_btm 0.281635f
C20512 a_15559_46634# a_16388_46812# 2.85e-19
C20513 a_12991_46634# a_765_45546# 1.31e-19
C20514 a_n881_46662# a_5210_46482# 0.002203f
C20515 a_n743_46660# a_14275_46494# 0.006268f
C20516 a_13747_46662# a_10809_44734# 0.045104f
C20517 a_19321_45002# a_6945_45028# 0.042647f
C20518 a_2107_46812# a_11133_46155# 7.92e-20
C20519 a_n1613_43370# a_5431_46482# 6.82e-22
C20520 a_5342_30871# a_n4064_37440# 0.028573f
C20521 a_4883_46098# a_12638_46436# 0.009375f
C20522 a_13507_46334# a_14371_46494# 0.001286f
C20523 a_16327_47482# a_18051_46116# 2.01e-20
C20524 a_17591_47464# a_16375_45002# 4.87e-19
C20525 a_n443_46116# a_2957_45546# 0.020365f
C20526 a_2063_45854# a_1609_45822# 0.035351f
C20527 a_17973_43940# a_18533_43940# 5.23e-19
C20528 a_17061_44734# a_16409_43396# 1.3e-20
C20529 a_9313_44734# a_4361_42308# 0.082952f
C20530 a_5883_43914# a_9127_43156# 3.96e-19
C20531 a_20193_45348# a_21195_42852# 1.43e-20
C20532 a_3905_42865# a_3626_43646# 0.036343f
C20533 a_18451_43940# a_18797_44260# 0.013377f
C20534 a_n1059_45260# a_5932_42308# 8.52e-19
C20535 a_n913_45002# a_6171_42473# 0.034189f
C20536 a_n2017_45002# a_6481_42558# 0.001353f
C20537 a_10193_42453# a_18799_45938# 3.31e-21
C20538 a_6194_45824# a_3357_43084# 0.004141f
C20539 a_11301_43218# a_10227_46804# 1.79e-19
C20540 a_5745_43940# a_5937_45572# 4.36e-20
C20541 a_11967_42832# a_n443_42852# 0.00555f
C20542 a_10765_43646# a_3090_45724# 6.96e-19
C20543 a_8952_43230# a_n2293_46634# 1.4e-20
C20544 a_14579_43548# a_15227_44166# 7.96e-19
C20545 a_5534_30871# a_5807_45002# 3.81e-20
C20546 a_15037_43940# a_3483_46348# 0.007725f
C20547 a_7754_40130# CAL_P 0.04831f
C20548 a_n3420_37984# EN_VIN_BSTR_P 0.031779f
C20549 a_12741_44636# VDD 0.988199f
C20550 a_7174_31319# a_n3420_37440# 0.002179f
C20551 a_4958_30871# a_11206_38545# 1.83e-20
C20552 a_9823_46155# a_2324_44458# 1.64e-20
C20553 a_10903_43370# a_13759_46122# 8.61e-19
C20554 a_12005_46116# a_13351_46090# 1.07e-19
C20555 a_1208_46090# a_1337_46436# 0.010132f
C20556 a_17339_46660# a_18243_46436# 0.001467f
C20557 a_17829_46910# a_13259_45724# 8.1e-20
C20558 a_22365_46825# a_8049_45260# 0.001257f
C20559 a_20835_44721# a_20753_42852# 5.18e-21
C20560 a_20974_43370# a_4361_42308# 0.122936f
C20561 a_n2293_43922# a_5379_42460# 0.4571f
C20562 a_n356_44636# a_11323_42473# 1.17e-19
C20563 a_17538_32519# a_13467_32519# 0.051209f
C20564 a_21381_43940# a_13678_32519# 5.1e-21
C20565 a_17737_43940# a_17701_42308# 1.13e-19
C20566 a_14401_32519# a_21855_43396# 0.00125f
C20567 a_n97_42460# a_17021_43396# 4.28e-19
C20568 a_11599_46634# DATA[5] 9.31e-19
C20569 a_17591_47464# RST_Z 2.7e-19
C20570 a_14311_47204# CLK 1.56e-19
C20571 a_16115_45572# a_11691_44458# 1.01e-20
C20572 a_15861_45028# a_11827_44484# 1.34e-19
C20573 a_10193_42453# a_16112_44458# 1.55e-19
C20574 a_11962_45724# a_8975_43940# 3.26e-21
C20575 a_16147_45260# a_16405_45348# 0.001516f
C20576 a_n1059_45260# a_1423_45028# 8.02e-22
C20577 a_2437_43646# a_2448_45028# 4.11e-19
C20578 a_6431_45366# a_5205_44484# 0.018787f
C20579 a_6171_45002# a_7276_45260# 0.00899f
C20580 a_3232_43370# a_7229_43940# 0.180766f
C20581 a_5111_44636# a_8191_45002# 1.43e-20
C20582 a_15279_43071# a_3483_46348# 5.23e-21
C20583 a_14543_43071# a_4185_45028# 9.15e-22
C20584 a_19511_42282# a_13661_43548# 4.91e-21
C20585 a_648_43396# a_n443_42852# 0.002995f
C20586 a_10083_42826# a_8953_45546# 8.07e-20
C20587 a_10835_43094# a_8199_44636# 4.6e-21
C20588 a_8037_42858# a_9290_44172# 2.48e-20
C20589 a_n3565_39304# a_n2312_39304# 0.104981f
C20590 a_17730_32519# VCM 0.068103f
C20591 a_19237_31679# VREF 0.046045f
C20592 a_2437_43646# a_14955_47212# 0.009063f
C20593 a_20623_45572# a_10227_46804# 4e-20
C20594 a_19365_45572# a_16327_47482# 4.87e-19
C20595 a_3357_43084# a_12861_44030# 3.68e-19
C20596 a_413_45260# a_3381_47502# 0.001239f
C20597 a_3065_45002# a_2063_45854# 4.37e-20
C20598 a_3232_43370# a_n237_47217# 7.83e-20
C20599 a_3429_45260# a_584_46384# 4.23e-21
C20600 a_327_44734# a_n1151_42308# 8.48e-19
C20601 a_18479_45785# a_11453_44696# 0.003588f
C20602 a_20273_45572# a_18479_47436# 0.028755f
C20603 a_8696_44636# a_n1613_43370# 5.83e-19
C20604 a_16680_45572# a_n881_46662# 0.051767f
C20605 a_13249_42308# a_n2293_46634# 0.027384f
C20606 a_11823_42460# a_n743_46660# 5.08e-19
C20607 a_5907_45546# a_4646_46812# 3.34e-21
C20608 a_n2661_45546# a_n1079_45724# 0.008911f
C20609 a_n2472_45546# a_n2293_45546# 0.171197f
C20610 a_13259_45724# a_n443_42852# 0.022577f
C20611 a_19478_44306# a_19647_42308# 2.55e-20
C20612 a_1568_43370# a_1755_42282# 7.17e-19
C20613 a_5649_42852# a_17333_42852# 1.49e-20
C20614 a_4361_42308# a_18599_43230# 9.24e-21
C20615 a_19862_44208# a_19511_42282# 1.12e-19
C20616 a_n1557_42282# a_n1630_35242# 0.865968f
C20617 a_14579_43548# a_14635_42282# 0.124652f
C20618 a_3080_42308# a_1184_42692# 1.44e-20
C20619 a_n4318_39768# a_n4064_39072# 2.48e-21
C20620 a_1756_43548# a_1606_42308# 3.46e-19
C20621 VDAC_Pi a_8912_37509# 1.57e-19
C20622 a_7754_38470# a_8530_39574# 0.143675f
C20623 a_7754_40130# CAL_N 0.050321f
C20624 a_7754_39964# VDAC_P 0.003276f
C20625 a_2903_42308# VDD 0.22017f
C20626 a_n452_47436# a_n971_45724# 0.330438f
C20627 a_n1741_47186# a_n785_47204# 0.026399f
C20628 a_n2109_47186# a_1209_47178# 0.226908f
C20629 a_n815_47178# a_n746_45260# 0.001861f
C20630 a_13777_45326# a_13857_44734# 8.93e-19
C20631 a_9482_43914# a_14815_43914# 0.024524f
C20632 a_2711_45572# a_19478_44056# 4.36e-19
C20633 a_n2017_45002# a_3422_30871# 2.49e-20
C20634 a_6481_42558# a_526_44458# 0.001415f
C20635 a_5932_42308# a_n1925_42282# 0.004062f
C20636 a_19511_42282# a_4185_45028# 9.41e-20
C20637 a_8791_45572# a_3483_46348# 5.57e-19
C20638 a_18175_45572# a_18280_46660# 1.14e-20
C20639 a_11691_44458# a_5807_45002# 0.117249f
C20640 a_11827_44484# a_19321_45002# 0.037739f
C20641 a_22959_45036# a_13747_46662# 4.74e-20
C20642 a_20205_45028# a_12549_44172# 7.43e-20
C20643 a_16321_45348# a_n743_46660# 7.66e-19
C20644 a_19113_45348# a_13661_43548# 0.003675f
C20645 a_3232_43370# a_8270_45546# 0.020859f
C20646 a_3357_43084# a_14180_46812# 1.32e-20
C20647 a_413_45260# a_15009_46634# 1.08e-20
C20648 a_7705_45326# a_7832_46660# 7.57e-21
C20649 a_n913_45002# a_19692_46634# 2.2e-20
C20650 a_11652_45724# a_10903_43370# 0.010404f
C20651 a_11823_42460# a_11189_46129# 1.55e-19
C20652 a_11322_45546# a_12594_46348# 1.17e-19
C20653 a_n1177_44458# a_n1613_43370# 0.332209f
C20654 a_13076_44458# a_12465_44636# 0.01224f
C20655 a_10341_42308# a_5742_30871# 0.031841f
C20656 a_13887_32519# a_21613_42308# 0.00157f
C20657 a_13467_32519# a_22465_38105# 0.076379f
C20658 a_n2293_42282# a_3581_42558# 0.001341f
C20659 a_3080_42308# C0_P_btm 0.018211f
C20660 a_12891_46348# a_13569_47204# 9.78e-20
C20661 a_n881_46662# a_13747_46662# 0.550574f
C20662 a_n310_47243# a_n2661_46634# 2.6e-19
C20663 a_n2312_39304# a_n1925_46634# 0.071018f
C20664 a_6575_47204# a_6540_46812# 1.87e-19
C20665 a_4915_47217# a_7411_46660# 4.06e-20
C20666 a_n1435_47204# a_4651_46660# 5.31e-20
C20667 a_2063_45854# a_10249_46116# 0.078073f
C20668 a_n1151_42308# a_10150_46912# 8.58e-20
C20669 a_18494_42460# a_15493_43940# 0.02195f
C20670 a_21101_45002# a_21115_43940# 3.47e-20
C20671 a_n356_44636# a_644_44056# 2.5e-19
C20672 a_11827_44484# a_20623_43914# 0.004538f
C20673 a_n2661_44458# a_10405_44172# 1.99e-20
C20674 a_11691_44458# a_19478_44306# 3.14e-20
C20675 a_2711_45572# a_17701_42308# 5.54e-20
C20676 a_7499_43078# a_8605_42826# 0.026478f
C20677 a_20193_45348# a_15493_43396# 3.33e-21
C20678 C9_N_btm VDD 0.345685f
C20679 a_13556_45296# VDD 0.569056f
C20680 a_n1630_35242# a_n83_35174# 7.97e-19
C20681 a_1209_43370# a_584_46384# 0.02923f
C20682 a_n1557_42282# a_n971_45724# 0.06901f
C20683 a_14021_43940# a_11453_44696# 8.33e-20
C20684 a_n2661_43370# a_2324_44458# 0.082794f
C20685 a_n2472_45002# a_n2661_45546# 0.004199f
C20686 a_n2840_45002# a_n2956_38216# 0.01122f
C20687 a_1423_45028# a_n1925_42282# 0.021671f
C20688 a_11963_45334# a_8049_45260# 1.58e-20
C20689 a_15682_43940# a_12549_44172# 0.058263f
C20690 a_n3674_39768# a_n2438_43548# 0.007137f
C20691 a_n1177_44458# a_n2293_46098# 1.38e-20
C20692 a_n2267_44484# a_n1991_46122# 7.99e-21
C20693 a_n2661_44458# a_n901_46420# 9.89e-21
C20694 a_3160_47472# VDD 0.256092f
C20695 a_n4318_38216# a_n4064_38528# 0.057645f
C20696 a_n3674_38216# a_n3420_38528# 0.152701f
C20697 a_n4318_37592# a_n3565_38502# 3.09e-20
C20698 a_5932_42308# a_n4315_30879# 6.05e-21
C20699 a_n1613_43370# a_4704_46090# 4.05e-20
C20700 a_12465_44636# a_12594_46348# 9.31e-21
C20701 a_n1435_47204# a_n1379_46482# 7.65e-21
C20702 a_4883_46098# a_13759_46122# 0.044004f
C20703 a_13507_46334# a_14493_46090# 0.001974f
C20704 a_16327_47482# a_19900_46494# 0.216811f
C20705 a_10227_46804# a_18819_46122# 2.52e-20
C20706 a_11599_46634# a_10809_44734# 0.06157f
C20707 a_15811_47375# a_6945_45028# 0.037131f
C20708 a_18597_46090# a_17583_46090# 4.74e-20
C20709 a_4791_45118# a_5431_46482# 0.001192f
C20710 a_n881_46662# a_4419_46090# 0.045203f
C20711 a_22612_30879# a_12741_44636# 1.68e-20
C20712 a_n2661_46634# a_11415_45002# 0.494836f
C20713 a_768_44030# a_1138_42852# 0.021091f
C20714 a_20916_46384# a_21076_30879# 9.97e-20
C20715 a_21588_30879# a_22959_46660# 0.001846f
C20716 a_n2661_46098# a_765_45546# 0.0407f
C20717 a_6755_46942# a_11901_46660# 0.587021f
C20718 a_10249_46116# a_12469_46902# 8.44e-20
C20719 a_n2661_43922# a_7112_43396# 3.6e-21
C20720 a_n2661_42834# a_8147_43396# 1.43e-20
C20721 a_11823_42460# a_15486_42560# 0.003207f
C20722 a_19721_31679# a_13467_32519# 0.051394f
C20723 a_2998_44172# a_3737_43940# 0.003753f
C20724 a_13249_42308# a_13249_42558# 0.003175f
C20725 a_10193_42453# a_11633_42308# 0.003739f
C20726 a_5891_43370# a_8229_43396# 1.73e-20
C20727 a_16112_44458# a_16137_43396# 2.27e-19
C20728 a_3422_30871# a_21845_43940# 4.36e-19
C20729 en_comp a_13291_42460# 4.34e-21
C20730 a_n1059_45260# a_17141_43172# 0.001223f
C20731 a_n2017_45002# a_18504_43218# 0.016191f
C20732 a_20362_44736# VDD 0.275577f
C20733 a_10193_42453# a_11962_45724# 0.044438f
C20734 a_10490_45724# a_11525_45546# 0.06936f
C20735 a_2711_45572# a_11136_45572# 0.002612f
C20736 a_8746_45002# a_11652_45724# 2.41e-21
C20737 a_4190_30871# a_5807_45002# 8.86e-22
C20738 a_21259_43561# a_13661_43548# 2.35e-20
C20739 a_n356_44636# a_n23_45546# 1.17e-20
C20740 a_2998_44172# a_2324_44458# 2.03e-19
C20741 a_n1991_42858# a_n1613_43370# 0.029351f
C20742 a_10796_42968# a_10227_46804# 0.024053f
C20743 a_8483_43230# a_n971_45724# 2.48e-19
C20744 a_413_45260# SINGLE_ENDED 0.037852f
C20745 a_13607_46688# VDD 0.209568f
C20746 a_n4064_39072# C1_P_btm 9.59e-21
C20747 a_5932_42308# a_n3420_37440# 5.13e-19
C20748 a_472_46348# a_167_45260# 0.001848f
C20749 a_1208_46090# a_1823_45246# 0.006027f
C20750 a_1176_45822# a_1138_42852# 0.41217f
C20751 a_1799_45572# a_n443_42852# 4.66e-20
C20752 a_11901_46660# a_8049_45260# 8.89e-20
C20753 a_6755_46942# a_15194_46482# 0.002244f
C20754 a_n2293_46098# a_4704_46090# 2.86e-20
C20755 a_11415_45002# a_8199_44636# 4.09e-20
C20756 a_19123_46287# a_17583_46090# 1.17e-20
C20757 a_765_45546# a_17957_46116# 0.133328f
C20758 a_18285_46348# a_17715_44484# 2.97e-20
C20759 a_13059_46348# a_6945_45028# 3.04e-19
C20760 a_17829_46910# a_18189_46348# 4.65e-19
C20761 a_5663_43940# a_5755_42852# 0.001147f
C20762 a_19478_44306# a_4190_30871# 2.22e-20
C20763 a_17737_43940# a_4361_42308# 1.14e-20
C20764 a_4699_43561# a_2982_43646# 1.91e-20
C20765 a_n97_42460# a_7287_43370# 0.004081f
C20766 a_14021_43940# a_17324_43396# 0.009103f
C20767 a_4093_43548# a_3626_43646# 0.011002f
C20768 a_19862_44208# a_21259_43561# 8.37e-19
C20769 a_n2661_42282# a_n1641_43230# 1.25e-20
C20770 a_20512_43084# a_18083_42858# 1.67e-21
C20771 a_3422_30871# a_19164_43230# 5.64e-20
C20772 a_458_43396# a_548_43396# 0.008441f
C20773 a_15493_43396# a_20301_43646# 2.14e-19
C20774 a_n699_43396# a_2903_42308# 1.29e-19
C20775 a_5883_43914# a_1755_42282# 2.89e-20
C20776 a_6293_42852# VDD 0.401011f
C20777 a_16855_45546# a_16751_45260# 4.68e-19
C20778 a_15861_45028# a_15595_45028# 0.072432f
C20779 a_8696_44636# a_16019_45002# 2.28e-19
C20780 a_3357_43084# a_n913_45002# 2.04e-19
C20781 a_20107_42308# a_12861_44030# 1.45e-21
C20782 a_n3420_38528# w_1575_34946# 5.84e-19
C20783 a_18907_42674# a_16327_47482# 0.001573f
C20784 a_4958_30871# a_10227_46804# 0.036177f
C20785 a_15681_43442# a_2324_44458# 0.006403f
C20786 a_4181_43396# a_n1925_42282# 1.15e-19
C20787 a_4156_43218# a_3090_45724# 2.05e-21
C20788 a_20922_43172# a_19692_46634# 5.29e-20
C20789 a_21259_43561# a_4185_45028# 4.43e-21
C20790 a_16375_45002# VDD 1.14948f
C20791 a_2711_45572# a_12891_46348# 0.027614f
C20792 a_6598_45938# a_n881_46662# 0.031336f
C20793 a_7227_45028# a_n1613_43370# 8.73e-21
C20794 a_11322_45546# a_12465_44636# 5.04e-19
C20795 a_10180_45724# a_11453_44696# 2.98e-19
C20796 a_11652_45724# a_4883_46098# 1.56e-19
C20797 a_8696_44636# a_4791_45118# 0.097007f
C20798 a_14579_43548# a_14543_43071# 0.032593f
C20799 a_21855_43396# a_22223_43396# 7.52e-19
C20800 a_13678_32519# a_5649_42852# 0.506367f
C20801 a_13467_32519# a_22591_43396# 4.5e-22
C20802 a_14205_43396# a_13635_43156# 0.002342f
C20803 a_743_42282# a_20749_43396# 0.09037f
C20804 a_4905_42826# a_4649_42852# 0.006342f
C20805 a_4361_42308# a_13887_32519# 2.22e-19
C20806 VDAC_N C10_N_btm 0.883474p
C20807 a_11554_42852# VDD 0.078978f
C20808 a_n143_45144# a_n23_44458# 0.001215f
C20809 a_n37_45144# a_n356_44636# 4.09e-19
C20810 a_8953_45002# a_10157_44484# 0.002321f
C20811 a_6171_45002# a_13720_44458# 3.19e-20
C20812 a_20447_31679# a_9313_44734# 1.21e-20
C20813 a_n967_45348# a_n998_44484# 0.001023f
C20814 a_4921_42308# a_4185_45028# 0.059648f
C20815 a_10518_42984# a_n443_42852# 1.45e-19
C20816 a_15279_43071# a_n357_42282# 0.007143f
C20817 a_17538_32519# VCM 0.0424f
C20818 a_22612_30879# C9_N_btm 0.003123f
C20819 a_21588_30879# C10_N_btm 0.002325f
C20820 a_4223_44672# a_n1151_42308# 1.31e-20
C20821 a_6298_44484# a_2063_45854# 5.31e-21
C20822 RST_Z VDD 4.72146f
C20823 a_21005_45260# a_16327_47482# 0.004367f
C20824 a_3357_43084# a_5894_47026# 1.88e-19
C20825 a_413_45260# a_2959_46660# 0.011261f
C20826 a_n1059_45260# a_4646_46812# 0.001886f
C20827 a_7705_45326# a_n743_46660# 4.03e-20
C20828 a_2274_45254# a_2443_46660# 9.71e-22
C20829 a_2437_43646# a_5257_43370# 7.48e-20
C20830 a_16223_45938# a_3090_45724# 0.002393f
C20831 a_16751_45260# a_13661_43548# 1.24e-19
C20832 a_13159_45002# a_n2661_46634# 0.062031f
C20833 a_1307_43914# a_13747_46662# 5.92e-20
C20834 a_16115_45572# a_15227_44166# 2.6e-21
C20835 a_1176_45572# a_1138_42852# 7.3e-19
C20836 a_1260_45572# a_1176_45822# 0.00411f
C20837 a_15781_43660# a_16104_42674# 4.99e-20
C20838 a_5649_42852# a_6123_31319# 0.062309f
C20839 a_4361_42308# a_8515_42308# 0.007572f
C20840 a_743_42282# a_8685_42308# 0.039566f
C20841 a_17595_43084# a_17665_42852# 0.011552f
C20842 a_3080_42308# comp_n 2.82e-19
C20843 a_n2860_38778# VDD 0.004252f
C20844 a_4915_47217# a_13661_43548# 3.51e-19
C20845 a_9313_45822# a_12891_46348# 2.26e-20
C20846 a_11459_47204# a_11309_47204# 0.183357f
C20847 a_11599_46634# a_n881_46662# 0.100714f
C20848 a_n785_47204# a_n743_46660# 7.46e-20
C20849 a_n1741_47186# a_2107_46812# 2.24e-19
C20850 a_n746_45260# a_171_46873# 0.120194f
C20851 a_n23_47502# a_n2438_43548# 3.57e-20
C20852 a_n237_47217# a_n133_46660# 6.22e-19
C20853 a_1209_47178# a_n1925_46634# 3.96e-20
C20854 a_n971_45724# a_33_46660# 5.37e-19
C20855 a_2553_47502# a_n2661_46634# 3.46e-20
C20856 a_4883_46098# a_22731_47423# 9.43e-21
C20857 a_13507_46334# a_11453_44696# 0.060476f
C20858 a_21811_47423# a_22223_47212# 0.031065f
C20859 a_11967_42832# CAL_N 0.001103f
C20860 a_5891_43370# a_9313_44734# 0.028253f
C20861 a_8696_44636# a_8791_43396# 3.5e-20
C20862 a_14537_43396# a_11341_43940# 0.032289f
C20863 a_10193_42453# a_17499_43370# 0.009503f
C20864 a_n2293_42834# a_3499_42826# 0.029158f
C20865 a_2711_45572# a_4361_42308# 0.031943f
C20866 a_11823_42460# a_13837_43396# 0.001813f
C20867 a_13720_44458# a_14673_44172# 2.95e-20
C20868 a_9482_43914# a_9248_44260# 5.36e-21
C20869 a_13258_32519# a_n357_42282# 0.022774f
C20870 a_21363_45546# VDD 0.36538f
C20871 a_1423_45028# a_2698_46116# 6.57e-22
C20872 a_2304_45348# a_167_45260# 6.8e-19
C20873 a_5009_45028# a_n2293_46098# 0.009429f
C20874 a_2903_45348# a_1823_45246# 1.47e-19
C20875 a_11827_44484# a_13059_46348# 0.495367f
C20876 a_18911_45144# a_17339_46660# 1.25e-21
C20877 a_18579_44172# a_13747_46662# 1.11e-20
C20878 a_8975_43940# a_8270_45546# 0.207334f
C20879 a_20512_43084# a_12549_44172# 0.002813f
C20880 a_949_44458# a_3090_45724# 3.71e-22
C20881 a_18681_44484# a_13661_43548# 6.47e-19
C20882 a_n2810_45028# a_n2956_39304# 0.042912f
C20883 a_9482_43914# a_8016_46348# 0.293982f
C20884 a_n1331_43914# a_n1613_43370# 0.16678f
C20885 a_6171_45002# a_13351_46090# 1.13e-20
C20886 a_8953_45002# a_10355_46116# 4.75e-20
C20887 a_413_45260# a_19335_46494# 1.78e-21
C20888 a_4574_45260# a_2324_44458# 9.08e-20
C20889 a_10555_44260# a_2063_45854# 0.001312f
C20890 a_3318_42354# a_5742_30871# 1.46e-20
C20891 a_6761_42308# a_8515_42308# 1.96e-20
C20892 a_6123_31319# a_7963_42308# 0.192155f
C20893 a_7227_42308# a_5934_30871# 5.66e-20
C20894 a_n443_46116# a_4419_46090# 0.20069f
C20895 a_5807_45002# a_15227_44166# 0.042586f
C20896 a_13661_43548# a_18834_46812# 0.1407f
C20897 a_4817_46660# a_5072_46660# 0.06121f
C20898 a_5167_46660# a_5732_46660# 7.99e-20
C20899 a_4955_46873# a_5275_47026# 7.88e-19
C20900 a_n2661_46634# a_12251_46660# 0.001121f
C20901 a_12891_46348# a_12513_46660# 3.56e-19
C20902 a_11453_44696# a_20623_46660# 0.029618f
C20903 a_18479_47436# a_20202_43084# 0.040227f
C20904 a_13507_46334# a_17639_46660# 0.005147f
C20905 a_n1435_47204# a_n1076_46494# 2.92e-21
C20906 a_n2497_47436# a_2324_44458# 0.796031f
C20907 a_4791_45118# a_4704_46090# 0.001482f
C20908 a_4700_47436# a_5068_46348# 1.09e-20
C20909 a_n1151_42308# a_6419_46155# 0.028969f
C20910 a_2063_45854# a_5937_45572# 0.012248f
C20911 a_n356_44636# a_104_43370# 0.001131f
C20912 a_n23_44458# a_n97_42460# 4.48e-19
C20913 a_20835_44721# a_11341_43940# 6.34e-20
C20914 a_20766_44850# a_21115_43940# 4.08e-19
C20915 a_20640_44752# a_15493_43940# 7.7e-20
C20916 a_18579_44172# a_20269_44172# 7.35e-20
C20917 a_19279_43940# a_20935_43940# 2.95e-19
C20918 a_4223_44672# a_6197_43396# 1.94e-19
C20919 a_11691_44458# a_13667_43396# 3.82e-21
C20920 a_1414_42308# a_2253_44260# 0.001444f
C20921 a_6453_43914# a_7542_44172# 2.4e-20
C20922 a_n2661_42834# a_10555_43940# 8.1e-20
C20923 a_5111_44636# a_7765_42852# 3.95e-20
C20924 a_3232_43370# a_5755_42852# 5.23e-21
C20925 a_n913_45002# a_5342_30871# 0.122483f
C20926 a_n1059_45260# a_15567_42826# 0.048229f
C20927 a_n2017_45002# a_16414_43172# 2.51e-19
C20928 a_n1190_44850# VDD 5.02e-19
C20929 a_n4315_30879# VREF 1.73216f
C20930 a_n4064_40160# VIN_P 0.06337f
C20931 a_n3565_39304# C10_P_btm 2.44e-19
C20932 a_n4209_39304# C8_P_btm 9.97e-19
C20933 CAL_N a_13259_45724# 0.005414f
C20934 a_743_42282# a_12861_44030# 6.92e-20
C20935 a_16855_43396# a_16327_47482# 1.79e-19
C20936 a_15125_43396# a_10227_46804# 1.54e-19
C20937 a_10617_44484# a_10809_44734# 0.014699f
C20938 a_20193_45348# a_n357_42282# 0.006712f
C20939 a_7640_43914# a_526_44458# 1.26e-20
C20940 a_11341_43940# a_3090_45724# 0.041393f
C20941 a_8685_43396# a_768_44030# 1.24e-19
C20942 a_n4209_39304# a_n4334_38528# 6.38e-20
C20943 a_n4334_39392# a_n4209_38502# 6.38e-20
C20944 a_n4209_39590# a_n3565_38216# 0.03183f
C20945 a_n3565_39590# a_n4209_38216# 0.0313f
C20946 a_n3420_39072# a_n2860_39072# 0.003211f
C20947 a_2609_46660# VDD 0.312974f
C20948 a_5742_30871# C10_N_btm 0.00237f
C20949 a_4651_46660# a_526_44458# 6.28e-21
C20950 a_2107_46812# a_10586_45546# 1.85e-19
C20951 a_n2661_46634# a_13259_45724# 0.009129f
C20952 a_13747_46662# a_19443_46116# 1.58e-20
C20953 a_19321_45002# a_20009_46494# 1.68e-19
C20954 a_n881_46662# a_1848_45724# 8.39e-20
C20955 a_7577_46660# a_6945_45028# 0.001401f
C20956 COMP_P a_2113_38308# 1.33e-19
C20957 a_19123_46287# a_20885_46660# 5.98e-21
C20958 a_10405_44172# a_9145_43396# 1.63e-19
C20959 a_13483_43940# a_8685_43396# 2.97e-20
C20960 a_20512_43084# a_21855_43396# 0.013929f
C20961 a_n2293_43922# a_12089_42308# 0.183316f
C20962 a_9313_44734# a_17595_43084# 0.006038f
C20963 a_n2293_42834# a_3318_42354# 4.09e-21
C20964 a_3422_30871# a_14209_32519# 0.031148f
C20965 a_21205_44306# a_21381_43940# 8.17e-20
C20966 a_n913_45002# a_20107_42308# 3.57e-19
C20967 a_n2017_45002# a_7174_31319# 2.34e-19
C20968 a_7499_43940# VDD 0.193884f
C20969 a_5263_45724# a_1423_45028# 5.02e-21
C20970 a_18341_45572# a_18596_45572# 0.056391f
C20971 a_18909_45814# a_19256_45572# 0.051162f
C20972 a_11652_45724# a_3232_43370# 0.009948f
C20973 a_11525_45546# a_6171_45002# 9.43e-19
C20974 a_13291_42460# a_13661_43548# 7.75e-21
C20975 a_17364_32525# a_19692_46634# 0.001936f
C20976 a_8333_44056# a_n755_45592# 1.1e-19
C20977 a_1568_43370# a_2324_44458# 0.001169f
C20978 a_n1329_42308# a_n2312_39304# 8.42e-20
C20979 a_n961_42308# a_n2312_40392# 2.36e-20
C20980 a_n3565_37414# VCM 0.03748f
C20981 a_8912_37509# RST_Z 0.082942f
C20982 a_n3420_37440# VREF 9.37e-19
C20983 a_n4064_37440# VIN_P 0.078489f
C20984 VDAC_P C2_P_btm 3.46245f
C20985 a_19721_31679# VCM 0.03544f
C20986 a_18985_46122# VDD 0.253642f
C20987 a_6194_45824# a_6151_47436# 0.227219f
C20988 a_12427_45724# a_n1741_47186# 1.48e-19
C20989 a_7227_45028# a_4791_45118# 0.288276f
C20990 a_n2293_46098# a_2957_45546# 0.00827f
C20991 a_472_46348# a_n863_45724# 1.63e-20
C20992 a_1823_45246# a_n2661_45546# 0.181403f
C20993 a_n901_46420# a_n1099_45572# 0.002063f
C20994 a_17583_46090# a_8049_45260# 5.45e-20
C20995 a_12005_46116# a_12005_46436# 0.009374f
C20996 a_10903_43370# a_12379_46436# 2.66e-19
C20997 a_9290_44172# a_11315_46155# 0.001284f
C20998 a_16243_43396# a_16759_43396# 0.106647f
C20999 a_15681_43442# a_15743_43084# 0.001131f
C21000 a_16137_43396# a_17499_43370# 1.55e-19
C21001 a_19319_43548# a_19339_43156# 0.006943f
C21002 a_n97_42460# a_12089_42308# 4.02e-19
C21003 a_9313_44734# a_21887_42336# 0.001765f
C21004 a_16547_43609# a_16977_43638# 6.72e-20
C21005 a_2982_43646# a_1847_42826# 4.13e-21
C21006 a_10341_43396# a_16855_43396# 8.56e-19
C21007 a_20916_46384# SINGLE_ENDED 0.020511f
C21008 a_16131_47204# CLK 3.58e-19
C21009 a_22612_30879# RST_Z 0.058603f
C21010 a_10991_42826# VDD 0.201891f
C21011 a_10775_45002# a_n2661_43370# 0.009126f
C21012 a_10907_45822# a_n2661_42834# 7.86e-20
C21013 a_16147_45260# a_16979_44734# 6.23e-20
C21014 a_11823_42460# a_12829_44484# 2.31e-19
C21015 a_22959_45572# a_19721_31679# 0.005929f
C21016 a_20447_31679# a_18114_32519# 0.051474f
C21017 a_3357_43084# a_n2661_44458# 0.027126f
C21018 a_17364_32525# a_20692_30879# 0.054134f
C21019 a_n4209_38502# a_n2312_38680# 0.095213f
C21020 a_10723_42308# a_3090_45724# 4.98e-22
C21021 a_13291_42460# a_4185_45028# 6.95e-20
C21022 a_22959_43948# RST_Z 0.001362f
C21023 a_8697_45822# a_8492_46660# 2.64e-20
C21024 a_16789_45572# a_n743_46660# 1.94e-19
C21025 a_10193_42453# a_8270_45546# 3e-20
C21026 a_1990_45572# a_3090_45724# 2.91e-20
C21027 a_2437_43646# a_5807_45002# 0.004842f
C21028 a_19610_45572# a_19594_46812# 5.07e-20
C21029 a_n967_45348# a_n1613_43370# 0.213625f
C21030 a_14537_43396# a_16327_47482# 3.85e-20
C21031 a_1307_43914# a_11599_46634# 3.42e-19
C21032 a_13348_45260# a_10227_46804# 6.18e-19
C21033 a_n2293_42834# a_n1151_42308# 0.051075f
C21034 a_5009_45028# a_4791_45118# 0.007533f
C21035 a_2809_45028# a_n443_46116# 5.61e-19
C21036 a_18083_42858# a_18249_42858# 0.699797f
C21037 a_2982_43646# a_15486_42560# 9.69e-20
C21038 a_3626_43646# a_14113_42308# 0.077829f
C21039 a_20974_43370# a_21887_42336# 8.61e-21
C21040 a_3935_42891# a_3863_42891# 6.64e-19
C21041 a_7227_42852# a_7309_43172# 0.003935f
C21042 a_3483_46348# CLK 0.408122f
C21043 a_17303_42282# VDD 0.379254f
C21044 a_n2288_47178# a_n2312_39304# 0.01565f
C21045 a_n2109_47186# a_n2312_40392# 0.005539f
C21046 a_7903_47542# a_9313_45822# 3.57e-20
C21047 a_6151_47436# a_12861_44030# 0.39397f
C21048 a_9067_47204# a_9863_47436# 0.007473f
C21049 a_6491_46660# a_n1435_47204# 7.35e-19
C21050 a_12883_44458# a_13076_44458# 0.142643f
C21051 a_949_44458# a_n356_44636# 0.009584f
C21052 a_12607_44458# a_13720_44458# 0.122704f
C21053 a_375_42282# a_n2065_43946# 2.58e-21
C21054 a_7499_43078# a_3626_43646# 0.002457f
C21055 a_n452_44636# a_n310_44811# 0.005572f
C21056 a_11827_44484# a_11649_44734# 5.76e-21
C21057 a_n2661_44458# a_5826_44734# 6.36e-19
C21058 a_n1059_45260# a_10405_44172# 2.46e-20
C21059 a_5205_44484# a_6453_43914# 7.72e-19
C21060 a_413_45260# a_3499_42826# 4.69e-19
C21061 a_7229_43940# a_5495_43940# 6.48e-21
C21062 a_7174_31319# a_526_44458# 4.88e-21
C21063 a_n4064_40160# a_n2956_38680# 6.27e-19
C21064 a_n2302_40160# a_n2956_39304# 4.04e-19
C21065 a_13070_42354# a_13259_45724# 6.28e-20
C21066 a_14209_32519# VREF_GND 0.034351f
C21067 a_17364_32525# VIN_N 0.039314f
C21068 a_20835_44721# a_16327_47482# 0.157393f
C21069 a_19789_44512# a_12861_44030# 2.27e-19
C21070 a_895_43940# a_584_46384# 0.025246f
C21071 a_n4318_39768# SMPL_ON_P 0.039185f
C21072 a_n875_44318# a_n2497_47436# 9.25e-20
C21073 a_17517_44484# a_4883_46098# 7.99e-22
C21074 a_9159_44484# a_n1613_43370# 3.29e-21
C21075 a_8696_44636# a_6945_45028# 4.49e-20
C21076 a_1609_45572# a_n2661_45546# 1.69e-19
C21077 a_11652_45724# a_11608_46482# 2.38e-19
C21078 a_12427_45724# a_10586_45546# 2.09e-19
C21079 a_13249_42308# a_8049_45260# 0.00179f
C21080 a_n967_45348# a_n2293_46098# 2.05e-20
C21081 a_15595_45028# a_13059_46348# 1.93e-20
C21082 a_14539_43914# a_n743_46660# 1.85e-19
C21083 a_413_45260# a_22959_46660# 0.018266f
C21084 a_n1059_45260# a_n901_46420# 2.16e-20
C21085 a_n2661_44458# a_3877_44458# 0.035165f
C21086 a_21356_42826# a_13258_32519# 6.82e-21
C21087 a_19164_43230# a_7174_31319# 3.33e-21
C21088 a_196_42282# a_1184_42692# 2.75e-19
C21089 a_n784_42308# a_1576_42282# 0.038241f
C21090 a_n473_42460# a_961_42354# 2.64e-21
C21091 a_n3674_37592# a_n1630_35242# 0.096752f
C21092 COMP_P a_1606_42308# 2.6775f
C21093 a_10752_42852# a_5742_30871# 5.4e-20
C21094 a_n4318_38680# a_n2860_38778# 1.77e-20
C21095 a_n881_46662# a_7411_46660# 0.025876f
C21096 a_n1613_43370# a_7715_46873# 8.67e-20
C21097 a_16327_47482# a_3090_45724# 1.00134f
C21098 a_11599_46634# a_17609_46634# 5.91e-20
C21099 a_10227_46804# a_12991_46634# 0.349162f
C21100 a_15811_47375# a_15559_46634# 0.018669f
C21101 a_15507_47210# a_16292_46812# 3.28e-19
C21102 a_13717_47436# a_19692_46634# 3.9e-20
C21103 a_6151_47436# a_14180_46812# 6.21e-19
C21104 a_12861_44030# a_19466_46812# 0.004139f
C21105 a_2553_47502# a_765_45546# 0.003113f
C21106 a_n1151_42308# a_14226_46660# 2.85e-20
C21107 a_n2956_39768# a_n2661_46098# 1.22e-20
C21108 a_n743_46660# a_2107_46812# 0.72755f
C21109 a_n2661_46634# a_1799_45572# 0.0082f
C21110 a_n2438_43548# a_948_46660# 0.054839f
C21111 a_n133_46660# a_1123_46634# 0.043619f
C21112 a_33_46660# a_601_46902# 0.17072f
C21113 a_n1925_46634# a_288_46660# 0.003365f
C21114 a_171_46873# a_383_46660# 3.12e-19
C21115 a_22315_44484# a_22591_44484# 0.001038f
C21116 a_14537_43396# a_10341_43396# 0.013753f
C21117 a_9313_44734# a_10807_43548# 0.033005f
C21118 a_n2293_42834# a_6197_43396# 1.31e-19
C21119 a_1307_43914# a_14358_43442# 1.45e-20
C21120 a_n2661_42834# a_n2661_42282# 0.019795f
C21121 a_3422_30871# a_17730_32519# 0.004485f
C21122 a_7499_43078# a_8649_43218# 5.01e-19
C21123 a_n913_45002# a_743_42282# 0.25834f
C21124 a_19963_31679# a_14209_32519# 0.051256f
C21125 a_20447_31679# a_13887_32519# 0.051465f
C21126 a_7754_39964# VDD 0.848281f
C21127 a_19778_44110# VDD 0.469922f
C21128 a_15433_44458# a_11415_45002# 1.94e-20
C21129 a_13857_44734# a_12741_44636# 0.003456f
C21130 a_5205_44734# a_3483_46348# 3.63e-20
C21131 a_21381_43940# a_12549_44172# 0.099617f
C21132 a_19237_31679# a_19692_46634# 4.44e-20
C21133 a_375_42282# a_n755_45592# 0.366231f
C21134 a_2304_45348# a_n863_45724# 0.091195f
C21135 a_17613_45144# a_8049_45260# 1.7e-20
C21136 a_501_45348# a_n357_42282# 1.02e-19
C21137 a_13017_45260# a_n443_42852# 2.72e-20
C21138 a_4185_45348# a_n2661_45546# 1.35e-19
C21139 a_13720_44458# a_10903_43370# 2.88e-20
C21140 a_5883_43914# a_2324_44458# 0.002714f
C21141 a_n1917_43396# a_n1613_43370# 0.153085f
C21142 a_14579_43548# a_4915_47217# 2.85e-21
C21143 a_21613_42308# a_21421_42336# 5.76e-19
C21144 a_n784_42308# C1_P_btm 0.027772f
C21145 a_15559_46634# a_13059_46348# 0.167936f
C21146 a_14084_46812# a_14226_46660# 0.007833f
C21147 a_12251_46660# a_765_45546# 0.001931f
C21148 a_n881_46662# a_4365_46436# 5.52e-19
C21149 a_n743_46660# a_14493_46090# 0.007037f
C21150 a_13661_43548# a_10809_44734# 0.043589f
C21151 a_19452_47524# a_6945_45028# 4.72e-19
C21152 a_2107_46812# a_11189_46129# 1.06e-20
C21153 a_11453_44696# a_10586_45546# 0.005294f
C21154 a_4883_46098# a_12379_46436# 0.007631f
C21155 a_13507_46334# a_14180_46482# 0.001677f
C21156 a_11599_46634# a_19443_46116# 0.026712f
C21157 a_584_46384# a_1609_45822# 1.57e-20
C21158 a_2063_45854# a_n443_42852# 8.99e-20
C21159 a_n443_46116# a_1848_45724# 0.041711f
C21160 a_2124_47436# a_2277_45546# 5.88e-21
C21161 a_20835_44721# a_10341_43396# 2.07e-20
C21162 a_3600_43914# a_3626_43646# 3.68e-19
C21163 a_17973_43940# a_19319_43548# 2.01e-22
C21164 a_20193_45348# a_21356_42826# 1.21e-20
C21165 a_5883_43914# a_8387_43230# 2.5e-20
C21166 a_18451_43940# a_18533_44260# 0.003935f
C21167 a_5841_44260# a_n97_42460# 6.63e-22
C21168 a_9313_44734# a_13467_32519# 0.057668f
C21169 a_3537_45260# a_1755_42282# 0.002095f
C21170 a_n1059_45260# a_6171_42473# 2.78e-20
C21171 a_n2017_45002# a_5932_42308# 0.005049f
C21172 a_n913_45002# a_5755_42308# 0.036226f
C21173 a_6511_45714# a_2437_43646# 2.64e-21
C21174 a_5907_45546# a_3357_43084# 0.023698f
C21175 a_11229_43218# a_10227_46804# 0.001903f
C21176 a_n3674_37592# a_n971_45724# 0.022388f
C21177 a_n3420_37984# a_n923_35174# 0.002459f
C21178 a_19237_31679# a_20692_30879# 0.051625f
C21179 a_18249_42858# a_12549_44172# 4.15e-20
C21180 a_9127_43156# a_n2293_46634# 1.56e-19
C21181 a_13460_43230# a_13661_43548# 7.36e-20
C21182 a_10341_43396# a_3090_45724# 0.07129f
C21183 a_13565_43940# a_3483_46348# 0.006953f
C21184 a_20820_30879# VDD 0.719502f
C21185 a_n4064_39072# a_n3420_37984# 0.045543f
C21186 a_n3420_39072# a_n4064_37984# 0.045827f
C21187 a_4958_30871# VDAC_P 0.017827f
C21188 a_765_45546# a_13259_45724# 0.036082f
C21189 a_17339_46660# a_18147_46436# 0.002157f
C21190 a_10903_43370# a_13351_46090# 0.181897f
C21191 a_9569_46155# a_2324_44458# 5.17e-20
C21192 a_12005_46116# a_12594_46348# 0.065075f
C21193 a_472_46348# a_1431_46436# 6.01e-19
C21194 a_17737_43940# a_17595_43084# 8.42e-21
C21195 a_11341_43940# a_12379_42858# 2.86e-20
C21196 a_10555_44260# a_10083_42826# 9.41e-22
C21197 a_n2661_42282# a_n2293_42282# 1.04835f
C21198 a_n2293_43922# a_5267_42460# 4.38e-20
C21199 a_5891_43370# a_8515_42308# 1.03e-19
C21200 a_n356_44636# a_10723_42308# 2.77e-19
C21201 a_14539_43914# a_15486_42560# 4.81e-21
C21202 a_20974_43370# a_13467_32519# 0.017399f
C21203 a_14401_32519# a_4361_42308# 8.07e-20
C21204 a_n97_42460# a_16855_43396# 8.47e-19
C21205 a_16588_47582# RST_Z 5.09e-20
C21206 a_13487_47204# CLK 7.51e-19
C21207 a_11652_45724# a_8975_43940# 1.25e-20
C21208 a_8696_44636# a_11827_44484# 0.039f
C21209 a_16333_45814# a_11691_44458# 3.71e-21
C21210 a_2711_45572# a_5891_43370# 8.73e-21
C21211 a_16147_45260# a_16321_45348# 0.002641f
C21212 a_n913_45002# a_626_44172# 7.19e-20
C21213 a_3357_43084# a_6125_45348# 0.001261f
C21214 a_6171_45002# a_5205_44484# 0.0168f
C21215 a_5691_45260# a_7229_43940# 2.13e-20
C21216 a_3232_43370# a_7276_45260# 0.027376f
C21217 a_5534_30871# a_3483_46348# 2.26e-20
C21218 a_4921_42308# a_5257_43370# 0.002713f
C21219 a_548_43396# a_n443_42852# 2.03e-19
C21220 a_8952_43230# a_8953_45546# 0.01883f
C21221 a_10518_42984# a_8199_44636# 7.84e-20
C21222 a_n4334_39392# a_n2312_39304# 3.7e-20
C21223 a_17730_32519# VREF_GND 0.241027f
C21224 a_19237_31679# VIN_N 0.029585f
C21225 a_20107_45572# a_18479_47436# 0.025968f
C21226 a_2437_43646# a_14311_47204# 0.00629f
C21227 a_20841_45814# a_10227_46804# 3.53e-19
C21228 a_20731_45938# a_16327_47482# 0.012637f
C21229 a_3357_43084# a_13717_47436# 0.024679f
C21230 a_413_45260# a_n1151_42308# 0.135643f
C21231 a_5691_45260# a_n237_47217# 2.17e-21
C21232 a_3065_45002# a_584_46384# 0.085314f
C21233 a_6171_45002# a_n971_45724# 0.030962f
C21234 a_18175_45572# a_11453_44696# 0.036949f
C21235 a_19256_45572# a_4883_46098# 1.02e-20
C21236 a_16855_45546# a_n881_46662# 0.052296f
C21237 a_12016_45572# a_12549_44172# 7.31e-20
C21238 a_2711_45572# a_4817_46660# 9.24e-20
C21239 a_10053_45546# a_2107_46812# 1.1e-19
C21240 a_12427_45724# a_n743_46660# 1.63e-20
C21241 a_5907_45546# a_3877_44458# 4.21e-21
C21242 a_n2472_45546# a_n2956_38216# 0.157892f
C21243 a_n2661_45546# a_n2293_45546# 0.077901f
C21244 a_21076_30879# a_22521_39511# 6.56e-20
C21245 a_20820_30879# a_22469_39537# 7.31e-20
C21246 a_14513_46634# CLK 2.54e-20
C21247 a_1568_43370# a_1606_42308# 0.007194f
C21248 a_4190_30871# a_21195_42852# 1.06e-20
C21249 a_3935_42891# a_4520_42826# 0.017436f
C21250 a_5649_42852# a_18083_42858# 4.21e-20
C21251 a_4361_42308# a_18817_42826# 1.3e-20
C21252 a_n1557_42282# a_564_42282# 0.003471f
C21253 a_15493_43940# a_17531_42308# 1.35e-21
C21254 a_11341_43940# a_18727_42674# 3.06e-21
C21255 a_14579_43548# a_13291_42460# 0.007999f
C21256 a_3080_42308# a_1576_42282# 1.7e-20
C21257 a_n3674_39768# a_n3420_39072# 2.58e-20
C21258 a_7754_39964# a_8912_37509# 0.003864f
C21259 a_7754_40130# a_11206_38545# 0.736866f
C21260 a_2713_42308# VDD 0.208275f
C21261 a_n815_47178# a_n971_45724# 0.013837f
C21262 a_n1741_47186# a_n23_47502# 0.007866f
C21263 a_n2109_47186# a_327_47204# 0.041762f
C21264 SMPL_ON_P a_n237_47217# 4.88e-23
C21265 a_n1920_47178# a_n785_47204# 1.29e-19
C21266 a_13556_45296# a_13857_44734# 0.01375f
C21267 a_626_44172# a_556_44484# 0.00387f
C21268 a_2711_45572# a_18533_43940# 0.004398f
C21269 a_9482_43914# a_14112_44734# 0.004038f
C21270 a_19963_31679# a_17730_32519# 0.054244f
C21271 a_13657_42308# a_9290_44172# 1.07e-19
C21272 a_5932_42308# a_526_44458# 3.79e-19
C21273 a_8697_45572# a_3483_46348# 7.8e-19
C21274 a_11787_45002# a_6755_46942# 9.54e-22
C21275 a_19113_45348# a_5807_45002# 9.15e-19
C21276 a_21359_45002# a_19321_45002# 4.39e-19
C21277 a_22223_45036# a_13747_46662# 2.35e-19
C21278 a_19929_45028# a_12549_44172# 3.72e-20
C21279 a_3357_43084# a_14035_46660# 2.73e-20
C21280 a_n2661_44458# a_8128_46384# 1.73e-21
C21281 a_11525_45546# a_10903_43370# 0.040993f
C21282 a_11823_42460# a_9290_44172# 0.864145f
C21283 a_8162_45546# a_2324_44458# 4.52e-20
C21284 a_7227_45028# a_6945_45028# 0.016808f
C21285 a_11652_45724# a_11387_46155# 1.9e-19
C21286 a_11322_45546# a_12005_46116# 2.36e-19
C21287 a_12427_45724# a_11189_46129# 1.25e-19
C21288 a_10490_45724# a_12594_46348# 9.79e-19
C21289 a_n1917_44484# a_n1613_43370# 0.153277f
C21290 a_10440_44484# a_11453_44696# 4.13e-20
C21291 a_12883_44458# a_12465_44636# 0.017889f
C21292 a_18287_44626# a_18597_46090# 6.68e-22
C21293 a_13467_32519# a_22397_42558# 5.38e-19
C21294 a_4361_42308# a_21421_42336# 6.95e-19
C21295 a_10922_42852# a_5742_30871# 7.65e-19
C21296 a_12089_42308# a_10533_42308# 8.19e-21
C21297 a_10341_42308# a_11323_42473# 1.11e-19
C21298 a_n2293_42282# a_3497_42558# 0.001879f
C21299 a_3080_42308# C1_P_btm 0.011373f
C21300 a_n881_46662# a_13661_43548# 3.79e-20
C21301 a_2747_46873# a_n2661_46634# 0.019513f
C21302 a_n2312_39304# a_n2312_38680# 0.082563f
C21303 a_11453_44696# a_n743_46660# 0.004481f
C21304 a_4915_47217# a_5257_43370# 8.75e-20
C21305 a_n1435_47204# a_4646_46812# 4.92e-20
C21306 a_n237_47217# a_8035_47026# 1.8e-20
C21307 a_2063_45854# a_10554_47026# 0.002948f
C21308 a_n1151_42308# a_9863_46634# 2.6e-19
C21309 a_4791_45118# a_7715_46873# 1.8e-19
C21310 C8_N_btm VDD 0.19922f
C21311 a_18184_42460# a_15493_43940# 0.022388f
C21312 a_21101_45002# a_20935_43940# 0.001207f
C21313 a_n356_44636# a_175_44278# 6.51e-20
C21314 a_15433_44458# a_11967_42832# 7e-22
C21315 a_9313_44734# a_22315_44484# 2.17e-21
C21316 a_n2661_44458# a_9672_43914# 4.07e-20
C21317 a_11691_44458# a_15493_43396# 1.33e-19
C21318 a_11827_44484# a_20365_43914# 0.0059f
C21319 a_14537_43396# a_n97_42460# 1.86e-20
C21320 a_7499_43078# a_8037_42858# 0.160087f
C21321 a_2711_45572# a_17595_43084# 2.52e-20
C21322 a_4574_45260# a_3539_42460# 5.02e-22
C21323 a_5111_44636# a_2982_43646# 1.32e-19
C21324 a_n913_45002# a_2813_43396# 5.93e-20
C21325 a_9482_43914# VDD 1.75061f
C21326 a_n1630_35242# EN_VIN_BSTR_P 0.009334f
C21327 CAL_N a_20202_43084# 0.002046f
C21328 a_15037_43940# a_12861_44030# 1.65e-19
C21329 a_458_43396# a_584_46384# 0.196763f
C21330 a_14021_43940# SMPL_ON_N 1.94e-20
C21331 a_11361_45348# a_2324_44458# 1.97e-19
C21332 a_n2661_45010# a_n2661_45546# 0.014492f
C21333 a_2437_43646# a_n755_45592# 0.017992f
C21334 a_1423_45028# a_526_44458# 0.133656f
C21335 a_n2293_43922# a_3090_45724# 0.02667f
C21336 a_14955_43940# a_12549_44172# 0.010132f
C21337 a_n4318_39768# a_n2438_43548# 6.52e-19
C21338 a_13483_43940# a_768_44030# 0.002743f
C21339 a_n2267_44484# a_n1853_46287# 1.43e-21
C21340 a_22959_45036# a_4185_45028# 0.17601f
C21341 a_n2129_44697# a_n1991_46122# 2.79e-21
C21342 a_n2661_44458# a_n1641_46494# 1.32e-20
C21343 a_11691_44458# a_3483_46348# 0.039125f
C21344 a_2905_45572# VDD 1.22598f
C21345 a_n1630_35242# a_n2302_39072# 5.02e-20
C21346 a_n784_42308# a_1736_39043# 1.49e-20
C21347 a_n3674_38216# a_n3690_38528# 4.64e-19
C21348 a_14113_42308# a_13921_42308# 2.46e-19
C21349 a_15890_42674# a_15720_42674# 2.6e-19
C21350 a_n4318_37592# a_n4334_38528# 7.61e-20
C21351 a_n881_46662# a_4185_45028# 0.001491f
C21352 a_11453_44696# a_11189_46129# 2.99e-20
C21353 a_n1435_47204# a_n1545_46494# 4.84e-20
C21354 a_4883_46098# a_13351_46090# 0.006426f
C21355 a_13507_46334# a_13925_46122# 0.003355f
C21356 a_16327_47482# a_20075_46420# 0.270434f
C21357 a_14955_47212# a_10809_44734# 9.82e-20
C21358 a_15507_47210# a_6945_45028# 0.04755f
C21359 a_18597_46090# a_15682_46116# 1.97e-20
C21360 a_18143_47464# a_18189_46348# 1.76e-19
C21361 a_n443_46116# a_4365_46436# 1.01e-19
C21362 a_4791_45118# a_5210_46482# 1.81e-19
C21363 a_2063_45854# a_6633_46155# 4.03e-21
C21364 a_n1613_43370# a_4419_46090# 2.2e-19
C21365 a_21588_30879# a_12741_44636# 0.001298f
C21366 a_22612_30879# a_20820_30879# 0.061094f
C21367 a_8035_47026# a_8270_45546# 7.91e-21
C21368 a_6755_46942# a_11813_46116# 0.028837f
C21369 a_10249_46116# a_11901_46660# 3.57e-19
C21370 a_1799_45572# a_765_45546# 0.225248f
C21371 a_22315_44484# a_20974_43370# 1.76e-21
C21372 a_n2661_42834# a_7112_43396# 3.36e-20
C21373 a_n2661_43922# a_7287_43370# 2.05e-21
C21374 a_20193_45348# a_20749_43396# 0.003298f
C21375 a_11823_42460# a_15051_42282# 0.367924f
C21376 a_18114_32519# a_13467_32519# 0.055508f
C21377 a_10193_42453# a_10149_42308# 0.002618f
C21378 a_13249_42308# a_14456_42282# 1.37e-19
C21379 a_3422_30871# a_17538_32519# 0.005569f
C21380 a_n356_44636# a_10341_43396# 1.27e-20
C21381 a_2998_44172# a_3353_43940# 3.09e-19
C21382 a_5111_44636# a_5837_42852# 7.13e-19
C21383 a_20159_44458# VDD 0.345429f
C21384 a_10490_45724# a_11322_45546# 0.246478f
C21385 a_6511_45714# a_8192_45572# 1.94e-20
C21386 a_10193_42453# a_11652_45724# 0.197229f
C21387 a_8746_45002# a_11525_45546# 3.44e-21
C21388 a_2711_45572# a_11064_45572# 2.3e-19
C21389 a_8333_44056# a_3483_46348# 5.87e-19
C21390 a_15493_43940# a_12741_44636# 2.5e-19
C21391 a_n97_42460# a_3090_45724# 0.001209f
C21392 a_19177_43646# a_13661_43548# 0.015951f
C21393 a_5649_42852# a_12549_44172# 9.86e-20
C21394 a_n356_44636# a_n356_45724# 0.001699f
C21395 a_15433_44458# a_13259_45724# 2.36e-21
C21396 a_n1853_43023# a_n1613_43370# 0.423772f
C21397 a_10835_43094# a_10227_46804# 0.295543f
C21398 a_n914_42852# a_n1151_42308# 1.43e-19
C21399 a_413_45260# START 0.035622f
C21400 a_12816_46660# VDD 0.293798f
C21401 a_1208_46090# a_1138_42852# 0.043831f
C21402 a_805_46414# a_1823_45246# 6.82e-20
C21403 a_472_46348# a_2202_46116# 3.26e-20
C21404 a_376_46348# a_167_45260# 1.16e-21
C21405 a_3524_46660# a_3503_45724# 8.08e-21
C21406 a_11813_46116# a_8049_45260# 0.00127f
C21407 a_6755_46942# a_14949_46494# 5.41e-19
C21408 a_17339_46660# a_17957_46116# 0.098952f
C21409 a_765_45546# a_18189_46348# 0.013467f
C21410 a_14543_46987# a_10809_44734# 4.31e-19
C21411 a_5742_30871# VDAC_Pi 1.57e-19
C21412 a_5934_30871# a_3754_38470# 1.86e-19
C21413 a_n2293_46098# a_4419_46090# 0.051687f
C21414 a_9313_44734# a_18695_43230# 5.53e-19
C21415 a_5495_43940# a_5755_42852# 8.96e-22
C21416 a_15493_43396# a_4190_30871# 6e-19
C21417 a_15682_43940# a_4361_42308# 1.15e-20
C21418 a_4235_43370# a_2982_43646# 7.35e-20
C21419 a_n97_42460# a_6547_43396# 8.98e-20
C21420 a_14021_43940# a_17499_43370# 0.011011f
C21421 a_n2661_42282# a_n1423_42826# 2.27e-20
C21422 a_3422_30871# a_19339_43156# 1.85e-21
C21423 a_6031_43396# VDD 0.47547f
C21424 a_8696_44636# a_15595_45028# 1.68e-20
C21425 a_21188_45572# a_413_45260# 2.54e-21
C21426 a_3357_43084# a_n1059_45260# 0.003773f
C21427 a_18727_42674# a_16327_47482# 0.003774f
C21428 a_16269_42308# a_10227_46804# 1.79e-19
C21429 a_13258_32519# a_12861_44030# 9.87e-21
C21430 a_1755_42282# a_n2293_46634# 7.99e-22
C21431 a_6123_31319# a_768_44030# 1.76e-21
C21432 a_19987_42826# a_19692_46634# 5.42e-19
C21433 a_4361_42308# a_1823_45246# 0.11884f
C21434 a_2711_45572# a_11309_47204# 1.1e-19
C21435 a_6667_45809# a_n881_46662# 0.006711f
C21436 a_6598_45938# a_n1613_43370# 0.009561f
C21437 a_11682_45822# a_11599_46634# 7.01e-19
C21438 a_n1533_46116# a_n2293_45546# 2.26e-19
C21439 a_3080_42308# a_4649_42852# 5.53e-20
C21440 a_9145_43396# a_5342_30871# 0.002082f
C21441 a_4361_42308# a_22223_43396# 9.86e-19
C21442 a_21855_43396# a_5649_42852# 0.057783f
C21443 a_10341_43396# a_12379_42858# 2.27e-19
C21444 a_14358_43442# a_13635_43156# 8.12e-19
C21445 a_14579_43548# a_13460_43230# 1.97e-19
C21446 a_9028_43914# a_8685_42308# 1.61e-21
C21447 a_13467_32519# a_13887_32519# 0.058303f
C21448 a_3539_42460# a_4743_43172# 8.63e-20
C21449 a_20512_43084# a_21613_42308# 2.76e-20
C21450 VDAC_N C9_N_btm 0.44188p
C21451 a_7715_46873# DATA[3] 7.9e-19
C21452 a_18341_45572# a_17517_44484# 1.28e-20
C21453 a_626_44172# a_n2661_44458# 0.031248f
C21454 a_375_42282# a_n2129_44697# 1.85e-20
C21455 a_n143_45144# a_n356_44636# 4.67e-19
C21456 a_8953_45002# a_9838_44484# 0.013986f
C21457 a_6171_45002# a_13076_44458# 2.44e-20
C21458 a_n467_45028# a_n23_44458# 0.038286f
C21459 a_4933_42558# a_4185_45028# 0.001444f
C21460 a_10083_42826# a_n443_42852# 5.44e-19
C21461 a_5534_30871# a_n357_42282# 0.04831f
C21462 a_17538_32519# VREF_GND 0.117023f
C21463 a_21588_30879# C9_N_btm 0.786375f
C21464 a_20567_45036# a_16327_47482# 0.009073f
C21465 a_n2661_44458# a_6151_47436# 3.69e-21
C21466 a_20193_45348# a_12861_44030# 0.680394f
C21467 C2_P_btm VDD 0.268945f
C21468 a_n2661_43370# a_n2312_39304# 1.64e-20
C21469 a_n2017_45002# a_4646_46812# 5.44e-19
C21470 a_5111_44636# a_2107_46812# 7.67e-20
C21471 a_8191_45002# a_n1925_46634# 9.69e-19
C21472 a_413_45260# a_3177_46902# 0.006595f
C21473 a_16751_45260# a_5807_45002# 0.001196f
C21474 a_16020_45572# a_3090_45724# 0.001921f
C21475 a_10951_45334# a_n2293_46634# 3.22e-21
C21476 a_1307_43914# a_13661_43548# 0.396211f
C21477 a_13017_45260# a_n2661_46634# 0.123713f
C21478 a_15143_45578# a_765_45546# 1.48e-21
C21479 a_16333_45814# a_15227_44166# 4.01e-21
C21480 a_6598_45938# a_n2293_46098# 8.22e-20
C21481 a_1176_45572# a_1176_45822# 0.001923f
C21482 a_791_42968# a_961_42354# 0.003403f
C21483 a_1847_42826# a_1184_42692# 0.001067f
C21484 a_4361_42308# a_5934_30871# 0.092304f
C21485 a_5649_42852# a_7227_42308# 1.31e-19
C21486 a_743_42282# a_8325_42308# 0.02734f
C21487 a_16759_43396# a_15803_42450# 8.82e-20
C21488 a_10341_43396# a_18727_42674# 1.72e-20
C21489 a_3080_42308# a_1736_39043# 1.41e-19
C21490 a_13678_32519# a_6123_31319# 0.00363f
C21491 a_18599_43230# a_18695_43230# 0.013793f
C21492 a_n2302_38778# VDD 0.35162f
C21493 a_4915_47217# a_5807_45002# 0.766023f
C21494 a_9313_45822# a_11309_47204# 0.027145f
C21495 a_14955_47212# a_n881_46662# 0.008266f
C21496 a_n1435_47204# a_9804_47204# 1.58e-19
C21497 a_n2109_47186# a_1983_46706# 9.03e-20
C21498 a_n1741_47186# a_948_46660# 1.63e-20
C21499 a_n785_47204# a_n1021_46688# 0.001633f
C21500 a_n23_47502# a_n743_46660# 1.99e-20
C21501 a_n237_47217# a_n2438_43548# 0.02231f
C21502 a_n746_45260# a_n133_46660# 0.042075f
C21503 a_327_47204# a_n1925_46634# 1.53e-19
C21504 a_n971_45724# a_171_46873# 0.002898f
C21505 a_2063_45854# a_n2661_46634# 1.75382f
C21506 a_21177_47436# a_11453_44696# 3.75e-20
C21507 a_4883_46098# a_22223_47212# 1.16e-19
C21508 a_21811_47423# a_12465_44636# 0.00101f
C21509 a_2711_45572# a_13467_32519# 2.9e-19
C21510 a_n23_44458# a_n2661_43922# 0.007348f
C21511 a_18114_32519# a_22315_44484# 0.017551f
C21512 a_10193_42453# a_16759_43396# 5.51e-19
C21513 a_13556_45296# a_15493_43940# 2.77e-19
C21514 a_11823_42460# a_13749_43396# 1.72e-20
C21515 a_8375_44464# a_9313_44734# 8.59e-20
C21516 a_n356_44636# a_n2293_43922# 0.025509f
C21517 a_3537_45260# a_3737_43940# 0.012872f
C21518 a_19963_31679# a_17538_32519# 0.051095f
C21519 a_20447_31679# a_14401_32519# 0.054145f
C21520 a_19647_42308# a_n357_42282# 7.07e-20
C21521 a_20623_45572# VDD 0.200978f
C21522 a_1307_43914# a_4185_45028# 0.025209f
C21523 a_2809_45348# a_1823_45246# 2.74e-19
C21524 a_20640_44752# a_20916_46384# 9.21e-22
C21525 a_18587_45118# a_17339_46660# 0.003347f
C21526 a_18579_44172# a_13661_43548# 0.229269f
C21527 a_19279_43940# a_19321_45002# 0.019898f
C21528 a_10057_43914# a_8270_45546# 3.3e-19
C21529 a_17478_45572# a_18051_46116# 6.12e-19
C21530 a_13385_45572# a_13259_45724# 8.8e-20
C21531 a_3357_43084# a_n1925_42282# 0.067793f
C21532 a_n1761_44111# a_n881_46662# 6.91e-21
C21533 a_n1899_43946# a_n1613_43370# 0.038349f
C21534 a_6171_45002# a_12594_46348# 4.26e-20
C21535 a_8953_45002# a_9823_46155# 5.32e-19
C21536 a_413_45260# a_19553_46090# 4.37e-21
C21537 a_3537_45260# a_2324_44458# 0.015845f
C21538 a_2903_42308# a_5742_30871# 2.87e-20
C21539 a_6761_42308# a_5934_30871# 1.73e-20
C21540 a_22821_38993# RST_Z 1.55e-20
C21541 a_4791_45118# a_4419_46090# 4.81e-19
C21542 a_13661_43548# a_17609_46634# 0.002022f
C21543 a_4651_46660# a_5275_47026# 9.73e-19
C21544 a_4955_46873# a_5072_46660# 0.17431f
C21545 a_5385_46902# a_5732_46660# 0.051162f
C21546 a_4817_46660# a_6540_46812# 2.48e-19
C21547 a_3877_44458# a_3878_46660# 8.89e-19
C21548 a_12891_46348# a_12347_46660# 4.22e-19
C21549 a_n2661_46634# a_12469_46902# 0.001353f
C21550 a_2107_46812# a_6086_46660# 2.62e-19
C21551 a_2747_46873# a_765_45546# 0.040029f
C21552 a_11453_44696# a_20841_46902# 0.0185f
C21553 a_12465_44636# a_22000_46634# 0.001537f
C21554 a_10227_46804# a_11415_45002# 0.139042f
C21555 a_n1435_47204# a_n901_46420# 4.38e-21
C21556 a_4700_47436# a_4704_46090# 1.44e-19
C21557 a_2063_45854# a_8199_44636# 0.037924f
C21558 a_n1151_42308# a_6165_46155# 0.055317f
C21559 a_n443_46116# a_4185_45028# 6.94e-20
C21560 a_20679_44626# a_11341_43940# 4.56e-20
C21561 a_20766_44850# a_20935_43940# 0.003556f
C21562 a_18579_44172# a_19862_44208# 0.091151f
C21563 a_19279_43940# a_20623_43914# 1.14e-19
C21564 a_20835_44721# a_21115_43940# 3.62e-19
C21565 a_n356_44636# a_n97_42460# 1.46232f
C21566 a_4223_44672# a_6293_42852# 2.53e-19
C21567 a_11827_44484# a_14205_43396# 5.23e-22
C21568 a_9313_44734# a_19319_43548# 1.9e-20
C21569 a_n2661_42834# a_9801_43940# 4.77e-19
C21570 a_1414_42308# a_1525_44260# 2.45e-19
C21571 a_453_43940# a_1241_44260# 5.21e-19
C21572 a_5663_43940# a_7542_44172# 7.37e-21
C21573 a_5111_44636# a_7871_42858# 2.52e-19
C21574 a_3537_45260# a_8387_43230# 3.75e-19
C21575 a_3232_43370# a_5111_42852# 1.6e-21
C21576 a_n1059_45260# a_5342_30871# 0.030512f
C21577 a_n2017_45002# a_15567_42826# 0.002448f
C21578 a_n913_45002# a_15279_43071# 2.22e-19
C21579 a_n1809_44850# VDD 0.132538f
C21580 a_n4209_39304# C9_P_btm 3.29e-19
C21581 a_n4209_37414# a_n2810_45572# 3.74e-21
C21582 a_15037_43396# a_10227_46804# 0.002187f
C21583 a_11691_44458# a_n357_42282# 2.63e-20
C21584 a_18287_44626# a_8049_45260# 1.03e-20
C21585 a_8685_43396# a_12549_44172# 3.53e-19
C21586 a_15493_43396# a_15227_44166# 0.046514f
C21587 a_18579_44172# a_4185_45028# 1.48e-22
C21588 a_n4209_39304# a_n4209_38502# 0.042459f
C21589 a_n3565_39304# a_n2216_39072# 0.003034f
C21590 a_2443_46660# VDD 0.413663f
C21591 a_5742_30871# C9_N_btm 0.003249f
C21592 a_20107_46660# a_19636_46660# 3.64e-21
C21593 a_19123_46287# a_20719_46660# 8.64e-21
C21594 a_3877_44458# a_n1925_42282# 0.034241f
C21595 a_4646_46812# a_526_44458# 0.020719f
C21596 a_n743_46660# a_14180_46482# 0.002131f
C21597 a_19321_45002# a_19597_46482# 5.66e-19
C21598 a_n881_46662# a_997_45618# 1.94e-19
C21599 a_6755_46942# a_15682_46116# 0.116442f
C21600 a_6969_46634# a_2324_44458# 7e-22
C21601 a_7715_46873# a_6945_45028# 0.001653f
C21602 a_3090_45724# a_5204_45822# 2.88e-19
C21603 a_n1613_43370# a_1848_45724# 6.13e-21
C21604 a_n784_42308# a_n3420_37984# 0.009139f
C21605 a_17339_46660# a_11415_45002# 0.025523f
C21606 a_15227_44166# a_3483_46348# 0.595533f
C21607 a_22315_44484# a_13887_32519# 2.2e-22
C21608 a_9672_43914# a_9145_43396# 1.12e-19
C21609 a_12429_44172# a_8685_43396# 2.43e-20
C21610 a_20512_43084# a_4361_42308# 0.02826f
C21611 a_n2293_43922# a_12379_42858# 0.030458f
C21612 a_9313_44734# a_16795_42852# 0.008194f
C21613 a_n2293_42834# a_2903_42308# 1.2e-20
C21614 a_18184_42460# a_22765_42852# 0.012194f
C21615 a_n913_45002# a_13258_32519# 0.025596f
C21616 a_19963_31679# a_22465_38105# 3.53e-19
C21617 a_6671_43940# VDD 0.227011f
C21618 a_4099_45572# a_1423_45028# 2.06e-20
C21619 a_18479_45785# a_18596_45572# 0.183223f
C21620 a_18175_45572# a_18799_45938# 9.73e-19
C21621 a_18341_45572# a_19256_45572# 0.116691f
C21622 a_11525_45546# a_3232_43370# 7.67e-19
C21623 a_11322_45546# a_6171_45002# 0.069025f
C21624 a_8568_45546# a_8953_45002# 0.001119f
C21625 a_7499_43078# a_8191_45002# 0.002543f
C21626 a_n3565_37414# VREF_GND 0.0061f
C21627 a_9396_43370# a_4185_45028# 7.23e-21
C21628 a_13291_42460# a_5807_45002# 5.69e-21
C21629 a_22959_43396# a_19692_46634# 9.22e-20
C21630 a_15953_42852# a_12549_44172# 9.14e-21
C21631 a_261_44278# a_n443_42852# 2.42e-19
C21632 a_8333_44056# a_n357_42282# 6.5e-22
C21633 a_n4318_39304# a_n2956_38680# 0.023179f
C21634 a_15493_43940# a_16375_45002# 2.37e-20
C21635 a_2982_43646# a_9290_44172# 0.001406f
C21636 VDAC_N RST_Z 0.154233f
C21637 COMP_P a_n2312_39304# 0.00156f
C21638 a_n1329_42308# a_n2312_40392# 4e-20
C21639 VDAC_P C3_P_btm 6.90991f
C21640 a_18114_32519# VCM 0.121302f
C21641 a_19721_31679# VREF_GND 0.001975f
C21642 a_18819_46122# VDD 0.453432f
C21643 a_6511_45714# a_4915_47217# 2.36e-21
C21644 a_6194_45824# a_5815_47464# 2.21e-20
C21645 a_5907_45546# a_6151_47436# 0.274247f
C21646 a_6598_45938# a_4791_45118# 3.84e-19
C21647 a_6428_45938# a_2063_45854# 3.74e-19
C21648 a_8746_45002# a_n971_45724# 9.8e-20
C21649 a_11962_45724# a_n1741_47186# 6.79e-20
C21650 a_n4064_38528# VDAC_P 2.4e-19
C21651 a_n3565_38216# a_n2216_37690# 1e-19
C21652 a_n2293_46098# a_1848_45724# 0.006569f
C21653 a_n1853_46287# a_n755_45592# 0.021472f
C21654 a_1138_42852# a_n2661_45546# 0.023338f
C21655 a_376_46348# a_n863_45724# 1.69e-21
C21656 a_n1641_46494# a_n1099_45572# 0.0023f
C21657 a_15682_46116# a_8049_45260# 0.015666f
C21658 a_4905_42826# a_5111_42852# 0.105155f
C21659 a_9145_43396# a_743_42282# 1.59e-19
C21660 a_16243_43396# a_16977_43638# 0.053479f
C21661 a_16547_43609# a_16409_43396# 0.206231f
C21662 a_16137_43396# a_16759_43396# 2.32e-19
C21663 a_2896_43646# a_1847_42826# 9.63e-20
C21664 a_n97_42460# a_12379_42858# 5.61e-19
C21665 a_11967_42832# a_12563_42308# 1.15e-20
C21666 a_9313_44734# a_21335_42336# 0.002222f
C21667 a_10341_43396# a_17486_43762# 1.07e-19
C21668 a_5807_45002# DATA[5] 3.78e-20
C21669 a_21588_30879# RST_Z 0.052092f
C21670 a_10796_42968# VDD 0.270235f
C21671 a_16147_45260# a_14539_43914# 4.45e-20
C21672 a_10193_42453# a_17517_44484# 4.26e-19
C21673 a_10544_45572# a_9313_44734# 5.83e-20
C21674 a_11823_42460# a_12553_44484# 1.28e-19
C21675 a_8953_45002# a_n2661_43370# 0.034058f
C21676 a_n913_45002# a_20193_45348# 0.224918f
C21677 a_19963_31679# a_19721_31679# 9.01086f
C21678 a_6171_45002# a_15060_45348# 2.19e-19
C21679 a_17364_32525# a_20205_31679# 0.053947f
C21680 a_4190_30871# a_n357_42282# 0.035963f
C21681 a_16664_43396# a_n443_42852# 2.07e-20
C21682 a_10533_42308# a_3090_45724# 5.9e-20
C21683 a_14635_42282# a_3483_46348# 1.83e-20
C21684 a_15493_43940# RST_Z 0.004544f
C21685 a_n3420_37984# SMPL_ON_P 6.62e-21
C21686 a_13904_45546# a_6755_46942# 2.1e-21
C21687 a_19610_45572# a_19321_45002# 7.05e-19
C21688 en_comp a_n1613_43370# 1.09e-19
C21689 a_413_45260# a_3315_47570# 7.08e-19
C21690 a_6171_45002# a_12465_44636# 0.03098f
C21691 a_5205_44484# a_4883_46098# 1.69e-20
C21692 a_16019_45002# a_11599_46634# 8.13e-20
C21693 a_13159_45002# a_10227_46804# 1.01e-20
C21694 a_7639_45394# a_n1151_42308# 0.004199f
C21695 a_2448_45028# a_n443_46116# 6.56e-19
C21696 a_10903_45394# a_2063_45854# 1.39e-19
C21697 a_18083_42858# a_17333_42852# 0.284837f
C21698 a_2982_43646# a_15051_42282# 6.3e-19
C21699 a_n97_42460# a_18727_42674# 3.76e-20
C21700 a_4190_30871# a_18707_42852# 0.006254f
C21701 a_17701_42308# a_18249_42858# 2.98e-20
C21702 a_4958_30871# VDD 1.06745f
C21703 a_6545_47178# a_n1435_47204# 9.45e-19
C21704 a_6151_47436# a_13717_47436# 0.17202f
C21705 a_n2288_47178# a_n2312_40392# 0.153632f
C21706 a_n2497_47436# a_n2312_39304# 0.061823f
C21707 a_n971_45724# a_4883_46098# 0.031452f
C21708 a_4915_47217# a_14311_47204# 0.001913f
C21709 a_742_44458# a_n356_44636# 0.207503f
C21710 a_12607_44458# a_13076_44458# 0.200168f
C21711 a_n2661_44458# a_5289_44734# 5.74e-19
C21712 a_21363_45546# a_15493_43940# 1.34e-22
C21713 a_n2017_45002# a_10405_44172# 1.01e-20
C21714 a_413_45260# a_2537_44260# 1.26e-19
C21715 a_3232_43370# a_7542_44172# 1.17e-20
C21716 a_4921_42308# a_n755_45592# 0.001431f
C21717 a_n4334_40480# a_n2956_38680# 4.16e-19
C21718 a_n4064_40160# a_n2956_39304# 6.96e-19
C21719 a_5934_30871# a_n2810_45572# 1.88e-21
C21720 a_13887_32519# VCM 0.011087f
C21721 a_14209_32519# VREF 2.95e-20
C21722 a_20679_44626# a_16327_47482# 0.318301f
C21723 a_11967_42832# a_10227_46804# 0.461417f
C21724 a_2479_44172# a_584_46384# 0.054912f
C21725 a_n1287_44306# a_n2497_47436# 8.39e-19
C21726 a_2127_44172# a_2063_45854# 5.29e-20
C21727 a_14673_44172# a_12465_44636# 0.101564f
C21728 a_1260_45572# a_n2661_45546# 7.47e-19
C21729 a_11962_45724# a_10586_45546# 0.137051f
C21730 a_13904_45546# a_8049_45260# 0.003111f
C21731 en_comp a_n2293_46098# 0.003369f
C21732 a_2437_43646# a_3483_46348# 4.71e-20
C21733 a_16112_44458# a_n743_46660# 0.001708f
C21734 a_15415_45028# a_13059_46348# 2.08e-20
C21735 a_413_45260# a_12741_44636# 0.009139f
C21736 a_19987_42826# a_20107_42308# 0.001063f
C21737 a_20922_43172# a_13258_32519# 7.84e-20
C21738 a_n473_42460# a_1184_42692# 1.41e-19
C21739 a_n784_42308# a_1067_42314# 0.064066f
C21740 a_n327_42558# a_n1630_35242# 0.053474f
C21741 a_n3674_37592# a_564_42282# 1.04e-19
C21742 a_11554_42852# a_5742_30871# 3.85e-19
C21743 a_n2840_46634# a_n2661_46098# 3.35e-19
C21744 a_n1925_46634# a_1983_46706# 0.007111f
C21745 a_n743_46660# a_948_46660# 0.038448f
C21746 a_n2438_43548# a_1123_46634# 0.075317f
C21747 a_n133_46660# a_383_46660# 0.105995f
C21748 a_171_46873# a_601_46902# 2.33e-20
C21749 a_n881_46662# a_5257_43370# 0.447042f
C21750 a_n1613_43370# a_7411_46660# 1.61e-20
C21751 a_3080_42308# a_n3420_37984# 0.002941f
C21752 a_11599_46634# a_16292_46812# 7.78e-19
C21753 a_10227_46804# a_12251_46660# 0.188053f
C21754 a_15507_47210# a_15559_46634# 0.011624f
C21755 a_15811_47375# a_15368_46634# 2.18e-19
C21756 a_6151_47436# a_14035_46660# 6.85e-19
C21757 a_13717_47436# a_19466_46812# 2.28e-20
C21758 a_4915_47217# a_14226_46987# 8.89e-19
C21759 a_2063_45854# a_765_45546# 1.71006f
C21760 a_14797_45144# a_14955_43396# 4.74e-21
C21761 a_15004_44636# a_14021_43940# 7.55e-21
C21762 a_22315_44484# a_22485_44484# 0.109468f
C21763 a_9313_44734# a_10949_43914# 3.03e-20
C21764 a_4223_44672# a_7499_43940# 0.030206f
C21765 a_n2293_42834# a_6293_42852# 0.008221f
C21766 a_7499_43078# a_7309_42852# 0.011818f
C21767 a_3422_30871# a_22591_44484# 8.92e-19
C21768 a_n2661_42834# a_6101_44260# 2.26e-19
C21769 a_n1059_45260# a_743_42282# 0.198704f
C21770 a_19479_31679# a_17364_32525# 0.05375f
C21771 a_6171_45002# a_16409_43396# 6.7e-20
C21772 a_18911_45144# VDD 0.218047f
C21773 a_5742_30871# RST_Z 0.003575f
C21774 a_14815_43914# a_11415_45002# 0.070306f
C21775 a_13468_44734# a_12741_44636# 9.06e-19
C21776 a_4181_44734# a_3483_46348# 6.14e-20
C21777 a_5891_43370# a_1823_45246# 5.34e-19
C21778 a_19741_43940# a_12549_44172# 0.001206f
C21779 a_11967_42832# a_17339_46660# 0.493072f
C21780 a_17023_45118# a_8049_45260# 1.03e-20
C21781 a_375_42282# a_n357_42282# 0.142311f
C21782 a_2232_45348# a_n863_45724# 0.002794f
C21783 a_13076_44458# a_10903_43370# 5.54e-19
C21784 a_12607_44458# a_12594_46348# 1.79e-19
C21785 a_8701_44490# a_2324_44458# 0.001089f
C21786 a_n1699_43638# a_n1613_43370# 0.160308f
C21787 a_7_47243# VDD 7.01e-19
C21788 a_5342_30871# a_n3420_37440# 0.030303f
C21789 a_5534_30871# a_n4064_37440# 0.041703f
C21790 a_3877_44458# a_2698_46116# 6.32e-21
C21791 a_10467_46802# a_11415_45002# 7.12e-22
C21792 a_15368_46634# a_13059_46348# 0.101997f
C21793 a_15559_46634# a_15227_46910# 7.75e-19
C21794 a_14976_45028# a_16388_46812# 4.43e-20
C21795 a_n881_46662# a_1337_46116# 0.043447f
C21796 a_n743_46660# a_13925_46122# 0.041274f
C21797 a_5807_45002# a_10809_44734# 0.065594f
C21798 a_13747_46662# a_6945_45028# 0.035381f
C21799 a_2107_46812# a_9290_44172# 0.091636f
C21800 a_n2293_46634# a_2324_44458# 0.021161f
C21801 a_13507_46334# a_12638_46436# 0.001374f
C21802 a_4883_46098# a_12005_46436# 1.01e-19
C21803 a_10227_46804# a_13259_45724# 0.335001f
C21804 a_16327_47482# a_19431_46494# 1.79e-19
C21805 a_11599_46634# a_20254_46482# 3.41e-19
C21806 a_3785_47178# a_3503_45724# 9.09e-22
C21807 a_584_46384# a_n443_42852# 1.36389f
C21808 a_n443_46116# a_997_45618# 0.080297f
C21809 a_13717_47436# a_20205_31679# 2.49e-20
C21810 a_20679_44626# a_10341_43396# 1.82e-20
C21811 a_3600_43914# a_3540_43646# 1.75e-19
C21812 a_n2661_42282# a_n1177_43370# 1.78e-22
C21813 a_3905_42865# a_2982_43646# 0.006358f
C21814 a_8701_44490# a_8387_43230# 1.48e-20
C21815 a_18326_43940# a_18533_44260# 6.08e-19
C21816 a_20193_45348# a_20922_43172# 7.72e-19
C21817 a_1414_42308# a_1512_43396# 8.62e-19
C21818 a_2998_44172# a_3626_43646# 1.65e-19
C21819 a_n1059_45260# a_5755_42308# 1.66e-19
C21820 a_n2017_45002# a_6171_42473# 0.003106f
C21821 a_3537_45260# a_1606_42308# 3.89e-20
C21822 a_n913_45002# a_5421_42558# 0.006411f
C21823 a_10907_45822# a_8696_44636# 0.001403f
C21824 a_13904_45546# a_14127_45572# 0.011458f
C21825 a_6472_45840# a_2437_43646# 3.74e-21
C21826 a_15785_43172# a_12861_44030# 4.72e-19
C21827 a_n327_42558# a_n971_45724# 0.01976f
C21828 a_19237_31679# a_20205_31679# 0.051574f
C21829 a_9885_43646# a_3090_45724# 0.003881f
C21830 a_14955_43396# a_14976_45028# 6.28e-20
C21831 a_17333_42852# a_12549_44172# 9.44e-21
C21832 a_8387_43230# a_n2293_46634# 4.77e-21
C21833 a_13635_43156# a_13661_43548# 0.004897f
C21834 a_22591_46660# VDD 0.251892f
C21835 a_472_46348# a_1337_46436# 9.76e-19
C21836 a_3090_45724# a_3503_45724# 0.006081f
C21837 a_17339_46660# a_13259_45724# 0.038367f
C21838 a_15227_44166# a_n357_42282# 0.023198f
C21839 a_16388_46812# a_18051_46116# 3.66e-19
C21840 a_10903_43370# a_12594_46348# 0.169312f
C21841 a_11387_46155# a_13351_46090# 5.76e-21
C21842 a_9625_46129# a_2324_44458# 0.002476f
C21843 a_1343_38525# a_2113_38308# 0.325474f
C21844 a_n3565_39304# a_n2302_37984# 1.31e-19
C21845 a_5244_44056# a_5193_42852# 3.06e-21
C21846 a_21381_43940# a_4361_42308# 0.195418f
C21847 a_n2293_43922# a_3823_42558# 4.58e-20
C21848 a_5891_43370# a_5934_30871# 0.027588f
C21849 a_n356_44636# a_10533_42308# 1.57e-19
C21850 a_14539_43914# a_15051_42282# 1.16e-20
C21851 a_14401_32519# a_13467_32519# 0.050489f
C21852 a_11341_43940# a_10341_42308# 3.2e-20
C21853 a_16763_47508# RST_Z 2.3e-19
C21854 a_12861_44030# CLK 4.17e-19
C21855 a_11525_45546# a_8975_43940# 1.35e-20
C21856 a_15765_45572# a_11691_44458# 3.92e-20
C21857 a_2711_45572# a_8375_44464# 1.54e-21
C21858 a_n1059_45260# a_626_44172# 2.24e-19
C21859 a_6171_45002# a_6431_45366# 0.017465f
C21860 a_3232_43370# a_5205_44484# 0.217288f
C21861 a_14543_43071# a_3483_46348# 5.23e-21
C21862 a_13635_43156# a_4185_45028# 7.46e-20
C21863 a_743_42282# a_n1925_42282# 0.052333f
C21864 a_n144_43396# a_n443_42852# 5.19e-20
C21865 a_9127_43156# a_8953_45546# 0.00897f
C21866 a_7871_42858# a_9290_44172# 2.35e-19
C21867 a_n4209_39304# a_n2312_39304# 0.19527f
C21868 a_17730_32519# VREF 1.53e-20
C21869 a_19431_45546# a_4883_46098# 5.31e-20
C21870 a_20528_45572# a_16327_47482# 0.011969f
C21871 a_3357_43084# a_n1435_47204# 1.08491f
C21872 a_2437_43646# a_13487_47204# 0.014506f
C21873 a_413_45260# a_3160_47472# 0.208121f
C21874 a_2382_45260# a_2063_45854# 5.84e-19
C21875 a_3232_43370# a_n971_45724# 0.058382f
C21876 a_n37_45144# a_n1151_42308# 4.16e-19
C21877 a_16147_45260# a_11453_44696# 0.026325f
C21878 a_20273_45572# a_10227_46804# 4.14e-20
C21879 a_16115_45572# a_n881_46662# 0.033547f
C21880 a_11778_45572# a_12549_44172# 1.09e-19
C21881 a_2711_45572# a_4955_46873# 2.02e-20
C21882 a_5263_45724# a_3877_44458# 3.55e-21
C21883 a_9049_44484# a_2107_46812# 0.240008f
C21884 a_11962_45724# a_n743_46660# 1.66e-20
C21885 a_n2661_45546# a_n2956_38216# 0.15505f
C21886 a_n2810_45572# a_n2293_45546# 4.68e-19
C21887 a_15493_43396# a_19511_42282# 1.63e-19
C21888 a_21259_43561# a_21195_42852# 7.25e-20
C21889 a_4190_30871# a_21356_42826# 0.011885f
C21890 a_5649_42852# a_17701_42308# 4.59e-20
C21891 a_4361_42308# a_18249_42858# 1.62e-19
C21892 a_19095_43396# a_18599_43230# 3.23e-19
C21893 a_743_42282# a_19987_42826# 0.009731f
C21894 a_n1557_42282# a_n3674_37592# 0.022251f
C21895 a_n97_42460# a_3823_42558# 4.7e-21
C21896 a_15493_43940# a_17303_42282# 7.91e-22
C21897 a_n3674_39768# a_n3690_39392# 3.4e-19
C21898 a_n4318_39768# a_n3420_39072# 2.16e-21
C21899 a_20820_30879# a_22821_38993# 1.52e-19
C21900 a_14180_46812# CLK 1.54e-20
C21901 a_3754_38470# a_8530_39574# 0.059662f
C21902 VDAC_Pi a_6886_37412# 0.259481f
C21903 a_7754_39964# VDAC_N 2.46e-19
C21904 a_7754_40130# VDAC_P 0.334598f
C21905 a_2725_42558# VDD 0.005543f
C21906 a_n815_47178# a_n452_47436# 0.107449f
C21907 a_n1605_47204# a_n971_45724# 3.64e-19
C21908 a_n1741_47186# a_n237_47217# 0.083957f
C21909 a_n2109_47186# a_n785_47204# 0.43597f
C21910 SMPL_ON_P a_n746_45260# 9.03e-22
C21911 a_9482_43914# a_13857_44734# 0.011887f
C21912 a_2711_45572# a_19319_43548# 0.225335f
C21913 a_19479_31679# a_19237_31679# 9.049419f
C21914 a_19963_31679# a_22591_44484# 8.88e-20
C21915 a_22591_45572# a_17730_32519# 7.45e-20
C21916 a_11897_42308# a_9290_44172# 7.06e-19
C21917 a_14635_42282# a_n357_42282# 0.010701f
C21918 a_6171_42473# a_526_44458# 4.56e-20
C21919 a_9803_43646# CLK 2.81e-19
C21920 a_10951_45334# a_6755_46942# 8.67e-21
C21921 a_11827_44484# a_13747_46662# 0.044822f
C21922 a_21101_45002# a_19321_45002# 0.005955f
C21923 a_1307_43914# a_5257_43370# 0.020655f
C21924 a_2437_43646# a_14513_46634# 2.95e-20
C21925 a_3357_43084# a_13885_46660# 2.28e-20
C21926 a_413_45260# a_13607_46688# 1.59e-20
C21927 a_7229_43940# a_7832_46660# 7.4e-21
C21928 a_6598_45938# a_6945_45028# 0.005236f
C21929 a_10490_45724# a_12005_46116# 6.17e-19
C21930 a_11322_45546# a_10903_43370# 0.313957f
C21931 a_11525_45546# a_11387_46155# 4.09e-19
C21932 a_11962_45724# a_11189_46129# 1.89e-19
C21933 a_10193_42453# a_13351_46090# 3.16e-21
C21934 a_n1699_44726# a_n1613_43370# 0.166123f
C21935 a_12607_44458# a_12465_44636# 0.186652f
C21936 a_10334_44484# a_11453_44696# 0.001021f
C21937 a_18248_44752# a_18597_46090# 8.18e-21
C21938 a_13467_32519# a_21421_42336# 6.18e-19
C21939 a_4361_42308# a_21125_42558# 2.86e-19
C21940 a_10991_42826# a_5742_30871# 0.002659f
C21941 a_10796_42968# a_11551_42558# 8.41e-19
C21942 a_10835_43094# a_11633_42558# 3.72e-19
C21943 a_10341_42308# a_10723_42308# 0.024028f
C21944 a_13678_32519# a_22775_42308# 0.024479f
C21945 a_5649_42852# a_21613_42308# 0.02466f
C21946 a_17364_32525# a_13258_32519# 0.053358f
C21947 a_12549_44172# a_768_44030# 0.490163f
C21948 a_n881_46662# a_5807_45002# 0.243322f
C21949 a_n2312_39304# a_n2104_46634# 0.018871f
C21950 a_n2312_40392# a_n2312_38680# 0.052461f
C21951 a_n1435_47204# a_3877_44458# 5.83e-20
C21952 a_n443_46116# a_5257_43370# 4.89e-19
C21953 a_n237_47217# a_7832_46660# 0.008175f
C21954 a_2063_45854# a_10623_46897# 0.009821f
C21955 a_n1151_42308# a_8492_46660# 1.89e-20
C21956 a_n1741_47186# a_8270_45546# 1.71e-19
C21957 a_19778_44110# a_15493_43940# 0.033844f
C21958 a_18494_42460# a_11341_43940# 0.025825f
C21959 a_21005_45260# a_20935_43940# 4.06e-20
C21960 a_9313_44734# a_3422_30871# 0.043499f
C21961 a_n2661_44458# a_9028_43914# 4.82e-21
C21962 a_11827_44484# a_20269_44172# 0.002504f
C21963 a_14815_43914# a_11967_42832# 5.37e-21
C21964 a_7499_43078# a_7765_42852# 0.008252f
C21965 a_14673_44172# a_16241_44734# 0.002281f
C21966 a_3537_45260# a_3539_42460# 0.264936f
C21967 C7_N_btm VDD 0.121904f
C21968 a_13348_45260# VDD 0.083657f
C21969 a_n784_42308# EN_VIN_BSTR_N 0.051272f
C21970 a_n1630_35242# a_n923_35174# 0.029967f
C21971 a_22765_42852# RST_Z 1.67e-19
C21972 VDAC_N a_20820_30879# 0.001867f
C21973 a_13565_43940# a_12861_44030# 1.02e-19
C21974 a_n229_43646# a_584_46384# 3.24e-19
C21975 a_8704_45028# a_2324_44458# 9.12e-20
C21976 a_2437_43646# a_n357_42282# 1.4e-19
C21977 a_n2840_45002# a_n2661_45546# 0.002083f
C21978 a_626_44172# a_n1925_42282# 4.51e-21
C21979 a_10951_45334# a_8049_45260# 1.03e-20
C21980 a_17061_44484# a_6755_46942# 9.81e-19
C21981 a_13483_43940# a_12549_44172# 0.007788f
C21982 a_12429_44172# a_768_44030# 0.007216f
C21983 a_18989_43940# a_17339_46660# 0.002356f
C21984 a_n2661_43922# a_3090_45724# 0.044809f
C21985 a_22223_45036# a_4185_45028# 0.002889f
C21986 a_2952_47436# VDD 0.089131f
C21987 a_1606_42308# a_1343_38525# 1.72e-20
C21988 a_n3674_38680# a_n4064_38528# 0.557806f
C21989 a_n4318_38216# a_n3420_38528# 0.31769f
C21990 a_n4318_37592# a_n4209_38502# 1.31e-19
C21991 a_n1630_35242# a_n4064_39072# 1.85e-20
C21992 a_14113_42308# a_13657_42308# 6.05e-20
C21993 COMP_P a_2112_39137# 1.26e-21
C21994 a_4190_30871# a_n4064_37440# 0.032722f
C21995 a_6755_46942# a_11735_46660# 0.61229f
C21996 a_10249_46116# a_11813_46116# 0.001399f
C21997 a_n743_46660# a_16655_46660# 0.004413f
C21998 a_n881_46662# a_3699_46348# 0.203393f
C21999 a_n1613_43370# a_4185_45028# 1.83e-19
C22000 a_12465_44636# a_10903_43370# 0.003556f
C22001 a_11453_44696# a_9290_44172# 0.064153f
C22002 a_4883_46098# a_12594_46348# 0.022174f
C22003 a_13507_46334# a_13759_46122# 0.004601f
C22004 a_16327_47482# a_19335_46494# 0.155998f
C22005 a_11599_46634# a_6945_45028# 0.04727f
C22006 a_14311_47204# a_10809_44734# 3.31e-20
C22007 a_10227_46804# a_18189_46348# 2.07e-20
C22008 a_n443_46116# a_1337_46116# 0.002343f
C22009 a_n1741_47186# a_12638_46436# 0.016323f
C22010 a_2063_45854# a_6347_46155# 2.92e-21
C22011 a_20916_46384# a_12741_44636# 0.023496f
C22012 a_21588_30879# a_20820_30879# 0.084472f
C22013 a_3422_30871# a_20974_43370# 0.020902f
C22014 a_22315_44484# a_14401_32519# 0.002016f
C22015 a_n2661_43922# a_6547_43396# 6.85e-21
C22016 a_n2661_42834# a_7287_43370# 1.79e-19
C22017 a_11823_42460# a_14113_42308# 0.103699f
C22018 a_2889_44172# a_3353_43940# 6.46e-21
C22019 a_13249_42308# a_13575_42558# 0.088907f
C22020 a_20193_45348# a_17364_32525# 1.2e-19
C22021 a_10193_42453# a_9885_42308# 2.33e-20
C22022 a_2998_44172# a_3052_44056# 3.81e-19
C22023 a_5111_44636# a_5193_42852# 0.018763f
C22024 a_n1059_45260# a_16328_43172# 0.009298f
C22025 a_19615_44636# VDD 0.203841f
C22026 a_10193_42453# a_11525_45546# 0.0979f
C22027 a_7499_43078# a_11823_42460# 0.002874f
C22028 a_8746_45002# a_11322_45546# 3.97e-21
C22029 a_2711_45572# a_10544_45572# 2.65e-19
C22030 a_15493_43940# a_20820_30879# 1.28e-20
C22031 a_13678_32519# a_12549_44172# 0.004825f
C22032 a_21845_43940# a_19692_46634# 0.014352f
C22033 a_15743_43084# a_n2293_46634# 8.65e-20
C22034 a_14815_43914# a_13259_45724# 0.001261f
C22035 a_2675_43914# a_2324_44458# 7.61e-20
C22036 a_n2157_42858# a_n1613_43370# 0.303592f
C22037 a_10518_42984# a_10227_46804# 0.225803f
C22038 a_413_45260# RST_Z 0.199496f
C22039 a_12991_46634# VDD 0.357655f
C22040 a_n3420_39072# C1_P_btm 6.64e-20
C22041 a_n2293_46098# a_4185_45028# 0.06423f
C22042 a_472_46348# a_1823_45246# 0.001742f
C22043 a_1208_46090# a_1176_45822# 0.141891f
C22044 a_805_46414# a_1138_42852# 2.41e-19
C22045 a_11735_46660# a_8049_45260# 8.52e-20
C22046 a_3699_46634# a_3503_45724# 6.06e-21
C22047 a_8270_45546# a_10586_45546# 3.82e-21
C22048 a_17339_46660# a_18189_46348# 0.170772f
C22049 a_765_45546# a_17715_44484# 0.117636f
C22050 a_14226_46987# a_10809_44734# 4.26e-19
C22051 a_19328_44172# a_4190_30871# 4.64e-22
C22052 a_15037_43940# a_9145_43396# 3.15e-19
C22053 a_14021_43940# a_16759_43396# 0.007414f
C22054 a_4093_43548# a_2982_43646# 1.2e-20
C22055 a_n2661_42282# a_n1991_42858# 7.14e-21
C22056 a_5495_43940# a_5111_42852# 5.29e-20
C22057 a_3422_30871# a_18599_43230# 6.68e-21
C22058 a_n229_43646# a_n144_43396# 1.48e-19
C22059 a_n2293_43922# a_12800_43218# 0.011493f
C22060 a_9313_44734# a_18504_43218# 0.002026f
C22061 a_n97_42460# a_6765_43638# 2.79e-19
C22062 a_n2956_37592# a_n3565_38216# 0.074137f
C22063 a_16115_45572# a_1307_43914# 0.001401f
C22064 a_8696_44636# a_15415_45028# 4.71e-20
C22065 a_3357_43084# a_n2017_45002# 3.91e-19
C22066 a_16197_42308# a_10227_46804# 0.001903f
C22067 a_3457_43396# a_526_44458# 0.002177f
C22068 a_6511_45714# a_n881_46662# 0.149116f
C22069 a_6667_45809# a_n1613_43370# 0.007328f
C22070 a_11322_45546# a_4883_46098# 9.36e-20
C22071 a_15143_45578# a_10227_46804# 0.010124f
C22072 a_2324_44458# a_2277_45546# 8.22e-19
C22073 a_4699_43561# a_4649_42852# 1.98e-20
C22074 a_4361_42308# a_5649_42852# 0.064476f
C22075 a_21855_43396# a_13678_32519# 0.17881f
C22076 a_13667_43396# a_13460_43230# 8.37e-20
C22077 a_12281_43396# a_10835_43094# 3.18e-20
C22078 a_19237_31679# a_13258_32519# 0.055803f
C22079 a_4190_30871# a_20749_43396# 0.018962f
C22080 a_14579_43548# a_13635_43156# 0.003436f
C22081 a_3080_42308# a_4149_42891# 0.001517f
C22082 a_3539_42460# a_4649_43172# 0.001762f
C22083 a_10341_43396# a_10341_42308# 9.26e-19
C22084 a_n97_42460# a_12800_43218# 4.03e-19
C22085 a_20512_43084# a_21887_42336# 1.58e-19
C22086 VDAC_N C8_N_btm 0.220913p
C22087 a_7411_46660# DATA[3] 7.26e-20
C22088 a_18479_45785# a_17517_44484# 0.023114f
C22089 a_9482_43914# a_4223_44672# 3.83e-21
C22090 a_8953_45002# a_5883_43914# 0.008516f
C22091 a_n467_45028# a_n356_44636# 0.052527f
C22092 a_3232_43370# a_13076_44458# 4.99e-21
C22093 a_8952_43230# a_n443_42852# 7.98e-19
C22094 a_14543_43071# a_n357_42282# 0.004653f
C22095 a_3080_42308# EN_VIN_BSTR_N 0.04304f
C22096 a_14401_32519# VCM 0.007907f
C22097 a_21588_30879# C8_N_btm 0.002806f
C22098 a_13490_45067# a_13507_46334# 6.13e-20
C22099 a_11827_44484# a_11599_46634# 1.7e-22
C22100 a_18494_42460# a_16327_47482# 0.083754f
C22101 a_16922_45042# a_18597_46090# 0.028931f
C22102 a_11691_44458# a_12861_44030# 0.196929f
C22103 C3_P_btm VDD 0.26836f
C22104 a_8975_43940# a_n971_45724# 7.38e-21
C22105 a_n2661_43370# a_n2312_40392# 1.34e-19
C22106 a_7229_43940# a_n743_46660# 6.59e-21
C22107 a_7705_45326# a_n1925_46634# 9.07e-21
C22108 a_5147_45002# a_2107_46812# 4.3e-20
C22109 a_413_45260# a_2609_46660# 0.022446f
C22110 a_8696_44636# a_15368_46634# 2.65e-20
C22111 a_2903_45348# a_768_44030# 0.001561f
C22112 a_15861_45028# a_14976_45028# 1.41e-19
C22113 a_16019_45002# a_13661_43548# 0.001206f
C22114 a_10775_45002# a_n2293_46634# 1.79e-21
C22115 a_1307_43914# a_5807_45002# 0.007287f
C22116 a_15595_45028# a_13747_46662# 3.1e-20
C22117 a_11963_45334# a_n2661_46634# 0.036874f
C22118 a_15765_45572# a_15227_44166# 2.32e-20
C22119 a_17478_45572# a_3090_45724# 0.128299f
C22120 a_6667_45809# a_n2293_46098# 1.01e-20
C22121 a_16977_43638# a_15803_42450# 9.29e-20
C22122 a_791_42968# a_1184_42692# 8.46e-19
C22123 a_5111_42852# a_n784_42308# 3.45e-21
C22124 a_5649_42852# a_6761_42308# 9.04e-20
C22125 a_4361_42308# a_7963_42308# 0.007925f
C22126 a_10341_43396# a_18057_42282# 5.97e-21
C22127 a_3080_42308# a_1239_39043# 1.03e-19
C22128 a_13467_32519# a_5934_30871# 0.003932f
C22129 a_16795_42852# a_16877_42852# 0.171361f
C22130 a_8292_43218# a_8483_43230# 4.61e-19
C22131 a_18599_43230# a_18504_43218# 0.049827f
C22132 a_18817_42826# a_18695_43230# 3.16e-19
C22133 a_1847_42826# a_1576_42282# 2.07e-19
C22134 a_743_42282# a_8337_42558# 4.14e-19
C22135 a_n4064_38528# VDD 1.69517f
C22136 a_11031_47542# a_11309_47204# 0.110775f
C22137 a_14311_47204# a_n881_46662# 0.037789f
C22138 a_9313_45822# a_11117_47542# 6.66e-19
C22139 a_n1435_47204# a_8128_46384# 9.08e-20
C22140 a_n2109_47186# a_2107_46812# 0.032545f
C22141 a_n1741_47186# a_1123_46634# 9.86e-20
C22142 a_n746_45260# a_n2438_43548# 0.031949f
C22143 a_n237_47217# a_n743_46660# 0.192378f
C22144 a_n971_45724# a_n133_46660# 0.011188f
C22145 a_584_46384# a_n2661_46634# 0.034039f
C22146 a_n785_47204# a_n1925_46634# 2.12e-19
C22147 a_20990_47178# a_11453_44696# 1.3e-19
C22148 a_4883_46098# a_12465_44636# 0.024607f
C22149 a_13777_45326# a_11341_43940# 3.2e-21
C22150 a_n356_44636# a_n2661_43922# 0.041936f
C22151 a_n23_44458# a_n2661_42834# 0.001339f
C22152 a_9482_43914# a_15493_43940# 1.42e-19
C22153 a_18114_32519# a_3422_30871# 0.001438f
C22154 a_13720_44458# a_13940_44484# 0.009965f
C22155 a_7640_43914# a_9313_44734# 0.001487f
C22156 a_10193_42453# a_16977_43638# 7.87e-19
C22157 a_3065_45002# a_3992_43940# 0.002689f
C22158 a_19511_42282# a_n357_42282# 0.056757f
C22159 a_7174_31319# a_n863_45724# 4.84e-21
C22160 a_20841_45814# VDD 0.209907f
C22161 a_1423_45028# a_167_45260# 0.123079f
C22162 a_2304_45348# a_1823_45246# 4.41e-19
C22163 a_18315_45260# a_17339_46660# 0.009833f
C22164 a_18579_44172# a_5807_45002# 0.003978f
C22165 a_20766_44850# a_19321_45002# 0.004119f
C22166 a_13249_42308# a_n443_42852# 0.033352f
C22167 a_13297_45572# a_13259_45724# 0.003457f
C22168 a_19418_45938# a_8049_45260# 1.68e-19
C22169 a_3357_43084# a_526_44458# 0.04478f
C22170 a_11963_45334# a_8199_44636# 8.83e-21
C22171 a_n1761_44111# a_n1613_43370# 0.148121f
C22172 a_6171_45002# a_12005_46116# 1.39e-20
C22173 a_8953_45002# a_9569_46155# 0.002046f
C22174 a_413_45260# a_18985_46122# 1.46e-21
C22175 a_3429_45260# a_2324_44458# 2.54e-20
C22176 a_2713_42308# a_5742_30871# 1.69e-20
C22177 a_6761_42308# a_7963_42308# 9.72e-20
C22178 a_7227_42308# a_6123_31319# 0.189956f
C22179 EN_VIN_BSTR_P a_n83_35174# 0.652984f
C22180 a_22545_38993# RST_Z 1.94e-21
C22181 a_n743_46660# a_8270_45546# 0.274248f
C22182 a_5807_45002# a_17609_46634# 2.45e-19
C22183 a_n2661_46634# a_11901_46660# 0.030789f
C22184 a_13747_46662# a_15559_46634# 1.73e-20
C22185 a_4817_46660# a_5732_46660# 0.118759f
C22186 a_4651_46660# a_5072_46660# 0.083408f
C22187 a_4646_46812# a_5275_47026# 8.49e-19
C22188 a_3877_44458# a_3633_46660# 2.14e-19
C22189 a_n1925_46634# a_8601_46660# 6.89e-21
C22190 a_12891_46348# a_12978_47026# 1.98e-19
C22191 a_2107_46812# a_5841_46660# 1.55e-19
C22192 a_12465_44636# a_21188_46660# 3.64e-21
C22193 a_11453_44696# a_20273_46660# 0.545219f
C22194 a_10227_46804# a_20202_43084# 0.022898f
C22195 a_4915_47217# a_3483_46348# 1.09e-19
C22196 a_n1435_47204# a_n1641_46494# 2.5e-20
C22197 a_18479_47436# a_20885_46660# 6.01e-19
C22198 a_n1151_42308# a_5497_46414# 0.089064f
C22199 a_4791_45118# a_4185_45028# 0.064362f
C22200 a_18494_42460# a_10341_43396# 0.030934f
C22201 a_20159_44458# a_15493_43940# 7.59e-20
C22202 a_20835_44721# a_20935_43940# 4.15e-19
C22203 a_20640_44752# a_11341_43940# 4.18e-22
C22204 a_20679_44626# a_21115_43940# 0.003825f
C22205 a_17517_44484# a_14021_43940# 6.77e-21
C22206 a_18579_44172# a_19478_44306# 0.040429f
C22207 a_19279_43940# a_20365_43914# 0.003068f
C22208 a_4223_44672# a_6031_43396# 1.22e-19
C22209 a_1414_42308# a_1241_44260# 9.75e-20
C22210 a_3537_45260# a_8605_42826# 2.91e-20
C22211 a_5111_44636# a_7227_42852# 1.22e-20
C22212 a_n913_45002# a_5534_30871# 0.274894f
C22213 a_n1059_45260# a_15279_43071# 0.021145f
C22214 a_n2017_45002# a_5342_30871# 0.038471f
C22215 a_n2012_44484# VDD 0.077632f
C22216 a_n4315_30879# VIN_P 0.187185f
C22217 a_n4209_39304# C10_P_btm 4.87e-19
C22218 a_15743_43084# a_18597_46090# 0.023066f
C22219 a_4190_30871# a_12861_44030# 6.78e-20
C22220 a_n1076_43230# a_n1151_42308# 0.00783f
C22221 a_18248_44752# a_8049_45260# 6.37e-21
C22222 a_20935_43940# a_3090_45724# 1.49e-20
C22223 a_3539_42460# a_n2293_46634# 0.003606f
C22224 a_8685_43396# a_12891_46348# 3.82e-20
C22225 a_n4209_39590# a_n4209_38216# 0.031951f
C22226 a_n4064_39072# a_n3607_39392# 4.68e-19
C22227 a_n3565_39304# a_n2860_39072# 0.001021f
C22228 a_n2661_46098# VDD 0.979859f
C22229 a_5742_30871# C8_N_btm 0.003514f
C22230 a_19551_46910# a_19636_46660# 1.48e-19
C22231 a_768_44030# a_n2661_45546# 0.07332f
C22232 a_3877_44458# a_526_44458# 0.017621f
C22233 a_5807_45002# a_19443_46116# 0.003665f
C22234 a_13747_46662# a_20009_46494# 9.03e-20
C22235 a_n881_46662# a_n755_45592# 0.077214f
C22236 a_6755_46942# a_2324_44458# 0.155169f
C22237 a_7411_46660# a_6945_45028# 0.004283f
C22238 a_3090_45724# a_5164_46348# 1.94e-19
C22239 a_n1613_43370# a_997_45618# 1.47e-20
C22240 a_n2661_43922# a_12379_42858# 2.39e-19
C22241 a_n2293_43922# a_10341_42308# 1.51e-20
C22242 a_9313_44734# a_16414_43172# 0.007521f
C22243 a_1307_43914# a_9223_42460# 3.82e-21
C22244 a_3422_30871# a_13887_32519# 0.031713f
C22245 a_18494_42460# a_20356_42852# 0.014237f
C22246 a_20512_43084# a_13467_32519# 0.021245f
C22247 a_18184_42460# a_20753_42852# 0.029113f
C22248 a_n2661_42834# a_12089_42308# 1.12e-20
C22249 a_n913_45002# a_19647_42308# 3.13e-19
C22250 a_n1059_45260# a_13258_32519# 4.14e-21
C22251 a_5829_43940# VDD 0.156797f
C22252 a_6511_45714# a_1307_43914# 9.73e-22
C22253 a_18175_45572# a_18596_45572# 0.086708f
C22254 a_18341_45572# a_19431_45546# 0.041762f
C22255 a_18909_45814# a_18691_45572# 0.209641f
C22256 a_18479_45785# a_19256_45572# 0.044595f
C22257 a_11322_45546# a_3232_43370# 4.14e-19
C22258 a_10490_45724# a_6171_45002# 3.24e-19
C22259 a_8568_45546# a_8191_45002# 9.41e-20
C22260 a_7499_43078# a_7705_45326# 2.7e-19
C22261 a_n4209_37414# VCM 0.03628f
C22262 a_8791_43396# a_4185_45028# 4.43e-22
C22263 a_5837_43396# a_1823_45246# 3.58e-21
C22264 a_14209_32519# a_19692_46634# 9.21e-20
C22265 a_13814_43218# a_13661_43548# 4.89e-20
C22266 a_n4318_39304# a_n2956_39304# 0.023717f
C22267 a_6886_37412# RST_Z 0.031637f
C22268 COMP_P a_n2312_40392# 0.035637f
C22269 a_n4318_37592# a_n2312_39304# 0.023445f
C22270 a_n3565_37414# VREF 0.046045f
C22271 a_n3420_37440# VIN_P 0.143165f
C22272 VDAC_P C4_P_btm 13.8049f
C22273 a_n2661_44458# CLK 2.88e-19
C22274 a_18114_32519# VREF_GND 0.493553f
C22275 a_19721_31679# VREF 0.057702f
C22276 a_17957_46116# VDD 0.138777f
C22277 a_6472_45840# a_4915_47217# 6.14e-21
C22278 a_2711_45572# a_6851_47204# 3.11e-21
C22279 a_5263_45724# a_6151_47436# 3e-19
C22280 a_6667_45809# a_4791_45118# 0.005119f
C22281 a_n2293_46098# a_997_45618# 0.003758f
C22282 a_1176_45822# a_n2661_45546# 0.004027f
C22283 a_n1076_46494# a_n863_45724# 1.04e-19
C22284 a_n901_46420# a_n452_45724# 0.004896f
C22285 a_n2956_38680# a_n1925_42282# 4.34e-20
C22286 a_2324_44458# a_8049_45260# 0.054166f
C22287 a_11189_46129# a_12638_46436# 1.22e-19
C22288 a_8685_43396# a_4361_42308# 1.36e-19
C22289 a_16243_43396# a_16409_43396# 0.575934f
C22290 a_16137_43396# a_16977_43638# 6.31e-20
C22291 a_18533_43940# a_18249_42858# 1.68e-20
C22292 a_4905_42826# a_4520_42826# 0.147708f
C22293 a_n97_42460# a_10341_42308# 0.005646f
C22294 a_895_43940# a_1755_42282# 3.72e-21
C22295 a_9313_44734# a_7174_31319# 1.37e-19
C22296 a_10341_43396# a_15940_43402# 4.63e-19
C22297 a_20843_47204# SINGLE_ENDED 0.007105f
C22298 a_5807_45002# DATA[4] 3.14e-21
C22299 a_20916_46384# RST_Z 3.17e-20
C22300 a_10835_43094# VDD 0.43308f
C22301 a_16147_45260# a_16112_44458# 7.04e-19
C22302 a_2711_45572# a_3422_30871# 1.83e-19
C22303 a_10193_42453# a_17061_44734# 0.012286f
C22304 a_8191_45002# a_n2661_43370# 0.013381f
C22305 a_n913_45002# a_11691_44458# 2.08e-20
C22306 a_19963_31679# a_18114_32519# 0.051445f
C22307 a_22591_45572# a_19721_31679# 0.001292f
C22308 a_6171_45002# a_14976_45348# 1.2e-19
C22309 a_9306_43218# a_8953_45546# 2.14e-19
C22310 a_14209_32519# a_20692_30879# 0.051612f
C22311 a_21259_43561# a_n357_42282# 1.65e-19
C22312 a_n2216_39072# a_n2312_38680# 3.1e-19
C22313 a_22223_43948# RST_Z 7.78e-20
C22314 a_13527_45546# a_6755_46942# 0.001323f
C22315 a_21363_45546# a_20916_46384# 2.9e-19
C22316 a_21350_45938# a_13747_46662# 1.02e-20
C22317 a_2437_43646# a_16942_47570# 3.81e-19
C22318 a_413_45260# a_3094_47570# 7.88e-19
C22319 a_3232_43370# a_12465_44636# 1.26e-20
C22320 a_15595_45028# a_11599_46634# 0.001416f
C22321 a_13017_45260# a_10227_46804# 9.45e-19
C22322 a_7418_45394# a_n1151_42308# 1.53e-19
C22323 a_9396_43370# a_9223_42460# 4.27e-20
C22324 a_17701_42308# a_17333_42852# 0.061051f
C22325 a_2982_43646# a_14113_42308# 2.12e-19
C22326 a_n97_42460# a_18057_42282# 2.69e-20
C22327 a_5755_42852# a_6101_43172# 0.013377f
C22328 a_17595_43084# a_18249_42858# 2.35e-19
C22329 a_4419_46090# DATA[2] 2.81e-19
C22330 a_2063_45854# a_10227_46804# 0.186188f
C22331 a_6151_47436# a_n1435_47204# 0.061966f
C22332 a_6575_47204# a_9067_47204# 0.210614f
C22333 a_4915_47217# a_13487_47204# 0.013601f
C22334 a_n2497_47436# a_n2312_40392# 0.194574f
C22335 a_n2833_47464# a_n2312_39304# 0.009425f
C22336 a_n1352_44484# a_n23_44458# 2.56e-20
C22337 a_n452_44636# a_n356_44636# 0.318214f
C22338 a_12607_44458# a_12883_44458# 0.11453f
C22339 a_7499_43078# a_2982_43646# 6.36e-19
C22340 a_n1699_44726# a_n1243_44484# 4.2e-19
C22341 a_n2661_44458# a_5205_44734# 2.45e-19
C22342 a_11827_44484# a_10617_44484# 1.33e-19
C22343 a_20623_45572# a_15493_43940# 1.03e-21
C22344 a_5205_44484# a_5495_43940# 4.22e-20
C22345 a_n913_45002# a_8333_44056# 3.9e-21
C22346 a_n1059_45260# a_9028_43914# 0.002455f
C22347 a_n967_45348# a_n2661_42282# 2.72e-19
C22348 a_413_45260# a_2253_44260# 1.2e-19
C22349 a_6171_45002# a_6453_43914# 1.38e-19
C22350 a_3232_43370# a_7281_43914# 0.001158f
C22351 a_5932_42308# a_n863_45724# 4.31e-21
C22352 a_4921_42308# a_n357_42282# 3.76e-19
C22353 a_n4315_30879# a_n2956_38680# 0.024632f
C22354 a_n4334_40480# a_n2956_39304# 2.77e-19
C22355 a_13887_32519# VREF_GND 0.047292f
C22356 a_14209_32519# VIN_N 0.044892f
C22357 a_14581_44484# a_12465_44636# 5.1e-19
C22358 a_17517_44484# a_13507_46334# 0.018934f
C22359 a_20640_44752# a_16327_47482# 0.044807f
C22360 a_18753_44484# a_12861_44030# 2.16e-19
C22361 a_2127_44172# a_584_46384# 8.16e-20
C22362 a_n1453_44318# a_n2497_47436# 0.001884f
C22363 a_14127_45572# a_2324_44458# 6.43e-19
C22364 a_1176_45572# a_n2661_45546# 5.5e-19
C22365 a_10193_42453# a_12005_46436# 2.62e-20
C22366 a_9241_45822# a_5066_45546# 2.98e-19
C22367 a_13527_45546# a_8049_45260# 0.001929f
C22368 a_11652_45724# a_10586_45546# 0.046802f
C22369 a_413_45260# a_20820_30879# 0.033659f
C22370 a_16922_45042# a_6755_46942# 6.22e-19
C22371 a_14797_45144# a_13059_46348# 0.066603f
C22372 a_n745_45366# a_n1853_46287# 0.002206f
C22373 a_2437_43646# a_3147_46376# 1.06e-20
C22374 a_n913_45002# a_n1991_46122# 2.75e-20
C22375 a_18599_43230# a_7174_31319# 2.71e-21
C22376 a_19987_42826# a_13258_32519# 2.93e-19
C22377 a_n4318_38680# a_n4064_38528# 0.047936f
C22378 a_n784_42308# a_n1630_35242# 0.063076f
C22379 a_11301_43218# a_5742_30871# 1.38e-19
C22380 a_n1925_46634# a_2107_46812# 1.12874f
C22381 a_n743_46660# a_1123_46634# 0.054493f
C22382 a_n2438_43548# a_383_46660# 0.0336f
C22383 a_171_46873# a_33_46660# 0.207108f
C22384 a_n133_46660# a_601_46902# 0.053479f
C22385 a_n881_46662# a_5429_46660# 3.91e-20
C22386 a_n1613_43370# a_5257_43370# 0.025984f
C22387 a_10227_46804# a_12469_46902# 0.181535f
C22388 a_11599_46634# a_15559_46634# 0.028826f
C22389 a_15811_47375# a_14976_45028# 2.33e-19
C22390 a_12861_44030# a_15227_44166# 0.810382f
C22391 a_6151_47436# a_13885_46660# 0.001762f
C22392 a_13717_47436# a_19333_46634# 1.58e-20
C22393 a_4915_47217# a_14513_46634# 2.71e-19
C22394 a_584_46384# a_765_45546# 0.086068f
C22395 a_14797_45144# a_15095_43370# 1.1e-20
C22396 a_9313_44734# a_10729_43914# 0.001217f
C22397 a_4223_44672# a_6671_43940# 0.03251f
C22398 a_14537_43396# a_14955_43396# 0.027267f
C22399 a_n2293_42834# a_6031_43396# 1.5e-19
C22400 a_n2293_43922# a_3499_42826# 8.88e-21
C22401 a_18494_42460# a_n97_42460# 2.68e-19
C22402 a_22315_44484# a_20512_43084# 0.004063f
C22403 a_3422_30871# a_22485_44484# 0.003365f
C22404 a_13720_44458# a_14021_43940# 8.41e-19
C22405 a_n2661_42834# a_5841_44260# 5.31e-20
C22406 a_n2017_45002# a_743_42282# 7.84646f
C22407 a_n913_45002# a_4190_30871# 0.061913f
C22408 a_19963_31679# a_13887_32519# 0.051213f
C22409 a_7754_40130# VDD 13.6809f
C22410 a_18587_45118# VDD 0.085535f
C22411 a_5742_30871# C2_P_btm 0.030783f
C22412 a_5934_30871# VCM 0.121361f
C22413 a_13213_44734# a_12741_44636# 0.00239f
C22414 a_14112_44734# a_11415_45002# 1.45e-20
C22415 a_19006_44850# a_17339_46660# 1.58e-20
C22416 a_3353_43940# a_n2293_46634# 5.23e-19
C22417 a_1307_43914# a_n755_45592# 0.007948f
C22418 a_1423_45028# a_n863_45724# 0.113534f
C22419 a_16922_45042# a_8049_45260# 8.87e-20
C22420 a_n2661_44458# a_n2956_39304# 1.51e-20
C22421 a_n4318_40392# a_n2956_38680# 0.024261f
C22422 a_375_42282# a_310_45028# 0.078376f
C22423 a_2304_45348# a_n2293_45546# 0.032829f
C22424 a_n2129_43609# a_n881_46662# 1.93e-21
C22425 a_12883_44458# a_10903_43370# 6.65e-20
C22426 a_n2267_43396# a_n1613_43370# 0.04778f
C22427 a_21335_42336# a_21421_42336# 0.006584f
C22428 a_n310_47243# VDD 2.4e-19
C22429 a_5257_43370# a_n2293_46098# 0.049293f
C22430 a_4955_46873# a_1823_45246# 0.001178f
C22431 a_3090_45724# a_16388_46812# 1.08e-19
C22432 a_15368_46634# a_15227_46910# 0.050747f
C22433 a_14976_45028# a_13059_46348# 0.209989f
C22434 a_11901_46660# a_765_45546# 0.007273f
C22435 a_12156_46660# a_12347_46660# 4.61e-19
C22436 a_n881_46662# a_835_46155# 2.99e-19
C22437 a_19321_45002# a_19900_46494# 0.002634f
C22438 a_n743_46660# a_13759_46122# 0.01783f
C22439 a_13661_43548# a_6945_45028# 0.015293f
C22440 a_20916_46384# a_18985_46122# 5.23e-20
C22441 a_2107_46812# a_10355_46116# 7.69e-19
C22442 a_4883_46098# a_10037_46155# 4.58e-19
C22443 a_13507_46334# a_12379_46436# 0.001281f
C22444 a_584_46384# a_509_45822# 3.94e-19
C22445 a_1431_47204# a_1609_45822# 9.46e-22
C22446 a_n443_46116# a_n755_45592# 0.651643f
C22447 a_n1151_42308# a_n356_45724# 4.29e-20
C22448 a_11599_46634# a_20009_46494# 2.17e-19
C22449 a_16327_47482# a_19240_46482# 2.52e-19
C22450 a_17591_47464# a_13259_45724# 3.28e-20
C22451 a_10227_46804# a_14383_46116# 0.01306f
C22452 a_n2661_42282# a_n1917_43396# 4.78e-21
C22453 a_9313_44734# a_21487_43396# 1.21e-19
C22454 a_11967_42832# a_12281_43396# 0.027232f
C22455 a_3499_42826# a_n97_42460# 0.019497f
C22456 a_5891_43370# a_5649_42852# 6.09e-19
C22457 a_1467_44172# a_1512_43396# 2.14e-20
C22458 a_20193_45348# a_19987_42826# 0.008117f
C22459 a_n2017_45002# a_5755_42308# 0.004115f
C22460 a_3065_45002# a_1755_42282# 4.51e-19
C22461 a_n913_45002# a_5337_42558# 0.006397f
C22462 a_13904_45546# a_14033_45572# 0.010132f
C22463 a_10793_43218# a_10227_46804# 2.95e-19
C22464 a_n784_42308# a_n971_45724# 0.006301f
C22465 a_n1630_35242# SMPL_ON_P 6.11548f
C22466 a_1606_42308# w_11334_34010# 0.001329f
C22467 a_17730_32519# a_20692_30879# 0.05146f
C22468 a_9672_43914# a_526_44458# 1.87e-19
C22469 a_18083_42858# a_12549_44172# 5.88e-21
C22470 a_14955_43396# a_3090_45724# 0.07523f
C22471 a_15743_43084# a_6755_46942# 7.96e-20
C22472 a_11415_45002# VDD 1.84504f
C22473 a_n2293_46098# a_1337_46116# 0.002811f
C22474 a_3090_45724# a_3316_45546# 0.04556f
C22475 a_3483_46348# a_10809_44734# 0.02965f
C22476 a_8953_45546# a_2324_44458# 0.047906f
C22477 a_10903_43370# a_12005_46116# 0.277468f
C22478 a_4958_30871# VDAC_N 0.021971f
C22479 a_n3565_39304# a_n4064_37984# 0.028081f
C22480 a_n3420_39072# a_n3420_37984# 0.046468f
C22481 a_15682_43940# a_16795_42852# 7.6e-20
C22482 a_2982_43646# a_15781_43660# 1.65e-20
C22483 a_20974_43370# a_21487_43396# 0.03755f
C22484 a_21381_43940# a_13467_32519# 0.002377f
C22485 a_n2293_43922# a_3318_42354# 4.38e-20
C22486 a_5891_43370# a_7963_42308# 0.036306f
C22487 a_3905_42865# a_5193_42852# 0.001894f
C22488 a_16023_47582# RST_Z 1.03e-19
C22489 a_13717_47436# CLK 0.057477f
C22490 a_16327_47482# START 4.67e-19
C22491 a_11322_45546# a_8975_43940# 2.88e-19
C22492 a_15903_45785# a_11691_44458# 4.76e-21
C22493 a_16855_45546# a_11827_44484# 7.23e-23
C22494 a_2711_45572# a_7640_43914# 3.03e-20
C22495 a_n2017_45002# a_626_44172# 1.24e-20
C22496 a_n913_45002# a_375_42282# 0.01541f
C22497 a_5691_45260# a_5205_44484# 9.01e-20
C22498 a_5111_44636# a_7229_43940# 4.19e-21
C22499 a_3537_45260# a_8953_45002# 2.96e-19
C22500 a_3232_43370# a_6431_45366# 0.005731f
C22501 a_13460_43230# a_3483_46348# 7.53e-19
C22502 a_12895_43230# a_4185_45028# 1.02e-20
C22503 a_743_42282# a_526_44458# 0.042759f
C22504 a_12281_43396# a_13259_45724# 3.97e-20
C22505 a_9127_43156# a_5937_45572# 5.33e-21
C22506 a_8952_43230# a_8199_44636# 1.83e-19
C22507 a_17730_32519# VIN_N 0.048461f
C22508 a_20107_45572# a_10227_46804# 2.37e-20
C22509 a_21188_45572# a_16327_47482# 0.227468f
C22510 a_3357_43084# a_13381_47204# 1.79e-19
C22511 a_2437_43646# a_12861_44030# 0.022753f
C22512 a_413_45260# a_2905_45572# 0.124898f
C22513 a_n143_45144# a_n1151_42308# 0.002247f
C22514 a_2274_45254# a_2063_45854# 2.23e-19
C22515 a_5111_44636# a_n237_47217# 6.91e-20
C22516 a_2382_45260# a_584_46384# 0.185451f
C22517 a_16333_45814# a_n881_46662# 0.04285f
C22518 a_11688_45572# a_12549_44172# 6.24e-20
C22519 a_3775_45552# a_3524_46660# 1.42e-20
C22520 a_2711_45572# a_4651_46660# 5.93e-20
C22521 a_4099_45572# a_3877_44458# 0.01632f
C22522 a_7499_43078# a_2107_46812# 6.63e-20
C22523 a_11652_45724# a_n743_46660# 2.53e-19
C22524 a_n2840_45546# a_n2293_45546# 2.81e-19
C22525 a_n2661_45546# a_n2472_45546# 0.040937f
C22526 a_n2810_45572# a_n2956_38216# 6.20057f
C22527 a_4190_30871# a_20922_43172# 8.66e-20
C22528 a_21259_43561# a_21356_42826# 3.61e-19
C22529 a_5649_42852# a_17595_43084# 9.42e-21
C22530 a_4361_42308# a_17333_42852# 3.75e-20
C22531 a_743_42282# a_19164_43230# 5.07e-20
C22532 a_11341_43940# a_17531_42308# 2.85e-21
C22533 a_19328_44172# a_19511_42282# 2.58e-21
C22534 a_14209_32519# a_5342_30871# 0.028644f
C22535 a_n1557_42282# a_n327_42558# 0.001953f
C22536 a_3080_42308# a_n1630_35242# 0.032975f
C22537 a_1209_43370# a_1606_42308# 1.26e-20
C22538 a_15493_43940# a_4958_30871# 4.56e-21
C22539 a_21076_30879# a_22459_39145# 3.89e-20
C22540 a_14035_46660# CLK 3.17e-20
C22541 a_7754_39964# a_6886_37412# 0.035115f
C22542 VDAC_Pi a_5700_37509# 2.20213f
C22543 a_7754_40130# a_8912_37509# 1.81084f
C22544 a_3754_38470# a_7754_38470# 3.02e-20
C22545 a_n39_42308# VDD 0.00143f
C22546 a_n1605_47204# a_n452_47436# 3.88e-21
C22547 SMPL_ON_P a_n971_45724# 2.75e-21
C22548 a_n1741_47186# a_n746_45260# 0.032595f
C22549 a_n2109_47186# a_n23_47502# 0.043455f
C22550 a_n2288_47178# a_n785_47204# 6.98e-20
C22551 a_1423_45028# a_9313_44734# 0.241551f
C22552 a_11691_44458# a_n2661_44458# 0.021716f
C22553 a_9482_43914# a_13468_44734# 0.00165f
C22554 a_11823_42460# a_12603_44260# 2.91e-20
C22555 a_6171_45002# a_14673_44172# 6.91e-20
C22556 a_19479_31679# a_22959_44484# 0.001721f
C22557 a_11633_42308# a_9290_44172# 0.001629f
C22558 a_13291_42460# a_n357_42282# 0.008613f
C22559 a_5755_42308# a_526_44458# 3.22e-19
C22560 a_9145_43396# CLK 2.67e-21
C22561 a_n2302_37984# a_n2312_38680# 1.26e-19
C22562 a_19778_44110# a_20916_46384# 2.1e-21
C22563 a_10775_45002# a_6755_46942# 6.89e-22
C22564 a_10951_45334# a_10249_46116# 8.11e-22
C22565 a_11827_44484# a_13661_43548# 0.120515f
C22566 a_21005_45260# a_19321_45002# 0.002433f
C22567 a_21359_45002# a_13747_46662# 0.060042f
C22568 a_5365_45348# a_3877_44458# 6.25e-22
C22569 a_2437_43646# a_14180_46812# 1.36e-20
C22570 a_413_45260# a_12816_46660# 4.83e-21
C22571 a_5111_44636# a_8270_45546# 0.035253f
C22572 a_n913_45002# a_15227_44166# 1.05e-19
C22573 a_n2129_44697# a_n881_46662# 1.78e-19
C22574 a_10490_45724# a_10903_43370# 0.057318f
C22575 a_11652_45724# a_11189_46129# 0.00549f
C22576 a_6667_45809# a_6945_45028# 0.015851f
C22577 a_10193_42453# a_12594_46348# 1.09e-19
C22578 a_11322_45546# a_11387_46155# 4.47e-19
C22579 a_n2267_44484# a_n1613_43370# 0.025052f
C22580 a_8975_43940# a_12465_44636# 3.06e-19
C22581 a_n2293_43922# a_n1151_42308# 1.39e-19
C22582 a_13467_32519# a_21125_42558# 1.91e-19
C22583 a_4361_42308# a_18997_42308# 1.34e-19
C22584 a_10796_42968# a_5742_30871# 0.003276f
C22585 a_10835_43094# a_11551_42558# 4.09e-19
C22586 a_10341_42308# a_10533_42308# 0.035479f
C22587 a_10922_42852# a_10723_42308# 0.001007f
C22588 a_10991_42826# a_11323_42473# 1.78e-19
C22589 a_5649_42852# a_21887_42336# 0.017243f
C22590 a_13678_32519# a_21613_42308# 0.024855f
C22591 a_13887_32519# a_7174_31319# 0.003259f
C22592 a_12891_46348# a_768_44030# 0.193145f
C22593 a_n1613_43370# a_5807_45002# 0.086053f
C22594 a_n2312_39304# a_n2293_46634# 0.021162f
C22595 a_2063_45854# a_10467_46802# 0.036614f
C22596 a_n971_45724# a_8035_47026# 8.58e-19
C22597 a_n1151_42308# a_8667_46634# 1.5e-19
C22598 a_4791_45118# a_5257_43370# 0.36404f
C22599 a_18911_45144# a_15493_43940# 2.89e-20
C22600 a_18184_42460# a_11341_43940# 0.029749f
C22601 a_n356_44636# a_n809_44244# 0.00336f
C22602 a_n2661_44458# a_8333_44056# 4.4e-20
C22603 a_11691_44458# a_18451_43940# 0.001358f
C22604 a_11827_44484# a_19862_44208# 0.015537f
C22605 a_7499_43078# a_7871_42858# 0.146369f
C22606 a_742_44458# a_3499_42826# 4.13e-19
C22607 a_2711_45572# a_16414_43172# 3.78e-19
C22608 a_16147_45260# a_17499_43370# 5.95e-20
C22609 a_3537_45260# a_3626_43646# 0.002395f
C22610 C6_N_btm VDD 0.210613f
C22611 a_13159_45002# VDD 0.321035f
C22612 COMP_P a_21589_35634# 7.17e-19
C22613 a_n784_42308# a_11530_34132# 0.006009f
C22614 a_n1630_35242# a_n1532_35090# 0.462421f
C22615 a_14485_44260# a_12465_44636# 0.009374f
C22616 a_n97_42460# a_n1151_42308# 8.22e-19
C22617 a_n2661_45010# a_n2840_45546# 3.35e-19
C22618 a_n2840_45002# a_n2810_45572# 4.88e-19
C22619 a_626_44172# a_526_44458# 0.180416f
C22620 a_10775_45002# a_8049_45260# 7.17e-20
C22621 a_16789_44484# a_6755_46942# 2.63e-19
C22622 a_12429_44172# a_12549_44172# 0.137881f
C22623 a_11750_44172# a_768_44030# 0.00229f
C22624 a_18374_44850# a_17339_46660# 0.009147f
C22625 a_n2661_42834# a_3090_45724# 0.164804f
C22626 a_18248_44752# a_18285_46348# 3.14e-21
C22627 a_13483_43940# a_12891_46348# 0.062818f
C22628 a_n2129_44697# a_n2157_46122# 8.63e-21
C22629 a_n2267_44484# a_n2293_46098# 2.71e-20
C22630 a_11827_44484# a_4185_45028# 0.03083f
C22631 a_n2661_44458# a_n1991_46122# 1.24e-22
C22632 a_2553_47502# VDD 0.150286f
C22633 a_15959_42545# a_15890_42674# 0.209641f
C22634 a_8515_42308# a_7174_31319# 4.88e-21
C22635 a_n3674_38216# a_n4334_38528# 2.59e-19
C22636 a_n3674_38680# a_n2946_38778# 4.03e-21
C22637 a_5742_30871# a_4958_30871# 0.032374f
C22638 a_21588_30879# a_22591_46660# 5.88e-20
C22639 a_5807_45002# a_n2293_46098# 2.61e-20
C22640 a_20916_46384# a_20820_30879# 4.91e-20
C22641 a_22612_30879# a_11415_45002# 1.26e-21
C22642 a_10249_46116# a_11735_46660# 7.95e-19
C22643 a_6755_46942# a_11186_47026# 0.014167f
C22644 a_n743_46660# a_16434_46660# 6.95e-19
C22645 a_n881_46662# a_3483_46348# 0.5947f
C22646 a_n1613_43370# a_3699_46348# 2.1e-19
C22647 a_6151_47436# a_526_44458# 3.76e-20
C22648 a_4883_46098# a_12005_46116# 0.012933f
C22649 a_13507_46334# a_13351_46090# 0.214666f
C22650 a_16327_47482# a_19553_46090# 0.172776f
C22651 a_14955_47212# a_6945_45028# 0.013254f
C22652 a_10227_46804# a_17715_44484# 1.63e-20
C22653 a_13487_47204# a_10809_44734# 1.49e-19
C22654 a_2063_45854# a_8034_45724# 0.034258f
C22655 a_n1741_47186# a_12379_46436# 0.067348f
C22656 a_5891_43370# a_8685_43396# 0.145735f
C22657 a_2998_44172# a_2455_43940# 1.95e-19
C22658 a_n2661_43922# a_6765_43638# 4.58e-22
C22659 a_n2661_42834# a_6547_43396# 2.31e-19
C22660 a_14539_43914# a_15781_43660# 1.8e-20
C22661 a_11823_42460# a_13657_42558# 0.009593f
C22662 a_n356_44636# a_14955_43396# 5.49e-21
C22663 a_13249_42308# a_13070_42354# 0.141799f
C22664 a_2711_45572# a_7174_31319# 0.008877f
C22665 a_3422_30871# a_14401_32519# 0.096501f
C22666 a_2889_44172# a_3052_44056# 0.004767f
C22667 a_2675_43914# a_3353_43940# 0.011812f
C22668 a_20512_43084# a_19319_43548# 1.25e-19
C22669 a_5147_45002# a_5193_42852# 4.91e-21
C22670 a_n913_45002# a_14635_42282# 0.332583f
C22671 a_n1059_45260# a_15785_43172# 3.54e-19
C22672 a_11967_42832# VDD 2.67441f
C22673 a_10193_42453# a_11322_45546# 0.024616f
C22674 a_8746_45002# a_10490_45724# 0.116339f
C22675 a_2711_45572# a_10306_45572# 7.5e-19
C22676 a_11341_43940# a_12741_44636# 9.61e-20
C22677 a_17538_32519# a_19692_46634# 0.002f
C22678 a_21855_43396# a_12549_44172# 0.001702f
C22679 a_14112_44734# a_13259_45724# 0.001601f
C22680 a_895_43940# a_2324_44458# 0.011941f
C22681 a_n2472_42826# a_n1613_43370# 6.43e-21
C22682 a_10083_42826# a_10227_46804# 0.292997f
C22683 a_12251_46660# VDD 0.195617f
C22684 a_n3565_39304# C0_P_btm 9.35e-21
C22685 a_5934_30871# VDAC_Ni 3.94e-19
C22686 a_6123_31319# a_3754_38470# 2.11e-19
C22687 a_n2293_46098# a_3699_46348# 3.53e-20
C22688 a_376_46348# a_1823_45246# 9.94e-21
C22689 a_472_46348# a_1138_42852# 0.028956f
C22690 a_805_46414# a_1176_45822# 0.024739f
C22691 a_8270_45546# a_8379_46155# 8.95e-21
C22692 a_3090_45724# a_5066_45546# 1.9e-19
C22693 a_17339_46660# a_17715_44484# 0.018672f
C22694 a_765_45546# a_17583_46090# 0.067337f
C22695 a_14513_46634# a_10809_44734# 0.002278f
C22696 a_9313_44734# a_17141_43172# 1.4e-19
C22697 a_18079_43940# a_743_42282# 3.93e-21
C22698 a_18451_43940# a_4190_30871# 3.13e-19
C22699 a_n97_42460# a_6197_43396# 0.003645f
C22700 a_14021_43940# a_16977_43638# 0.005856f
C22701 a_n2661_42282# a_n1853_43023# 4.23e-20
C22702 a_5013_44260# a_5111_42852# 2.02e-21
C22703 a_3422_30871# a_18817_42826# 1.01e-20
C22704 a_15493_43396# a_19177_43646# 0.001461f
C22705 a_1756_43548# a_2982_43646# 7.54e-20
C22706 a_13565_43940# a_9145_43396# 0.001581f
C22707 a_n2810_45028# a_n3565_38216# 0.349341f
C22708 a_648_43396# VDD 9.68e-19
C22709 a_15765_45572# a_16751_45260# 8.52e-20
C22710 a_11823_42460# a_n2661_43370# 0.006541f
C22711 a_8696_44636# a_14797_45144# 7.63e-21
C22712 a_16333_45814# a_1307_43914# 6.14e-21
C22713 a_15861_45028# a_14537_43396# 2.27e-20
C22714 a_17531_42308# a_16327_47482# 7.43e-19
C22715 a_15761_42308# a_10227_46804# 2.95e-19
C22716 a_9223_42460# a_n1613_43370# 0.007135f
C22717 a_2813_43396# a_526_44458# 0.013054f
C22718 a_17538_32519# a_20692_30879# 0.05141f
C22719 a_n1630_35242# a_n2438_43548# 1.24e-19
C22720 a_13259_45724# VDD 2.41738f
C22721 a_6472_45840# a_n881_46662# 0.179318f
C22722 a_6511_45714# a_n1613_43370# 0.017587f
C22723 a_7499_43078# a_11453_44696# 0.02227f
C22724 a_10490_45724# a_4883_46098# 7.84e-20
C22725 a_14495_45572# a_10227_46804# 0.001891f
C22726 a_8049_45260# a_12839_46116# 0.004724f
C22727 a_8333_44056# a_8325_42308# 1.23e-22
C22728 a_13667_43396# a_13635_43156# 0.006368f
C22729 a_4361_42308# a_13678_32519# 0.048617f
C22730 a_21259_43561# a_20749_43396# 7.22e-19
C22731 a_9145_43396# a_5534_30871# 2.86e-19
C22732 a_20512_43084# a_21335_42336# 1.26e-21
C22733 a_13467_32519# a_5649_42852# 0.042596f
C22734 a_4190_30871# a_17364_32525# 1.46e-20
C22735 a_3080_42308# a_3863_42891# 9.93e-20
C22736 a_3422_30871# a_21421_42336# 5.28e-19
C22737 VDAC_N C7_N_btm 0.11042p
C22738 a_5257_43370# DATA[3] 9.23e-21
C22739 a_9114_42852# VDD 4.6e-19
C22740 a_18175_45572# a_17517_44484# 1.07e-20
C22741 a_375_42282# a_n2661_44458# 0.025194f
C22742 a_8191_45002# a_5883_43914# 4.94e-22
C22743 a_8953_45002# a_8701_44490# 0.005993f
C22744 a_6171_45002# a_12607_44458# 5.85e-20
C22745 a_3232_43370# a_12883_44458# 1.44e-20
C22746 a_9127_43156# a_n443_42852# 0.001064f
C22747 a_13460_43230# a_n357_42282# 0.007447f
C22748 a_3080_42308# a_11530_34132# 0.001927f
C22749 a_14401_32519# VREF_GND 0.066097f
C22750 a_17538_32519# VIN_N 0.041176f
C22751 a_14309_45348# a_12465_44636# 1.46e-20
C22752 a_18184_42460# a_16327_47482# 0.168018f
C22753 a_19113_45348# a_12861_44030# 0.003723f
C22754 C4_P_btm VDD 0.265463f
C22755 a_2779_44458# a_2905_45572# 7.14e-20
C22756 a_4743_44484# a_2063_45854# 3.42e-21
C22757 a_1667_45002# a_1799_45572# 1.16e-19
C22758 a_8953_45002# a_n2293_46634# 4.11e-20
C22759 a_4558_45348# a_2107_46812# 1.43e-21
C22760 a_327_44734# a_n2661_46098# 1.48e-20
C22761 a_413_45260# a_2443_46660# 0.020902f
C22762 a_2809_45348# a_768_44030# 0.001559f
C22763 a_16680_45572# a_15368_46634# 2.35e-20
C22764 a_8696_44636# a_14976_45028# 2.84e-19
C22765 a_11787_45002# a_n2661_46634# 0.004953f
C22766 a_15595_45028# a_13661_43548# 0.214904f
C22767 a_15415_45028# a_13747_46662# 2.47e-20
C22768 a_15861_45028# a_3090_45724# 0.125763f
C22769 a_15903_45785# a_15227_44166# 0.005114f
C22770 a_6511_45714# a_n2293_46098# 7.32e-20
C22771 a_743_42282# a_4169_42308# 4.3e-19
C22772 a_16409_43396# a_15803_42450# 9.67e-20
C22773 a_4520_42826# a_n784_42308# 4.32e-21
C22774 a_4361_42308# a_6123_31319# 0.065399f
C22775 a_16243_43396# a_15890_42674# 1.41e-20
C22776 a_13887_32519# a_5932_42308# 0.003117f
C22777 a_18249_42858# a_18695_43230# 2.28e-19
C22778 a_n2946_38778# VDD 0.383009f
C22779 a_6151_47436# a_13759_47204# 0.00136f
C22780 a_11031_47542# a_11117_47542# 0.006584f
C22781 a_9313_45822# a_10037_47542# 0.00168f
C22782 a_13487_47204# a_n881_46662# 0.108977f
C22783 a_4791_45118# a_5807_45002# 0.129041f
C22784 a_n2109_47186# a_948_46660# 5.02e-20
C22785 a_n1741_47186# a_383_46660# 4.76e-20
C22786 a_n23_47502# a_n1925_46634# 4.04e-20
C22787 a_n746_45260# a_n743_46660# 0.068305f
C22788 a_n971_45724# a_n2438_43548# 0.038673f
C22789 a_2124_47436# a_n2661_46634# 1.6e-20
C22790 a_13507_46334# a_22223_47212# 0.001502f
C22791 a_20894_47436# a_11453_44696# 7.99e-20
C22792 a_21496_47436# a_12465_44636# 2.84e-19
C22793 a_4883_46098# a_21811_47423# 0.054014f
C22794 a_10951_45334# a_10555_44260# 5.79e-20
C22795 a_n356_44636# a_n2661_42834# 0.024765f
C22796 a_13556_45296# a_11341_43940# 0.001133f
C22797 a_11823_42460# a_15681_43442# 6.78e-20
C22798 a_10193_42453# a_16409_43396# 2.72e-19
C22799 a_12607_44458# a_14673_44172# 2.97e-21
C22800 a_1307_43914# a_15493_43396# 2.1e-19
C22801 a_18114_32519# a_21398_44850# 4.06e-20
C22802 a_n1655_44484# a_n2661_43922# 6.56e-19
C22803 a_19963_31679# a_14401_32519# 0.053905f
C22804 a_3065_45002# a_3737_43940# 0.005754f
C22805 a_22465_38105# a_20692_30879# 5.07e-19
C22806 a_20273_45572# VDD 0.571099f
C22807 a_1307_43914# a_3483_46348# 0.095243f
C22808 a_1145_45348# a_167_45260# 5.7e-19
C22809 a_17719_45144# a_17339_46660# 8.89e-19
C22810 a_11691_44458# a_14035_46660# 4.42e-21
C22811 a_17613_45144# a_765_45546# 1.04e-21
C22812 a_19279_43940# a_13747_46662# 0.048937f
C22813 a_20835_44721# a_19321_45002# 7.19e-19
C22814 a_19721_31679# a_19692_46634# 5.55e-20
C22815 a_16922_45042# a_18285_46348# 4.22e-21
C22816 a_20637_44484# a_12549_44172# 8.68e-20
C22817 a_16223_45938# a_16375_45002# 3.86e-20
C22818 a_n2017_45002# a_n2956_38680# 7.75e-22
C22819 a_11787_45002# a_8199_44636# 2.96e-20
C22820 a_n2065_43946# a_n1613_43370# 0.30437f
C22821 a_6171_45002# a_10903_43370# 0.041534f
C22822 a_8953_45002# a_9625_46129# 0.004507f
C22823 a_413_45260# a_18819_46122# 1.56e-20
C22824 a_3065_45002# a_2324_44458# 0.017588f
C22825 a_6761_42308# a_6123_31319# 0.187371f
C22826 a_1606_42308# a_14456_42282# 3.31e-20
C22827 a_n923_35174# a_n83_35174# 0.480251f
C22828 a_13661_43548# a_15559_46634# 8.86e-22
C22829 a_13747_46662# a_15368_46634# 0.110984f
C22830 a_n2661_46634# a_11813_46116# 0.162517f
C22831 a_5807_45002# a_16292_46812# 0.202526f
C22832 a_4651_46660# a_6540_46812# 7.72e-21
C22833 a_5385_46902# a_5167_46660# 0.209641f
C22834 a_4817_46660# a_5907_46634# 0.042415f
C22835 a_19321_45002# a_3090_45724# 0.163821f
C22836 a_4646_46812# a_5072_46660# 0.013764f
C22837 a_n881_46662# a_14513_46634# 0.017832f
C22838 a_11453_44696# a_20411_46873# 0.020751f
C22839 a_12465_44636# a_21363_46634# 5.44e-20
C22840 a_4883_46098# a_22000_46634# 0.004514f
C22841 a_16327_47482# a_12741_44636# 0.074082f
C22842 a_13507_46334# a_20731_47026# 8.28e-19
C22843 a_2063_45854# a_8016_46348# 8.48e-19
C22844 a_n1151_42308# a_5204_45822# 0.487224f
C22845 a_n1741_47186# a_13351_46090# 7.57e-20
C22846 a_n443_46116# a_3483_46348# 0.009289f
C22847 a_18479_47436# a_20719_46660# 8e-19
C22848 a_n1435_47204# a_n1423_46090# 2.49e-19
C22849 a_10227_46804# a_22365_46825# 2.64e-20
C22850 a_19615_44636# a_15493_43940# 4.39e-21
C22851 a_20835_44721# a_20623_43914# 2.27e-19
C22852 a_20640_44752# a_21115_43940# 7.54e-19
C22853 a_11691_44458# a_9145_43396# 4.24e-19
C22854 a_5663_43940# a_6453_43914# 0.017005f
C22855 a_18579_44172# a_15493_43396# 0.070538f
C22856 a_19279_43940# a_20269_44172# 0.002186f
C22857 a_20679_44626# a_20935_43940# 7.96e-20
C22858 a_n699_43396# a_648_43396# 3.48e-19
C22859 a_11827_44484# a_14579_43548# 9.5e-23
C22860 a_18184_42460# a_10341_43396# 0.034231f
C22861 a_1115_44172# a_1525_44260# 0.007617f
C22862 a_453_43940# a_261_44278# 5.76e-19
C22863 a_5495_43940# a_7281_43914# 1.28e-20
C22864 a_14673_44172# a_14761_44260# 1.45e-19
C22865 a_n2661_42834# a_9165_43940# 3.03e-20
C22866 a_3232_43370# a_3935_42891# 2.51e-20
C22867 a_5111_44636# a_5755_42852# 0.002818f
C22868 a_3537_45260# a_8037_42858# 0.010068f
C22869 a_n913_45002# a_14543_43071# 0.036401f
C22870 a_n1059_45260# a_5534_30871# 0.025423f
C22871 a_n2017_45002# a_15279_43071# 0.002198f
C22872 a_18989_43940# VDD 0.342796f
C22873 a_n4064_39616# C2_P_btm 4.56e-20
C22874 a_16664_43396# a_10227_46804# 5.15e-19
C22875 a_21259_43561# a_12861_44030# 3.06e-20
C22876 a_n901_43156# a_n1151_42308# 0.01984f
C22877 a_19721_31679# a_20692_30879# 0.051673f
C22878 a_20623_43914# a_3090_45724# 4.66e-20
C22879 a_3626_43646# a_n2293_46634# 0.012347f
C22880 a_18579_44172# a_3483_46348# 2.2e-21
C22881 a_1343_38525# a_2112_39137# 0.22564f
C22882 a_n4064_39072# a_n4251_39392# 4.37e-19
C22883 a_n4209_39304# a_n2216_39072# 0.001412f
C22884 a_1799_45572# VDD 0.381212f
C22885 a_5742_30871# C7_N_btm 0.04157f
C22886 a_21188_46660# a_22000_46634# 2.08e-19
C22887 a_20623_46660# a_20731_47026# 0.057222f
C22888 a_19123_46287# a_19636_46660# 1.03e-19
C22889 a_n743_46660# a_12379_46436# 1.32e-19
C22890 a_2107_46812# a_10044_46482# 2.82e-19
C22891 a_n881_46662# a_n357_42282# 7.4e-19
C22892 a_6755_46942# a_14840_46494# 0.021842f
C22893 a_8270_45546# a_9290_44172# 0.433963f
C22894 a_5257_43370# a_6945_45028# 6.65e-21
C22895 a_n1613_43370# a_n755_45592# 0.052236f
C22896 a_3422_30871# a_22223_43396# 2.47e-20
C22897 a_10807_43548# a_8685_43396# 0.029811f
C22898 a_n2293_43922# a_10922_42852# 1.19e-20
C22899 a_9313_44734# a_15567_42826# 0.01457f
C22900 a_18184_42460# a_20356_42852# 0.008384f
C22901 a_n356_44636# a_n2293_42282# 1.10197f
C22902 a_18494_42460# a_20256_42852# 0.001548f
C22903 a_20512_43084# a_19095_43396# 1.93e-19
C22904 a_n913_45002# a_19511_42282# 0.120073f
C22905 a_n1059_45260# a_19647_42308# 2.95e-20
C22906 a_5745_43940# VDD 0.144352f
C22907 a_18175_45572# a_19256_45572# 0.102355f
C22908 a_18341_45572# a_18691_45572# 0.206455f
C22909 a_18479_45785# a_19431_45546# 0.009466f
C22910 a_2711_45572# a_1423_45028# 6.59e-21
C22911 a_16147_45260# a_18596_45572# 9.29e-20
C22912 a_8746_45002# a_6171_45002# 0.069475f
C22913 a_8162_45546# a_8191_45002# 0.003007f
C22914 a_9049_44484# a_7229_43940# 4.55e-21
C22915 a_10490_45724# a_3232_43370# 9.93e-20
C22916 a_n4209_37414# VREF_GND 0.00198f
C22917 a_10341_43396# a_12741_44636# 4.16e-20
C22918 a_22591_43396# a_19692_46634# 2.85e-19
C22919 a_3499_42826# a_3503_45724# 9.02e-22
C22920 a_11341_43940# a_16375_45002# 4.26e-20
C22921 a_5700_37509# RST_Z 0.051902f
C22922 a_n1736_42282# a_n2312_39304# 3.28e-20
C22923 a_n4318_37592# a_n2312_40392# 0.025292f
C22924 VDAC_P C5_P_btm 27.6071f
C22925 a_18114_32519# VREF 1.12e-19
C22926 a_19721_31679# VIN_N 0.029175f
C22927 a_18189_46348# VDD 0.211855f
C22928 a_6194_45824# a_4915_47217# 1.57e-22
C22929 a_2711_45572# a_6491_46660# 1.46e-21
C22930 a_6511_45714# a_4791_45118# 0.034343f
C22931 a_9049_44484# a_n237_47217# 0.001811f
C22932 a_3775_45552# a_3785_47178# 7.52e-20
C22933 a_n3420_38528# VDAC_P 2.69e-19
C22934 a_n2293_46098# a_n755_45592# 0.086057f
C22935 a_1208_46090# a_n2661_45546# 4.43e-20
C22936 a_n1076_46494# a_n1079_45724# 8.64e-19
C22937 a_376_46348# a_n2293_45546# 1.03e-21
C22938 a_n901_46420# a_n863_45724# 0.00998f
C22939 a_n1991_46122# a_n1099_45572# 5.38e-19
C22940 a_n2956_39304# a_n1925_42282# 5.53e-20
C22941 a_14840_46494# a_8049_45260# 0.002948f
C22942 a_11189_46129# a_12379_46436# 1.91e-20
C22943 a_n3565_38216# a_n2302_37690# 0.002384f
C22944 a_20843_47204# START 1.11e-19
C22945 a_5807_45002# DATA[3] 4.68e-21
C22946 a_2479_44172# a_1755_42282# 6.04e-21
C22947 a_3080_42308# a_4520_42826# 4.7e-19
C22948 a_16243_43396# a_16547_43609# 0.165289f
C22949 a_16137_43396# a_16409_43396# 0.011989f
C22950 a_19319_43548# a_18249_42858# 7.61e-19
C22951 a_n97_42460# a_10922_42852# 3.12e-20
C22952 a_11967_42832# a_11551_42558# 6.75e-19
C22953 a_9313_44734# a_20712_42282# 6.9e-20
C22954 a_3422_30871# a_5934_30871# 0.02193f
C22955 a_10341_43396# a_15868_43402# 7.33e-20
C22956 a_10518_42984# VDD 0.273357f
C22957 a_10193_42453# a_16241_44734# 8.94e-19
C22958 a_7705_45326# a_n2661_43370# 0.00431f
C22959 a_n2017_45002# a_20193_45348# 1.2e-20
C22960 a_2437_43646# a_n2661_44458# 0.036499f
C22961 a_n1059_45260# a_11691_44458# 4.15e-20
C22962 a_6171_45002# a_14403_45348# 3.44e-19
C22963 a_3357_43084# a_19721_31679# 5.18e-19
C22964 a_9061_43230# a_8953_45546# 3.71e-19
C22965 a_14209_32519# a_20205_31679# 0.051418f
C22966 a_2113_38308# w_1575_34946# 6.01e-20
C22967 a_9049_44484# a_8270_45546# 0.006099f
C22968 a_13163_45724# a_6755_46942# 6.64e-21
C22969 a_3775_45552# a_3090_45724# 0.001359f
C22970 a_20623_45572# a_20916_46384# 0.006579f
C22971 a_2437_43646# a_16697_47582# 1.94e-19
C22972 a_n745_45366# a_n881_46662# 0.152998f
C22973 a_15415_45028# a_11599_46634# 0.013635f
C22974 a_6171_45002# a_4883_46098# 0.020043f
C22975 a_11963_45334# a_10227_46804# 7.17e-21
C22976 a_1423_45028# a_9313_45822# 1.31e-20
C22977 a_17595_43084# a_17333_42852# 0.057438f
C22978 a_21381_43940# a_21335_42336# 0.002309f
C22979 a_n97_42460# a_17531_42308# 1.1e-21
C22980 a_5755_42852# a_5837_43172# 0.003935f
C22981 a_17701_42308# a_18083_42858# 2.35e-19
C22982 a_4190_30871# a_19273_43230# 5.82e-21
C22983 a_4185_45028# DATA[2] 0.002615f
C22984 a_5815_47464# a_n1435_47204# 0.001005f
C22985 a_4915_47217# a_12861_44030# 0.025257f
C22986 a_6151_47436# a_13381_47204# 0.014822f
C22987 a_n2833_47464# a_n2312_40392# 0.064992f
C22988 a_n1352_44484# a_n356_44636# 0.003615f
C22989 a_n2267_44484# a_n1243_44484# 2.36e-20
C22990 a_n2661_44458# a_4181_44734# 5.47e-19
C22991 a_6171_45002# a_5663_43940# 7.76e-21
C22992 a_5205_44484# a_5013_44260# 4e-20
C22993 a_3232_43370# a_6453_43914# 0.001417f
C22994 a_5111_44636# a_7845_44172# 0.063408f
C22995 en_comp a_n2661_42282# 0.103098f
C22996 a_1755_42282# a_n443_42852# 0.055323f
C22997 a_3905_42558# a_n755_45592# 4.35e-20
C22998 a_n4315_30879# a_n2956_39304# 0.024812f
C22999 a_15143_45578# VDD 0.12071f
C23000 a_13887_32519# VREF 3.68e-19
C23001 a_13940_44484# a_12465_44636# 1.26e-19
C23002 a_20362_44736# a_16327_47482# 0.213851f
C23003 a_18681_44484# a_12861_44030# 1.24e-19
C23004 a_n984_44318# a_n1151_42308# 0.009157f
C23005 a_453_43940# a_584_46384# 0.125447f
C23006 a_n1644_44306# a_n2497_47436# 0.008707f
C23007 a_14033_45572# a_2324_44458# 6.09e-19
C23008 a_8697_45822# a_5066_45546# 0.033513f
C23009 a_13163_45724# a_8049_45260# 0.008063f
C23010 a_11525_45546# a_10586_45546# 0.115475f
C23011 a_9838_44484# a_2107_46812# 5.07e-20
C23012 a_5891_43370# a_768_44030# 0.050862f
C23013 a_n913_45002# a_n1853_46287# 1.34e-20
C23014 a_n1059_45260# a_n1991_46122# 3.7e-20
C23015 a_413_45260# a_22591_46660# 1.37e-20
C23016 a_n2661_45010# a_376_46348# 7.98e-23
C23017 a_14537_43396# a_13059_46348# 0.30244f
C23018 a_18817_42826# a_7174_31319# 8.9e-21
C23019 a_20922_43172# a_19511_42282# 2.35e-19
C23020 a_196_42282# a_n1630_35242# 0.032791f
C23021 a_n784_42308# a_564_42282# 0.003938f
C23022 a_n327_42558# a_n3674_37592# 3.94e-19
C23023 a_11229_43218# a_5742_30871# 8.46e-20
C23024 a_n4318_38680# a_n2946_38778# 3.13e-20
C23025 a_n1925_46634# a_948_46660# 0.006613f
C23026 a_n743_46660# a_383_46660# 0.035839f
C23027 a_n2438_43548# a_601_46902# 0.043115f
C23028 a_n133_46660# a_33_46660# 0.580914f
C23029 a_n2661_46634# a_1110_47026# 1.44e-19
C23030 a_n881_46662# a_5263_46660# 2.48e-19
C23031 a_n1613_43370# a_5429_46660# 0.001925f
C23032 a_10227_46804# a_11901_46660# 0.055248f
C23033 a_11599_46634# a_15368_46634# 0.320705f
C23034 a_15811_47375# a_3090_45724# 1.43e-19
C23035 a_4915_47217# a_14180_46812# 0.017902f
C23036 a_13717_47436# a_15227_44166# 2.25e-20
C23037 a_12861_44030# a_18834_46812# 4.27e-19
C23038 a_2124_47436# a_765_45546# 0.003536f
C23039 a_3422_30871# a_20512_43084# 0.125955f
C23040 a_9313_44734# a_10405_44172# 0.009407f
C23041 a_14537_43396# a_15095_43370# 0.019641f
C23042 a_1307_43914# a_10695_43548# 6.81e-19
C23043 a_n2661_43922# a_3499_42826# 0.001904f
C23044 a_4223_44672# a_5829_43940# 0.037008f
C23045 a_18184_42460# a_n97_42460# 4.22e-19
C23046 a_n2661_42834# a_3820_44260# 5.39e-19
C23047 a_n913_45002# a_21259_43561# 1.9e-20
C23048 a_n1059_45260# a_4190_30871# 0.133926f
C23049 en_comp a_16823_43084# 6.51e-22
C23050 a_19479_31679# a_14209_32519# 0.051176f
C23051 a_20447_31679# a_13678_32519# 0.051589f
C23052 a_6171_45002# a_16243_43396# 1.07e-19
C23053 a_18315_45260# VDD 0.12623f
C23054 a_5742_30871# C3_P_btm 0.030866f
C23055 a_5934_30871# VREF_GND 0.002663f
C23056 a_n2293_43922# a_12741_44636# 0.114756f
C23057 a_13857_44734# a_11415_45002# 1.47e-20
C23058 a_18588_44850# a_17339_46660# 0.00201f
C23059 a_19478_44056# a_12549_44172# 2.21e-20
C23060 a_375_42282# a_n1099_45572# 8.14e-19
C23061 a_1307_43914# a_n357_42282# 0.044512f
C23062 a_2232_45348# a_n2293_45546# 0.004093f
C23063 a_n4318_40392# a_n2956_39304# 0.023379f
C23064 a_1145_45348# a_n863_45724# 4.99e-20
C23065 a_2903_45348# a_n2661_45546# 4.28e-19
C23066 a_12607_44458# a_10903_43370# 0.004073f
C23067 a_6298_44484# a_2324_44458# 0.315008f
C23068 a_n2129_43609# a_n1613_43370# 0.44294f
C23069 a_3626_43646# a_18597_46090# 1.01e-19
C23070 a_6511_45714# DATA[3] 1.62e-21
C23071 a_21613_42308# a_22775_42308# 0.225363f
C23072 a_5742_30871# a_n4064_38528# 0.005505f
C23073 a_2747_46873# VDD 0.626468f
C23074 a_3877_44458# a_167_45260# 5.06e-20
C23075 a_4651_46660# a_1823_45246# 0.001115f
C23076 a_14976_45028# a_15227_46910# 0.060892f
C23077 a_3090_45724# a_13059_46348# 0.167043f
C23078 a_15009_46634# a_16388_46812# 3.35e-20
C23079 a_11813_46116# a_765_45546# 0.003083f
C23080 a_n881_46662# a_518_46155# 3.47e-19
C23081 a_13747_46662# a_20708_46348# 2.93e-21
C23082 a_19321_45002# a_20075_46420# 9.9e-20
C23083 a_20916_46384# a_18819_46122# 7.33e-21
C23084 a_2107_46812# a_9823_46155# 0.002289f
C23085 a_n743_46660# a_13351_46090# 0.008315f
C23086 a_19594_46812# a_19335_46494# 2.8e-19
C23087 a_5807_45002# a_6945_45028# 0.057813f
C23088 a_5534_30871# a_n3420_37440# 0.04166f
C23089 a_4791_45118# a_n755_45592# 0.001705f
C23090 a_n443_46116# a_n357_42282# 0.153614f
C23091 a_10227_46804# a_15194_46482# 0.002224f
C23092 a_16327_47482# a_16375_45002# 0.032962f
C23093 a_13507_46334# a_12005_46436# 7.68e-21
C23094 a_4883_46098# a_9751_46155# 3.69e-19
C23095 a_2998_44172# a_2982_43646# 7.48e-19
C23096 a_5883_43914# a_7765_42852# 2.76e-21
C23097 a_11827_44484# a_21671_42860# 3.44e-21
C23098 a_8701_44490# a_8037_42858# 1.63e-21
C23099 a_20193_45348# a_19164_43230# 3.76e-21
C23100 a_16241_44734# a_16137_43396# 7.77e-20
C23101 a_3065_45002# a_1606_42308# 1.43e-20
C23102 a_n913_45002# a_4921_42308# 0.169235f
C23103 a_n2017_45002# a_5421_42558# 0.001147f
C23104 a_n822_43940# VDD 5.19e-19
C23105 a_10193_42453# a_18691_45572# 6.6e-21
C23106 a_10553_43218# a_10227_46804# 0.001965f
C23107 a_1606_42308# w_1575_34946# 0.001337f
C23108 a_17730_32519# a_20205_31679# 0.051307f
C23109 a_18579_44172# a_n357_42282# 2.1e-19
C23110 a_9028_43914# a_526_44458# 3.93e-21
C23111 a_17701_42308# a_12549_44172# 3.43e-21
C23112 a_8037_42858# a_n2293_46634# 1.56e-20
C23113 a_14205_43396# a_14976_45028# 4.75e-21
C23114 a_15095_43370# a_3090_45724# 0.00771f
C23115 a_9145_43396# a_15227_44166# 0.001689f
C23116 a_n97_42460# a_12741_44636# 3.68e-21
C23117 a_20202_43084# VDD 0.987622f
C23118 a_n4209_39304# a_n2302_37984# 1.04e-19
C23119 a_17124_42282# CAL_N 0.001755f
C23120 a_n2293_46098# a_835_46155# 2.73e-19
C23121 a_3090_45724# a_3218_45724# 0.100752f
C23122 a_13059_46348# a_15002_46116# 1.85e-19
C23123 a_5937_45572# a_2324_44458# 0.407894f
C23124 a_15682_43940# a_16414_43172# 3.58e-19
C23125 a_20974_43370# a_20556_43646# 0.076332f
C23126 a_n2293_43922# a_2903_42308# 8.6e-20
C23127 a_5891_43370# a_6123_31319# 0.028865f
C23128 a_3905_42865# a_4649_42852# 0.04156f
C23129 a_3499_42826# a_3445_43172# 2.31e-19
C23130 a_11341_43940# a_10991_42826# 2.93e-19
C23131 a_14401_32519# a_21487_43396# 6.94e-19
C23132 a_n1435_47204# CLK 1.41989f
C23133 a_13717_47436# EN_OFFSET_CAL 0.002392f
C23134 a_16327_47482# RST_Z 1.85e-19
C23135 a_16867_43762# VDD 0.132317f
C23136 a_15599_45572# a_11691_44458# 1.35e-20
C23137 a_10490_45724# a_8975_43940# 7.33e-22
C23138 a_2711_45572# a_6109_44484# 3.03e-20
C23139 a_n1059_45260# a_375_42282# 0.0165f
C23140 a_5691_45260# a_6431_45366# 0.005044f
C23141 a_3537_45260# a_8191_45002# 0.00226f
C23142 a_5147_45002# a_7229_43940# 1.65e-22
C23143 a_4927_45028# a_5205_44484# 9.25e-21
C23144 a_3232_43370# a_6171_45002# 0.314056f
C23145 a_13635_43156# a_3483_46348# 1.81e-20
C23146 a_13113_42826# a_4185_45028# 3.91e-21
C23147 a_9396_43370# a_n357_42282# 1.13e-19
C23148 a_10341_43396# a_16375_45002# 1.23e-20
C23149 a_9127_43156# a_8199_44636# 0.01079f
C23150 a_10083_42826# a_8016_46348# 1.33e-19
C23151 a_8605_42826# a_8953_45546# 3.03e-19
C23152 a_18909_45814# a_4883_46098# 1.42e-21
C23153 a_19431_45546# a_13507_46334# 2.47e-20
C23154 a_21363_45546# a_16327_47482# 0.276554f
C23155 a_3357_43084# a_11459_47204# 5.7e-19
C23156 a_2437_43646# a_13717_47436# 0.085485f
C23157 a_21513_45002# a_12861_44030# 2.48e-20
C23158 a_413_45260# a_2952_47436# 0.026401f
C23159 a_5147_45002# a_n237_47217# 5.93e-20
C23160 a_2274_45254# a_584_46384# 3.31e-21
C23161 a_n467_45028# a_n1151_42308# 0.406349f
C23162 a_15765_45572# a_n881_46662# 0.58719f
C23163 a_11136_45572# a_12549_44172# 1.78e-21
C23164 a_3775_45552# a_3699_46634# 5.03e-19
C23165 a_2711_45572# a_4646_46812# 0.053113f
C23166 a_8568_45546# a_2107_46812# 2.03e-20
C23167 a_11525_45546# a_n743_46660# 1.75e-21
C23168 a_n2840_45546# a_n2956_38216# 0.019918f
C23169 a_n2810_45572# a_n2472_45546# 0.002308f
C23170 a_19095_43396# a_18249_42858# 6.34e-19
C23171 a_4190_30871# a_19987_42826# 3.95e-19
C23172 a_5649_42852# a_16795_42852# 4.02e-21
C23173 a_4361_42308# a_18083_42858# 2.01e-19
C23174 a_743_42282# a_19339_43156# 2.4e-20
C23175 a_n1557_42282# a_n784_42308# 0.058812f
C23176 a_9145_43396# a_14635_42282# 3.74e-20
C23177 a_21076_30879# a_22521_40055# 2.11e-20
C23178 a_20820_30879# a_22521_39511# 5.7e-20
C23179 a_13885_46660# CLK 2.64e-20
C23180 VDAC_Pi a_5088_37509# 0.391059f
C23181 a_7754_40130# VDAC_N 0.434929f
C23182 a_7754_39964# a_5700_37509# 0.095724f
C23183 VDAC_Ni a_8530_39574# 1.72e-20
C23184 a_n327_42308# VDD 1.42e-19
C23185 a_n1741_47186# a_n971_45724# 0.157081f
C23186 a_n1605_47204# a_n815_47178# 2.38e-19
C23187 a_n2109_47186# a_n237_47217# 0.730469f
C23188 a_n2497_47436# a_n785_47204# 4.85e-19
C23189 SMPL_ON_P a_n452_47436# 3.73e-21
C23190 a_1307_43914# a_3363_44484# 5.2e-19
C23191 a_9482_43914# a_13213_44734# 0.003145f
C23192 a_13556_45296# a_n2293_43922# 1.07e-20
C23193 a_375_42282# a_484_44484# 8.95e-19
C23194 a_11823_42460# a_12495_44260# 9.96e-20
C23195 a_3357_43084# a_22591_44484# 7.11e-20
C23196 a_22591_45572# a_22485_44484# 1.77e-19
C23197 a_19479_31679# a_17730_32519# 0.052745f
C23198 a_10149_42308# a_9290_44172# 0.001223f
C23199 a_9306_43218# a_n443_42852# 3.58e-20
C23200 a_13003_42852# a_n357_42282# 0.002208f
C23201 a_7174_31319# a_1823_45246# 1.97e-20
C23202 a_10341_43396# RST_Z 2.8e-19
C23203 a_10775_45002# a_10249_46116# 1.35e-22
C23204 a_10951_45334# a_10554_47026# 2.81e-22
C23205 a_20567_45036# a_19321_45002# 0.205038f
C23206 a_11827_44484# a_5807_45002# 0.022597f
C23207 a_21101_45002# a_13747_46662# 0.081818f
C23208 a_5105_45348# a_3877_44458# 9.23e-22
C23209 a_n2661_43370# a_2107_46812# 0.02614f
C23210 a_413_45260# a_12991_46634# 4.46e-20
C23211 a_8953_45002# a_6755_46942# 6.77e-20
C23212 a_n1059_45260# a_15227_44166# 0.099892f
C23213 a_2437_43646# a_14035_46660# 1.31e-19
C23214 a_6511_45714# a_6945_45028# 0.028815f
C23215 a_10490_45724# a_11387_46155# 1.07e-20
C23216 a_11525_45546# a_11189_46129# 0.085926f
C23217 a_11322_45546# a_11133_46155# 0.001455f
C23218 a_11652_45724# a_9290_44172# 0.020364f
C23219 a_10193_42453# a_12005_46116# 0.016165f
C23220 a_8746_45002# a_10903_43370# 1.84e-19
C23221 a_n2129_44697# a_n1613_43370# 0.026334f
C23222 a_n2661_43922# a_n1151_42308# 0.056653f
C23223 a_21855_43396# a_21613_42308# 2.52e-21
C23224 a_10835_43094# a_5742_30871# 0.011953f
C23225 a_10796_42968# a_11323_42473# 8.05e-20
C23226 a_5649_42852# a_21335_42336# 6.37e-20
C23227 a_13678_32519# a_21887_42336# 0.012293f
C23228 a_14209_32519# a_13258_32519# 0.051594f
C23229 a_n2293_42282# a_3823_42558# 3.04e-21
C23230 a_10341_42308# a_10545_42558# 0.002951f
C23231 a_1793_42852# a_1755_42282# 3.44e-19
C23232 a_1848_45724# DATA[1] 9.34e-21
C23233 a_12891_46348# a_12549_44172# 0.309821f
C23234 a_n2312_40392# a_n2293_46634# 4.37e-19
C23235 a_n2312_39304# a_n2442_46660# 0.15211f
C23236 a_4791_45118# a_5429_46660# 6.03e-19
C23237 a_2063_45854# a_10428_46928# 0.04306f
C23238 a_n971_45724# a_7832_46660# 0.013782f
C23239 a_n1151_42308# a_7927_46660# 5.63e-20
C23240 a_6491_46660# a_6540_46812# 0.079263f
C23241 a_18587_45118# a_15493_43940# 4.11e-22
C23242 a_19778_44110# a_11341_43940# 0.004296f
C23243 a_20567_45036# a_20623_43914# 4.97e-21
C23244 a_21359_45002# a_19862_44208# 0.001254f
C23245 a_11827_44484# a_19478_44306# 0.002282f
C23246 a_18184_42460# a_21115_43940# 1.01e-21
C23247 a_7499_43078# a_7227_42852# 0.126148f
C23248 a_14581_44484# a_14673_44172# 7.47e-20
C23249 a_2711_45572# a_15567_42826# 6.6e-20
C23250 a_15861_45028# a_17486_43762# 5.8e-21
C23251 a_3537_45260# a_3540_43646# 2.04e-20
C23252 a_3065_45002# a_3539_42460# 0.300764f
C23253 a_n913_45002# a_6452_43396# 1.57e-20
C23254 C5_N_btm VDD 0.267489f
C23255 a_13017_45260# VDD 0.263701f
C23256 COMP_P a_19864_35138# 3.57e-19
C23257 a_n1630_35242# a_n1386_35608# 0.019114f
C23258 a_14021_43940# a_12465_44636# 0.015806f
C23259 a_n447_43370# a_n1151_42308# 1.85e-19
C23260 a_n1557_42282# SMPL_ON_P 2.98e-20
C23261 a_3357_43084# a_n863_45724# 0.003254f
C23262 a_8953_45002# a_8049_45260# 7.24e-19
C23263 a_n2840_45002# a_n2840_45546# 0.026152f
C23264 a_375_42282# a_n1925_42282# 2.07e-19
C23265 a_n3674_39768# a_n2312_38680# 0.023176f
C23266 a_9313_44734# a_19692_46634# 3.49e-20
C23267 a_10807_43548# a_768_44030# 0.001051f
C23268 a_18443_44721# a_17339_46660# 0.006967f
C23269 a_2063_45854# VDD 3.60498f
C23270 a_5934_30871# a_7174_31319# 0.473128f
C23271 a_15803_42450# a_15890_42674# 0.07009f
C23272 a_n3674_38680# a_n3420_38528# 0.07337f
C23273 a_n3674_38216# a_n4209_38502# 4.47e-20
C23274 a_15764_42576# a_15720_42674# 1.46e-19
C23275 a_n3674_37592# a_n4064_39072# 0.019349f
C23276 a_21588_30879# a_11415_45002# 2.68e-19
C23277 a_10467_46802# a_11901_46660# 0.001328f
C23278 a_10249_46116# a_11186_47026# 0.172467f
C23279 a_7832_46660# a_8023_46660# 4.61e-19
C23280 a_1110_47026# a_765_45546# 2.11e-20
C23281 a_n881_46662# a_3147_46376# 0.073958f
C23282 a_n1613_43370# a_3483_46348# 0.029573f
C23283 a_4190_30871# a_n3420_37440# 0.034998f
C23284 a_13507_46334# a_12594_46348# 3.5e-19
C23285 a_4883_46098# a_10903_43370# 0.025531f
C23286 a_16327_47482# a_18985_46122# 0.051538f
C23287 a_10227_46804# a_17583_46090# 8.3e-22
C23288 a_14311_47204# a_6945_45028# 0.008982f
C23289 a_17591_47464# a_17715_44484# 0.001482f
C23290 a_11599_46634# a_20708_46348# 1.58e-20
C23291 a_12861_44030# a_10809_44734# 0.156561f
C23292 a_n1741_47186# a_12005_46436# 5.93e-20
C23293 a_n443_46116# a_518_46155# 0.001648f
C23294 a_n237_47217# a_8062_46155# 1.73e-19
C23295 a_11750_44172# a_12429_44172# 1.03e-20
C23296 a_2998_44172# a_2253_43940# 2.08e-19
C23297 a_n2661_42834# a_6765_43638# 4.91e-21
C23298 a_n2661_43922# a_6197_43396# 1.61e-20
C23299 a_14539_43914# a_15681_43442# 4.94e-20
C23300 a_20980_44850# a_20974_43370# 4.87e-21
C23301 a_3422_30871# a_21381_43940# 0.006676f
C23302 a_10193_42453# a_15890_42674# 8.41e-20
C23303 a_2711_45572# a_20712_42282# 4.18e-19
C23304 a_2675_43914# a_3052_44056# 7.61e-19
C23305 a_13249_42308# a_12563_42308# 1.64e-19
C23306 a_11823_42460# a_13333_42558# 0.003508f
C23307 a_n2293_43922# a_6293_42852# 9.77e-21
C23308 a_20193_45348# a_14209_32519# 5.6e-19
C23309 a_n913_45002# a_13291_42460# 0.070562f
C23310 a_n1059_45260# a_14635_42282# 0.063373f
C23311 a_3537_45260# a_7309_42852# 4.49e-19
C23312 a_19006_44850# VDD 0.077608f
C23313 a_10193_42453# a_10490_45724# 0.062365f
C23314 a_2711_45572# a_10216_45572# 9.36e-19
C23315 a_n2661_42282# a_4185_45028# 0.833759f
C23316 a_15493_43940# a_11415_45002# 1.15e-19
C23317 a_4361_42308# a_12549_44172# 8.96e-19
C23318 a_20974_43370# a_19692_46634# 0.012779f
C23319 a_16823_43084# a_13661_43548# 7.25e-19
C23320 a_13857_44734# a_13259_45724# 0.03212f
C23321 a_9313_44734# a_20692_30879# 1.31e-20
C23322 a_2479_44172# a_2324_44458# 0.010173f
C23323 a_8952_43230# a_10227_46804# 7.54e-21
C23324 a_12469_46902# VDD 0.203316f
C23325 a_n3565_39304# C1_P_btm 1.3e-20
C23326 a_5742_30871# a_7754_40130# 0.005581f
C23327 a_n2293_46098# a_3483_46348# 0.044283f
C23328 a_805_46414# a_1208_46090# 0.002746f
C23329 a_472_46348# a_1176_45822# 0.146555f
C23330 a_376_46348# a_1138_42852# 3.05e-21
C23331 a_2959_46660# a_3316_45546# 5.39e-21
C23332 a_3877_44458# a_n863_45724# 4.38e-21
C23333 a_8270_45546# a_8062_46155# 8.57e-21
C23334 a_17339_46660# a_17583_46090# 0.004328f
C23335 a_765_45546# a_15682_46116# 0.005634f
C23336 a_14180_46812# a_10809_44734# 0.012862f
C23337 a_9313_44734# a_16877_43172# 5.07e-19
C23338 a_5244_44056# a_5111_42852# 9.76e-21
C23339 a_12429_44172# a_4361_42308# 1.84e-21
C23340 a_n97_42460# a_6293_42852# 0.018467f
C23341 a_14021_43940# a_16409_43396# 0.025204f
C23342 a_n2661_42282# a_n2157_42858# 4.07e-20
C23343 a_742_44458# a_2903_42308# 0.0077f
C23344 a_3422_30871# a_18249_42858# 1.45e-20
C23345 a_1568_43370# a_2982_43646# 0.002246f
C23346 a_n2956_37592# a_n4209_38216# 0.104159f
C23347 a_548_43396# VDD 4.01e-19
C23348 a_15765_45572# a_1307_43914# 9.23e-20
C23349 a_8696_44636# a_14537_43396# 0.024289f
C23350 a_15903_45785# a_16751_45260# 2.12e-20
C23351 a_17303_42282# a_16327_47482# 4.29e-19
C23352 a_15521_42308# a_10227_46804# 0.001965f
C23353 a_8791_42308# a_n1613_43370# 6.28e-21
C23354 a_17538_32519# a_20205_31679# 0.051233f
C23355 a_16823_43084# a_4185_45028# 6.8e-21
C23356 a_n2293_43922# RST_Z 4.75e-21
C23357 a_14383_46116# VDD 0.132317f
C23358 a_2711_45572# a_9804_47204# 2.39e-19
C23359 a_6194_45824# a_n881_46662# 0.063172f
C23360 a_6472_45840# a_n1613_43370# 0.017909f
C23361 a_8746_45002# a_4883_46098# 0.032616f
C23362 a_13249_42308# a_10227_46804# 0.064815f
C23363 a_n1379_46482# a_n2293_45546# 1.3e-20
C23364 a_8049_45260# a_11601_46155# 6.51e-19
C23365 a_2324_44458# a_n443_42852# 2.42e-19
C23366 a_4361_42308# a_21855_43396# 0.167446f
C23367 a_10341_43396# a_10991_42826# 7.08e-20
C23368 a_15095_43370# a_12379_42858# 1.62e-21
C23369 a_13467_32519# a_13678_32519# 10.9526f
C23370 a_17730_32519# a_13258_32519# 0.05785f
C23371 a_3422_30871# a_21125_42558# 2.49e-20
C23372 VDAC_N C6_N_btm 55.2142f
C23373 a_16147_45260# a_17517_44484# 8.68e-20
C23374 a_6171_45002# a_8975_43940# 0.175346f
C23375 a_3232_43370# a_12607_44458# 1.04e-20
C23376 a_5932_42308# a_1823_45246# 8.68e-21
C23377 a_8387_43230# a_n443_42852# 0.006907f
C23378 a_13635_43156# a_n357_42282# 0.008746f
C23379 a_n97_42460# RST_Z 2.62e-20
C23380 a_n2661_43370# a_11453_44696# 0.002123f
C23381 a_19778_44110# a_16327_47482# 0.037655f
C23382 a_16922_45042# a_18479_47436# 6.1e-20
C23383 C5_P_btm VDD 0.267489f
C23384 a_n452_44636# a_n1151_42308# 0.238824f
C23385 a_6517_45366# a_n881_46662# 5.23e-19
C23386 a_7229_43940# a_n1925_46634# 3.86e-21
C23387 a_5205_44484# a_n743_46660# 2.07e-20
C23388 a_4574_45260# a_2107_46812# 3.63e-20
C23389 a_413_45260# a_n2661_46098# 1.23e-20
C23390 a_16855_45546# a_15368_46634# 6.26e-21
C23391 a_15415_45028# a_13661_43548# 0.133591f
C23392 a_10951_45334# a_n2661_46634# 9.5e-21
C23393 a_8696_44636# a_3090_45724# 0.038457f
C23394 a_13904_45546# a_765_45546# 7.77e-22
C23395 a_15599_45572# a_15227_44166# 4.09e-21
C23396 a_6472_45840# a_n2293_46098# 6.84e-21
C23397 a_743_42282# a_3905_42308# 3.67e-19
C23398 a_16547_43609# a_15803_42450# 1.5e-20
C23399 a_16243_43396# a_15959_42545# 6.33e-20
C23400 a_16409_43396# a_15764_42576# 6.83e-20
C23401 a_791_42968# a_1067_42314# 2.04e-19
C23402 a_18249_42858# a_18504_43218# 0.05936f
C23403 a_4361_42308# a_7227_42308# 0.01047f
C23404 a_16137_43396# a_15890_42674# 2.67e-21
C23405 a_10341_43396# a_17303_42282# 1.21e-20
C23406 a_13467_32519# a_6123_31319# 2.49e-19
C23407 a_16414_43172# a_16245_42852# 0.08213f
C23408 a_n3420_38528# VDD 0.522772f
C23409 a_3422_30871# a_8530_39574# 1.13e-19
C23410 a_6151_47436# a_13675_47204# 0.002433f
C23411 a_9313_45822# a_9804_47204# 0.171044f
C23412 a_12861_44030# a_n881_46662# 0.135351f
C23413 a_n746_45260# a_n1021_46688# 8.61e-21
C23414 a_n2109_47186# a_1123_46634# 3.71e-19
C23415 a_n452_47436# a_n2438_43548# 3.48e-19
C23416 a_n237_47217# a_n1925_46634# 0.079348f
C23417 a_1431_47204# a_n2661_46634# 0.001833f
C23418 a_n971_45724# a_n743_46660# 0.122713f
C23419 a_13507_46334# a_12465_44636# 0.029101f
C23420 a_21496_47436# a_21811_47423# 3.73e-19
C23421 a_19787_47423# a_11453_44696# 1.96e-19
C23422 a_10775_45002# a_10555_44260# 2.44e-20
C23423 a_9482_43914# a_11341_43940# 0.037822f
C23424 a_13076_44458# a_13296_44484# 0.009965f
C23425 a_700_44734# a_556_44484# 6.84e-19
C23426 a_8375_44464# a_8783_44734# 5.23e-21
C23427 a_n2661_43370# a_n3674_39768# 0.144159f
C23428 a_12607_44458# a_14581_44484# 3.05e-21
C23429 a_n1821_44484# a_n2661_43922# 0.001334f
C23430 a_n1655_44484# a_n2661_42834# 5.04e-19
C23431 a_19479_31679# a_17538_32519# 0.051112f
C23432 a_2382_45260# a_3992_43940# 4.5e-19
C23433 a_22465_38105# a_20205_31679# 3.95e-19
C23434 a_20107_45572# VDD 0.458237f
C23435 a_626_44172# a_167_45260# 0.04273f
C23436 a_1423_45028# a_1823_45246# 0.024089f
C23437 a_20679_44626# a_19321_45002# 0.023087f
C23438 a_19279_43940# a_13661_43548# 6.72e-19
C23439 a_18114_32519# a_19692_46634# 5.21e-19
C23440 a_20397_44484# a_12549_44172# 1.48e-19
C23441 a_20766_44850# a_13747_46662# 1.67e-19
C23442 a_n2017_45002# a_n2956_39304# 9.09e-22
C23443 a_2437_43646# a_n1925_42282# 2.49e-20
C23444 a_10951_45334# a_8199_44636# 0.237774f
C23445 a_10775_45002# a_5937_45572# 1.83e-20
C23446 a_n2472_43914# a_n1613_43370# 1.2e-19
C23447 a_8953_45002# a_8953_45546# 0.023516f
C23448 a_2680_45002# a_2324_44458# 9e-20
C23449 a_3232_43370# a_10903_43370# 0.114259f
C23450 a_n913_45002# a_10809_44734# 0.0025f
C23451 a_6761_42308# a_7227_42308# 0.173849f
C23452 a_5932_42308# a_5934_30871# 1.37963f
C23453 a_1606_42308# a_13575_42558# 1.77e-20
C23454 a_n1532_35090# a_n83_35174# 0.558402f
C23455 a_n923_35174# EN_VIN_BSTR_P 1.02927f
C23456 a_n1925_46634# a_8270_45546# 0.109762f
C23457 a_5807_45002# a_15559_46634# 0.006621f
C23458 a_13747_46662# a_14976_45028# 0.016638f
C23459 a_n2661_46634# a_11735_46660# 0.044956f
C23460 a_16131_47204# a_16292_46812# 2.31e-19
C23461 a_4817_46660# a_5167_46660# 0.218775f
C23462 a_4646_46812# a_6540_46812# 0.029952f
C23463 a_4651_46660# a_5732_46660# 0.102355f
C23464 a_3877_44458# a_5072_46660# 0.021873f
C23465 a_13661_43548# a_15368_46634# 3.74e-20
C23466 a_n881_46662# a_14180_46812# 0.028137f
C23467 a_11453_44696# a_20107_46660# 0.050203f
C23468 a_12465_44636# a_20623_46660# 4.37e-20
C23469 a_n1741_47186# a_12594_46348# 0.150956f
C23470 a_2063_45854# a_7920_46348# 3.54e-19
C23471 a_n1151_42308# a_5164_46348# 0.110485f
C23472 a_n237_47217# a_10355_46116# 1.06e-20
C23473 a_4007_47204# a_4185_45028# 7.03e-19
C23474 a_n443_46116# a_3147_46376# 0.002662f
C23475 a_4791_45118# a_3483_46348# 0.088998f
C23476 a_18597_46090# a_18900_46660# 0.00136f
C23477 a_10227_46804# a_20885_46660# 0.001925f
C23478 a_n1435_47204# a_n1991_46122# 1.76e-20
C23479 a_4883_46098# a_21188_46660# 0.012559f
C23480 a_21811_47423# a_21363_46634# 0.010128f
C23481 a_13507_46334# a_20528_46660# 0.00277f
C23482 a_11967_42832# a_15493_43940# 0.299734f
C23483 a_20159_44458# a_11341_43940# 6.61e-20
C23484 a_20679_44626# a_20623_43914# 0.009865f
C23485 a_19279_43940# a_19862_44208# 0.012567f
C23486 a_20640_44752# a_20935_43940# 4.13e-20
C23487 a_18579_44172# a_19328_44172# 0.053539f
C23488 a_1115_44172# a_1241_44260# 0.013015f
C23489 a_5495_43940# a_6453_43914# 5.83e-20
C23490 a_n699_43396# a_548_43396# 2.06e-19
C23491 a_n1761_44111# a_n2661_42282# 5.46e-20
C23492 a_19778_44110# a_10341_43396# 1.31e-19
C23493 a_n2661_42834# a_8487_44056# 1.89e-21
C23494 a_n2017_45002# a_5534_30871# 0.025363f
C23495 a_n1059_45260# a_14543_43071# 0.002239f
C23496 a_n913_45002# a_13460_43230# 0.04239f
C23497 a_3232_43370# a_3681_42891# 0.005411f
C23498 a_5111_44636# a_5111_42852# 0.148196f
C23499 a_3537_45260# a_7765_42852# 2.41e-19
C23500 a_18374_44850# VDD 0.203584f
C23501 a_n4064_39616# C3_P_btm 5.52e-20
C23502 a_n4064_39072# EN_VIN_BSTR_P 0.959329f
C23503 a_15743_43084# a_18479_47436# 4.35e-20
C23504 a_n1641_43230# a_n1151_42308# 9.41e-19
C23505 a_4181_44734# a_n1925_42282# 6.6e-19
C23506 a_18114_32519# a_20692_30879# 0.051555f
C23507 a_19721_31679# a_20205_31679# 0.052217f
C23508 a_17767_44458# a_8049_45260# 9.2e-21
C23509 a_20365_43914# a_3090_45724# 1.09e-19
C23510 a_18326_43940# a_15227_44166# 5.29e-20
C23511 a_3540_43646# a_n2293_46634# 0.003694f
C23512 a_n2472_43914# a_n2293_46098# 5.06e-21
C23513 a_n4064_39072# a_n2302_39072# 0.250408f
C23514 a_n4064_40160# a_n3565_38216# 0.02828f
C23515 a_n4064_39616# a_n4064_38528# 0.05063f
C23516 a_n3420_39072# a_n3607_39392# 8.36e-19
C23517 a_5742_30871# C6_N_btm 0.170624f
C23518 a_20841_46902# a_20731_47026# 0.097745f
C23519 a_21363_46634# a_22000_46634# 0.017308f
C23520 a_20623_46660# a_20528_46660# 0.049827f
C23521 a_19123_46287# a_18900_46660# 0.001018f
C23522 a_2107_46812# a_9823_46482# 2.17e-19
C23523 a_n881_46662# a_310_45028# 7.88e-19
C23524 a_6755_46942# a_15015_46420# 0.133517f
C23525 a_3090_45724# a_4704_46090# 4.99e-19
C23526 a_8270_45546# a_10355_46116# 2.83e-19
C23527 a_n1613_43370# a_n357_42282# 0.030838f
C23528 a_10949_43914# a_8685_43396# 4.56e-21
C23529 a_2253_43940# a_1568_43370# 3.94e-19
C23530 a_18579_44172# a_20749_43396# 5.9e-20
C23531 a_20512_43084# a_21487_43396# 0.003816f
C23532 a_n2293_43922# a_10991_42826# 2.64e-20
C23533 a_9313_44734# a_5342_30871# 0.026413f
C23534 a_1307_43914# a_8685_42308# 1.98e-21
C23535 a_18184_42460# a_20256_42852# 0.01674f
C23536 a_19319_43548# a_19741_43940# 0.048788f
C23537 a_3422_30871# a_5649_42852# 0.291966f
C23538 a_n1059_45260# a_19511_42282# 3.28e-19
C23539 a_n2017_45002# a_19647_42308# 1.94e-19
C23540 en_comp a_19332_42282# 4.59e-20
C23541 a_20447_31679# a_22775_42308# 4.98e-21
C23542 a_19479_31679# a_22465_38105# 2.87e-19
C23543 a_5326_44056# VDD 0.001151f
C23544 a_18341_45572# a_18909_45814# 0.170692f
C23545 a_18479_45785# a_18691_45572# 0.036486f
C23546 a_18175_45572# a_19431_45546# 0.043567f
C23547 a_16147_45260# a_19256_45572# 2.79e-20
C23548 a_8746_45002# a_3232_43370# 0.439467f
C23549 a_7499_43078# a_7229_43940# 9.29e-21
C23550 a_10193_42453# a_6171_45002# 0.411891f
C23551 a_8791_43396# a_3483_46348# 4.38e-23
C23552 a_19700_43370# a_17339_46660# 3.22e-19
C23553 a_13887_32519# a_19692_46634# 2.91e-19
C23554 a_15493_43940# a_13259_45724# 0.019228f
C23555 a_7584_44260# a_n357_42282# 7.22e-20
C23556 a_3626_43646# a_8953_45546# 0.005746f
C23557 a_n1736_42282# a_n2312_40392# 4.5e-20
C23558 a_n3674_38216# a_n2312_39304# 0.023615f
C23559 a_5088_37509# RST_Z 0.059771f
C23560 a_n4209_37414# VREF 0.056254f
C23561 a_n3565_37414# VIN_P 0.029764f
C23562 VDAC_P C6_P_btm 55.214397f
C23563 a_18114_32519# VIN_N 0.063295f
C23564 a_17715_44484# VDD 0.526119f
C23565 a_5907_45546# a_4915_47217# 4.1e-22
C23566 a_2711_45572# a_6545_47178# 8.4e-19
C23567 a_7499_43078# a_n237_47217# 4.22e-20
C23568 a_6194_45824# a_n443_46116# 8.96e-21
C23569 a_6472_45840# a_4791_45118# 0.025301f
C23570 a_11322_45546# a_n1741_47186# 0.003846f
C23571 a_n3565_38216# a_n4064_37440# 0.032797f
C23572 a_n2293_46098# a_n357_42282# 0.014918f
C23573 a_n1076_46494# a_n2293_45546# 7.13e-22
C23574 a_805_46414# a_n2661_45546# 7.52e-20
C23575 a_n901_46420# a_n1079_45724# 1.93e-20
C23576 a_n1853_46287# a_n1099_45572# 0.067343f
C23577 a_15015_46420# a_8049_45260# 0.002448f
C23578 a_12594_46348# a_10586_45546# 8.27e-20
C23579 a_4699_43561# a_4520_42826# 1.02e-19
C23580 a_16137_43396# a_16547_43609# 0.151161f
C23581 a_3080_42308# a_3935_42891# 0.017131f
C23582 a_n97_42460# a_10991_42826# 6.43e-20
C23583 a_9313_44734# a_20107_42308# 8.02e-20
C23584 a_14579_43548# a_16823_43084# 3.51e-21
C23585 a_10341_43396# a_15231_43396# 1.63e-19
C23586 a_19321_45002# SINGLE_ENDED 1.12e-19
C23587 a_19594_46812# START 0.020669f
C23588 a_10083_42826# VDD 0.461256f
C23589 a_13249_42308# a_14815_43914# 4.82e-21
C23590 a_3357_43084# a_18114_32519# 8.45e-21
C23591 a_6709_45028# a_n2661_43370# 0.041021f
C23592 a_19479_31679# a_19721_31679# 9.039419f
C23593 a_8191_45002# a_8704_45028# 8.88e-19
C23594 a_n2017_45002# a_11691_44458# 4.56e-21
C23595 a_6171_45002# a_14309_45348# 3.25e-19
C23596 a_4361_42308# a_n2661_45546# 1.97e-21
C23597 a_13887_32519# a_20692_30879# 0.051577f
C23598 a_743_42282# a_n863_45724# 0.05133f
C23599 a_15743_43084# a_n443_42852# 0.034562f
C23600 a_14097_32519# a_21076_30879# 0.054945f
C23601 a_12791_45546# a_6755_46942# 4.95e-22
C23602 a_7499_43078# a_8270_45546# 0.063428f
C23603 a_2711_45572# a_19692_46634# 4.14e-20
C23604 a_20841_45814# a_20916_46384# 1.18e-19
C23605 a_20528_45572# a_19321_45002# 7.43e-20
C23606 a_2437_43646# a_16285_47570# 7.17e-19
C23607 a_n913_45002# a_n881_46662# 0.00874f
C23608 a_n745_45366# a_n1613_43370# 0.012092f
C23609 a_3232_43370# a_4883_46098# 0.017979f
C23610 a_11787_45002# a_10227_46804# 1.63e-21
C23611 a_1307_43914# a_12861_44030# 0.038753f
C23612 a_16795_42852# a_17333_42852# 0.108694f
C23613 a_17595_43084# a_18083_42858# 0.046381f
C23614 a_3626_43646# a_14456_42282# 0.005342f
C23615 a_n97_42460# a_17303_42282# 2.32e-20
C23616 a_17538_32519# a_13258_32519# 0.054578f
C23617 a_4190_30871# a_18861_43218# 9.99e-19
C23618 a_n1741_47186# a_12465_44636# 4.19e-22
C23619 a_5129_47502# a_n1435_47204# 4.12e-19
C23620 a_7227_47204# a_9067_47204# 3.76e-21
C23621 a_7903_47542# a_6575_47204# 0.046223f
C23622 a_6151_47436# a_11459_47204# 0.034818f
C23623 a_4915_47217# a_13717_47436# 4.05e-19
C23624 a_n1177_44458# a_n356_44636# 1.98e-19
C23625 a_8975_43940# a_12607_44458# 0.004748f
C23626 a_n2661_44458# a_700_44734# 5e-19
C23627 a_n2956_37592# a_n2661_42282# 1.91e-20
C23628 a_n2017_45002# a_8333_44056# 1.11e-21
C23629 a_5111_44636# a_7542_44172# 0.039468f
C23630 a_5205_44484# a_5244_44056# 1.29e-20
C23631 a_3232_43370# a_5663_43940# 0.090892f
C23632 a_20623_45572# a_11341_43940# 1.76e-21
C23633 a_1606_42308# a_n443_42852# 0.003624f
C23634 a_3581_42558# a_n755_45592# 2.25e-19
C23635 a_14495_45572# VDD 0.238674f
C23636 a_13678_32519# VCM 0.014539f
C23637 a_13887_32519# VIN_N 0.061374f
C23638 a_13296_44484# a_12465_44636# 1.43e-19
C23639 a_20159_44458# a_16327_47482# 0.270426f
C23640 a_18579_44172# a_12861_44030# 0.221909f
C23641 a_n809_44244# a_n1151_42308# 0.02481f
C23642 a_1414_42308# a_584_46384# 0.321387f
C23643 a_n3674_39768# a_n2497_47436# 5.96e-20
C23644 a_15903_45785# a_10809_44734# 2.74e-20
C23645 a_8336_45822# a_5066_45546# 8.57e-20
C23646 a_12791_45546# a_8049_45260# 0.005799f
C23647 a_11322_45546# a_10586_45546# 0.220166f
C23648 a_n2017_45002# a_n1991_46122# 5.3e-19
C23649 a_5883_43914# a_2107_46812# 0.009818f
C23650 a_5009_45028# a_3090_45724# 0.008714f
C23651 a_8375_44464# a_768_44030# 0.001943f
C23652 a_13076_44458# a_n743_46660# 9.1e-21
C23653 a_14180_45002# a_13059_46348# 0.073427f
C23654 a_n1059_45260# a_n1853_46287# 0.006746f
C23655 a_413_45260# a_11415_45002# 0.063143f
C23656 a_2437_43646# a_2698_46116# 6.23e-21
C23657 a_n2293_45010# a_n1641_46494# 2.7e-19
C23658 a_n2661_45010# a_n1076_46494# 1.72e-21
C23659 a_18249_42858# a_7174_31319# 1.28e-20
C23660 a_19987_42826# a_19511_42282# 1.28e-19
C23661 a_196_42282# a_564_42282# 7.52e-19
C23662 a_n473_42460# a_n1630_35242# 0.049561f
C23663 a_n4318_38680# a_n3420_38528# 0.001905f
C23664 a_n784_42308# a_n3674_37592# 0.254719f
C23665 a_n1925_46634# a_1123_46634# 0.018809f
C23666 a_n743_46660# a_601_46902# 0.022066f
C23667 a_n2438_43548# a_33_46660# 0.588568f
C23668 a_n133_46660# a_171_46873# 0.163873f
C23669 a_n1613_43370# a_5263_46660# 7.38e-19
C23670 a_11599_46634# a_14976_45028# 0.020184f
C23671 a_10227_46804# a_11813_46116# 0.094518f
C23672 a_15811_47375# a_15009_46634# 2.23e-19
C23673 a_4915_47217# a_14035_46660# 0.075669f
C23674 a_12861_44030# a_17609_46634# 0.183853f
C23675 a_1431_47204# a_765_45546# 0.00505f
C23676 a_9482_43914# a_10341_43396# 7.76e-20
C23677 a_18989_43940# a_15493_43940# 0.025737f
C23678 a_9313_44734# a_9672_43914# 1.48e-19
C23679 a_1307_43914# a_9803_43646# 9.06e-20
C23680 a_14537_43396# a_14205_43396# 0.080783f
C23681 a_n2661_42834# a_3499_42826# 0.009315f
C23682 a_4223_44672# a_5745_43940# 0.040431f
C23683 a_3422_30871# a_21145_44484# 6.39e-20
C23684 a_20193_45348# a_17538_32519# 2.12e-19
C23685 a_n2661_43922# a_2537_44260# 1.23e-19
C23686 a_n2293_42834# a_648_43396# 6.38e-19
C23687 a_n2293_45010# a_743_42282# 1.96e-21
C23688 a_n2017_45002# a_4190_30871# 0.025499f
C23689 a_3754_39964# VDD 0.033808f
C23690 a_17719_45144# VDD 0.1297f
C23691 a_5742_30871# C4_P_btm 0.03103f
C23692 a_6123_31319# VCM 0.144585f
C23693 a_n3565_37414# a_n2956_38680# 9.9e-21
C23694 a_n2661_43922# a_12741_44636# 0.00322f
C23695 a_n2661_42282# a_5257_43370# 0.01339f
C23696 a_22485_44484# a_19692_46634# 1.22e-19
C23697 a_375_42282# a_380_45546# 3.56e-19
C23698 a_626_44172# a_n863_45724# 0.097275f
C23699 a_1423_45028# a_n2293_45546# 0.06244f
C23700 a_2809_45348# a_n2661_45546# 9.78e-19
C23701 a_8975_43940# a_10903_43370# 0.043009f
C23702 a_5518_44484# a_2324_44458# 0.112753f
C23703 a_13720_44458# a_9290_44172# 2.01e-19
C23704 a_n2661_44458# a_10809_44734# 0.033319f
C23705 a_n2433_43396# a_n1613_43370# 0.299968f
C23706 a_6472_45840# DATA[3] 2.3e-21
C23707 a_13258_32519# a_22465_38105# 0.056749f
C23708 a_4646_46812# a_1823_45246# 8.67e-19
C23709 a_15009_46634# a_13059_46348# 0.054389f
C23710 a_11735_46660# a_765_45546# 0.006002f
C23711 a_3090_45724# a_15227_46910# 0.010657f
C23712 a_n881_46662# a_3873_46454# 0.003191f
C23713 a_13747_46662# a_19900_46494# 0.001247f
C23714 a_n743_46660# a_12594_46348# 0.0427f
C23715 a_19321_45002# a_19335_46494# 0.006071f
C23716 a_2107_46812# a_9569_46155# 0.018199f
C23717 a_19594_46812# a_19553_46090# 8.61e-19
C23718 a_16131_47204# a_6945_45028# 0.003013f
C23719 a_n2661_46634# a_2324_44458# 0.0278f
C23720 a_n1151_42308# a_3316_45546# 5.6e-21
C23721 a_4791_45118# a_n357_42282# 0.020355f
C23722 a_n443_46116# a_310_45028# 0.06667f
C23723 a_10227_46804# a_14949_46494# 6.03e-19
C23724 a_11599_46634# a_18051_46116# 0.03664f
C23725 a_4883_46098# a_11608_46482# 5.79e-19
C23726 a_n23_44458# a_n1853_43023# 4.42e-21
C23727 a_8103_44636# a_8037_42858# 2.12e-21
C23728 a_20159_44458# a_10341_43396# 3.98e-20
C23729 a_2998_44172# a_2896_43646# 0.001865f
C23730 a_n2661_42282# a_n2267_43396# 5.11e-21
C23731 a_9313_44734# a_743_42282# 0.024013f
C23732 a_n2017_45002# a_5337_42558# 0.001525f
C23733 en_comp a_5379_42460# 1.81e-20
C23734 a_n913_45002# a_4933_42558# 0.005299f
C23735 a_n1059_45260# a_4921_42308# 6.43e-19
C23736 a_2382_45260# a_1755_42282# 4.8e-19
C23737 a_261_44278# VDD 2.43e-19
C23738 a_8697_45822# a_8696_44636# 1.69e-20
C23739 a_2711_45572# a_3357_43084# 0.037825f
C23740 a_13003_42852# a_12861_44030# 6.07e-20
C23741 a_n473_42460# a_n971_45724# 0.094491f
C23742 a_1184_42692# a_n2497_47436# 3.5e-22
C23743 a_n3674_37592# SMPL_ON_P 0.051746f
C23744 a_15493_43940# a_18189_46348# 1.31e-20
C23745 a_8333_44056# a_526_44458# 1.1e-21
C23746 a_12545_42858# a_13661_43548# 1.24e-19
C23747 a_17595_43084# a_12549_44172# 2.6e-20
C23748 a_7765_42852# a_n2293_46634# 6.5e-21
C23749 a_14205_43396# a_3090_45724# 0.040425f
C23750 a_22365_46825# VDD 0.193587f
C23751 a_1736_39587# a_2113_38308# 0.100626f
C23752 a_n4209_39304# a_n4064_37984# 0.029462f
C23753 a_n3565_39304# a_n3420_37984# 0.028129f
C23754 a_16522_42674# CAL_N 2.6e-20
C23755 a_n1076_46494# a_n914_46116# 0.006453f
C23756 a_n2293_46098# a_518_46155# 3.23e-19
C23757 a_3090_45724# a_2957_45546# 0.167712f
C23758 a_3483_46348# a_6945_45028# 0.002307f
C23759 a_11189_46129# a_12594_46348# 0.001927f
C23760 a_11387_46155# a_10903_43370# 7.72e-19
C23761 a_8199_44636# a_2324_44458# 0.412215f
C23762 a_15682_43940# a_15567_42826# 1.02e-19
C23763 a_21381_43940# a_21487_43396# 0.007531f
C23764 a_3499_42826# a_n2293_42282# 0.058548f
C23765 a_5891_43370# a_7227_42308# 8.82e-19
C23766 a_n2293_43922# a_2713_42308# 4.97e-20
C23767 a_20193_45348# a_22465_38105# 7.48e-20
C23768 a_19721_31679# a_13258_32519# 0.054727f
C23769 a_9396_43370# a_9803_43646# 9.33e-19
C23770 a_20974_43370# a_743_42282# 1.42e-19
C23771 a_3905_42865# a_4149_42891# 0.002034f
C23772 a_11341_43940# a_10796_42968# 4.28e-19
C23773 a_14401_32519# a_20556_43646# 2.02e-19
C23774 a_13381_47204# CLK 2.37e-19
C23775 a_16241_47178# RST_Z 5.18e-20
C23776 a_16664_43396# VDD 0.077608f
C23777 a_16333_45814# a_11827_44484# 3.46e-21
C23778 a_10490_45724# a_10057_43914# 4.22e-20
C23779 a_8746_45002# a_8975_43940# 0.016889f
C23780 a_5691_45260# a_6171_45002# 0.057463f
C23781 a_5111_44636# a_5205_44484# 0.200189f
C23782 a_n2661_45010# a_1423_45028# 4.66e-19
C23783 a_n2017_45002# a_375_42282# 0.03181f
C23784 a_n913_45002# a_1307_43914# 0.298747f
C23785 a_n2293_45010# a_626_44172# 0.024201f
C23786 a_12545_42858# a_4185_45028# 3.65e-20
C23787 a_19332_42282# a_13661_43548# 1.85e-21
C23788 a_8147_43396# a_n755_45592# 0.134231f
C23789 a_8791_43396# a_n357_42282# 1.18e-21
C23790 a_2813_43396# a_n863_45724# 1.63e-19
C23791 a_3539_42460# a_n443_42852# 0.02291f
C23792 a_8387_43230# a_8199_44636# 9.49e-20
C23793 a_8037_42858# a_8953_45546# 0.017317f
C23794 w_11334_34010# C0_dummy_N_btm 3.87e-21
C23795 a_18341_45572# a_4883_46098# 1.94e-20
C23796 a_18691_45572# a_13507_46334# 6.86e-21
C23797 a_20623_45572# a_16327_47482# 0.168593f
C23798 a_3357_43084# a_9313_45822# 2.85e-19
C23799 a_2437_43646# a_n1435_47204# 0.191468f
C23800 a_1667_45002# a_584_46384# 3.89e-20
C23801 a_5111_44636# a_n971_45724# 0.381443f
C23802 a_n913_45002# a_n443_46116# 0.002757f
C23803 a_n955_45028# a_n1151_42308# 2.98e-19
C23804 a_413_45260# a_2553_47502# 0.004176f
C23805 a_15903_45785# a_n881_46662# 0.032602f
C23806 a_11823_42460# a_n2293_46634# 0.072996f
C23807 a_2711_45572# a_3877_44458# 0.099631f
C23808 a_11322_45546# a_n743_46660# 3.68e-19
C23809 a_n2810_45572# a_n2661_45546# 0.006676f
C23810 a_n2840_45546# a_n2472_45546# 7.52e-19
C23811 a_1568_43370# a_1184_42692# 2.36e-19
C23812 a_1756_43548# a_1576_42282# 1e-20
C23813 a_4190_30871# a_19164_43230# 0.005605f
C23814 a_4361_42308# a_17701_42308# 0.004927f
C23815 a_743_42282# a_18599_43230# 1.85e-20
C23816 a_n1557_42282# a_196_42282# 0.031105f
C23817 a_1049_43396# a_961_42354# 1.08e-19
C23818 a_14021_43940# a_15890_42674# 3.09e-21
C23819 a_n4318_39768# a_n4334_39392# 3.4e-19
C23820 a_13887_32519# a_5342_30871# 0.028465f
C23821 a_14209_32519# a_5534_30871# 0.057361f
C23822 a_9145_43396# a_13291_42460# 6.23e-20
C23823 a_11341_43940# a_4958_30871# 2.27e-20
C23824 VDAC_Ni a_7754_38470# 0.005657f
C23825 VDAC_Pi a_4338_37500# 1.92369f
C23826 a_7754_40130# a_6886_37412# 0.006212f
C23827 a_7754_39964# a_5088_37509# 0.392826f
C23828 a_16721_46634# RST_Z 5.46e-22
C23829 a_2351_42308# VDD 0.188239f
C23830 a_n1741_47186# a_n452_47436# 0.013149f
C23831 a_n1920_47178# a_n971_45724# 1.39e-20
C23832 a_n2109_47186# a_n746_45260# 0.295988f
C23833 SMPL_ON_P a_n815_47178# 0.002605f
C23834 a_n2833_47464# a_n785_47204# 5.95e-22
C23835 a_13348_45260# a_13213_44734# 1.03e-19
C23836 a_1423_45028# a_8855_44734# 1.81e-20
C23837 a_9482_43914# a_n2293_43922# 0.018115f
C23838 a_413_45260# a_11967_42832# 4.85e-22
C23839 a_n913_45002# a_18579_44172# 7.45e-21
C23840 a_19479_31679# a_22591_44484# 0.00246f
C23841 a_21513_45002# a_19237_31679# 4.7e-20
C23842 a_9061_43230# a_n443_42852# 1.22e-20
C23843 a_4921_42308# a_n1925_42282# 1.23e-19
C23844 a_19332_42282# a_4185_45028# 1.64e-19
C23845 a_10775_45002# a_10554_47026# 2.81e-22
C23846 a_10951_45334# a_10623_46897# 4.99e-21
C23847 a_18494_42460# a_19321_45002# 0.084551f
C23848 a_21005_45260# a_13747_46662# 0.058269f
C23849 a_4640_45348# a_3877_44458# 1.44e-20
C23850 a_2437_43646# a_13885_46660# 1.22e-20
C23851 a_8953_45002# a_10249_46116# 9.14e-20
C23852 a_n2017_45002# a_15227_44166# 0.005144f
C23853 a_n2661_44458# a_n881_46662# 0.001141f
C23854 a_11525_45546# a_9290_44172# 0.001224f
C23855 a_10193_42453# a_10903_43370# 0.402091f
C23856 a_6472_45840# a_6945_45028# 0.034109f
C23857 a_11322_45546# a_11189_46129# 0.05577f
C23858 a_10490_45724# a_11133_46155# 3.4e-20
C23859 a_n2433_44484# a_n1613_43370# 0.29864f
C23860 a_8975_43940# a_4883_46098# 0.018394f
C23861 a_n2661_42834# a_n1151_42308# 0.038196f
C23862 a_21855_43396# a_21887_42336# 1.39e-19
C23863 a_22591_43396# a_13258_32519# 1.79e-20
C23864 a_10796_42968# a_10723_42308# 0.003077f
C23865 a_10835_43094# a_11323_42473# 3.74e-19
C23866 a_13467_32519# a_22775_42308# 0.016923f
C23867 a_n2293_42282# a_3318_42354# 0.01699f
C23868 a_10341_42308# a_9885_42558# 0.003164f
C23869 a_4361_42308# a_21613_42308# 0.001002f
C23870 a_5649_42852# a_7174_31319# 0.025928f
C23871 a_1793_42852# a_1606_42308# 2.01e-20
C23872 a_10518_42984# a_5742_30871# 0.001042f
C23873 a_n2312_39304# a_n2472_46634# 0.016291f
C23874 a_n2312_40392# a_n2442_46660# 5.91846f
C23875 a_12465_44636# a_n743_46660# 0.026136f
C23876 a_4791_45118# a_5263_46660# 0.001102f
C23877 a_2063_45854# a_10150_46912# 0.008885f
C23878 a_n1151_42308# a_8145_46902# 3.91e-20
C23879 a_6545_47178# a_6540_46812# 0.013617f
C23880 a_6491_46660# a_5732_46660# 6.78e-19
C23881 a_18911_45144# a_11341_43940# 2.97e-20
C23882 a_21101_45002# a_19862_44208# 0.00117f
C23883 a_11691_44458# a_18079_43940# 4.05e-20
C23884 a_11827_44484# a_15493_43396# 0.00117f
C23885 a_7499_43078# a_5755_42852# 2.12e-20
C23886 C4_N_btm VDD 0.265463f
C23887 a_3065_45002# a_3626_43646# 0.480498f
C23888 a_n913_45002# a_9396_43370# 9.91e-20
C23889 a_3232_43370# a_4905_42826# 4.37e-21
C23890 a_3537_45260# a_2982_43646# 7.1e-19
C23891 a_11963_45334# VDD 0.229584f
C23892 a_1606_42308# CAL_P 0.00911f
C23893 a_n1630_35242# a_n1838_35608# 0.00968f
C23894 a_n784_42308# EN_VIN_BSTR_P 0.051272f
C23895 a_8191_45002# a_8049_45260# 0.084237f
C23896 a_10903_45394# a_2324_44458# 3.37e-19
C23897 a_375_42282# a_526_44458# 0.007075f
C23898 a_16241_44484# a_6755_46942# 9.75e-20
C23899 a_n2661_42282# a_5807_45002# 1.81e-19
C23900 a_n4318_39768# a_n2312_38680# 0.023285f
C23901 a_10949_43914# a_768_44030# 0.007821f
C23902 a_18287_44626# a_17339_46660# 0.018815f
C23903 a_n2433_44484# a_n2293_46098# 1.34e-21
C23904 a_11827_44484# a_3483_46348# 0.060892f
C23905 a_584_46384# VDD 2.50905f
C23906 a_15803_42450# a_15959_42545# 0.110532f
C23907 a_15764_42576# a_15890_42674# 0.181217f
C23908 a_7963_42308# a_7174_31319# 4.88e-21
C23909 a_1606_42308# a_1736_39587# 1.72e-20
C23910 a_n3674_38680# a_n3690_38528# 0.071909f
C23911 a_n4318_38216# a_n4334_38528# 5.87e-19
C23912 a_15486_42560# a_15720_42674# 0.006453f
C23913 COMP_P comp_n 0.033828f
C23914 a_20916_46384# a_11415_45002# 7.86e-20
C23915 a_19594_46812# a_12741_44636# 6.75e-20
C23916 a_10467_46802# a_11813_46116# 2.89e-19
C23917 a_10249_46116# a_10768_47026# 0.027091f
C23918 a_6755_46942# a_8846_46660# 8.14e-19
C23919 a_10428_46928# a_11901_46660# 0.004685f
C23920 a_n881_46662# a_2804_46116# 0.050669f
C23921 a_n1613_43370# a_3147_46376# 0.004069f
C23922 a_4883_46098# a_11387_46155# 0.010865f
C23923 a_13507_46334# a_12005_46116# 2.73e-19
C23924 a_16327_47482# a_18819_46122# 0.324239f
C23925 a_10227_46804# a_15682_46116# 0.001531f
C23926 a_11599_46634# a_19900_46494# 0.055271f
C23927 a_17591_47464# a_17583_46090# 6.37e-19
C23928 a_13717_47436# a_10809_44734# 0.004969f
C23929 a_13487_47204# a_6945_45028# 0.015556f
C23930 a_n1151_42308# a_5066_45546# 0.5423f
C23931 a_2998_44172# a_1443_43940# 7.55e-21
C23932 a_n2661_42834# a_6197_43396# 1.61e-19
C23933 a_n356_44636# a_14205_43396# 6.46e-21
C23934 a_10193_42453# a_15959_42545# 1.6e-19
C23935 a_2711_45572# a_20107_42308# 0.164316f
C23936 a_2675_43914# a_2455_43940# 0.007392f
C23937 a_2479_44172# a_3353_43940# 4.3e-20
C23938 a_7499_43078# a_10149_42308# 3.73e-19
C23939 a_11823_42460# a_13249_42558# 0.004086f
C23940 a_20193_45348# a_22591_43396# 0.001393f
C23941 a_n1059_45260# a_13291_42460# 0.03043f
C23942 a_n2017_45002# a_14635_42282# 0.025779f
C23943 a_3537_45260# a_5837_42852# 0.042825f
C23944 a_n913_45002# a_13003_42852# 0.026478f
C23945 a_18588_44850# VDD 0.132317f
C23946 a_7499_43078# a_11652_45724# 1.11e-20
C23947 a_7227_45028# a_8697_45822# 3.36e-20
C23948 a_10193_42453# a_8746_45002# 0.11003f
C23949 a_2711_45572# a_9159_45572# 0.003753f
C23950 a_10180_45724# a_10490_45724# 7.31e-21
C23951 a_15493_43940# a_20202_43084# 0.02138f
C23952 a_22223_43948# a_11415_45002# 9.62e-19
C23953 a_13467_32519# a_12549_44172# 3.15e-20
C23954 a_14401_32519# a_19692_46634# 4.68e-19
C23955 a_9313_44734# a_20205_31679# 1.02e-20
C23956 a_13468_44734# a_13259_45724# 0.004213f
C23957 a_2127_44172# a_2324_44458# 0.00237f
C23958 a_n2293_42282# a_n1151_42308# 3.68e-19
C23959 a_11901_46660# VDD 0.57548f
C23960 a_1606_42308# CAL_N 0.006757f
C23961 a_376_46348# a_1176_45822# 0.001135f
C23962 a_n2293_46098# a_3147_46376# 1.09e-19
C23963 a_472_46348# a_1208_46090# 0.088629f
C23964 a_2609_46660# a_3503_45724# 2.66e-19
C23965 a_2959_46660# a_3218_45724# 1.15e-19
C23966 a_765_45546# a_2324_44458# 5.17e-20
C23967 a_14035_46660# a_10809_44734# 0.00805f
C23968 a_14513_46634# a_6945_45028# 3.51e-20
C23969 a_17339_46660# a_15682_46116# 2.86e-19
C23970 a_6123_31319# VDAC_Ni 4.39e-19
C23971 a_9313_44734# a_16328_43172# 1.1e-19
C23972 a_3905_42865# a_5111_42852# 0.079376f
C23973 a_18079_43940# a_4190_30871# 4.22e-21
C23974 a_11750_44172# a_4361_42308# 1.32e-21
C23975 a_17737_43940# a_743_42282# 9.59e-21
C23976 a_n97_42460# a_6031_43396# 0.002248f
C23977 a_14021_43940# a_16547_43609# 0.005885f
C23978 a_3422_30871# a_17333_42852# 1.02e-20
C23979 a_742_44458# a_2713_42308# 7.64e-19
C23980 a_1756_43548# a_1987_43646# 0.004999f
C23981 a_15493_43940# a_16867_43762# 6.77e-19
C23982 a_n2810_45028# a_n4209_38216# 0.063751f
C23983 SMPL_ON_P EN_VIN_BSTR_P 1.58e-19
C23984 a_n144_43396# VDD 3.23e-19
C23985 a_15765_45572# a_16019_45002# 0.001223f
C23986 a_15599_45572# a_16751_45260# 0.012353f
C23987 a_8696_44636# a_14180_45002# 5.97e-21
C23988 a_2711_45572# a_16237_45028# 0.001569f
C23989 a_16680_45572# a_14537_43396# 3.12e-20
C23990 a_11652_45724# a_11915_45394# 6.1e-19
C23991 a_15903_45785# a_1307_43914# 8.62e-19
C23992 a_4958_30871# a_16327_47482# 2.84e-19
C23993 a_17124_42282# a_10227_46804# 1.7e-20
C23994 a_n2302_39072# SMPL_ON_P 5.6e-20
C23995 a_9145_43396# a_10809_44734# 4.72e-20
C23996 a_8685_42308# a_n1613_43370# 0.002002f
C23997 a_14401_32519# a_20692_30879# 0.054254f
C23998 a_n3674_37592# a_n2438_43548# 0.001205f
C23999 a_5907_45546# a_n881_46662# 0.070761f
C24000 a_2711_45572# a_8128_46384# 1.58e-19
C24001 a_6194_45824# a_n1613_43370# 2.79e-20
C24002 a_10193_42453# a_4883_46098# 0.040505f
C24003 a_13904_45546# a_10227_46804# 5.42e-19
C24004 a_9159_45572# a_9313_45822# 0.051702f
C24005 a_n1545_46494# a_n2293_45546# 8.21e-20
C24006 a_8049_45260# a_11315_46155# 1.74e-19
C24007 a_13467_32519# a_21855_43396# 0.003525f
C24008 a_21487_43396# a_5649_42852# 8.4e-20
C24009 a_10341_43396# a_10796_42968# 9.03e-20
C24010 a_9145_43396# a_13460_43230# 0.002473f
C24011 a_20512_43084# a_20712_42282# 2.86e-20
C24012 a_4190_30871# a_14209_32519# 0.031783f
C24013 VDAC_N C5_N_btm 27.606901f
C24014 a_1307_43914# a_n2661_44458# 0.007888f
C24015 a_7499_43078# a_7845_44172# 0.112307f
C24016 a_6171_45002# a_10057_43914# 1.53e-19
C24017 a_3232_43370# a_8975_43940# 0.620589f
C24018 a_n967_45348# a_n356_44636# 2.16e-20
C24019 a_8191_45002# a_8103_44636# 2.19e-19
C24020 a_5379_42460# a_4185_45028# 0.189676f
C24021 a_8605_42826# a_n443_42852# 0.001815f
C24022 a_12895_43230# a_n357_42282# 0.00578f
C24023 a_1606_42308# a_8199_44636# 2.7e-20
C24024 a_n784_42308# a_10903_43370# 1.58e-20
C24025 a_3080_42308# EN_VIN_BSTR_P 0.043903f
C24026 a_14401_32519# VIN_N 0.03172f
C24027 a_21588_30879# C5_N_btm 5.07e-20
C24028 a_18911_45144# a_16327_47482# 3.79e-19
C24029 C6_P_btm VDD 0.210613f
C24030 a_n2661_44458# a_n443_46116# 0.034876f
C24031 a_n1352_44484# a_n1151_42308# 0.001499f
C24032 a_4223_44672# a_2063_45854# 1.1e-20
C24033 a_n699_43396# a_584_46384# 0.632931f
C24034 a_7276_45260# a_n1925_46634# 8.36e-22
C24035 a_3537_45260# a_2107_46812# 1.32e-20
C24036 a_n37_45144# a_n2661_46098# 1.2e-20
C24037 a_413_45260# a_1799_45572# 7.25e-20
C24038 a_3357_43084# a_6540_46812# 0.001035f
C24039 a_16115_45572# a_15368_46634# 6.95e-20
C24040 a_15415_45028# a_5807_45002# 1.7e-21
C24041 a_14797_45144# a_13661_43548# 0.116989f
C24042 a_10775_45002# a_n2661_46634# 3.04e-22
C24043 a_16680_45572# a_3090_45724# 0.009229f
C24044 a_13527_45546# a_765_45546# 2.42e-21
C24045 a_14537_43396# a_13747_46662# 0.006836f
C24046 a_6194_45824# a_n2293_46098# 2.86e-19
C24047 a_16547_43609# a_15764_42576# 2.95e-21
C24048 a_16243_43396# a_15803_42450# 2.1e-20
C24049 a_3681_42891# a_n784_42308# 1.66e-21
C24050 a_17333_42852# a_18504_43218# 0.157683f
C24051 a_16137_43396# a_15959_42545# 0.001471f
C24052 a_5649_42852# a_5932_42308# 0.126438f
C24053 a_4361_42308# a_6761_42308# 0.042179f
C24054 a_743_42282# a_8515_42308# 0.005514f
C24055 a_15567_42826# a_16245_42852# 0.03084f
C24056 a_18083_42858# a_18695_43230# 0.001881f
C24057 a_10341_43396# a_4958_30871# 4.26e-20
C24058 a_n3690_38528# VDD 0.363159f
C24059 a_3422_30871# a_7754_38470# 6.77e-20
C24060 a_6151_47436# a_13569_47204# 0.004336f
C24061 a_9863_47436# a_10037_47542# 0.006584f
C24062 a_13717_47436# a_n881_46662# 0.039579f
C24063 a_9313_45822# a_8128_46384# 0.013269f
C24064 a_n452_47436# a_n743_46660# 6.22e-21
C24065 a_n971_45724# a_n1021_46688# 0.002801f
C24066 a_n2109_47186# a_383_46660# 2.96e-20
C24067 a_n1741_47186# a_33_46660# 4.45e-20
C24068 a_n815_47178# a_n2438_43548# 1.87e-19
C24069 a_n746_45260# a_n1925_46634# 0.036469f
C24070 a_1239_47204# a_n2661_46634# 0.002062f
C24071 a_21177_47436# a_12465_44636# 2.23e-19
C24072 a_19386_47436# a_11453_44696# 1.38e-19
C24073 a_21496_47436# a_4883_46098# 0.257837f
C24074 a_13507_46334# a_21811_47423# 4.35e-19
C24075 a_13348_45260# a_11341_43940# 1.4e-21
C24076 a_22959_45036# a_19237_31679# 0.005799f
C24077 a_10193_42453# a_16243_43396# 2.07e-19
C24078 a_13249_42308# a_12281_43396# 1.91e-19
C24079 a_2711_45572# a_743_42282# 0.039036f
C24080 a_8375_44464# a_8333_44734# 7.47e-21
C24081 a_12883_44458# a_13296_44484# 5.31e-19
C24082 a_12607_44458# a_13940_44484# 5.31e-19
C24083 a_5891_43370# a_8238_44734# 9.85e-19
C24084 a_n2661_43370# a_n4318_39768# 0.068386f
C24085 a_n1821_44484# a_n2661_42834# 0.001026f
C24086 a_2382_45260# a_3737_43940# 0.027805f
C24087 a_6171_45002# a_14021_43940# 5.61e-20
C24088 a_1307_43914# a_2804_46116# 3.01e-21
C24089 a_1423_45028# a_1138_42852# 7.83e-19
C24090 a_16922_45042# a_765_45546# 6.35e-21
C24091 a_19279_43940# a_5807_45002# 4.49e-20
C24092 a_20640_44752# a_19321_45002# 0.034599f
C24093 a_16979_44734# a_6755_46942# 0.00119f
C24094 a_20835_44721# a_13747_46662# 0.006757f
C24095 a_9838_44484# a_8270_45546# 4.89e-20
C24096 a_17478_45572# a_16375_45002# 0.009252f
C24097 a_2437_43646# a_526_44458# 0.005693f
C24098 a_10775_45002# a_8199_44636# 0.064568f
C24099 a_n2840_43914# a_n1613_43370# 6.54e-20
C24100 a_8953_45002# a_5937_45572# 0.062333f
C24101 a_6171_45002# a_11133_46155# 4.63e-21
C24102 a_2382_45260# a_2324_44458# 0.044897f
C24103 a_3232_43370# a_11387_46155# 3.73e-20
C24104 a_1443_43940# a_n2497_47436# 1.71e-19
C24105 a_6171_42473# a_5934_30871# 1.01e-20
C24106 a_1606_42308# a_13070_42354# 1.69e-20
C24107 a_n1386_35608# a_n83_35174# 0.081924f
C24108 a_n1532_35090# EN_VIN_BSTR_P 0.340449f
C24109 a_3785_47178# a_4419_46090# 2.07e-20
C24110 a_5807_45002# a_15368_46634# 0.029781f
C24111 a_13747_46662# a_3090_45724# 0.139869f
C24112 a_2107_46812# a_6969_46634# 2.09e-19
C24113 a_3877_44458# a_6540_46812# 0.244975f
C24114 a_4646_46812# a_5732_46660# 0.050752f
C24115 a_4651_46660# a_5907_46634# 0.043482f
C24116 a_4817_46660# a_5385_46902# 0.170485f
C24117 a_13661_43548# a_14976_45028# 0.162789f
C24118 a_4955_46873# a_5167_46660# 0.003269f
C24119 a_n2661_46634# a_11186_47026# 0.002094f
C24120 a_12891_46348# a_12359_47026# 0.002172f
C24121 a_n1925_46634# a_8189_46660# 1.2e-19
C24122 a_n881_46662# a_14035_46660# 9.06e-20
C24123 a_2063_45854# a_6419_46155# 1.49e-19
C24124 a_3160_47472# a_5164_46348# 9.48e-21
C24125 a_n1741_47186# a_12005_46116# 0.174477f
C24126 a_n1151_42308# a_5068_46348# 0.089946f
C24127 a_n237_47217# a_9823_46155# 4.34e-20
C24128 a_n443_46116# a_2804_46116# 0.018109f
C24129 a_n1435_47204# a_n1853_46287# 2.54e-20
C24130 a_10227_46804# a_20719_46660# 3.17e-19
C24131 a_18597_46090# a_18280_46660# 3.97e-19
C24132 a_21496_47436# a_21188_46660# 2.45e-19
C24133 a_4883_46098# a_21363_46634# 0.066909f
C24134 a_20990_47178# a_20731_47026# 6.38e-19
C24135 a_13507_46334# a_22000_46634# 0.183978f
C24136 a_11453_44696# a_19551_46910# 0.047386f
C24137 a_12465_44636# a_20841_46902# 3.04e-20
C24138 a_5111_44636# a_4520_42826# 1.98e-19
C24139 a_n1059_45260# a_13460_43230# 0.004971f
C24140 a_n913_45002# a_13635_43156# 0.036742f
C24141 a_3537_45260# a_7871_42858# 8.33e-19
C24142 a_3232_43370# a_2905_42968# 0.008509f
C24143 a_5147_45002# a_5111_42852# 1.57e-20
C24144 a_n2661_42834# a_8415_44056# 1.54e-35
C24145 a_20766_44850# a_19862_44208# 1.08e-19
C24146 a_n699_43396# a_n144_43396# 1.99e-19
C24147 a_n2661_44458# a_9396_43370# 1.17e-21
C24148 a_19279_43940# a_19478_44306# 0.03583f
C24149 a_18579_44172# a_18451_43940# 0.147572f
C24150 a_14673_44172# a_14021_43940# 4.52e-19
C24151 a_5495_43940# a_5663_43940# 0.227135f
C24152 a_20640_44752# a_20623_43914# 0.003088f
C24153 a_19615_44636# a_11341_43940# 2.34e-21
C24154 a_18911_45144# a_10341_43396# 2.05e-21
C24155 a_18443_44721# VDD 0.193515f
C24156 a_n4064_39616# C4_P_btm 6.79e-20
C24157 a_n3420_39616# C2_P_btm 2.28e-20
C24158 a_n4064_39072# a_n923_35174# 0.007158f
C24159 a_15433_44458# a_2324_44458# 0.021739f
C24160 a_11827_44484# a_n357_42282# 1.01e-20
C24161 a_18114_32519# a_20205_31679# 0.051478f
C24162 a_20269_44172# a_3090_45724# 1.17e-19
C24163 a_2982_43646# a_n2293_46634# 0.015801f
C24164 a_479_46660# VDD 1.63e-19
C24165 a_n4064_40160# a_n4334_38304# 0.013157f
C24166 a_n2946_39072# a_n2302_39072# 6.68e-19
C24167 a_n3690_39392# a_n3607_39392# 0.007692f
C24168 a_5742_30871# C5_N_btm 0.089375f
C24169 a_21363_46634# a_21188_46660# 0.233657f
C24170 a_18285_46348# a_18900_46660# 0.004259f
C24171 a_20273_46660# a_20731_47026# 0.027606f
C24172 a_19123_46287# a_18280_46660# 8.18e-20
C24173 a_5807_45002# a_19597_46482# 1.86e-20
C24174 a_2107_46812# a_9241_46436# 2.55e-19
C24175 a_n743_46660# a_10037_46155# 3.34e-19
C24176 a_n881_46662# a_n1099_45572# 0.088565f
C24177 a_6755_46942# a_14275_46494# 1.11e-19
C24178 a_10623_46897# a_2324_44458# 1.46e-20
C24179 a_8270_45546# a_9823_46155# 3.17e-19
C24180 a_n1613_43370# a_310_45028# 1.46e-20
C24181 a_n4318_37592# a_n4064_37984# 0.050508f
C24182 a_n3674_38216# a_n4251_38304# 8.42e-19
C24183 a_3090_45724# a_4419_46090# 0.001764f
C24184 a_10729_43914# a_8685_43396# 5.97e-22
C24185 a_1443_43940# a_1568_43370# 4.63e-19
C24186 a_n2293_43922# a_10796_42968# 2.47e-20
C24187 a_9313_44734# a_15279_43071# 0.007423f
C24188 a_3422_30871# a_13678_32519# 0.452533f
C24189 a_20512_43084# a_20556_43646# 9.96e-19
C24190 a_18184_42460# a_19326_42852# 1.25e-20
C24191 a_n2017_45002# a_19511_42282# 6.66e-20
C24192 en_comp a_18907_42674# 1.94e-20
C24193 a_n1059_45260# a_18548_42308# 0.001247f
C24194 a_5025_43940# VDD 0.004306f
C24195 a_10180_45724# a_6171_45002# 0.03378f
C24196 a_10193_42453# a_3232_43370# 0.016241f
C24197 a_18479_45785# a_18909_45814# 0.023226f
C24198 a_18175_45572# a_18691_45572# 0.105995f
C24199 a_5907_45546# a_1307_43914# 2.22e-20
C24200 a_8147_43396# a_3483_46348# 2.1e-21
C24201 a_14955_43396# a_12741_44636# 6.28e-23
C24202 a_7287_43370# a_4185_45028# 1.18e-21
C24203 a_3457_43396# a_1823_45246# 9.91e-20
C24204 a_19268_43646# a_17339_46660# 0.003554f
C24205 a_22223_43396# a_19692_46634# 0.001051f
C24206 a_n2661_42282# a_n755_45592# 0.025718f
C24207 a_n2104_42282# a_n2312_39304# 3.28e-20
C24208 a_n3674_38216# a_n2312_40392# 0.025514f
C24209 COMP_P SMPL_ON_N 2.13516f
C24210 a_4338_37500# RST_Z 0.01719f
C24211 VDAC_P C7_P_btm 0.11042p
C24212 a_17583_46090# VDD 0.23578f
C24213 a_2711_45572# a_6151_47436# 0.050517f
C24214 a_9049_44484# a_n971_45724# 1.51e-21
C24215 a_8568_45546# a_n237_47217# 1.04e-19
C24216 a_6194_45824# a_4791_45118# 0.004919f
C24217 a_3260_45572# a_2063_45854# 5.14e-21
C24218 a_n3565_38216# a_n2946_37690# 0.001566f
C24219 a_n4209_38216# a_n2302_37690# 0.001686f
C24220 a_n4334_38304# a_n4064_37440# 7.84e-19
C24221 a_n2293_46098# a_310_45028# 0.017313f
C24222 a_472_46348# a_n2661_45546# 2.09e-20
C24223 a_n901_46420# a_n2293_45546# 1.79e-20
C24224 a_n2157_46122# a_n1099_45572# 1.52e-19
C24225 a_14275_46494# a_8049_45260# 0.001971f
C24226 a_11387_46155# a_11608_46482# 0.007833f
C24227 a_10341_43396# a_15125_43396# 7.22e-20
C24228 a_9313_44734# a_13258_32519# 0.003166f
C24229 a_3422_30871# a_6123_31319# 0.021957f
C24230 a_n3674_39768# a_n4318_37592# 0.023075f
C24231 a_14401_32519# a_5342_30871# 0.062032f
C24232 a_n97_42460# a_10796_42968# 3.04e-19
C24233 a_3080_42308# a_3681_42891# 5.97e-19
C24234 a_4235_43370# a_4520_42826# 0.001794f
C24235 a_16137_43396# a_16243_43396# 0.182209f
C24236 a_19321_45002# START 0.10793f
C24237 a_19594_46812# RST_Z 3.35e-20
C24238 a_8952_43230# VDD 0.273404f
C24239 a_10775_45002# a_10903_45394# 0.004764f
C24240 a_7229_43940# a_n2661_43370# 0.040132f
C24241 a_19479_31679# a_18114_32519# 0.182316f
C24242 a_22223_45572# a_19721_31679# 8.73e-19
C24243 a_6171_45002# a_13711_45394# 9.69e-20
C24244 a_13887_32519# a_20205_31679# 0.051379f
C24245 a_22400_42852# a_21076_30879# 1.76e-19
C24246 a_20273_45572# a_20916_46384# 9.09e-20
C24247 a_8568_45546# a_8270_45546# 0.015327f
C24248 a_11823_42460# a_6755_46942# 3.55e-19
C24249 a_20731_45938# a_13747_46662# 2.78e-19
C24250 a_19365_45572# a_13661_43548# 9.66e-20
C24251 a_19610_45572# a_5807_45002# 7.29e-19
C24252 a_2437_43646# a_13759_47204# 8.24e-20
C24253 a_n1059_45260# a_n881_46662# 0.121542f
C24254 a_n913_45002# a_n1613_43370# 0.686014f
C24255 a_413_45260# a_2747_46873# 0.038809f
C24256 a_5691_45260# a_4883_46098# 5.88e-21
C24257 a_10951_45334# a_10227_46804# 0.001109f
C24258 a_14537_43396# a_11599_46634# 6.07e-21
C24259 a_6171_45002# a_13507_46334# 5.79e-20
C24260 a_n2661_43370# a_n237_47217# 3.56e-19
C24261 a_5093_45028# a_n1151_42308# 1.96e-21
C24262 a_8791_43396# a_8685_42308# 1.69e-21
C24263 a_20974_43370# a_13258_32519# 7.54e-21
C24264 a_17595_43084# a_17701_42308# 0.141211f
C24265 a_n97_42460# a_4958_30871# 0.069553f
C24266 a_16795_42852# a_18083_42858# 6.33e-21
C24267 a_3626_43646# a_13575_42558# 0.008305f
C24268 a_5111_42852# a_5457_43172# 0.013377f
C24269 a_16414_43172# a_17333_42852# 2.98e-20
C24270 a_3483_46348# DATA[2] 6.68e-19
C24271 a_4915_47217# a_n1435_47204# 0.038318f
C24272 a_7227_47204# a_6575_47204# 0.028925f
C24273 a_6151_47436# a_9313_45822# 0.032544f
C24274 a_n1151_42308# a_15811_47375# 1.38e-21
C24275 a_n2810_45028# a_n2661_42282# 2.09e-20
C24276 a_20528_45572# a_20365_43914# 4.03e-21
C24277 a_3232_43370# a_5495_43940# 0.060353f
C24278 a_5691_45260# a_5663_43940# 4.64e-21
C24279 a_n2129_44697# a_7_44811# 1.23e-19
C24280 a_n2433_44484# a_n1243_44484# 2.56e-19
C24281 a_20193_45348# a_9313_44734# 0.056112f
C24282 a_n1917_44484# a_n356_44636# 1.7e-20
C24283 a_15037_45618# a_15037_43940# 1.4e-21
C24284 a_3497_42558# a_n755_45592# 2.25e-19
C24285 a_13678_32519# VREF_GND 0.047887f
C24286 a_13249_42308# VDD 0.653917f
C24287 a_11541_44484# a_11453_44696# 0.004713f
C24288 a_12829_44484# a_12465_44636# 3.05e-19
C24289 a_19615_44636# a_16327_47482# 6.71e-19
C24290 a_n1549_44318# a_n1151_42308# 5.94e-21
C24291 a_1467_44172# a_584_46384# 0.005691f
C24292 a_n4318_39768# a_n2497_47436# 3e-20
C24293 a_11823_42460# a_8049_45260# 0.046281f
C24294 a_10490_45724# a_10586_45546# 0.235237f
C24295 a_556_44484# a_n1613_43370# 3.24e-20
C24296 a_n2293_45010# a_n1423_46090# 1.94e-19
C24297 a_413_45260# a_20202_43084# 3.33e-20
C24298 a_3357_43084# a_1823_45246# 0.062163f
C24299 a_14539_43914# a_n2293_46634# 0.045317f
C24300 a_7640_43914# a_768_44030# 0.036222f
C24301 a_949_44458# a_n2661_46098# 4.97e-22
C24302 a_13777_45326# a_13059_46348# 0.00155f
C24303 a_n1059_45260# a_n2157_46122# 8.24e-19
C24304 a_n2661_45010# a_n901_46420# 8.48e-21
C24305 a_n2661_43370# a_8270_45546# 0.022558f
C24306 a_n4318_38680# a_n3690_38528# 1.96e-19
C24307 a_10793_43218# a_5742_30871# 4.83e-21
C24308 a_n784_42308# a_n327_42558# 5.3e-19
C24309 a_n961_42308# a_n1630_35242# 0.028868f
C24310 a_196_42282# a_n3674_37592# 0.1528f
C24311 a_19164_43230# a_19511_42282# 0.001746f
C24312 a_19339_43156# a_19647_42308# 0.009735f
C24313 a_17333_42852# a_7174_31319# 7.1e-21
C24314 a_n1925_46634# a_383_46660# 0.009919f
C24315 a_n743_46660# a_33_46660# 0.025563f
C24316 a_n2438_43548# a_171_46873# 0.029723f
C24317 a_n2661_46634# a_491_47026# 0.003523f
C24318 a_n2293_46634# a_2107_46812# 3.61e-19
C24319 a_n1613_43370# a_5894_47026# 5.16e-19
C24320 a_10227_46804# a_11735_46660# 0.54163f
C24321 a_11599_46634# a_3090_45724# 0.133107f
C24322 a_15811_47375# a_14084_46812# 7.3e-20
C24323 a_4915_47217# a_13885_46660# 0.179458f
C24324 a_12861_44030# a_16292_46812# 0.059827f
C24325 a_n1151_42308# a_13059_46348# 0.003065f
C24326 a_1239_47204# a_765_45546# 9.93e-19
C24327 a_9482_43914# a_9885_43646# 7.99e-20
C24328 a_13556_45296# a_14955_43396# 8.22e-21
C24329 a_18374_44850# a_15493_43940# 4.07e-21
C24330 a_1423_45028# a_8685_43396# 1.34e-21
C24331 a_1307_43914# a_9145_43396# 0.003867f
C24332 a_14537_43396# a_14358_43442# 0.1418f
C24333 a_20193_45348# a_20974_43370# 0.026944f
C24334 a_21398_44850# a_21145_44484# 4.61e-19
C24335 a_3422_30871# a_21073_44484# 3.97e-20
C24336 a_4223_44672# a_5326_44056# 4.3e-19
C24337 a_n2661_43922# a_2253_44260# 3.34e-19
C24338 a_n2661_42834# a_2537_44260# 1.37e-19
C24339 a_n2293_42834# a_548_43396# 2.62e-19
C24340 a_19479_31679# a_13887_32519# 0.051118f
C24341 a_19963_31679# a_13678_32519# 0.051335f
C24342 a_n2216_37984# VDD 0.003985f
C24343 a_17613_45144# VDD 0.094022f
C24344 a_5934_30871# VIN_N 0.009408f
C24345 a_5742_30871# C5_P_btm 0.089375f
C24346 a_6123_31319# VREF_GND 0.00207f
C24347 a_n2661_42834# a_12741_44636# 5.02e-19
C24348 a_19319_43548# a_12549_44172# 0.024381f
C24349 a_20512_43084# a_19692_46634# 0.387138f
C24350 a_501_45348# a_n863_45724# 2.59e-19
C24351 a_2304_45348# a_n2661_45546# 0.004487f
C24352 a_8953_45002# a_n443_42852# 2.1e-20
C24353 a_5343_44458# a_2324_44458# 0.255488f
C24354 a_10057_43914# a_10903_43370# 0.052284f
C24355 a_n4318_39304# a_n1613_43370# 3.19e-20
C24356 a_2982_43646# a_18597_46090# 0.239147f
C24357 a_21887_42336# a_21613_42308# 0.071168f
C24358 a_5742_30871# a_n3420_38528# 0.004679f
C24359 a_19511_42282# a_21973_42336# 1.79e-19
C24360 a_3877_44458# a_1823_45246# 0.231164f
C24361 a_15559_46634# a_14513_46634# 2.81e-20
C24362 a_14084_46812# a_13059_46348# 5.17e-19
C24363 a_15009_46634# a_15227_46910# 0.08213f
C24364 a_11186_47026# a_765_45546# 5.79e-19
C24365 a_n881_46662# a_n1925_42282# 0.041426f
C24366 a_19321_45002# a_19553_46090# 0.008717f
C24367 a_13747_46662# a_20075_46420# 1.64e-20
C24368 a_n743_46660# a_12005_46116# 0.024033f
C24369 a_2107_46812# a_9625_46129# 0.184645f
C24370 a_19594_46812# a_18985_46122# 9.08e-20
C24371 a_16942_47570# a_6945_45028# 1.33e-19
C24372 a_5807_45002# a_20708_46348# 1.89e-19
C24373 a_3160_47472# a_3316_45546# 0.003495f
C24374 a_n1151_42308# a_3218_45724# 5.24e-20
C24375 a_2905_45572# a_3503_45724# 0.001385f
C24376 a_n443_46116# a_n1099_45572# 0.368941f
C24377 a_11599_46634# a_15002_46116# 4.2e-19
C24378 a_10227_46804# a_14537_46482# 0.001903f
C24379 a_4883_46098# a_11387_46482# 2.91e-19
C24380 a_n913_45002# a_3905_42558# 0.047606f
C24381 a_2382_45260# a_1606_42308# 1.35e-20
C24382 a_n2017_45002# a_4921_42308# 0.006208f
C24383 a_2479_44172# a_3626_43646# 3.71e-20
C24384 a_5891_43370# a_4361_42308# 0.028094f
C24385 a_11827_44484# a_21356_42826# 5.05e-21
C24386 a_5495_43940# a_4905_42826# 0.001789f
C24387 a_2889_44172# a_2896_43646# 0.001151f
C24388 a_644_44056# a_648_43396# 2.15e-19
C24389 a_19615_44636# a_10341_43396# 2.09e-21
C24390 a_8103_44636# a_7765_42852# 4.51e-20
C24391 a_n1441_43940# VDD 0.142719f
C24392 a_10193_42453# a_18341_45572# 6.23e-22
C24393 a_11064_45572# a_11136_45572# 0.003395f
C24394 a_13163_45724# a_13485_45572# 0.001367f
C24395 a_11823_42460# a_14127_45572# 3.38e-19
C24396 a_n961_42308# a_n971_45724# 3.58e-20
C24397 a_22485_44484# a_20205_31679# 2.08e-20
C24398 a_15493_43940# a_17715_44484# 0.005403f
C24399 a_14021_43940# a_10903_43370# 2.56e-21
C24400 a_7871_42858# a_n2293_46634# 6.83e-20
C24401 a_5649_42852# a_4646_46812# 1.19e-20
C24402 a_14358_43442# a_3090_45724# 6.05e-19
C24403 a_16104_42674# CAL_N 1.8e-20
C24404 a_376_46348# a_518_46482# 0.007833f
C24405 a_16388_46812# a_16375_45002# 0.039999f
C24406 a_3090_45724# a_1848_45724# 3.59e-19
C24407 a_11189_46129# a_12005_46116# 0.00104f
C24408 a_11133_46155# a_10903_43370# 2.09e-20
C24409 a_9290_44172# a_12594_46348# 1.22e-21
C24410 a_9396_43370# a_9145_43396# 0.030617f
C24411 a_11341_43940# a_10835_43094# 1.05e-19
C24412 a_5891_43370# a_6761_42308# 0.010358f
C24413 a_18114_32519# a_13258_32519# 0.059438f
C24414 a_20974_43370# a_20301_43646# 9.11e-21
C24415 a_3905_42865# a_3863_42891# 1.54e-19
C24416 a_17538_32519# a_4190_30871# 1.16e-20
C24417 a_20193_45348# a_22397_42558# 0.00176f
C24418 a_11459_47204# CLK 7.93e-19
C24419 a_n1435_47204# DATA[5] 0.031859f
C24420 a_15673_47210# RST_Z 1.57e-19
C24421 a_19700_43370# VDD 0.28578f
C24422 a_4927_45028# a_6171_45002# 8.82e-20
C24423 a_3537_45260# a_6709_45028# 5.94e-20
C24424 a_5147_45002# a_5205_44484# 0.018671f
C24425 a_5691_45260# a_3232_43370# 0.123939f
C24426 a_n1059_45260# a_1307_43914# 0.016622f
C24427 a_8746_45002# a_10057_43914# 0.003098f
C24428 a_15765_45572# a_11827_44484# 1.86e-20
C24429 a_10193_42453# a_8975_43940# 0.023559f
C24430 a_12089_42308# a_4185_45028# 3.84e-20
C24431 a_5379_42460# a_5257_43370# 7.23e-20
C24432 a_17749_42852# a_15227_44166# 0.00177f
C24433 a_8147_43396# a_n357_42282# 8.81e-19
C24434 a_3626_43646# a_n443_42852# 0.027303f
C24435 a_8605_42826# a_8199_44636# 1.4e-21
C24436 a_7765_42852# a_8953_45546# 3.74e-21
C24437 a_16147_45260# a_12465_44636# 2.41e-21
C24438 a_18479_45785# a_4883_46098# 8.72e-20
C24439 a_20841_45814# a_16327_47482# 0.161808f
C24440 a_3357_43084# a_11031_47542# 1.35e-19
C24441 a_2437_43646# a_13381_47204# 0.005327f
C24442 a_413_45260# a_2063_45854# 0.031952f
C24443 a_327_44734# a_584_46384# 0.040089f
C24444 a_4574_45260# a_n237_47217# 3.04e-20
C24445 a_n1059_45260# a_n443_46116# 3.62e-19
C24446 a_n913_45002# a_4791_45118# 0.254334f
C24447 a_15599_45572# a_n881_46662# 0.601034f
C24448 a_10490_45724# a_n743_46660# 2.02e-20
C24449 a_n2840_45546# a_n2661_45546# 0.175179f
C24450 a_n2661_42282# a_n2302_40160# 1.84e-20
C24451 a_14021_43940# a_15959_42545# 4.7e-21
C24452 a_1049_43396# a_1184_42692# 3.77e-21
C24453 a_n1557_42282# a_n473_42460# 0.077371f
C24454 a_743_42282# a_18817_42826# 1.5e-20
C24455 a_4361_42308# a_17595_43084# 3.75e-20
C24456 a_5649_42852# a_15567_42826# 8.45e-21
C24457 a_4905_42826# a_n784_42308# 3.17e-21
C24458 a_4190_30871# a_19339_43156# 0.002519f
C24459 a_19095_43396# a_18083_42858# 2.56e-19
C24460 a_1568_43370# a_1576_42282# 9.29e-19
C24461 a_20820_30879# a_22459_39145# 3.4e-20
C24462 a_16388_46812# RST_Z 3.56e-20
C24463 a_7754_38636# a_7754_38470# 0.296258f
C24464 a_7754_40130# a_5700_37509# 0.037095f
C24465 VDAC_Pi a_3726_37500# 1.17174f
C24466 a_7754_39964# a_4338_37500# 0.021449f
C24467 a_2123_42473# VDD 0.1936f
C24468 a_n2497_47436# a_n237_47217# 4.7e-20
C24469 SMPL_ON_P a_n1605_47204# 0.194856f
C24470 a_n1741_47186# a_n815_47178# 0.031488f
C24471 a_n2109_47186# a_n971_45724# 1.21934f
C24472 a_13159_45002# a_13213_44734# 2.87e-19
C24473 a_9482_43914# a_n2661_43922# 0.036658f
C24474 a_11136_45572# a_10807_43548# 5.02e-21
C24475 a_19479_31679# a_22485_44484# 0.001111f
C24476 a_3357_43084# a_20512_43084# 3.36e-21
C24477 a_4921_42308# a_526_44458# 0.002257f
C24478 a_8649_43218# a_n443_42852# 6.31e-19
C24479 a_18907_42674# a_4185_45028# 7.14e-20
C24480 a_10907_45822# a_3483_46348# 0.140023f
C24481 a_15861_45028# a_12741_44636# 0.075863f
C24482 a_n2661_43370# a_1123_46634# 3.92e-21
C24483 a_10775_45002# a_10623_46897# 3.09e-22
C24484 a_10951_45334# a_10467_46802# 2.26e-21
C24485 a_18184_42460# a_19321_45002# 0.094476f
C24486 a_20567_45036# a_13747_46662# 0.026034f
C24487 a_4185_45348# a_3877_44458# 7.28e-19
C24488 a_6709_45028# a_6969_46634# 9.02e-22
C24489 a_7705_45326# a_6755_46942# 1.11e-20
C24490 a_11322_45546# a_9290_44172# 0.077646f
C24491 a_10193_42453# a_11387_46155# 0.050391f
C24492 a_10490_45724# a_11189_46129# 0.03271f
C24493 a_10180_45724# a_10903_43370# 7.78e-20
C24494 a_n2661_44458# a_n1613_43370# 0.05666f
C24495 a_10057_43914# a_4883_46098# 2.16e-19
C24496 a_10083_42826# a_5742_30871# 2.48e-19
C24497 a_10835_43094# a_10723_42308# 0.006083f
C24498 a_10796_42968# a_10533_42308# 8.22e-19
C24499 a_n2293_42282# a_2903_42308# 0.005938f
C24500 a_5649_42852# a_20712_42282# 1.31e-19
C24501 a_13467_32519# a_21613_42308# 0.053076f
C24502 a_13887_32519# a_13258_32519# 0.054157f
C24503 a_5342_30871# a_5934_30871# 0.018148f
C24504 a_13678_32519# a_7174_31319# 7.78e-20
C24505 a_1709_42852# a_1606_42308# 4.98e-19
C24506 a_11309_47204# a_12891_46348# 9.04e-21
C24507 a_n2312_39304# a_n2661_46634# 0.105298f
C24508 a_n2312_40392# a_n2472_46634# 3.86e-20
C24509 a_2063_45854# a_9863_46634# 0.10786f
C24510 a_n1151_42308# a_7577_46660# 0.001579f
C24511 a_6491_46660# a_5907_46634# 0.002903f
C24512 a_6151_47436# a_6540_46812# 0.043688f
C24513 a_6545_47178# a_5732_46660# 1.97e-20
C24514 C3_N_btm VDD 0.26836f
C24515 a_3065_45002# a_3540_43646# 9.54e-20
C24516 a_n1059_45260# a_9396_43370# 1.51e-19
C24517 a_3232_43370# a_3080_42308# 0.001461f
C24518 a_2382_45260# a_3539_42460# 0.110439f
C24519 a_16147_45260# a_16409_43396# 1.28e-21
C24520 a_18184_42460# a_20623_43914# 4.99e-21
C24521 a_18494_42460# a_20365_43914# 0.003336f
C24522 a_11827_44484# a_19328_44172# 0.001549f
C24523 a_11691_44458# a_17973_43940# 3.47e-19
C24524 a_16237_45028# a_15682_43940# 1.42e-19
C24525 a_21005_45260# a_19862_44208# 6.37e-19
C24526 a_18587_45118# a_11341_43940# 1.05e-21
C24527 a_11787_45002# VDD 0.153399f
C24528 COMP_P a_18194_35068# 5.47e-19
C24529 a_n784_42308# a_n923_35174# 0.003268f
C24530 a_n1177_43370# a_n1151_42308# 3.34e-19
C24531 a_1307_43914# a_n1925_42282# 0.03653f
C24532 a_6171_45002# a_10586_45546# 0.001629f
C24533 a_7705_45326# a_8049_45260# 0.032872f
C24534 a_8560_45348# a_2324_44458# 0.070986f
C24535 a_10949_43914# a_12549_44172# 0.052089f
C24536 a_10729_43914# a_768_44030# 0.004644f
C24537 a_10617_44484# a_3090_45724# 0.003583f
C24538 a_18248_44752# a_17339_46660# 0.019889f
C24539 a_n2661_44458# a_n2293_46098# 0.026753f
C24540 a_n2433_44484# a_n2472_46090# 5.65e-21
C24541 a_2124_47436# VDD 0.086403f
C24542 a_n3674_37592# a_n3420_39072# 0.019892f
C24543 a_15486_42560# a_15890_42674# 0.051162f
C24544 a_13575_42558# a_13921_42308# 0.013377f
C24545 a_n1630_35242# a_n3565_39304# 2.9e-19
C24546 COMP_P a_1736_39043# 6.78e-21
C24547 a_n3674_38680# a_n3565_38502# 0.128677f
C24548 a_1606_42308# a_1239_39587# 9.67e-20
C24549 a_15764_42576# a_15959_42545# 0.21686f
C24550 a_6123_31319# a_7174_31319# 13.9919f
C24551 a_19321_45002# a_12741_44636# 0.113088f
C24552 a_20916_46384# a_20202_43084# 0.181561f
C24553 a_491_47026# a_765_45546# 1.57e-19
C24554 a_21588_30879# a_22365_46825# 5.32e-19
C24555 a_10428_46928# a_11813_46116# 1.23e-19
C24556 a_10467_46802# a_11735_46660# 0.096658f
C24557 a_10554_47026# a_10768_47026# 0.097745f
C24558 a_10623_46897# a_11186_47026# 0.049827f
C24559 a_6755_46942# a_8601_46660# 5.59e-19
C24560 a_n881_46662# a_2698_46116# 0.058407f
C24561 a_12465_44636# a_9290_44172# 7.82e-20
C24562 a_13507_46334# a_10903_43370# 0.016027f
C24563 a_4883_46098# a_11133_46155# 0.007956f
C24564 a_16327_47482# a_17957_46116# 6.07e-20
C24565 a_11599_46634# a_20075_46420# 0.021805f
C24566 a_10227_46804# a_2324_44458# 0.051051f
C24567 a_n1435_47204# a_10809_44734# 9.93e-19
C24568 a_12861_44030# a_6945_45028# 0.108969f
C24569 a_n443_46116# a_n1925_42282# 0.001452f
C24570 a_n1151_42308# a_5431_46482# 0.004507f
C24571 a_3160_47472# a_5066_45546# 1.83e-20
C24572 a_2063_45854# a_5527_46155# 8.53e-21
C24573 a_19615_44636# a_n97_42460# 5.97e-21
C24574 a_895_43940# a_2455_43940# 0.01899f
C24575 a_10949_43914# a_12429_44172# 0.156922f
C24576 a_2998_44172# a_1241_43940# 1.39e-20
C24577 a_n2661_42834# a_6293_42852# 1.51e-19
C24578 a_n2661_43922# a_6031_43396# 1.84e-20
C24579 a_n356_44636# a_14358_43442# 3.91e-21
C24580 a_11823_42460# a_14456_42282# 0.004505f
C24581 a_10193_42453# a_15803_42450# 3.64e-19
C24582 a_2711_45572# a_13258_32519# 0.02914f
C24583 a_20193_45348# a_13887_32519# 0.277027f
C24584 a_7499_43078# a_9885_42308# 0.00284f
C24585 a_2479_44172# a_3052_44056# 9.94e-20
C24586 a_n2017_45002# a_13291_42460# 0.042872f
C24587 a_3537_45260# a_5193_42852# 0.012016f
C24588 a_n1059_45260# a_13003_42852# 0.004401f
C24589 a_5111_44636# a_8483_43230# 1.96e-19
C24590 a_2711_45572# a_8791_45572# 6.36e-19
C24591 a_10180_45724# a_8746_45002# 0.304016f
C24592 a_10053_45546# a_10490_45724# 0.084842f
C24593 a_7499_43078# a_11525_45546# 1.14e-21
C24594 a_11341_43940# a_11415_45002# 6.83e-19
C24595 a_21381_43940# a_19692_46634# 0.022586f
C24596 a_8685_43396# a_4646_46812# 7.39e-20
C24597 a_13213_44734# a_13259_45724# 0.020051f
C24598 a_n310_44811# a_n755_45592# 0.001544f
C24599 a_12895_43230# a_12861_44030# 3e-19
C24600 a_11813_46116# VDD 0.434656f
C24601 a_1606_42308# a_11206_38545# 3.98e-20
C24602 a_376_46348# a_1208_46090# 5.21e-19
C24603 a_n2293_46098# a_2804_46116# 1.46e-20
C24604 a_472_46348# a_805_46414# 0.360492f
C24605 a_288_46660# a_n443_42852# 2.55e-21
C24606 a_2107_46812# a_2277_45546# 4.99e-20
C24607 a_2959_46660# a_2957_45546# 1.67e-20
C24608 a_2443_46660# a_3503_45724# 3.68e-20
C24609 a_13885_46660# a_10809_44734# 0.026009f
C24610 a_14180_46812# a_6945_45028# 4.2e-20
C24611 a_16388_46812# a_18985_46122# 5.62e-21
C24612 w_11334_34010# a_19864_35138# 0.005843f
C24613 SMPL_ON_P a_n923_35174# 2.32e-19
C24614 a_9313_44734# a_15785_43172# 7.07e-19
C24615 a_15493_43940# a_16664_43396# 9.17e-19
C24616 a_5343_44458# a_1606_42308# 1.12e-20
C24617 a_1756_43548# a_1891_43646# 0.008678f
C24618 a_n2661_42282# a_n2840_42826# 0.001572f
C24619 a_3422_30871# a_18083_42858# 2.69e-20
C24620 a_3905_42865# a_4520_42826# 0.054799f
C24621 a_15493_43396# a_16823_43084# 0.029968f
C24622 a_14021_43940# a_16243_43396# 0.017079f
C24623 a_3080_42308# a_4905_42826# 0.005659f
C24624 a_10807_43548# a_4361_42308# 0.006525f
C24625 a_15682_43940# a_743_42282# 3.41e-20
C24626 a_n998_43396# VDD 6.7e-20
C24627 a_15903_45785# a_16019_45002# 0.139976f
C24628 a_15765_45572# a_15595_45028# 1.18e-19
C24629 a_15599_45572# a_1307_43914# 1.34e-19
C24630 a_8696_44636# a_13777_45326# 5.73e-20
C24631 a_11652_45724# a_n2661_43370# 0.028174f
C24632 a_11322_45546# a_13105_45348# 6.34e-21
C24633 a_2711_45572# a_20193_45348# 5.96e-20
C24634 a_16522_42674# a_10227_46804# 2.46e-19
C24635 a_n4064_39072# SMPL_ON_P 1.17e-20
C24636 a_14401_32519# a_20205_31679# 0.054064f
C24637 a_6452_43396# a_526_44458# 9.65e-19
C24638 a_8325_42308# a_n1613_43370# 2.95e-20
C24639 a_743_42282# a_1823_45246# 0.06422f
C24640 a_16823_43084# a_3483_46348# 8.97e-20
C24641 a_9313_44734# CLK 9.52e-20
C24642 a_5263_45724# a_n881_46662# 0.180025f
C24643 a_5907_45546# a_n1613_43370# 2.13e-20
C24644 a_10180_45724# a_4883_46098# 0.001751f
C24645 a_13527_45546# a_10227_46804# 6.04e-19
C24646 a_8696_44636# a_n1151_42308# 5.67e-21
C24647 a_13467_32519# a_4361_42308# 0.121732f
C24648 a_21487_43396# a_13678_32519# 7.05e-19
C24649 a_10341_43396# a_10835_43094# 1.26e-19
C24650 a_9145_43396# a_13635_43156# 0.001181f
C24651 VDAC_N C4_N_btm 13.8047f
C24652 a_8495_42852# VDD 0.132018f
C24653 en_comp a_n356_44636# 3.08e-20
C24654 a_7229_43940# a_5883_43914# 0.026061f
C24655 a_3232_43370# a_10057_43914# 0.025371f
C24656 a_7499_43078# a_7542_44172# 0.069089f
C24657 a_5267_42460# a_4185_45028# 9.17e-19
C24658 a_8037_42858# a_n443_42852# 0.007515f
C24659 a_13113_42826# a_n357_42282# 0.008588f
C24660 a_3080_42308# a_n923_35174# 0.006061f
C24661 a_18587_45118# a_16327_47482# 0.002342f
C24662 a_11827_44484# a_12861_44030# 0.466435f
C24663 C7_P_btm VDD 0.121904f
C24664 a_n2661_44458# a_4791_45118# 0.095212f
C24665 a_n1177_44458# a_n1151_42308# 0.021669f
C24666 a_2779_44458# a_2063_45854# 1.24e-20
C24667 a_12607_44458# a_n1741_47186# 1.63e-22
C24668 a_4223_44672# a_584_46384# 0.044788f
C24669 a_6171_45002# a_n743_46660# 0.140224f
C24670 a_3357_43084# a_5732_46660# 0.017659f
C24671 a_3429_45260# a_2107_46812# 3.88e-21
C24672 a_5205_44484# a_n1925_46634# 3.1e-21
C24673 a_8953_45002# a_n2661_46634# 2.39e-20
C24674 a_n143_45144# a_n2661_46098# 2.28e-22
C24675 a_3232_43370# a_n2438_43548# 8.07e-21
C24676 a_16333_45814# a_15368_46634# 3.38e-20
C24677 a_14537_43396# a_13661_43548# 0.505634f
C24678 a_16855_45546# a_3090_45724# 0.007982f
C24679 a_1423_45028# a_768_44030# 0.096238f
C24680 a_13163_45724# a_765_45546# 4.54e-21
C24681 a_14180_45002# a_13747_46662# 5.33e-19
C24682 a_5907_45546# a_n2293_46098# 4.2e-19
C24683 a_17333_42852# a_17141_43172# 1.97e-19
C24684 a_15567_42826# a_15953_42852# 0.006406f
C24685 a_4743_43172# a_4649_42852# 1.26e-19
C24686 a_13678_32519# a_5932_42308# 1.17e-19
C24687 a_5649_42852# a_6171_42473# 0.00196f
C24688 a_743_42282# a_5934_30871# 0.020602f
C24689 a_5342_30871# a_16245_42852# 8.35e-20
C24690 a_18083_42858# a_18504_43218# 0.088127f
C24691 a_16137_43396# a_15803_42450# 0.002599f
C24692 a_2905_42968# a_n784_42308# 4.32e-21
C24693 a_16243_43396# a_15764_42576# 2.19e-20
C24694 a_n3565_38502# VDD 0.762011f
C24695 a_9863_47436# a_9804_47204# 0.109361f
C24696 a_n1435_47204# a_n881_46662# 0.068194f
C24697 a_n1741_47186# a_171_46873# 3.56e-20
C24698 a_n815_47178# a_n743_46660# 0.001755f
C24699 a_1209_47178# a_n2661_46634# 0.001337f
C24700 a_n971_45724# a_n1925_46634# 0.163523f
C24701 a_20990_47178# a_12465_44636# 3.04e-19
C24702 a_13507_46334# a_4883_46098# 4.09671f
C24703 a_18597_46090# a_11453_44696# 0.022871f
C24704 a_15415_45028# a_15493_43396# 2.36e-21
C24705 a_22959_45036# a_22959_44484# 0.025171f
C24706 a_10193_42453# a_16137_43396# 0.329316f
C24707 a_12607_44458# a_13296_44484# 0.002675f
C24708 a_20193_45348# a_22485_44484# 0.027057f
C24709 a_n2012_44484# a_n2293_43922# 9.53e-19
C24710 a_22223_45036# a_19237_31679# 7.18e-19
C24711 a_19479_31679# a_14401_32519# 0.053843f
C24712 a_1307_43914# a_2698_46116# 2.53e-20
C24713 a_375_42282# a_167_45260# 0.017297f
C24714 a_15415_45028# a_3483_46348# 5.74e-21
C24715 a_626_44172# a_1823_45246# 2.16e-20
C24716 a_1145_45348# a_1138_42852# 1.86e-19
C24717 a_16922_45042# a_17339_46660# 0.02918f
C24718 a_20362_44736# a_19321_45002# 0.009631f
C24719 a_5883_43914# a_8270_45546# 0.20967f
C24720 a_14539_43914# a_6755_46942# 0.094724f
C24721 a_20679_44626# a_13747_46662# 0.030878f
C24722 a_3422_30871# a_12549_44172# 0.148646f
C24723 a_14673_44172# a_n743_46660# 3.65e-21
C24724 a_15861_45028# a_16375_45002# 0.029833f
C24725 a_6171_45002# a_11189_46129# 7.06e-21
C24726 a_8953_45002# a_8199_44636# 0.12099f
C24727 a_8191_45002# a_5937_45572# 0.180306f
C24728 a_2274_45254# a_2324_44458# 0.007089f
C24729 a_413_45260# a_17715_44484# 4.56e-21
C24730 a_9028_43914# a_9313_45822# 3.91e-20
C24731 a_1241_43940# a_n2497_47436# 5.31e-20
C24732 a_4921_42308# a_4169_42308# 9.83e-20
C24733 a_2351_42308# a_5742_30871# 1.16e-20
C24734 a_5755_42308# a_5934_30871# 2.52e-20
C24735 a_5932_42308# a_6123_31319# 1.49414f
C24736 a_1606_42308# a_12563_42308# 3.31e-20
C24737 a_6773_42558# a_6761_42308# 0.01129f
C24738 a_n1532_35090# a_n923_35174# 0.400297f
C24739 a_n1386_35608# EN_VIN_BSTR_P 0.573134f
C24740 a_3626_43646# CAL_N 0.00204f
C24741 a_13661_43548# a_3090_45724# 0.177565f
C24742 a_5807_45002# a_14976_45028# 0.026261f
C24743 a_13747_46662# a_15009_46634# 6.01e-21
C24744 a_2107_46812# a_6755_46942# 0.002513f
C24745 a_3877_44458# a_5732_46660# 0.040487f
C24746 a_4646_46812# a_5907_46634# 0.037052f
C24747 a_4651_46660# a_5167_46660# 0.102946f
C24748 a_n2661_46634# a_10768_47026# 0.002208f
C24749 a_n1925_46634# a_8023_46660# 2.21e-19
C24750 a_n881_46662# a_13885_46660# 2.09e-19
C24751 a_2063_45854# a_6165_46155# 8.02e-20
C24752 a_n1741_47186# a_10903_43370# 0.066687f
C24753 a_n1151_42308# a_4704_46090# 0.001193f
C24754 a_n237_47217# a_9569_46155# 6.37e-20
C24755 a_3785_47178# a_4185_45028# 2.07e-20
C24756 a_4007_47204# a_3483_46348# 1.93e-19
C24757 a_n443_46116# a_2698_46116# 0.012019f
C24758 a_n1435_47204# a_n2157_46122# 1.63e-20
C24759 a_6151_47436# a_1823_45246# 3.85e-20
C24760 a_20894_47436# a_20731_47026# 2.28e-19
C24761 a_13507_46334# a_21188_46660# 0.03408f
C24762 a_21496_47436# a_21363_46634# 4.81e-20
C24763 a_4883_46098# a_20623_46660# 3.47e-20
C24764 a_16327_47482# a_11415_45002# 0.94171f
C24765 a_12465_44636# a_20273_46660# 3.92e-21
C24766 a_11453_44696# a_19123_46287# 0.021733f
C24767 a_n2017_45002# a_13460_43230# 2.95e-21
C24768 a_n913_45002# a_12895_43230# 0.029875f
C24769 a_n1059_45260# a_13635_43156# 0.006041f
C24770 a_3537_45260# a_7227_42852# 0.002978f
C24771 a_n2661_42834# a_7499_43940# 5.15e-19
C24772 a_10193_42453# a_n784_42308# 1.64e-19
C24773 a_n2661_44458# a_8791_43396# 2.51e-20
C24774 a_19279_43940# a_15493_43396# 0.003821f
C24775 a_5013_44260# a_5663_43940# 0.083171f
C24776 a_20362_44736# a_20623_43914# 0.001795f
C24777 a_18579_44172# a_18326_43940# 0.096332f
C24778 a_20835_44721# a_19862_44208# 0.00122f
C24779 a_11967_42832# a_11341_43940# 0.046075f
C24780 a_18287_44626# VDD 0.389383f
C24781 a_n4064_39616# C5_P_btm 8.54e-20
C24782 a_n3420_39616# C3_P_btm 2.76e-20
C24783 a_n4064_39072# a_n1532_35090# 9.45e-20
C24784 a_n3420_39072# EN_VIN_BSTR_P 0.772414f
C24785 a_15743_43084# a_10227_46804# 0.002448f
C24786 a_n1991_42858# a_n1151_42308# 2.39e-19
C24787 a_685_42968# a_n971_45724# 4.15e-21
C24788 a_17973_43940# a_15227_44166# 4.09e-19
C24789 a_19862_44208# a_3090_45724# 0.004983f
C24790 a_2896_43646# a_n2293_46634# 7.64e-19
C24791 a_14539_43914# a_8049_45260# 1.59e-36
C24792 a_14815_43914# a_2324_44458# 1.05e-20
C24793 a_9145_43396# a_n1613_43370# 7e-20
C24794 a_1110_47026# VDD 4.6e-19
C24795 a_n3420_39072# a_n2302_39072# 2.77e-19
C24796 a_1736_39587# a_2112_39137# 0.269796f
C24797 a_n3565_39304# a_n3607_39392# 0.001003f
C24798 a_n3420_39616# a_n4064_38528# 0.048102f
C24799 a_n4064_39616# a_n3420_38528# 0.052176f
C24800 a_n4064_40160# a_n4209_38216# 0.047163f
C24801 a_n4315_30879# a_n3565_38216# 0.043307f
C24802 a_1343_38525# comp_n 0.004961f
C24803 a_n2946_39072# a_n4064_39072# 0.053263f
C24804 a_5742_30871# C4_N_btm 0.03103f
C24805 a_n4318_38216# a_n3607_38304# 7.49e-20
C24806 a_13059_46348# a_12741_44636# 0.02008f
C24807 a_3090_45724# a_4185_45028# 0.770164f
C24808 a_15368_46634# a_3483_46348# 1.42e-21
C24809 a_18285_46348# a_18280_46660# 0.089884f
C24810 a_20273_46660# a_20528_46660# 0.056391f
C24811 a_20623_46660# a_21188_46660# 7.99e-20
C24812 a_2107_46812# a_8049_45260# 0.029889f
C24813 a_5807_45002# a_18051_46116# 0.006001f
C24814 a_19321_45002# a_16375_45002# 8.59e-21
C24815 a_n743_46660# a_9751_46155# 3.19e-19
C24816 a_13747_46662# a_19431_46494# 1.74e-19
C24817 a_n881_46662# a_380_45546# 0.001604f
C24818 a_6755_46942# a_14493_46090# 1.15e-20
C24819 a_8846_46660# a_5937_45572# 2.62e-19
C24820 a_8270_45546# a_9569_46155# 1.61e-19
C24821 a_n1613_43370# a_n1099_45572# 0.025553f
C24822 a_6298_44484# a_7309_42852# 1.49e-22
C24823 a_10405_44172# a_8685_43396# 4.99e-20
C24824 a_1241_43940# a_1568_43370# 1.38e-20
C24825 a_3422_30871# a_21855_43396# 0.005365f
C24826 a_n2661_42834# a_10991_42826# 1.88e-20
C24827 a_20512_43084# a_743_42282# 0.082751f
C24828 a_n2293_43922# a_10835_43094# 1.05e-20
C24829 a_9313_44734# a_5534_30871# 0.039673f
C24830 a_18184_42460# a_14097_32519# 9.17e-19
C24831 a_5829_43940# a_n97_42460# 7.1e-20
C24832 en_comp a_18727_42674# 3.94e-20
C24833 a_19963_31679# a_22775_42308# 4.22e-21
C24834 a_n1059_45260# a_18310_42308# 0.006864f
C24835 a_3992_43940# VDD 0.004127f
C24836 a_10180_45724# a_3232_43370# 1.58e-19
C24837 a_10053_45546# a_6171_45002# 5.53e-21
C24838 a_16147_45260# a_18691_45572# 9.71e-20
C24839 a_18479_45785# a_18341_45572# 0.21997f
C24840 a_18175_45572# a_18909_45814# 0.053479f
C24841 a_2813_43396# a_1823_45246# 5.33e-20
C24842 a_15743_43084# a_17339_46660# 0.450316f
C24843 a_5649_42852# a_19692_46634# 0.01341f
C24844 a_11341_43940# a_13259_45724# 0.045479f
C24845 a_n2661_42282# a_n357_42282# 0.055806f
C24846 a_3626_43646# a_8199_44636# 0.001453f
C24847 a_3726_37500# RST_Z 1.60318f
C24848 a_n2104_42282# a_n2312_40392# 4.5e-20
C24849 a_n4318_38216# a_n2312_39304# 0.023429f
C24850 VDAC_P C8_P_btm 0.220914p
C24851 a_n4209_37414# VIN_P 0.029528f
C24852 a_19721_31679# EN_OFFSET_CAL 3.03e-20
C24853 a_15682_46116# VDD 1.25004f
C24854 a_7227_45028# a_n1151_42308# 0.00514f
C24855 a_5907_45546# a_4791_45118# 0.02288f
C24856 a_7499_43078# a_n971_45724# 0.857375f
C24857 a_2211_45572# a_2063_45854# 0.006085f
C24858 a_n4209_38216# a_n4064_37440# 0.028219f
C24859 a_n3565_38216# a_n3420_37440# 0.038559f
C24860 a_n2293_46098# a_n1099_45572# 0.069723f
C24861 a_n1423_46090# a_n1079_45724# 1.85e-19
C24862 a_n1853_46287# a_n452_45724# 0.080546f
C24863 a_376_46348# a_n2661_45546# 4.24e-21
C24864 a_n1641_46494# a_n2293_45546# 1.27e-19
C24865 a_2324_44458# a_8034_45724# 1.84e-19
C24866 a_10903_43370# a_10586_45546# 0.238199f
C24867 a_14493_46090# a_8049_45260# 0.001687f
C24868 a_10341_43396# a_15037_43396# 1.71e-21
C24869 a_14955_43396# a_15231_43396# 0.00119f
C24870 a_n4318_39768# a_n4318_37592# 0.023201f
C24871 a_9313_44734# a_19647_42308# 9.5e-20
C24872 a_895_43940# a_961_42354# 7.76e-22
C24873 a_n97_42460# a_10835_43094# 7.73e-20
C24874 a_3080_42308# a_2905_42968# 3.9e-20
C24875 a_4093_43548# a_4520_42826# 0.077799f
C24876 a_n1557_42282# a_791_42968# 0.002272f
C24877 a_4235_43370# a_3935_42891# 0.082011f
C24878 a_1414_42308# a_1755_42282# 7.59e-19
C24879 a_453_43940# a_1606_42308# 2.97e-21
C24880 a_19452_47524# START 0.003297f
C24881 a_19321_45002# RST_Z 1.28e-19
C24882 a_9127_43156# VDD 0.468721f
C24883 a_22223_45572# a_18114_32519# 4.88e-19
C24884 a_7276_45260# a_n2661_43370# 0.007354f
C24885 a_n913_45002# a_11827_44484# 1.54e-19
C24886 a_2437_43646# a_19721_31679# 3.14e-19
C24887 a_6171_45002# a_13490_45394# 1.03e-19
C24888 a_16823_43084# a_n357_42282# 0.016884f
C24889 a_20753_42852# a_20202_43084# 8.28e-19
C24890 a_8162_45546# a_8270_45546# 0.170838f
C24891 a_20107_45572# a_20916_46384# 6.04e-21
C24892 a_20528_45572# a_13747_46662# 2.86e-19
C24893 a_2437_43646# a_13675_47204# 6.63e-20
C24894 a_n1059_45260# a_n1613_43370# 0.202724f
C24895 a_4927_45028# a_4883_46098# 2.86e-20
C24896 a_10775_45002# a_10227_46804# 0.006025f
C24897 a_15595_45028# a_12861_44030# 0.012748f
C24898 a_n2293_42834# a_584_46384# 0.049322f
C24899 a_n2661_43370# a_n746_45260# 0.060205f
C24900 a_3626_43646# a_13070_42354# 0.001839f
C24901 a_2982_43646# a_14456_42282# 2.19e-19
C24902 a_14401_32519# a_13258_32519# 0.053694f
C24903 a_5111_42852# a_5193_43172# 0.003935f
C24904 a_16795_42852# a_17701_42308# 2.09e-19
C24905 a_17124_42282# VDD 0.28176f
C24906 a_n2293_43922# a_7754_40130# 6.5e-19
C24907 a_7227_47204# a_7903_47542# 0.002513f
C24908 a_4915_47217# a_13381_47204# 0.045103f
C24909 a_6851_47204# a_6575_47204# 0.027563f
C24910 a_6151_47436# a_11031_47542# 0.03901f
C24911 a_n1741_47186# a_4883_46098# 0.031761f
C24912 a_n443_46116# a_n1435_47204# 8.31e-19
C24913 a_5111_44636# a_6453_43914# 2.3e-20
C24914 a_3232_43370# a_5013_44260# 0.081759f
C24915 a_5691_45260# a_5495_43940# 3.68e-21
C24916 a_20623_45572# a_20935_43940# 1.84e-19
C24917 a_11691_44458# a_9313_44734# 5.15e-20
C24918 a_n2129_44697# a_n310_44811# 8.5e-19
C24919 a_n1917_44484# a_n1655_44484# 0.001705f
C24920 a_n1352_44484# a_n1190_44850# 0.006453f
C24921 a_10057_43914# a_8975_43940# 0.069663f
C24922 a_n1699_44726# a_n356_44636# 1.11e-20
C24923 a_5379_42460# a_n755_45592# 0.038776f
C24924 a_1149_42558# a_n443_42852# 1.56e-19
C24925 a_13904_45546# VDD 0.135068f
C24926 a_13678_32519# VREF 1.33e-19
C24927 a_484_44484# a_n1613_43370# 1.49e-20
C24928 a_12553_44484# a_12465_44636# 3.52e-19
C24929 a_11967_42832# a_16327_47482# 0.241578f
C24930 a_3600_43914# a_n971_45724# 1.64e-20
C24931 a_1115_44172# a_584_46384# 0.174981f
C24932 a_13556_45296# a_13059_46348# 0.274813f
C24933 a_2437_43646# a_167_45260# 0.025008f
C24934 a_n2661_45010# a_n1641_46494# 2.26e-19
C24935 a_n2293_45010# a_n1991_46122# 4.53e-20
C24936 a_n1059_45260# a_n2293_46098# 2.7e-19
C24937 a_949_44458# a_1799_45572# 4.76e-19
C24938 a_12607_44458# a_n743_46660# 2.46e-22
C24939 a_6109_44484# a_768_44030# 0.04198f
C24940 a_n2017_45002# a_n2157_46122# 2.07e-20
C24941 en_comp a_21076_30879# 3.62e-19
C24942 a_12427_45724# a_8049_45260# 0.012343f
C24943 a_8746_45002# a_10586_45546# 0.001538f
C24944 a_n4318_38680# a_n3565_38502# 5.19e-20
C24945 a_n473_42460# a_n3674_37592# 0.054584f
C24946 a_n1329_42308# a_n1630_35242# 0.043579f
C24947 a_19339_43156# a_19511_42282# 4.61e-19
C24948 a_18083_42858# a_7174_31319# 1.26e-20
C24949 a_n1925_46634# a_601_46902# 0.004874f
C24950 a_n743_46660# a_171_46873# 0.075858f
C24951 a_n2438_43548# a_n133_46660# 0.848709f
C24952 a_768_44030# a_4646_46812# 0.047094f
C24953 a_n2661_46634# a_288_46660# 0.002871f
C24954 a_n1021_46688# a_33_46660# 1.18e-19
C24955 a_n1613_43370# a_3878_46660# 0.002879f
C24956 a_11453_44696# a_6755_46942# 0.026496f
C24957 a_11599_46634# a_15009_46634# 6.85e-19
C24958 a_14955_47212# a_3090_45724# 0.009113f
C24959 a_10227_46804# a_11186_47026# 0.018916f
C24960 a_12861_44030# a_15559_46634# 0.066578f
C24961 a_13717_47436# a_16292_46812# 1.08e-20
C24962 a_1209_47178# a_765_45546# 0.003605f
C24963 a_9482_43914# a_14955_43396# 5.1e-21
C24964 a_18443_44721# a_15493_43940# 1.61e-20
C24965 a_18989_43940# a_11341_43940# 0.004444f
C24966 a_14537_43396# a_14579_43548# 0.046172f
C24967 a_5837_45028# a_6031_43396# 5.01e-21
C24968 a_13556_45296# a_15095_43370# 6.47e-22
C24969 a_20193_45348# a_14401_32519# 0.175398f
C24970 a_4223_44672# a_5025_43940# 0.002864f
C24971 a_5891_43370# a_10807_43548# 1.3e-19
C24972 a_n2661_43922# a_1525_44260# 1.65e-19
C24973 a_n2661_42834# a_2253_44260# 3.6e-19
C24974 a_n2293_42834# a_n144_43396# 3.51e-19
C24975 a_20447_31679# a_13467_32519# 0.051601f
C24976 a_n2860_37984# VDD 0.004232f
C24977 a_17023_45118# VDD 0.086861f
C24978 a_5934_30871# VIN_P 0.009408f
C24979 a_5742_30871# C6_P_btm 0.170624f
C24980 a_n4209_37414# a_n2956_38680# 1.36e-21
C24981 a_n356_44636# a_4185_45028# 1.54308f
C24982 a_11649_44734# a_12741_44636# 3.54e-20
C24983 a_5841_44260# a_5257_43370# 3.99e-19
C24984 a_19808_44306# a_12549_44172# 6.88e-19
C24985 a_375_42282# a_n863_45724# 0.451905f
C24986 a_626_44172# a_n2293_45546# 0.150062f
C24987 a_19721_31679# a_22959_46124# 5.11e-20
C24988 a_2232_45348# a_n2661_45546# 7.5e-19
C24989 a_8191_45002# a_n443_42852# 3.74e-21
C24990 a_4743_44484# a_2324_44458# 0.042685f
C24991 a_n2661_44458# a_6945_45028# 1.65e-19
C24992 a_n2840_43370# a_n1613_43370# 2.32e-21
C24993 a_2711_45572# CLK 0.032985f
C24994 a_n89_47570# VDD 4.63e-19
C24995 a_21335_42336# a_21613_42308# 0.110671f
C24996 a_13258_32519# a_21421_42336# 7.85e-19
C24997 a_5342_30871# a_8530_39574# 1.55e-19
C24998 a_3067_47026# a_3147_46376# 2.75e-19
C24999 a_3524_46660# a_3699_46348# 4.06e-19
C25000 a_13607_46688# a_13059_46348# 9.43e-19
C25001 a_15559_46634# a_14180_46812# 0.001017f
C25002 a_n881_46662# a_526_44458# 0.060324f
C25003 a_13747_46662# a_19335_46494# 0.005102f
C25004 a_19321_45002# a_18985_46122# 0.019556f
C25005 a_n743_46660# a_10903_43370# 0.080542f
C25006 a_2107_46812# a_8953_45546# 0.007676f
C25007 a_19594_46812# a_18819_46122# 1.63e-19
C25008 a_16697_47582# a_6945_45028# 1.16e-19
C25009 a_5807_45002# a_19900_46494# 0.00115f
C25010 a_n1613_43370# a_n1925_42282# 1.08e-19
C25011 a_2905_45572# a_3316_45546# 0.004332f
C25012 a_n443_46116# a_380_45546# 0.073277f
C25013 a_327_47204# a_n443_42852# 3.15e-21
C25014 a_n237_47217# a_1990_45899# 8.97e-19
C25015 a_16327_47482# a_13259_45724# 0.584328f
C25016 a_10227_46804# a_12839_46116# 8.43e-21
C25017 a_4883_46098# a_10586_45546# 0.006953f
C25018 a_11453_44696# a_8049_45260# 0.032046f
C25019 a_n2017_45002# a_4933_42558# 0.00112f
C25020 a_n913_45002# a_3581_42558# 0.003935f
C25021 a_2479_44172# a_3540_43646# 5.31e-20
C25022 a_18184_42460# a_22959_42860# 0.004934f
C25023 a_5883_43914# a_5755_42852# 6.14e-21
C25024 a_9313_44734# a_4190_30871# 0.02726f
C25025 a_5013_44260# a_4905_42826# 3.52e-20
C25026 a_n2661_42282# a_n2433_43396# 1.4e-20
C25027 a_11967_42832# a_10341_43396# 0.076124f
C25028 a_n630_44306# VDD 1.8e-19
C25029 a_10193_42453# a_18479_45785# 1.12e-19
C25030 a_13163_45724# a_13385_45572# 0.001684f
C25031 a_11341_43940# a_18189_46348# 2.49e-20
C25032 a_n784_42308# SMPL_ON_P 0.001291f
C25033 a_14579_43548# a_3090_45724# 0.074713f
C25034 a_12379_42858# a_13661_43548# 1.34e-19
C25035 a_19279_43940# a_n357_42282# 3.11e-20
C25036 a_9801_43940# a_3483_46348# 0.027985f
C25037 a_n2293_46098# a_n1925_42282# 0.020467f
C25038 a_16388_46812# a_18243_46436# 0.004535f
C25039 a_11189_46129# a_10903_43370# 0.151119f
C25040 a_8016_46348# a_2324_44458# 0.048711f
C25041 a_9290_44172# a_12005_46116# 1.48e-19
C25042 a_n4209_39304# a_n3420_37984# 0.029539f
C25043 a_14539_43914# a_14456_42282# 5.4e-20
C25044 a_8791_43396# a_9145_43396# 0.092458f
C25045 a_20974_43370# a_4190_30871# 0.214288f
C25046 a_14955_43940# a_5342_30871# 1.82e-19
C25047 a_21381_43940# a_743_42282# 4.2e-21
C25048 a_n356_44636# a_9803_42558# 1.46e-19
C25049 a_9313_45822# CLK 0.027301f
C25050 a_n1435_47204# DATA[4] 0.033859f
C25051 a_15811_47375# RST_Z 1.42e-19
C25052 SMPL_ON_N a_22609_37990# 2.01e-20
C25053 a_19268_43646# VDD 0.237793f
C25054 a_4927_45028# a_3232_43370# 1.34e-20
C25055 a_3537_45260# a_7229_43940# 1.13e-19
C25056 a_5111_44636# a_6171_45002# 3.76e-19
C25057 a_n2293_45010# a_375_42282# 0.021456f
C25058 a_n2017_45002# a_1307_43914# 0.001015f
C25059 a_n2661_45010# a_626_44172# 0.0195f
C25060 a_10180_45724# a_8975_43940# 6.79e-20
C25061 a_8746_45002# a_10440_44484# 0.027688f
C25062 a_15903_45785# a_11827_44484# 3.96e-21
C25063 a_10193_42453# a_10057_43914# 4.92e-20
C25064 a_15037_45618# a_11691_44458# 1.37e-19
C25065 a_12379_42858# a_4185_45028# 6.62e-20
C25066 a_18727_42674# a_13661_43548# 1.61e-19
C25067 a_5267_42460# a_5257_43370# 9.2e-19
C25068 a_6123_31319# a_4646_46812# 0.004637f
C25069 a_10341_43396# a_13259_45724# 0.08137f
C25070 a_7287_43370# a_n755_45592# 1.51e-19
C25071 a_5565_43396# a_n2661_45546# 7.68e-21
C25072 a_7871_42858# a_8953_45546# 0.017048f
C25073 a_8037_42858# a_8199_44636# 2.18e-20
C25074 w_1575_34946# C0_dummy_P_btm 3.87e-21
C25075 a_20273_45572# a_16327_47482# 0.050306f
C25076 a_18175_45572# a_4883_46098# 6.22e-20
C25077 a_18341_45572# a_13507_46334# 7.32e-21
C25078 a_18799_45938# a_18597_46090# 1.88e-19
C25079 a_20528_45572# a_11599_46634# 1.32e-20
C25080 a_3357_43084# a_9863_47436# 1.35e-19
C25081 a_2437_43646# a_11459_47204# 0.004348f
C25082 a_413_45260# a_584_46384# 0.164383f
C25083 a_3537_45260# a_n237_47217# 3.39e-20
C25084 a_4558_45348# a_n971_45724# 1.27e-19
C25085 a_n2017_45002# a_n443_46116# 1.32e-19
C25086 a_n967_45348# a_n1151_42308# 0.170453f
C25087 a_n1059_45260# a_4791_45118# 0.020789f
C25088 a_8746_45002# a_n743_46660# 1.81e-19
C25089 a_1990_45572# a_1799_45572# 2.88e-19
C25090 a_15297_45822# a_n881_46662# 0.001288f
C25091 a_n2840_45546# a_n2810_45572# 0.162234f
C25092 a_15493_43940# a_15521_42308# 2.45e-20
C25093 a_1847_42826# a_3681_42891# 8.84e-21
C25094 a_n97_42460# a_n39_42308# 0.001449f
C25095 a_2075_43172# a_2905_42968# 0.023236f
C25096 a_13887_32519# a_5534_30871# 0.047233f
C25097 a_3080_42308# a_n784_42308# 0.170007f
C25098 a_n2661_42282# a_n4064_40160# 4.6e-21
C25099 a_14021_43940# a_15803_42450# 1.55e-20
C25100 a_n1557_42282# a_n961_42308# 0.041329f
C25101 a_743_42282# a_18249_42858# 4.69e-20
C25102 a_4361_42308# a_16795_42852# 2.38e-20
C25103 a_5649_42852# a_5342_30871# 0.091782f
C25104 a_4190_30871# a_18599_43230# 0.008694f
C25105 a_1209_43370# a_1184_42692# 0.001053f
C25106 a_458_43396# a_961_42354# 4.08e-20
C25107 a_15493_43396# a_19332_42282# 3.15e-19
C25108 a_20820_30879# a_22521_40055# 1.31e-20
C25109 a_13059_46348# RST_Z 0.002761f
C25110 VDAC_Ni a_3754_38470# 0.911632f
C25111 a_7754_40130# a_5088_37509# 0.036831f
C25112 a_7754_39964# a_3726_37500# 0.030605f
C25113 a_1755_42282# VDD 0.215277f
C25114 a_n1920_47178# a_n815_47178# 6.26e-20
C25115 a_n2497_47436# a_n746_45260# 0.046973f
C25116 a_n2109_47186# a_n452_47436# 0.039314f
C25117 a_n1741_47186# a_n1605_47204# 0.011722f
C25118 a_9482_43914# a_n2661_42834# 0.076592f
C25119 a_10193_42453# a_14021_43940# 0.033291f
C25120 a_20193_45348# a_20205_45028# 0.012189f
C25121 a_11827_44484# a_n2661_44458# 0.003582f
C25122 a_n2017_45002# a_18579_44172# 3.84e-19
C25123 a_11136_42852# a_n357_42282# 0.002171f
C25124 a_3905_42558# a_n1925_42282# 8.24e-19
C25125 a_5934_30871# a_n2956_38680# 4.1e-21
C25126 a_18727_42674# a_4185_45028# 1.37e-19
C25127 a_8696_44636# a_12741_44636# 2.20704f
C25128 a_16020_45572# a_11415_45002# 9.68e-19
C25129 a_10951_45334# a_10428_46928# 1.28e-19
C25130 a_10775_45002# a_10467_46802# 1.67e-22
C25131 a_19778_44110# a_19321_45002# 0.568668f
C25132 a_18494_42460# a_13747_46662# 0.004606f
C25133 a_3602_45348# a_3877_44458# 1.19e-19
C25134 a_17568_45572# a_765_45546# 2.41e-21
C25135 a_3537_45260# a_8270_45546# 0.002418f
C25136 a_413_45260# a_11901_46660# 4.96e-20
C25137 a_10193_42453# a_11133_46155# 0.039441f
C25138 a_10490_45724# a_9290_44172# 0.022805f
C25139 a_8746_45002# a_11189_46129# 6.97e-20
C25140 a_10053_45546# a_10903_43370# 4.05e-19
C25141 a_n4318_40392# a_n1613_43370# 4.23e-20
C25142 a_10440_44484# a_4883_46098# 3.27e-21
C25143 a_18989_43940# a_16327_47482# 0.100946f
C25144 a_743_42282# a_21125_42558# 3.76e-20
C25145 a_n2293_42282# a_2713_42308# 0.002882f
C25146 a_10518_42984# a_10723_42308# 6.75e-19
C25147 a_4361_42308# a_21335_42336# 0.013772f
C25148 a_13467_32519# a_21887_42336# 0.011781f
C25149 a_5649_42852# a_20107_42308# 1.31e-19
C25150 a_16328_43172# a_16245_42852# 1.48e-19
C25151 a_n755_45592# DATA[0] 1.08e-20
C25152 a_n881_46662# a_13759_47204# 2.74e-19
C25153 a_n1151_42308# a_7715_46873# 0.09029f
C25154 a_n237_47217# a_6969_46634# 1.13e-19
C25155 a_2063_45854# a_8492_46660# 0.005635f
C25156 a_n971_45724# a_6999_46987# 0.005614f
C25157 a_6151_47436# a_5732_46660# 0.002133f
C25158 a_4883_46098# a_n743_46660# 5.6639f
C25159 a_n2312_39304# a_n2956_39768# 5.91067f
C25160 a_n2312_40392# a_n2661_46634# 1.45e-20
C25161 C2_N_btm VDD 0.268945f
C25162 a_n2017_45002# a_9396_43370# 3.4e-20
C25163 a_n1059_45260# a_8791_43396# 0.196029f
C25164 a_n913_45002# a_8147_43396# 7.89e-20
C25165 a_3232_43370# a_4699_43561# 9.73e-20
C25166 a_2382_45260# a_3626_43646# 0.041715f
C25167 a_3065_45002# a_2982_43646# 0.026494f
C25168 a_19778_44110# a_20623_43914# 3.52e-20
C25169 a_n2293_43922# a_11967_42832# 0.022597f
C25170 a_18184_42460# a_20365_43914# 2.05e-19
C25171 a_5883_43914# a_7845_44172# 0.02286f
C25172 a_11827_44484# a_18451_43940# 0.006619f
C25173 a_11691_44458# a_17737_43940# 1.76e-19
C25174 a_18494_42460# a_20269_44172# 0.017863f
C25175 a_17613_45144# a_15493_43940# 4.03e-21
C25176 a_10951_45334# VDD 0.226705f
C25177 COMP_P EN_VIN_BSTR_N 0.004364f
C25178 a_14097_32519# RST_Z 0.051182f
C25179 a_8488_45348# a_2324_44458# 0.003185f
C25180 a_11173_44260# a_11453_44696# 3.43e-20
C25181 a_17970_44736# a_17339_46660# 0.002841f
C25182 a_10405_44172# a_768_44030# 0.001056f
C25183 a_9313_44734# a_15227_44166# 0.06548f
C25184 a_n3674_39768# a_n2442_46660# 0.023663f
C25185 a_10729_43914# a_12549_44172# 4.26e-20
C25186 a_1307_43914# a_526_44458# 0.467539f
C25187 a_3232_43370# a_10586_45546# 8.27e-19
C25188 a_2437_43646# a_n863_45724# 0.071802f
C25189 a_6709_45028# a_8049_45260# 4.7e-19
C25190 a_1431_47204# VDD 0.423871f
C25191 a_15486_42560# a_15959_42545# 7.99e-20
C25192 a_13575_42558# a_13657_42308# 0.003935f
C25193 a_5934_30871# a_13258_32519# 7.32e-19
C25194 a_n3674_38680# a_n4334_38528# 0.05024f
C25195 COMP_P a_1239_39043# 0.001354f
C25196 a_7227_42308# a_7174_31319# 9.76e-21
C25197 a_15764_42576# a_15803_42450# 0.901878f
C25198 a_10428_46928# a_11735_46660# 0.001328f
C25199 a_10467_46802# a_11186_47026# 0.082642f
C25200 a_5257_43370# a_3090_45724# 0.020885f
C25201 a_10623_46897# a_10768_47026# 0.057222f
C25202 a_288_46660# a_765_45546# 1.47e-21
C25203 a_n881_46662# a_2521_46116# 0.050613f
C25204 a_n1613_43370# a_2698_46116# 2.5e-20
C25205 a_4883_46098# a_11189_46129# 0.008441f
C25206 a_11599_46634# a_19335_46494# 0.030852f
C25207 a_10227_46804# a_14840_46494# 0.275527f
C25208 a_16588_47582# a_15682_46116# 0.00115f
C25209 a_16327_47482# a_18189_46348# 0.029513f
C25210 a_13381_47204# a_10809_44734# 1.08e-19
C25211 a_13717_47436# a_6945_45028# 0.038878f
C25212 a_n443_46116# a_526_44458# 0.366438f
C25213 a_4791_45118# a_n1925_42282# 1.87e-19
C25214 a_n237_47217# a_9241_46436# 2.14e-19
C25215 a_n1151_42308# a_5210_46482# 7.81e-19
C25216 a_2063_45854# a_5210_46155# 1.39e-19
C25217 a_18989_43940# a_10341_43396# 2.68e-19
C25218 a_11967_42832# a_n97_42460# 0.489711f
C25219 a_2479_44172# a_2455_43940# 0.025354f
C25220 a_895_43940# a_2253_43940# 0.053882f
C25221 a_10949_43914# a_11750_44172# 0.05299f
C25222 a_1414_42308# a_3737_43940# 1.01e-19
C25223 a_n2661_42834# a_6031_43396# 1.34e-19
C25224 a_11823_42460# a_13575_42558# 0.075921f
C25225 a_n356_44636# a_14579_43548# 5.95e-21
C25226 a_20193_45348# a_22223_43396# 0.020364f
C25227 a_10193_42453# a_15764_42576# 2.52e-19
C25228 a_2711_45572# a_19647_42308# 0.046367f
C25229 a_10729_43914# a_12429_44172# 1.01e-19
C25230 a_5891_43370# a_5837_43396# 1.86e-19
C25231 a_n2293_42834# a_8952_43230# 1.55e-19
C25232 a_3537_45260# a_4649_42852# 0.065656f
C25233 a_2711_45572# a_8697_45572# 3.48e-19
C25234 a_9049_44484# a_10490_45724# 1.71e-20
C25235 a_10180_45724# a_10193_42453# 0.145672f
C25236 a_10053_45546# a_8746_45002# 0.075884f
C25237 a_7499_43078# a_11322_45546# 8.22e-21
C25238 a_20365_43914# a_12741_44636# 3.64e-19
C25239 a_11341_43940# a_20202_43084# 0.033215f
C25240 a_21487_43396# a_12549_44172# 2.13e-19
C25241 a_n23_44458# a_n755_45592# 8.98e-19
C25242 a_n2293_43922# a_13259_45724# 2.67e-19
C25243 a_1414_42308# a_2324_44458# 2.25e-19
C25244 a_20447_31679# VCM 0.035344f
C25245 a_11735_46660# VDD 0.407307f
C25246 a_1606_42308# VDAC_P 0.006313f
C25247 a_n2293_46098# a_2698_46116# 6.74e-20
C25248 a_21076_30879# a_4185_45028# 2.52e-19
C25249 a_n901_46420# a_1176_45822# 1.16e-19
C25250 a_3524_46660# a_n755_45592# 5.56e-20
C25251 a_4651_46660# a_n2661_45546# 2.36e-20
C25252 a_16388_46812# a_18819_46122# 1.15e-19
C25253 a_765_45546# a_15015_46420# 4.38e-20
C25254 a_14035_46660# a_6945_45028# 4.05e-19
C25255 en_comp a_1177_38525# 0.205977f
C25256 a_4699_43561# a_4905_42826# 1.43e-19
C25257 a_1568_43370# a_1891_43646# 7.4e-19
C25258 a_9313_44734# a_14635_42282# 0.005265f
C25259 a_n97_42460# a_648_43396# 0.00481f
C25260 a_3422_30871# a_17701_42308# 2.82e-20
C25261 a_3905_42865# a_3935_42891# 0.240349f
C25262 a_18579_44172# a_19164_43230# 5.37e-20
C25263 a_14021_43940# a_16137_43396# 0.002723f
C25264 a_15493_43940# a_19700_43370# 5.37e-20
C25265 a_14955_43940# a_743_42282# 1.64e-22
C25266 a_19279_43940# a_21356_42826# 2.54e-19
C25267 w_11334_34010# a_19120_35138# 0.001523f
C25268 SMPL_ON_P a_n1532_35090# 4.33e-19
C25269 a_n1243_43396# VDD 4.56e-20
C25270 a_15599_45572# a_16019_45002# 0.001742f
C25271 a_16115_45572# a_14537_43396# 3.42e-21
C25272 a_15903_45785# a_15595_45028# 0.003784f
C25273 a_8696_44636# a_13556_45296# 0.022968f
C25274 a_2711_45572# a_11691_44458# 0.058464f
C25275 a_11322_45546# a_11915_45394# 3.21e-19
C25276 a_16147_45260# a_6171_45002# 0.072853f
C25277 a_22959_45572# a_20447_31679# 0.154273f
C25278 a_16104_42674# a_10227_46804# 0.012196f
C25279 a_n1630_35242# a_n2312_38680# 8.58e-19
C25280 a_9396_43370# a_526_44458# 2.4e-19
C25281 a_n97_42460# a_13259_45724# 0.182889f
C25282 a_743_42282# a_1138_42852# 8.9e-20
C25283 a_4099_45572# a_n881_46662# 7.8e-20
C25284 a_5263_45724# a_n1613_43370# 5.35e-21
C25285 a_10053_45546# a_4883_46098# 0.008211f
C25286 a_10193_42453# a_13507_46334# 0.008059f
C25287 a_13163_45724# a_10227_46804# 2.33e-19
C25288 a_15143_45578# a_16327_47482# 8.76e-21
C25289 a_8049_45260# a_14180_46482# 9.26e-19
C25290 a_8685_43396# a_5342_30871# 0.001246f
C25291 a_21487_43396# a_21855_43396# 7.52e-19
C25292 a_10341_43396# a_10518_42984# 5.04e-20
C25293 a_14579_43548# a_12379_42858# 2.62e-21
C25294 a_20512_43084# a_13258_32519# 2.41e-19
C25295 a_3422_30871# a_21613_42308# 0.027998f
C25296 a_4190_30871# a_13887_32519# 0.032018f
C25297 a_743_42282# a_5649_42852# 0.030921f
C25298 VDAC_N C3_N_btm 6.907279f
C25299 a_n467_45028# a_n2012_44484# 9.72e-23
C25300 a_3232_43370# a_10440_44484# 0.042872f
C25301 a_7705_45326# a_6298_44484# 0.004597f
C25302 a_7499_43078# a_7281_43914# 6.26e-21
C25303 a_8162_45546# a_7845_44172# 1.27e-21
C25304 a_3823_42558# a_4185_45028# 1.01e-19
C25305 a_7765_42852# a_n443_42852# 0.004527f
C25306 a_12545_42858# a_n357_42282# 0.042417f
C25307 a_3080_42308# a_n1532_35090# 6.43e-20
C25308 a_16501_45348# a_10227_46804# 4.16e-20
C25309 a_18315_45260# a_16327_47482# 4.78e-19
C25310 a_21359_45002# a_12861_44030# 1.13e-20
C25311 C8_P_btm VDD 0.19922f
C25312 a_949_44458# a_2063_45854# 9.64e-19
C25313 a_2779_44458# a_584_46384# 2.06e-20
C25314 a_n1917_44484# a_n1151_42308# 2.05e-19
C25315 a_16115_45572# a_3090_45724# 0.00765f
C25316 a_13777_45326# a_13747_46662# 1.16e-21
C25317 a_14537_43396# a_5807_45002# 0.001298f
C25318 a_15765_45572# a_15368_46634# 3.33e-19
C25319 a_14180_45002# a_13661_43548# 1.37e-19
C25320 a_3357_43084# a_5907_46634# 0.013466f
C25321 a_3065_45002# a_2107_46812# 2.48e-20
C25322 a_3232_43370# a_n743_46660# 7.45e-20
C25323 a_413_45260# a_479_46660# 2.29e-20
C25324 a_5365_45348# a_n881_46662# 2.78e-19
C25325 a_5263_45724# a_n2293_46098# 0.002594f
C25326 a_5342_30871# a_15953_42852# 5.76e-19
C25327 a_4649_43172# a_4649_42852# 6.96e-20
C25328 a_16409_43396# a_14113_42308# 1.57e-21
C25329 a_743_42282# a_7963_42308# 0.008222f
C25330 a_5649_42852# a_5755_42308# 0.008092f
C25331 a_16137_43396# a_15764_42576# 0.008757f
C25332 a_15567_42826# a_15597_42852# 0.025037f
C25333 a_685_42968# a_564_42282# 3.6e-19
C25334 a_n4334_38528# VDD 0.385889f
C25335 a_6151_47436# a_15928_47570# 2.62e-20
C25336 a_9067_47204# a_9804_47204# 0.001602f
C25337 a_13381_47204# a_n881_46662# 0.025748f
C25338 a_n1435_47204# a_n1613_43370# 2.68e-19
C25339 a_n237_47217# a_n2293_46634# 0.003267f
C25340 SMPL_ON_P a_n2438_43548# 0.003035f
C25341 a_n1151_42308# a_13747_46662# 0.050569f
C25342 a_n2109_47186# a_33_46660# 6.32e-20
C25343 a_n1741_47186# a_n133_46660# 4.48e-20
C25344 a_n815_47178# a_n1021_46688# 0.003455f
C25345 a_327_47204# a_n2661_46634# 0.004931f
C25346 a_20894_47436# a_12465_44636# 2.12e-19
C25347 a_21177_47436# a_4883_46098# 5.42e-19
C25348 a_13507_46334# a_21496_47436# 0.167302f
C25349 a_18780_47178# a_11453_44696# 2.2e-19
C25350 a_8375_44464# a_5891_43370# 0.094782f
C25351 a_20193_45348# a_20512_43084# 0.160912f
C25352 a_2711_45572# a_4190_30871# 0.051595f
C25353 a_n2012_44484# a_n2661_43922# 0.00414f
C25354 a_12607_44458# a_12829_44484# 5.19e-19
C25355 a_11827_44484# a_19237_31679# 3.81e-19
C25356 a_n2293_42834# a_n1441_43940# 0.001195f
C25357 a_19332_42282# a_n357_42282# 1.1e-19
C25358 a_19418_45938# VDD 4.6e-19
C25359 a_22959_42860# RST_Z 0.001357f
C25360 a_14797_45144# a_3483_46348# 2.2e-21
C25361 a_626_44172# a_1138_42852# 0.010739f
C25362 a_1145_45348# a_1176_45822# 5.36e-22
C25363 a_20159_44458# a_19321_45002# 0.065041f
C25364 a_8701_44490# a_8270_45546# 0.015888f
C25365 a_16112_44458# a_6755_46942# 0.023983f
C25366 a_20640_44752# a_13747_46662# 0.027627f
C25367 a_n356_44636# a_5257_43370# 1.18e-20
C25368 a_19929_45028# a_19466_46812# 0.012303f
C25369 a_16020_45572# a_13259_45724# 0.024851f
C25370 a_8696_44636# a_16375_45002# 0.043034f
C25371 a_11823_42460# a_n443_42852# 0.356965f
C25372 a_18799_45938# a_8049_45260# 0.004297f
C25373 a_8191_45002# a_8199_44636# 0.234072f
C25374 a_3232_43370# a_11189_46129# 3.91e-20
C25375 a_6171_45002# a_9290_44172# 0.028032f
C25376 a_413_45260# a_17583_46090# 1.29e-21
C25377 a_7705_45326# a_5937_45572# 0.070066f
C25378 a_5111_44636# a_10903_43370# 3.25e-20
C25379 a_11341_43940# a_2063_45854# 0.001102f
C25380 a_4921_42308# a_3905_42308# 6.09e-20
C25381 a_2123_42473# a_5742_30871# 1.16e-20
C25382 a_5932_42308# a_7227_42308# 1.68e-20
C25383 a_6171_42473# a_6123_31319# 8.95e-21
C25384 CAL_P a_21589_35634# 0.00593f
C25385 a_n1386_35608# a_n923_35174# 0.201937f
C25386 a_n1838_35608# EN_VIN_BSTR_P 2.62e-19
C25387 a_n237_47217# a_9625_46129# 2.69e-19
C25388 a_2063_45854# a_5497_46414# 1.5e-19
C25389 a_n1741_47186# a_11387_46155# 4.53e-19
C25390 a_n1151_42308# a_4419_46090# 2.82e-19
C25391 a_5807_45002# a_3090_45724# 0.032418f
C25392 a_13747_46662# a_14084_46812# 0.038349f
C25393 a_3877_44458# a_5907_46634# 0.073504f
C25394 a_4646_46812# a_5167_46660# 0.033486f
C25395 a_4955_46873# a_4817_46660# 0.318259f
C25396 a_4651_46660# a_5385_46902# 0.053479f
C25397 a_n2293_46634# a_8270_45546# 0.030248f
C25398 a_2107_46812# a_10249_46116# 4.12e-19
C25399 a_11309_47204# a_12156_46660# 4.26e-19
C25400 a_3815_47204# a_3483_46348# 2.65e-20
C25401 a_3785_47178# a_3699_46348# 4.8e-20
C25402 a_n443_46116# a_2521_46116# 0.00999f
C25403 a_18479_47436# a_18280_46660# 4.42e-20
C25404 a_16327_47482# a_20202_43084# 0.475502f
C25405 a_21177_47436# a_21188_46660# 5.06e-21
C25406 a_13507_46334# a_21363_46634# 0.029223f
C25407 a_4883_46098# a_20841_46902# 7.76e-20
C25408 a_12465_44636# a_20411_46873# 2.37e-20
C25409 a_11453_44696# a_18285_46348# 0.236771f
C25410 a_n1059_45260# a_12895_43230# 0.003645f
C25411 a_n913_45002# a_13113_42826# 0.018663f
C25412 a_n2017_45002# a_13635_43156# 4.66e-19
C25413 a_3537_45260# a_5755_42852# 0.088502f
C25414 a_5343_44458# a_3626_43646# 0.001955f
C25415 a_18579_44172# a_18079_43940# 3.67e-19
C25416 a_n2661_42834# a_6671_43940# 6.64e-19
C25417 a_11827_44484# a_9145_43396# 6.87e-20
C25418 a_19279_43940# a_19328_44172# 0.120319f
C25419 a_5244_44056# a_5663_43940# 7.46e-20
C25420 a_5013_44260# a_5495_43940# 0.251039f
C25421 a_20159_44458# a_20623_43914# 0.005333f
C25422 a_20679_44626# a_19862_44208# 0.001682f
C25423 a_20362_44736# a_20365_43914# 0.012553f
C25424 a_18989_43940# a_n97_42460# 1.52e-19
C25425 a_742_44458# a_648_43396# 6.39e-22
C25426 a_18248_44752# VDD 0.251171f
C25427 a_n4064_39616# C6_P_btm 1.1e-19
C25428 a_n3420_39616# C4_P_btm 3.39e-20
C25429 a_n3420_39072# a_n923_35174# 0.004736f
C25430 a_16137_43396# a_13507_46334# 1.52e-19
C25431 a_16867_43762# a_16327_47482# 0.012196f
C25432 a_16823_43084# a_12861_44030# 6.87e-21
C25433 a_n1853_43023# a_n1151_42308# 0.021207f
C25434 a_17737_43940# a_15227_44166# 0.013191f
C25435 a_19478_44306# a_3090_45724# 0.027139f
C25436 a_3457_43396# a_768_44030# 3.04e-20
C25437 a_1987_43646# a_n2293_46634# 5.42e-20
C25438 a_8975_43940# a_10586_45546# 2.76e-20
C25439 a_n935_46688# VDD 2.29e-19
C25440 a_n4064_40160# a_n3607_38528# 5.58e-20
C25441 a_n3565_39590# a_n2302_38778# 8.95e-20
C25442 a_n3420_39072# a_n4064_39072# 4.93427f
C25443 a_1343_38525# a_1736_39043# 0.310247f
C25444 a_5742_30871# C3_N_btm 0.030866f
C25445 a_n3674_38216# a_n4064_37984# 0.65176f
C25446 a_n4318_37592# a_n3420_37984# 0.404896f
C25447 a_n4318_38216# a_n4251_38304# 2.47e-19
C25448 a_14976_45028# a_3483_46348# 3.99e-20
C25449 a_20107_46660# a_20731_47026# 9.73e-19
C25450 a_20411_46873# a_20528_46660# 0.170785f
C25451 a_20841_46902# a_21188_46660# 0.051162f
C25452 a_20273_46660# a_22000_46634# 2.02e-19
C25453 a_18285_46348# a_17639_46660# 0.003315f
C25454 a_13747_46662# a_19240_46482# 0.012097f
C25455 a_2107_46812# a_8781_46436# 2.53e-19
C25456 a_n881_46662# a_n452_45724# 0.005284f
C25457 a_8270_45546# a_9625_46129# 0.001176f
C25458 a_6755_46942# a_13925_46122# 4.42e-19
C25459 a_10428_46928# a_2324_44458# 7.92e-21
C25460 a_8846_46660# a_8199_44636# 6.28e-20
C25461 a_9672_43914# a_8685_43396# 3.33e-20
C25462 a_1241_43940# a_1049_43396# 3.88e-19
C25463 a_3422_30871# a_4361_42308# 0.096125f
C25464 a_n2293_43922# a_10518_42984# 5.88e-21
C25465 a_n2661_42834# a_10796_42968# 6.58e-21
C25466 a_9313_44734# a_14543_43071# 0.00414f
C25467 a_20512_43084# a_20301_43646# 2.11e-20
C25468 a_18184_42460# a_22400_42852# 0.16156f
C25469 a_19319_43548# a_18533_43940# 2.47e-20
C25470 a_n2661_43370# a_n1630_35242# 2.37e-20
C25471 a_5745_43940# a_n97_42460# 8.52e-20
C25472 en_comp a_18057_42282# 2.2e-20
C25473 a_n1059_45260# a_18220_42308# 0.00103f
C25474 a_3737_43940# VDD 0.18423f
C25475 a_9049_44484# a_6171_45002# 0.026882f
C25476 a_16147_45260# a_18909_45814# 3.16e-20
C25477 a_18175_45572# a_18341_45572# 0.577068f
C25478 a_4099_45572# a_1307_43914# 1.48e-22
C25479 a_7287_43370# a_3483_46348# 3.53e-21
C25480 a_10341_43396# a_20202_43084# 0.037863f
C25481 a_18783_43370# a_17339_46660# 0.02025f
C25482 a_13678_32519# a_19692_46634# 0.004218f
C25483 a_6101_44260# a_n357_42282# 4.36e-20
C25484 a_n2472_42282# a_n2312_39304# 3.28e-20
C25485 a_n4318_38216# a_n2312_40392# 0.025276f
C25486 VDAC_P C9_P_btm 0.441881p
C25487 a_2324_44458# VDD 2.73366f
C25488 a_10193_42453# a_n1741_47186# 6.98e-20
C25489 a_8568_45546# a_n971_45724# 0.009964f
C25490 a_6598_45938# a_n1151_42308# 9.17e-20
C25491 a_5263_45724# a_4791_45118# 0.021183f
C25492 a_4099_45572# a_n443_46116# 1e-20
C25493 a_n2293_46098# a_380_45546# 0.007518f
C25494 a_n1853_46287# a_n863_45724# 0.019522f
C25495 a_n1423_46090# a_n2293_45546# 0.001036f
C25496 a_n1076_46494# a_n2661_45546# 1.51e-20
C25497 a_n1991_46122# a_n1079_45724# 0.001345f
C25498 a_13925_46122# a_8049_45260# 0.009027f
C25499 a_11387_46155# a_10586_45546# 7.66e-19
C25500 a_n4209_38216# a_n2946_37690# 5.11e-19
C25501 a_n3565_38216# a_n3690_37440# 7.25e-19
C25502 a_10341_43396# a_16867_43762# 0.001683f
C25503 a_4235_43370# a_3681_42891# 7.84e-21
C25504 a_15095_43370# a_15231_43396# 0.001002f
C25505 a_15781_43660# a_16409_43396# 2.7e-19
C25506 a_n3674_39768# a_n3674_38216# 0.02323f
C25507 a_1414_42308# a_1606_42308# 0.056716f
C25508 a_14955_43396# a_15125_43396# 0.001675f
C25509 a_14401_32519# a_5534_30871# 0.339008f
C25510 a_9313_44734# a_19511_42282# 0.001387f
C25511 a_895_43940# a_1184_42692# 2.55e-21
C25512 a_n97_42460# a_10518_42984# 1.55e-20
C25513 a_n1557_42282# a_685_42968# 0.003946f
C25514 a_8685_43396# a_743_42282# 1.88e-19
C25515 a_4093_43548# a_3935_42891# 0.00342f
C25516 a_13747_46662# START 0.062289f
C25517 a_16119_47582# CLK 2.67e-19
C25518 a_8387_43230# VDD 0.200672f
C25519 a_13904_45546# a_13857_44734# 4.52e-21
C25520 a_11652_45724# a_11541_44484# 1.11e-20
C25521 a_13249_42308# a_13468_44734# 2.67e-20
C25522 a_5205_44484# a_n2661_43370# 0.033807f
C25523 a_8953_45002# a_8560_45348# 0.001921f
C25524 en_comp a_18494_42460# 6.64e-20
C25525 a_21513_45002# a_19721_31679# 9.71e-20
C25526 a_n1059_45260# a_11827_44484# 9.98e-20
C25527 a_6171_45002# a_13105_45348# 5.33e-20
C25528 a_14097_32519# a_20820_30879# 0.052932f
C25529 a_20356_42852# a_20202_43084# 0.003203f
C25530 a_9223_42460# a_3090_45724# 1.31e-21
C25531 a_13678_32519# a_20692_30879# 0.051702f
C25532 a_n4064_37984# w_1575_34946# 3.17e-19
C25533 a_6511_45714# a_3090_45724# 1.98e-21
C25534 a_2711_45572# a_15227_44166# 0.113396f
C25535 a_7499_43078# a_8654_47026# 5.36e-21
C25536 a_21188_45572# a_13747_46662# 9.45e-19
C25537 a_20623_45572# a_19321_45002# 0.001031f
C25538 a_3357_43084# a_768_44030# 0.09747f
C25539 a_2437_43646# a_13569_47204# 5.26e-20
C25540 a_n2017_45002# a_n1613_43370# 0.015448f
C25541 a_13777_45326# a_11599_46634# 8.08e-19
C25542 a_5111_44636# a_4883_46098# 0.048482f
C25543 a_8953_45002# a_10227_46804# 0.017713f
C25544 a_5837_45348# a_4791_45118# 1.43e-20
C25545 a_n2661_43370# a_n971_45724# 0.064346f
C25546 a_8147_43396# a_8325_42308# 8.68e-22
C25547 a_20974_43370# a_19511_42282# 1.07e-21
C25548 a_16795_42852# a_17595_43084# 0.010079f
C25549 a_21381_43940# a_13258_32519# 1.65e-19
C25550 a_12281_43396# a_1606_42308# 1.94e-20
C25551 a_3626_43646# a_12563_42308# 0.005049f
C25552 a_2982_43646# a_13575_42558# 1.36e-19
C25553 a_4520_42826# a_5193_43172# 1.24e-19
C25554 a_n97_42460# a_16197_42308# 3.2e-21
C25555 a_6491_46660# a_6575_47204# 0.029984f
C25556 a_4915_47217# a_11459_47204# 0.03966f
C25557 a_6151_47436# a_9863_47436# 0.030884f
C25558 a_n1151_42308# a_11599_46634# 0.116147f
C25559 a_4791_45118# a_n1435_47204# 5.92e-19
C25560 a_16522_42674# VDD 0.077608f
C25561 a_n913_45002# a_n2661_42282# 0.054259f
C25562 a_20841_45814# a_20935_43940# 6.15e-21
C25563 a_3232_43370# a_5244_44056# 0.017099f
C25564 a_3537_45260# a_7845_44172# 0.001398f
C25565 a_5111_44636# a_5663_43940# 0.001818f
C25566 a_5691_45260# a_5013_44260# 9.29e-19
C25567 a_n2661_44458# a_7_44811# 3.19e-19
C25568 a_n2267_44484# a_n356_44636# 1.82e-20
C25569 a_n2129_44697# a_n23_44458# 2.23e-19
C25570 a_18479_45785# a_14021_43940# 0.025329f
C25571 a_n1699_44726# a_n1655_44484# 3.69e-19
C25572 a_n1917_44484# a_n1821_44484# 0.013793f
C25573 a_10440_44484# a_8975_43940# 0.045841f
C25574 a_5379_42460# a_n357_42282# 0.007085f
C25575 a_961_42354# a_n443_42852# 0.002615f
C25576 a_5267_42460# a_n755_45592# 1.87e-19
C25577 a_13527_45546# VDD 0.1902f
C25578 a_13467_32519# VCM 0.020152f
C25579 a_13678_32519# VIN_N 0.069898f
C25580 a_17478_45572# a_17957_46116# 1.77e-19
C25581 a_16335_44484# a_10227_46804# 4.36e-20
C25582 a_19006_44850# a_16327_47482# 0.028858f
C25583 a_19279_43940# a_12861_44030# 0.152657f
C25584 a_2998_44172# a_n971_45724# 2.34e-20
C25585 a_n1899_43946# a_n1151_42308# 2.4e-19
C25586 a_644_44056# a_584_46384# 0.004876f
C25587 a_9482_43914# a_13059_46348# 0.448068f
C25588 a_2437_43646# a_2202_46116# 0.022869f
C25589 a_n2109_45247# a_n2157_46122# 1.34e-21
C25590 a_6298_44484# a_2107_46812# 4.34e-21
C25591 a_8975_43940# a_n743_46660# 7.99e-22
C25592 a_n2017_45002# a_n2293_46098# 1.65e-19
C25593 a_n2293_45010# a_n1853_46287# 2.07e-20
C25594 a_742_44458# a_1799_45572# 1.46e-20
C25595 a_11962_45724# a_8049_45260# 0.019556f
C25596 a_10193_42453# a_10586_45546# 0.380236f
C25597 a_n473_42460# a_n327_42558# 0.171361f
C25598 a_n4318_38680# a_n4334_38528# 0.08371f
C25599 a_196_42282# a_n784_42308# 0.00268f
C25600 a_n961_42308# a_n3674_37592# 0.005438f
C25601 COMP_P a_n1630_35242# 2.45645f
C25602 a_17701_42308# a_7174_31319# 2.14e-20
C25603 a_n2661_46634# a_1983_46706# 0.005467f
C25604 a_n2293_46634# a_1123_46634# 6.6e-21
C25605 a_n743_46660# a_n133_46660# 0.205551f
C25606 a_n1925_46634# a_33_46660# 0.0095f
C25607 a_n1021_46688# a_171_46873# 1.98e-19
C25608 a_768_44030# a_3877_44458# 0.012394f
C25609 a_n1613_43370# a_3633_46660# 6.03e-19
C25610 a_10227_46804# a_10768_47026# 0.012196f
C25611 a_14955_47212# a_15009_46634# 0.001517f
C25612 a_13717_47436# a_15559_46634# 2.06e-21
C25613 a_12861_44030# a_15368_46634# 0.066698f
C25614 a_327_47204# a_765_45546# 8.96e-19
C25615 a_n1151_42308# a_13693_46688# 2.97e-19
C25616 a_9482_43914# a_15095_43370# 1.57e-19
C25617 a_18287_44626# a_15493_43940# 1.79e-20
C25618 a_13556_45296# a_14205_43396# 0.012255f
C25619 a_14180_45002# a_14579_43548# 9.2e-22
C25620 a_20193_45348# a_21381_43940# 0.01388f
C25621 a_4223_44672# a_3992_43940# 1.9e-19
C25622 a_5891_43370# a_10949_43914# 0.005033f
C25623 a_14537_43396# a_13667_43396# 2.79e-19
C25624 a_7499_43078# a_8483_43230# 8.28e-19
C25625 a_n2661_43922# a_1241_44260# 3.45e-19
C25626 a_n2661_42834# a_1525_44260# 1.72e-19
C25627 a_n2293_42834# a_n998_43396# 1.67e-19
C25628 a_n913_45002# a_16823_43084# 1.15e-20
C25629 a_2113_38308# VDD 0.004903f
C25630 a_16922_45042# VDD 1.54713f
C25631 a_6123_31319# VIN_N 0.01057f
C25632 a_5742_30871# C7_P_btm 0.04157f
C25633 a_n2661_43922# a_11415_45002# 2.28e-19
C25634 a_18797_44260# a_12549_44172# 5.67e-19
C25635 a_1423_45028# a_n2661_45546# 0.020024f
C25636 a_n699_43396# a_2324_44458# 0.070009f
C25637 a_12607_44458# a_9290_44172# 3.67e-20
C25638 a_3626_43646# a_10227_46804# 0.011826f
C25639 a_10341_43396# a_2063_45854# 1e-19
C25640 a_21335_42336# a_21887_42336# 0.001613f
C25641 a_13258_32519# a_21125_42558# 0.002663f
C25642 a_5742_30871# a_n3565_38502# 4.45e-21
C25643 a_n310_47570# VDD 3.35e-19
C25644 a_5342_30871# a_7754_38470# 1.06e-19
C25645 a_3699_46634# a_3699_46348# 0.005275f
C25646 a_3524_46660# a_3483_46348# 6.03e-20
C25647 a_15368_46634# a_14180_46812# 4.62e-20
C25648 a_12816_46660# a_13059_46348# 3.67e-19
C25649 a_n881_46662# a_2981_46116# 0.026038f
C25650 a_13747_46662# a_19553_46090# 3.31e-20
C25651 a_19321_45002# a_18819_46122# 0.018323f
C25652 a_n743_46660# a_11387_46155# 0.007599f
C25653 a_2107_46812# a_5937_45572# 0.027091f
C25654 a_16285_47570# a_6945_45028# 1.12e-19
C25655 a_5807_45002# a_20075_46420# 4.74e-19
C25656 a_n1613_43370# a_526_44458# 0.826565f
C25657 a_2905_45572# a_3218_45724# 0.021505f
C25658 a_n237_47217# a_2277_45546# 0.104529f
C25659 a_n1151_42308# a_1848_45724# 7.61e-21
C25660 a_n443_46116# a_n452_45724# 0.188857f
C25661 a_327_47204# a_509_45822# 1.76e-20
C25662 a_3785_47178# a_n755_45592# 8.67e-21
C25663 a_11599_46634# a_19240_46482# 0.016662f
C25664 SMPL_ON_N a_8049_45260# 1.15e-19
C25665 a_n913_45002# a_3497_42558# 0.004643f
C25666 a_n2017_45002# a_3905_42558# 0.006025f
C25667 a_5343_44458# a_8037_42858# 0.019942f
C25668 a_14955_43940# a_15037_43940# 0.171361f
C25669 a_18184_42460# a_22223_42860# 0.03037f
C25670 a_11827_44484# a_19987_42826# 2.96e-20
C25671 a_9313_44734# a_21259_43561# 1.06e-19
C25672 a_1414_42308# a_3539_42460# 5.28e-20
C25673 a_2479_44172# a_2982_43646# 0.019219f
C25674 a_5244_44056# a_4905_42826# 0.002354f
C25675 a_n875_44318# VDD 4.97e-20
C25676 a_10193_42453# a_18175_45572# 5.07e-21
C25677 a_13163_45724# a_13297_45572# 0.001089f
C25678 a_11341_43940# a_17715_44484# 0.001541f
C25679 a_13565_44260# a_10903_43370# 3.14e-19
C25680 a_12603_44260# a_12594_46348# 1e-20
C25681 a_n1630_35242# a_n2497_47436# 2.73e-20
C25682 COMP_P a_n971_45724# 8.93e-21
C25683 a_15567_42826# a_12549_44172# 1.56e-19
C25684 a_13667_43396# a_3090_45724# 1.98e-20
C25685 a_5755_42852# a_n2293_46634# 4.15e-20
C25686 a_3626_43646# a_17339_46660# 3.03e-20
C25687 a_21350_47026# VDD 4.6e-19
C25688 a_n2293_46098# a_526_44458# 0.053029f
C25689 a_n1423_46090# a_n914_46116# 2.6e-19
C25690 a_3090_45724# a_n755_45592# 0.051041f
C25691 a_16388_46812# a_18147_46436# 0.004345f
C25692 a_9290_44172# a_10903_43370# 0.340316f
C25693 a_7920_46348# a_2324_44458# 6.6e-21
C25694 a_11189_46129# a_11387_46155# 0.320331f
C25695 a_7174_31319# a_3754_38470# 2.41e-19
C25696 a_20974_43370# a_21259_43561# 0.049502f
C25697 a_n97_42460# a_16867_43762# 1.22e-19
C25698 a_n356_44636# a_9223_42460# 1.4e-19
C25699 a_14401_32519# a_4190_30871# 0.10855f
C25700 a_8147_43396# a_9145_43396# 1.64e-19
C25701 a_11599_46634# START 2.57e-19
C25702 a_11031_47542# CLK 4.33e-19
C25703 a_11459_47204# DATA[5] 0.370451f
C25704 a_n1435_47204# DATA[3] 0.02843f
C25705 a_15507_47210# RST_Z 2.28e-19
C25706 a_15743_43084# VDD 0.572249f
C25707 a_5147_45002# a_6171_45002# 3.36e-19
C25708 a_5111_44636# a_3232_43370# 0.134191f
C25709 a_4927_45028# a_5691_45260# 0.018415f
C25710 a_10180_45724# a_10057_43914# 0.002709f
C25711 a_8746_45002# a_10334_44484# 0.019787f
C25712 a_10907_45822# a_n2661_44458# 3.96e-19
C25713 a_15599_45572# a_11827_44484# 4.86e-21
C25714 a_10341_42308# a_4185_45028# 1.48e-20
C25715 a_20712_42282# a_12549_44172# 3.18e-19
C25716 a_7227_42308# a_4646_46812# 1.62e-20
C25717 a_6547_43396# a_n755_45592# 7.25e-21
C25718 a_7287_43370# a_n357_42282# 0.002031f
C25719 a_2982_43646# a_n443_42852# 0.037773f
C25720 a_4181_43396# a_n2661_45546# 0.009936f
C25721 a_7765_42852# a_8199_44636# 1.98e-19
C25722 a_18479_45785# a_13507_46334# 8.2e-20
C25723 a_20107_45572# a_16327_47482# 0.674639f
C25724 a_18596_45572# a_18597_46090# 8.84e-19
C25725 a_19256_45572# a_19386_47436# 6.77e-21
C25726 a_18799_45938# a_18780_47178# 9.94e-22
C25727 a_3357_43084# a_9067_47204# 5.7e-19
C25728 a_2437_43646# a_9313_45822# 0.045826f
C25729 a_n37_45144# a_584_46384# 9.32e-20
C25730 a_3429_45260# a_n237_47217# 7.06e-21
C25731 a_n2017_45002# a_4791_45118# 0.023951f
C25732 a_6171_45002# a_n2109_47186# 1.79e-19
C25733 en_comp a_n1151_42308# 8.03e-21
C25734 a_11823_42460# a_n2661_46634# 0.331717f
C25735 a_10193_42453# a_n743_46660# 0.25279f
C25736 a_9145_43396# a_13569_43230# 1.23e-19
C25737 a_13678_32519# a_5342_30871# 0.028488f
C25738 a_19328_44172# a_19332_42282# 1.13e-21
C25739 a_15493_43940# a_17124_42282# 1.54e-21
C25740 a_9165_43940# a_9223_42460# 4.51e-21
C25741 a_n1557_42282# a_n1329_42308# 0.075734f
C25742 a_4190_30871# a_18817_42826# 0.011301f
C25743 a_743_42282# a_17333_42852# 8.08e-20
C25744 a_1847_42826# a_2905_42968# 0.097535f
C25745 a_458_43396# a_1184_42692# 1.51e-20
C25746 a_7754_40130# a_4338_37500# 0.030623f
C25747 a_7754_38636# a_3754_38470# 0.037604f
C25748 a_1606_42308# VDD 0.631207f
C25749 a_n1920_47178# a_n1605_47204# 0.08571f
C25750 a_n2109_47186# a_n815_47178# 0.160027f
C25751 a_n2497_47436# a_n971_45724# 0.229429f
C25752 a_n1741_47186# SMPL_ON_P 0.178214f
C25753 a_22959_45036# a_19721_31679# 0.156264f
C25754 a_11136_45572# a_10729_43914# 1.39e-20
C25755 a_20193_45348# a_19929_45028# 4.23e-19
C25756 a_11691_44458# a_20205_45028# 2.19e-19
C25757 a_1423_45028# a_8238_44734# 2.37e-19
C25758 a_n1059_45260# a_18005_44484# 5.53e-20
C25759 a_18057_42282# a_4185_45028# 7.92e-20
C25760 a_3905_42558# a_526_44458# 0.006254f
C25761 a_5934_30871# a_n2956_39304# 5.05e-21
C25762 a_22469_40625# SMPL_ON_N 0.03403f
C25763 a_16680_45572# a_12741_44636# 5.61e-19
C25764 a_17478_45572# a_11415_45002# 0.002665f
C25765 a_9241_45822# a_3483_46348# 3e-19
C25766 a_10775_45002# a_10428_46928# 2.17e-22
C25767 a_18911_45144# a_19321_45002# 0.050257f
C25768 a_18184_42460# a_13747_46662# 0.123281f
C25769 a_18494_42460# a_13661_43548# 0.049953f
C25770 a_3495_45348# a_3877_44458# 1.26e-19
C25771 a_7229_43940# a_6755_46942# 6.9e-21
C25772 a_413_45260# a_11813_46116# 1.63e-20
C25773 a_9049_44484# a_10903_43370# 2.44e-20
C25774 a_10193_42453# a_11189_46129# 0.123385f
C25775 a_8746_45002# a_9290_44172# 0.004141f
C25776 a_10490_45724# a_10355_46116# 0.01084f
C25777 a_11823_42460# a_8199_44636# 0.00368f
C25778 a_n2840_44458# a_n1613_43370# 1.2e-19
C25779 a_10334_44484# a_4883_46098# 3.73e-21
C25780 a_18374_44850# a_16327_47482# 0.16003f
C25781 a_9313_44734# a_4915_47217# 1.84e-22
C25782 a_21487_43396# a_21613_42308# 9.66e-20
C25783 a_10083_42826# a_10723_42308# 0.001074f
C25784 a_10518_42984# a_10533_42308# 0.001423f
C25785 a_10341_42308# a_9803_42558# 0.108853f
C25786 a_13467_32519# a_21335_42336# 0.005979f
C25787 a_4361_42308# a_7174_31319# 0.024432f
C25788 a_5649_42852# a_13258_32519# 0.040931f
C25789 a_5342_30871# a_6123_31319# 0.018227f
C25790 a_5534_30871# a_5934_30871# 0.018227f
C25791 a_n2293_42282# a_2725_42558# 1.65e-19
C25792 a_11117_47542# a_11309_47204# 5.76e-19
C25793 a_n881_46662# a_13675_47204# 0.001593f
C25794 a_n1151_42308# a_7411_46660# 2.81e-19
C25795 a_n237_47217# a_6755_46942# 0.073038f
C25796 a_2063_45854# a_8667_46634# 0.00593f
C25797 a_n971_45724# a_6682_46987# 0.006879f
C25798 a_6151_47436# a_5907_46634# 9.7e-19
C25799 a_5815_47464# a_5732_46660# 0.002408f
C25800 a_4915_47217# a_5072_46660# 1.11e-19
C25801 a_6575_47204# a_4646_46812# 1.71e-19
C25802 a_n2312_40392# a_n2956_39768# 0.056063f
C25803 a_n2312_39304# a_n2840_46634# 0.018018f
C25804 C1_N_btm VDD 0.264503f
C25805 a_3232_43370# a_4235_43370# 6.06e-20
C25806 a_n2017_45002# a_8791_43396# 2.77e-21
C25807 a_n1059_45260# a_8147_43396# 4.32e-21
C25808 a_2382_45260# a_3540_43646# 0.006906f
C25809 a_3065_45002# a_2896_43646# 6.3e-21
C25810 a_5111_44636# a_4905_42826# 0.128918f
C25811 a_n2661_43922# a_11967_42832# 1.74e-20
C25812 a_5883_43914# a_7542_44172# 0.187537f
C25813 a_19778_44110# a_20365_43914# 1.6e-19
C25814 a_18184_42460# a_20269_44172# 0.002397f
C25815 a_11827_44484# a_18326_43940# 0.001776f
C25816 a_11691_44458# a_15682_43940# 0.013321f
C25817 a_18494_42460# a_19862_44208# 0.019692f
C25818 a_10775_45002# VDD 0.148349f
C25819 COMP_P a_11530_34132# 0.018284f
C25820 a_22400_42852# RST_Z 0.059674f
C25821 a_7229_43940# a_8049_45260# 0.014199f
C25822 a_8137_45348# a_2324_44458# 4.79e-19
C25823 a_14021_43940# a_13507_46334# 0.01995f
C25824 a_104_43370# a_584_46384# 0.001171f
C25825 a_1427_43646# a_n2497_47436# 8.12e-20
C25826 a_18494_42460# a_4185_45028# 2.49e-19
C25827 a_9672_43914# a_768_44030# 0.006402f
C25828 a_7845_44172# a_n2293_46634# 3.2e-20
C25829 a_n4318_39768# a_n2442_46660# 0.023739f
C25830 a_17767_44458# a_17339_46660# 9.16e-19
C25831 a_1239_47204# VDD 0.278979f
C25832 a_n784_42308# a_n3420_39072# 0.003982f
C25833 a_n1630_35242# a_n4209_39304# 4.66e-19
C25834 a_n3674_37592# a_n3565_39304# 6.52e-20
C25835 a_n3674_38680# a_n4209_38502# 0.04481f
C25836 a_6761_42308# a_7174_31319# 4.88e-21
C25837 a_14113_42308# a_15890_42674# 0.022182f
C25838 a_15486_42560# a_15803_42450# 0.102355f
C25839 a_13747_46662# a_12741_44636# 0.099721f
C25840 a_19594_46812# a_11415_45002# 2.74e-20
C25841 a_6755_46942# a_8270_45546# 0.045608f
C25842 a_10428_46928# a_11186_47026# 0.055625f
C25843 a_10467_46802# a_10768_47026# 9.73e-19
C25844 a_1983_46706# a_765_45546# 9.01e-19
C25845 a_10249_46116# a_10384_47026# 5.86e-19
C25846 a_n881_46662# a_167_45260# 0.108232f
C25847 a_n1613_43370# a_2521_46116# 8.1e-20
C25848 a_4883_46098# a_9290_44172# 0.055265f
C25849 a_11599_46634# a_19553_46090# 0.021903f
C25850 a_16327_47482# a_17715_44484# 0.03083f
C25851 a_10227_46804# a_15015_46420# 0.287571f
C25852 a_16763_47508# a_15682_46116# 0.001945f
C25853 a_n1435_47204# a_6945_45028# 0.030745f
C25854 a_n237_47217# a_8049_45260# 0.109887f
C25855 a_4791_45118# a_526_44458# 0.042209f
C25856 a_n443_46116# a_2981_46116# 0.017561f
C25857 a_18374_44850# a_10341_43396# 3.04e-21
C25858 a_2479_44172# a_2253_43940# 0.010537f
C25859 a_10729_43914# a_11750_44172# 0.144893f
C25860 a_10949_43914# a_10807_43548# 0.034945f
C25861 a_20193_45348# a_5649_42852# 0.052027f
C25862 a_11823_42460# a_13070_42354# 0.077142f
C25863 a_10193_42453# a_15486_42560# 8.28e-20
C25864 a_2711_45572# a_19511_42282# 0.234026f
C25865 a_2127_44172# a_2455_43940# 0.096132f
C25866 a_895_43940# a_1443_43940# 0.016028f
C25867 a_n2293_42834# a_9127_43156# 4.88e-19
C25868 a_n913_45002# a_11136_42852# 0.026537f
C25869 a_3537_45260# a_4149_42891# 2.78e-19
C25870 a_9049_44484# a_8746_45002# 0.025877f
C25871 a_2711_45572# a_8192_45572# 0.005217f
C25872 a_6598_45938# a_6977_45572# 3.16e-19
C25873 a_7499_43078# a_10490_45724# 4.9e-20
C25874 a_10053_45546# a_10193_42453# 0.086012f
C25875 a_20269_44172# a_12741_44636# 3.52e-20
C25876 a_21115_43940# a_20202_43084# 1.71e-19
C25877 a_743_42282# a_768_44030# 1.92e-19
C25878 a_20556_43646# a_12549_44172# 0.125209f
C25879 a_15743_43084# a_22612_30879# 4.17e-20
C25880 a_n356_44636# a_n755_45592# 2.42652f
C25881 a_n23_44458# a_n357_42282# 4.49e-20
C25882 a_14539_43914# a_n443_42852# 7.29e-19
C25883 a_8037_42858# a_10227_46804# 1.91e-20
C25884 a_12545_42858# a_12861_44030# 1.63e-20
C25885 a_20447_31679# VREF_GND 0.00199f
C25886 a_11186_47026# VDD 0.077608f
C25887 a_5932_42308# a_3754_38470# 2.78e-19
C25888 a_n2293_46098# a_2521_46116# 1.28e-20
C25889 a_376_46348# a_472_46348# 0.318161f
C25890 a_8270_45546# a_8049_45260# 0.321896f
C25891 a_4646_46812# a_n2661_45546# 7e-20
C25892 a_3699_46634# a_n755_45592# 3.16e-20
C25893 a_2609_46660# a_2957_45546# 7.62e-19
C25894 a_2107_46812# a_n443_42852# 1.15e-19
C25895 a_16388_46812# a_17957_46116# 0.140894f
C25896 a_13885_46660# a_6945_45028# 7.75e-21
C25897 a_12925_46660# a_10809_44734# 7.99e-21
C25898 a_n97_42460# a_548_43396# 9.03e-19
C25899 a_4235_43370# a_4905_42826# 8.27e-21
C25900 a_1756_43548# a_n1557_42282# 1.14e-20
C25901 a_9313_44734# a_13291_42460# 0.003344f
C25902 a_18579_44172# a_19339_43156# 3.57e-20
C25903 a_3422_30871# a_17595_43084# 6.38e-21
C25904 a_3905_42865# a_3681_42891# 0.101054f
C25905 a_2998_44172# a_4520_42826# 5.74e-20
C25906 a_15493_43940# a_19268_43646# 9.38e-20
C25907 a_15037_43940# a_8685_43396# 6.84e-19
C25908 a_1568_43370# a_1427_43646# 0.046825f
C25909 a_4699_43561# a_3080_42308# 0.223965f
C25910 a_13483_43940# a_743_42282# 4.27e-21
C25911 a_20679_44626# a_21671_42860# 3.31e-21
C25912 w_11334_34010# a_18194_35068# 0.796644f
C25913 SMPL_ON_P a_n1386_35608# 0.012082f
C25914 a_3539_42460# VDD 0.363092f
C25915 a_15599_45572# a_15595_45028# 2.01e-19
C25916 a_11322_45546# a_n2661_43370# 0.01285f
C25917 a_16333_45814# a_14537_43396# 4.99e-21
C25918 a_8696_44636# a_9482_43914# 0.042504f
C25919 a_19963_31679# a_20447_31679# 0.069779f
C25920 a_10341_43396# a_17715_44484# 1.37e-19
C25921 a_n3420_39072# SMPL_ON_P 1.03e-20
C25922 a_8791_43396# a_526_44458# 1.78e-20
C25923 a_12839_46116# VDD 0.347766f
C25924 a_4099_45572# a_n1613_43370# 1.78e-20
C25925 a_9049_44484# a_4883_46098# 0.001404f
C25926 a_12791_45546# a_10227_46804# 1.59e-20
C25927 a_15037_45618# a_4915_47217# 2.32e-22
C25928 a_9159_45572# a_9067_47204# 6.28e-22
C25929 a_n2956_38680# a_n2956_38216# 0.10753f
C25930 a_8685_43396# a_15279_43071# 0.011343f
C25931 a_21487_43396# a_4361_42308# 0.077645f
C25932 a_10341_43396# a_10083_42826# 0.002266f
C25933 a_8333_44056# a_5934_30871# 2.88e-21
C25934 a_3422_30871# a_21887_42336# 0.003456f
C25935 VDAC_N C2_N_btm 3.46253f
C25936 a_5205_44484# a_5883_43914# 0.003713f
C25937 a_5111_44636# a_8975_43940# 5.4e-19
C25938 a_3232_43370# a_10334_44484# 0.040395f
C25939 a_6171_45002# a_10157_44484# 4.27e-20
C25940 a_8191_45002# a_5343_44458# 1.33e-19
C25941 a_6709_45028# a_6298_44484# 0.006607f
C25942 a_7871_42858# a_n443_42852# 0.013386f
C25943 a_12089_42308# a_n357_42282# 0.027195f
C25944 a_16405_45348# a_10227_46804# 5.83e-20
C25945 a_18184_42460# a_11599_46634# 0.018223f
C25946 a_17719_45144# a_16327_47482# 2.77e-19
C25947 a_21101_45002# a_12861_44030# 1.67e-20
C25948 C9_P_btm VDD 0.345685f
C25949 a_949_44458# a_584_46384# 0.011926f
C25950 a_5883_43914# a_n971_45724# 0.027317f
C25951 a_n1699_44726# a_n1151_42308# 2.55e-19
C25952 a_4099_45572# a_n2293_46098# 0.00692f
C25953 a_16333_45814# a_3090_45724# 0.007872f
C25954 a_15903_45785# a_15368_46634# 6.84e-19
C25955 a_11823_42460# a_765_45546# 2.37e-20
C25956 a_15599_45572# a_15559_46634# 6.99e-21
C25957 a_14180_45002# a_5807_45002# 0.005192f
C25958 a_13777_45326# a_13661_43548# 0.001317f
C25959 a_626_44172# a_768_44030# 0.186913f
C25960 a_15765_45572# a_14976_45028# 1.08e-20
C25961 a_2437_43646# a_6540_46812# 5.76e-21
C25962 a_5691_45260# a_n743_46660# 3.07e-20
C25963 a_6171_45002# a_n1925_46634# 0.005306f
C25964 a_3357_43084# a_5167_46660# 2.88e-19
C25965 a_5342_30871# a_15597_42852# 0.003587f
C25966 a_4190_30871# a_5934_30871# 0.020923f
C25967 a_4361_42308# a_5932_42308# 0.072603f
C25968 a_743_42282# a_6123_31319# 0.018532f
C25969 a_1847_42826# a_n784_42308# 0.001475f
C25970 a_16547_43609# a_14113_42308# 6.85e-19
C25971 a_15781_43660# a_15890_42674# 2.11e-20
C25972 a_n1925_42282# DATA[2] 9.03e-20
C25973 a_6151_47436# a_768_44030# 0.096889f
C25974 a_4915_47217# a_13569_47204# 4.96e-19
C25975 a_6575_47204# a_9804_47204# 3.95e-20
C25976 a_11459_47204# a_n881_46662# 0.0707f
C25977 a_9067_47204# a_8128_46384# 4.87e-19
C25978 a_n2109_47186# a_171_46873# 7.56e-20
C25979 a_n815_47178# a_n1925_46634# 9.48e-20
C25980 a_n1741_47186# a_n2438_43548# 6.62e-19
C25981 a_n785_47204# a_n2661_46634# 0.006981f
C25982 a_n746_45260# a_n2293_46634# 0.048005f
C25983 a_20990_47178# a_4883_46098# 2.39e-20
C25984 a_19787_47423# a_12465_44636# 2.07e-19
C25985 a_18479_47436# a_11453_44696# 0.018416f
C25986 a_n4209_38502# VDD 0.811731f
C25987 a_11963_45334# a_11341_43940# 1.74e-20
C25988 a_7640_43914# a_5891_43370# 0.011186f
C25989 a_12607_44458# a_12553_44484# 6.75e-20
C25990 a_14537_43396# a_15493_43396# 5.06e-19
C25991 a_21359_45002# a_19237_31679# 8.84e-20
C25992 a_n2012_44484# a_n2661_42834# 0.001285f
C25993 a_18907_42674# a_n357_42282# 3.94e-20
C25994 a_22775_42308# a_20692_30879# 5.45e-21
C25995 a_17668_45572# VDD 9.68e-19
C25996 a_22223_42860# RST_Z 5.92e-20
C25997 a_14537_43396# a_3483_46348# 0.087339f
C25998 a_626_44172# a_1176_45822# 1.95e-19
C25999 a_5365_45348# a_n2293_46098# 4.09e-19
C26000 a_15004_44636# a_6755_46942# 5.2e-19
C26001 a_19615_44636# a_19321_45002# 0.035767f
C26002 a_20362_44736# a_13747_46662# 5.6e-20
C26003 a_n2661_43922# a_1799_45572# 3.03e-20
C26004 a_17478_45572# a_13259_45724# 0.048668f
C26005 a_16680_45572# a_16375_45002# 5.99e-20
C26006 a_18596_45572# a_8049_45260# 0.001924f
C26007 a_n2661_45010# a_n2956_39304# 1.05e-20
C26008 a_3232_43370# a_9290_44172# 0.087744f
C26009 a_6171_45002# a_10355_46116# 3.21e-22
C26010 a_8191_45002# a_8349_46414# 5.23e-21
C26011 a_413_45260# a_15682_46116# 3.05e-20
C26012 a_8953_45002# a_8016_46348# 0.016464f
C26013 a_6709_45028# a_5937_45572# 0.629301f
C26014 a_7229_43940# a_8953_45546# 7.78e-21
C26015 a_7705_45326# a_8199_44636# 8.08e-19
C26016 a_1755_42282# a_5742_30871# 3.99e-20
C26017 a_5932_42308# a_6761_42308# 0.001757f
C26018 a_5755_42308# a_6123_31319# 2.22e-20
C26019 a_1606_42308# a_11551_42558# 1.77e-20
C26020 a_14097_32519# a_4958_30871# 0.030871f
C26021 a_22400_42852# a_17303_42282# 0.004332f
C26022 a_2982_43646# CAL_N 0.181412f
C26023 CAL_P a_19864_35138# 0.003641f
C26024 a_n1386_35608# a_n1532_35090# 0.045378f
C26025 a_2063_45854# a_5204_45822# 0.174206f
C26026 a_n1741_47186# a_11133_46155# 1.23e-20
C26027 a_n237_47217# a_8953_45546# 0.090521f
C26028 a_5807_45002# a_15009_46634# 0.006271f
C26029 a_13747_46662# a_13607_46688# 0.168294f
C26030 a_3877_44458# a_5167_46660# 0.032716f
C26031 a_4646_46812# a_5385_46902# 0.042888f
C26032 a_4651_46660# a_4817_46660# 0.57393f
C26033 a_12549_44172# a_19692_46634# 0.491923f
C26034 a_n1925_46634# a_6903_46660# 7.98e-20
C26035 a_n1151_42308# a_4185_45028# 7.97e-20
C26036 a_n443_46116# a_167_45260# 0.794635f
C26037 a_3785_47178# a_3483_46348# 2.62e-20
C26038 a_4883_46098# a_20273_46660# 2.98e-19
C26039 a_13507_46334# a_20623_46660# 0.005302f
C26040 a_21177_47436# a_21363_46634# 2.52e-20
C26041 a_11599_46634# a_12741_44636# 0.183316f
C26042 a_11453_44696# a_17829_46910# 0.013408f
C26043 a_12465_44636# a_20107_46660# 2.35e-20
C26044 a_n2017_45002# a_12895_43230# 1.47e-19
C26045 a_n1059_45260# a_13113_42826# 0.002702f
C26046 a_n913_45002# a_12545_42858# 0.548984f
C26047 a_3537_45260# a_5111_42852# 0.123919f
C26048 a_n984_44318# a_n822_43940# 0.006453f
C26049 a_175_44278# a_261_44278# 0.006584f
C26050 a_19279_43940# a_18451_43940# 3.9e-19
C26051 a_18579_44172# a_17973_43940# 5.34e-19
C26052 a_5244_44056# a_5495_43940# 0.107037f
C26053 a_11967_42832# a_20935_43940# 9.08e-20
C26054 a_20640_44752# a_19862_44208# 0.001675f
C26055 a_20159_44458# a_20365_43914# 0.003347f
C26056 a_20362_44736# a_20269_44172# 2.05e-20
C26057 a_18374_44850# a_n97_42460# 1.3e-21
C26058 a_17970_44736# VDD 0.27753f
C26059 a_n4064_39616# C7_P_btm 1.47e-19
C26060 a_n3420_39616# C5_P_btm 4.27e-20
C26061 a_n3565_39304# EN_VIN_BSTR_P 2.04e-19
C26062 a_9313_44734# a_10809_44734# 0.001335f
C26063 a_16664_43396# a_16327_47482# 2.45e-19
C26064 a_n2157_42858# a_n1151_42308# 5.83e-19
C26065 a_15682_43940# a_15227_44166# 0.072383f
C26066 a_15493_43396# a_3090_45724# 0.134629f
C26067 a_2813_43396# a_768_44030# 4.65e-19
C26068 a_n1557_42282# a_n2312_38680# 1.6e-20
C26069 a_1891_43646# a_n2293_46634# 8.05e-20
C26070 a_10057_43914# a_10586_45546# 1.37e-19
C26071 a_491_47026# VDD 0.132552f
C26072 a_n4064_40160# a_n4251_38528# 0.001069f
C26073 a_n4209_39304# a_n3607_39392# 0.002352f
C26074 a_n4334_39392# a_n4251_39392# 0.007692f
C26075 a_n3420_39616# a_n3420_38528# 0.049464f
C26076 a_n4064_39616# a_n3565_38502# 0.02802f
C26077 a_n3565_39590# a_n4064_38528# 0.031177f
C26078 a_n4315_30879# a_n4209_38216# 0.053149f
C26079 a_1343_38525# a_1239_39043# 0.01446f
C26080 a_n3565_39304# a_n2302_39072# 0.066757f
C26081 a_n3690_39392# a_n4064_39072# 0.085872f
C26082 a_n3420_39072# a_n2946_39072# 0.238708f
C26083 a_5742_30871# C2_N_btm 0.030783f
C26084 a_n3674_38216# a_n2946_37984# 4.03e-21
C26085 a_3090_45724# a_3483_46348# 0.060766f
C26086 a_20273_46660# a_21188_46660# 0.118759f
C26087 a_20107_46660# a_20528_46660# 0.083408f
C26088 a_13747_46662# a_16375_45002# 0.021583f
C26089 a_5807_45002# a_19431_46494# 1.86e-20
C26090 a_n881_46662# a_n863_45724# 0.023273f
C26091 a_6755_46942# a_13759_46122# 9.15e-19
C26092 a_8270_45546# a_8953_45546# 1.06716f
C26093 a_n1613_43370# a_n452_45724# 6.53e-20
C26094 a_11453_44696# a_n443_42852# 4.16e-20
C26095 a_9028_43914# a_8685_43396# 1.97e-20
C26096 a_1241_43940# a_1209_43370# 3.49e-19
C26097 a_20512_43084# a_4190_30871# 0.006642f
C26098 a_n2293_43922# a_10083_42826# 2.45e-20
C26099 a_9313_44734# a_13460_43230# 0.004332f
C26100 a_375_42282# a_5934_30871# 1.48e-20
C26101 a_n2293_42834# a_1755_42282# 1.34e-19
C26102 a_3422_30871# a_13467_32519# 0.421402f
C26103 en_comp a_17531_42308# 1.87e-20
C26104 a_n1059_45260# a_18214_42558# 0.020063f
C26105 a_n913_45002# a_19332_42282# 2.77e-19
C26106 a_3353_43940# VDD 0.005542f
C26107 a_9049_44484# a_3232_43370# 0.17048f
C26108 a_7230_45938# a_7276_45260# 4.28e-19
C26109 a_7499_43078# a_6171_45002# 0.029896f
C26110 a_16147_45260# a_18341_45572# 0.001545f
C26111 a_18175_45572# a_18479_45785# 0.280208f
C26112 a_6197_43396# a_4185_45028# 7.89e-21
C26113 a_18525_43370# a_17339_46660# 0.060382f
C26114 a_21855_43396# a_19692_46634# 0.016876f
C26115 a_n97_42460# a_17715_44484# 8.03e-20
C26116 a_2982_43646# a_8199_44636# 3.15e-19
C26117 a_n2472_42282# a_n2312_40392# 4.5e-20
C26118 a_n3674_38680# a_n2312_39304# 0.023326f
C26119 VDAC_P C10_P_btm 0.883474p
C26120 a_14840_46494# VDD 0.275785f
C26121 a_2711_45572# a_4915_47217# 0.265557f
C26122 a_6667_45809# a_n1151_42308# 9.3e-20
C26123 a_8162_45546# a_n971_45724# 0.015463f
C26124 a_3175_45822# a_n443_46116# 0.002277f
C26125 a_n2293_46098# a_n452_45724# 0.007729f
C26126 a_n1853_46287# a_n1079_45724# 0.02186f
C26127 a_n901_46420# a_n2661_45546# 1.05e-19
C26128 a_n1991_46122# a_n2293_45546# 1.19e-19
C26129 a_n4209_38216# a_n3420_37440# 0.035706f
C26130 a_n3565_38216# a_n3565_37414# 0.046412f
C26131 a_9823_46155# a_10037_46155# 0.005572f
C26132 a_11133_46155# a_10586_45546# 0.006738f
C26133 a_13759_46122# a_8049_45260# 0.002564f
C26134 a_1467_44172# a_1606_42308# 2.54e-20
C26135 a_n1557_42282# a_421_43172# 3.1e-19
C26136 a_3080_42308# a_1847_42826# 2.31e-19
C26137 a_15681_43442# a_16409_43396# 3.1e-20
C26138 a_10341_43396# a_16664_43396# 0.005311f
C26139 a_15095_43370# a_15125_43396# 0.007578f
C26140 a_14955_43396# a_15037_43396# 0.005781f
C26141 a_n4318_39768# a_n3674_38216# 0.023361f
C26142 a_5891_43370# a_7174_31319# 9.47e-21
C26143 a_n97_42460# a_10083_42826# 6.2e-20
C26144 a_15781_43660# a_16547_43609# 5.24e-19
C26145 a_14673_44172# a_14113_42308# 2.36e-21
C26146 a_13661_43548# START 0.012406f
C26147 a_13747_46662# RST_Z 0.001276f
C26148 a_8605_42826# VDD 0.204898f
C26149 a_11525_45546# a_11541_44484# 2.97e-20
C26150 a_2232_45348# a_2304_45348# 0.003395f
C26151 a_10306_45572# a_5891_43370# 2.85e-21
C26152 a_13249_42308# a_13213_44734# 1.19e-20
C26153 a_6431_45366# a_n2661_43370# 0.009143f
C26154 a_21513_45002# a_18114_32519# 9.32e-20
C26155 en_comp a_18184_42460# 2.88e-20
C26156 a_7229_43940# a_7735_45067# 0.005614f
C26157 a_8191_45002# a_8560_45348# 0.03364f
C26158 a_6709_45028# a_7418_45067# 0.001659f
C26159 a_6171_45002# a_11915_45394# 7.98e-19
C26160 a_n2017_45002# a_11827_44484# 2.08e-20
C26161 a_22400_42852# a_20820_30879# 1.3e-19
C26162 a_20256_42852# a_20202_43084# 0.001339f
C26163 a_17324_43396# a_n443_42852# 1.63e-21
C26164 a_13678_32519# a_20205_31679# 0.051502f
C26165 a_6472_45840# a_3090_45724# 1.07e-21
C26166 a_11652_45724# a_6755_46942# 1.83e-20
C26167 a_3357_43084# a_12549_44172# 0.001325f
C26168 a_21363_45546# a_13747_46662# 0.001465f
C26169 a_2437_43646# a_16119_47582# 0.001405f
C26170 a_n2293_45010# a_n881_46662# 9.84e-21
C26171 a_5147_45002# a_4883_46098# 5.63e-20
C26172 a_13556_45296# a_11599_46634# 5.22e-21
C26173 a_5365_45348# a_4791_45118# 0.001047f
C26174 a_2982_43646# a_13070_42354# 7.37e-20
C26175 a_4520_42826# a_4743_43172# 0.011458f
C26176 a_16104_42674# VDD 0.134357f
C26177 a_6851_47204# a_7227_47204# 0.241208f
C26178 a_6545_47178# a_6575_47204# 0.11927f
C26179 a_6151_47436# a_9067_47204# 3.94e-19
C26180 a_4915_47217# a_9313_45822# 0.366722f
C26181 a_6491_46660# a_7903_47542# 5.79e-21
C26182 a_n2109_47186# a_4883_46098# 0.029241f
C26183 a_n1741_47186# a_13507_46334# 8.99e-20
C26184 a_4700_47436# a_n1435_47204# 2.1e-19
C26185 a_n1059_45260# a_n2661_42282# 0.028862f
C26186 a_3537_45260# a_7542_44172# 1.57e-19
C26187 a_3232_43370# a_3905_42865# 0.027169f
C26188 a_5147_45002# a_5663_43940# 0.019985f
C26189 a_5111_44636# a_5495_43940# 0.037006f
C26190 a_21188_45572# a_19862_44208# 1.49e-19
C26191 a_n2661_44458# a_n310_44811# 3.72e-19
C26192 a_n1699_44726# a_n1821_44484# 3.16e-19
C26193 a_10334_44484# a_8975_43940# 0.044798f
C26194 a_n2129_44697# a_n356_44636# 0.009952f
C26195 a_n2433_44484# a_n23_44458# 2.38e-21
C26196 a_10440_44484# a_10057_43914# 0.026774f
C26197 a_1184_42692# a_n443_42852# 0.003744f
C26198 a_5267_42460# a_n357_42282# 1.81e-20
C26199 a_3823_42558# a_n755_45592# 0.001851f
C26200 a_13163_45724# VDD 0.322298f
C26201 a_13467_32519# VREF_GND 0.048151f
C26202 a_11652_45724# a_8049_45260# 0.002134f
C26203 a_10180_45724# a_10586_45546# 7.02e-19
C26204 a_15037_45618# a_10809_44734# 4.19e-21
C26205 a_17478_45572# a_18189_46348# 0.002791f
C26206 a_12649_45572# a_2324_44458# 4.41e-19
C26207 a_16241_44484# a_10227_46804# 4.52e-20
C26208 a_18588_44850# a_16327_47482# 0.012252f
C26209 a_17517_44484# a_18597_46090# 0.021693f
C26210 a_20766_44850# a_12861_44030# 5.26e-19
C26211 a_175_44278# a_584_46384# 0.001131f
C26212 a_n1761_44111# a_n1151_42308# 0.642214f
C26213 a_2437_43646# a_1823_45246# 0.324477f
C26214 a_14537_43396# a_14513_46634# 1.12e-21
C26215 a_13348_45260# a_13059_46348# 0.010157f
C26216 a_10057_43914# a_n743_46660# 2.57e-20
C26217 a_n2661_45010# a_n1991_46122# 2.05e-19
C26218 a_n2293_45010# a_n2157_46122# 1.83e-20
C26219 a_n4318_37592# a_n1630_35242# 0.847279f
C26220 a_n3674_39304# a_n4334_38528# 6.7e-20
C26221 a_n4318_38680# a_n4209_38502# 0.105064f
C26222 a_n473_42460# a_n784_42308# 0.020033f
C26223 a_n1329_42308# a_n3674_37592# 0.005224f
C26224 a_22223_42860# a_17303_42282# 4.73e-19
C26225 a_17595_43084# a_7174_31319# 2.85e-21
C26226 a_n2661_46634# a_2107_46812# 0.00917f
C26227 a_n1021_46688# a_n133_46660# 1.36e-19
C26228 a_n1925_46634# a_171_46873# 0.027689f
C26229 a_n743_46660# a_n2438_43548# 0.426835f
C26230 a_n1613_43370# a_5275_47026# 0.039193f
C26231 a_11599_46634# a_13607_46688# 3.8e-19
C26232 a_12861_44030# a_14976_45028# 0.007077f
C26233 a_13717_47436# a_15368_46634# 3.91e-20
C26234 a_n785_47204# a_765_45546# 1.18e-19
C26235 a_18248_44752# a_15493_43940# 8.91e-20
C26236 a_18443_44721# a_11341_43940# 2.01e-20
C26237 a_3422_30871# a_22315_44484# 0.19914f
C26238 a_9482_43914# a_14205_43396# 1.91e-22
C26239 a_4223_44672# a_3737_43940# 1.52e-19
C26240 a_19279_43940# a_19237_31679# 5.63e-21
C26241 a_5891_43370# a_10729_43914# 0.001943f
C26242 a_7499_43078# a_8292_43218# 7.98e-20
C26243 a_11827_44484# a_21845_43940# 1.08e-19
C26244 a_n2661_42834# a_1241_44260# 3.84e-19
C26245 a_n2293_42834# a_n1243_43396# 1.39e-19
C26246 a_n1059_45260# a_16823_43084# 0.318918f
C26247 a_19479_31679# a_13678_32519# 0.051236f
C26248 a_19963_31679# a_13467_32519# 0.051345f
C26249 a_n3607_38304# VDD 2.79e-20
C26250 a_6123_31319# VIN_P 0.01057f
C26251 a_5742_30871# C8_P_btm 0.003514f
C26252 a_n2661_42834# a_11415_45002# 3.35e-20
C26253 a_9895_44260# a_2107_46812# 6.01e-19
C26254 a_18533_44260# a_12549_44172# 3.67e-19
C26255 a_1307_43914# a_n863_45724# 0.050349f
C26256 a_14537_43396# a_n357_42282# 7.25e-21
C26257 a_375_42282# a_n2293_45546# 0.104283f
C26258 a_1145_45348# a_n2661_45546# 1.22e-19
C26259 a_8975_43940# a_9290_44172# 0.114958f
C26260 a_4223_44672# a_2324_44458# 0.56408f
C26261 a_19511_42282# a_21421_42336# 8.32e-19
C26262 a_n2312_39304# VDD 0.587668f
C26263 a_14097_32519# C7_N_btm 7.66e-20
C26264 a_3699_46634# a_3483_46348# 3.01e-19
C26265 a_14976_45028# a_14180_46812# 1.12e-19
C26266 a_12991_46634# a_13059_46348# 0.003295f
C26267 a_13607_46688# a_13693_46688# 0.006584f
C26268 a_14084_46812# a_14543_46987# 6.64e-19
C26269 a_15559_46634# a_13885_46660# 8.64e-20
C26270 a_3090_45724# a_14513_46634# 6.29e-19
C26271 a_15368_46634# a_14035_46660# 5.28e-22
C26272 a_n881_46662# a_1431_46436# 5.43e-19
C26273 a_n743_46660# a_11133_46155# 0.006423f
C26274 a_13747_46662# a_18985_46122# 0.035795f
C26275 a_2107_46812# a_8199_44636# 0.022874f
C26276 a_5807_45002# a_19335_46494# 0.005114f
C26277 a_13759_47204# a_6945_45028# 7.25e-19
C26278 a_n237_47217# a_1609_45822# 0.141985f
C26279 a_n1151_42308# a_997_45618# 9.32e-22
C26280 a_n443_46116# a_n863_45724# 0.055503f
C26281 a_584_46384# a_n356_45724# 0.00412f
C26282 a_2063_45854# a_3503_45724# 0.002656f
C26283 a_2905_45572# a_2957_45546# 0.137248f
C26284 a_12861_44030# a_18051_46116# 2.97e-19
C26285 a_11599_46634# a_16375_45002# 0.407484f
C26286 a_5534_30871# a_8530_39574# 1.75e-19
C26287 a_n2017_45002# a_3581_42558# 0.001947f
C26288 a_n913_45002# a_5379_42460# 0.179494f
C26289 a_5111_44636# a_n784_42308# 2.01e-20
C26290 a_13829_44260# a_14021_43940# 1.97e-19
C26291 a_18184_42460# a_22165_42308# 0.026631f
C26292 a_11827_44484# a_19164_43230# 1.08e-21
C26293 a_11691_44458# a_18249_42858# 5.39e-21
C26294 a_5343_44458# a_7765_42852# 0.010279f
C26295 a_11967_42832# a_14955_43396# 2.03e-19
C26296 a_1414_42308# a_3626_43646# 0.015112f
C26297 a_2479_44172# a_2896_43646# 0.026857f
C26298 a_4223_44672# a_8387_43230# 4.84e-21
C26299 a_3905_42865# a_4905_42826# 0.404829f
C26300 a_6298_44484# a_7227_42852# 2.52e-20
C26301 a_n1287_44306# VDD 1.78e-19
C26302 a_10193_42453# a_16147_45260# 0.193225f
C26303 a_11823_42460# a_13385_45572# 1.28e-19
C26304 a_7845_44172# a_8049_45260# 7.46e-20
C26305 a_20835_44721# a_n357_42282# 8.73e-21
C26306 a_n2661_42282# a_n1925_42282# 2.27741f
C26307 a_15493_43940# a_2324_44458# 0.061147f
C26308 a_12710_44260# a_10903_43370# 0.001775f
C26309 a_564_42282# a_n2497_47436# 3.52e-21
C26310 a_4361_42308# a_4646_46812# 9.53e-20
C26311 a_10695_43548# a_3090_45724# 0.005861f
C26312 a_1847_42826# a_n2438_43548# 3.92e-21
C26313 a_5342_30871# a_12549_44172# 4.48e-20
C26314 a_16759_43396# a_6755_46942# 5.96e-19
C26315 a_n1991_46122# a_n914_46116# 1.46e-19
C26316 a_3090_45724# a_n357_42282# 0.002409f
C26317 a_16388_46812# a_13259_45724# 0.030634f
C26318 a_9290_44172# a_11387_46155# 0.008277f
C26319 a_6419_46155# a_2324_44458# 2.12e-20
C26320 a_11189_46129# a_11133_46155# 0.203074f
C26321 a_5891_43370# a_5932_42308# 0.001048f
C26322 a_21381_43940# a_4190_30871# 0.023285f
C26323 a_19319_43548# a_19095_43396# 0.006369f
C26324 a_n2293_43922# a_2351_42308# 3.54e-20
C26325 a_n356_44636# a_8791_42308# 2.77e-19
C26326 a_3626_43646# a_12281_43396# 0.001712f
C26327 a_8147_43396# a_8423_43396# 0.00119f
C26328 a_14401_32519# a_21259_43561# 2.5e-19
C26329 a_n97_42460# a_16664_43396# 0.002303f
C26330 SMPL_ON_N a_22609_38406# 9.53e-21
C26331 a_9863_47436# CLK 0.00103f
C26332 a_9313_45822# DATA[5] 0.055804f
C26333 a_11599_46634# RST_Z 2.3e-19
C26334 a_n1435_47204# DATA[2] 0.028258f
C26335 a_18783_43370# VDD 0.289099f
C26336 a_5147_45002# a_3232_43370# 0.253159f
C26337 a_5111_44636# a_5691_45260# 0.130044f
C26338 a_3537_45260# a_5205_44484# 7.92e-19
C26339 a_n2661_45010# a_375_42282# 0.017053f
C26340 a_n2293_45010# a_1307_43914# 0.008547f
C26341 a_9049_44484# a_8975_43940# 0.001423f
C26342 a_10180_45724# a_10440_44484# 8.08e-21
C26343 a_8746_45002# a_10157_44484# 0.003462f
C26344 a_10922_42852# a_4185_45028# 1.72e-20
C26345 a_6761_42308# a_4646_46812# 2.07e-21
C26346 a_17531_42308# a_13661_43548# 1.49e-21
C26347 a_20107_42308# a_12549_44172# 3.8e-21
C26348 a_3457_43396# a_n2661_45546# 0.030099f
C26349 a_7871_42858# a_8199_44636# 1.17e-20
C26350 a_n2216_39866# a_n2312_40392# 5.49e-20
C26351 a_3422_30871# VCM 1.12142f
C26352 a_15037_45618# a_n881_46662# 0.044816f
C26353 a_18175_45572# a_13507_46334# 3.67e-20
C26354 a_19431_45546# a_19386_47436# 8.77e-20
C26355 a_19256_45572# a_18597_46090# 0.001301f
C26356 a_18953_45572# a_16327_47482# 0.002336f
C26357 a_3357_43084# a_6575_47204# 8.41e-19
C26358 a_2437_43646# a_11031_47542# 0.003672f
C26359 a_3537_45260# a_n971_45724# 0.266743f
C26360 a_3065_45002# a_n237_47217# 2.45e-20
C26361 a_3232_43370# a_n2109_47186# 3.24e-19
C26362 a_12427_45724# a_n2661_46634# 4.09e-20
C26363 a_10180_45724# a_n743_46660# 2.31e-19
C26364 a_5649_42852# a_5534_30871# 0.234793f
C26365 a_15493_43396# a_18727_42674# 1.59e-21
C26366 a_14021_43940# a_15486_42560# 6.52e-22
C26367 a_n1557_42282# COMP_P 0.123881f
C26368 a_743_42282# a_18083_42858# 1.7e-19
C26369 a_4361_42308# a_15567_42826# 3.24e-20
C26370 a_4190_30871# a_18249_42858# 0.029356f
C26371 a_1847_42826# a_2075_43172# 0.103349f
C26372 a_1209_43370# a_1067_42314# 4.05e-20
C26373 a_7754_40130# a_3726_37500# 0.021358f
C26374 a_1221_42558# VDD 2.13e-19
C26375 a_n2288_47178# a_n815_47178# 6.95e-21
C26376 a_n2109_47186# a_n1605_47204# 0.041602f
C26377 a_n1920_47178# SMPL_ON_P 0.007059f
C26378 a_22959_45036# a_18114_32519# 0.004401f
C26379 a_1423_45028# a_5891_43370# 0.301629f
C26380 a_13249_42308# a_11341_43940# 0.032308f
C26381 a_22223_45036# a_19721_31679# 2.55e-19
C26382 a_11691_44458# a_19929_45028# 5.24e-19
C26383 a_1307_43914# a_9313_44734# 0.021168f
C26384 a_2437_43646# a_20512_43084# 3.76e-21
C26385 a_6123_31319# a_n2956_38680# 3.8e-21
C26386 a_14113_42308# a_10903_43370# 1.69e-20
C26387 a_17531_42308# a_4185_45028# 6.87e-20
C26388 a_22521_40599# SMPL_ON_N 1.14e-19
C26389 a_8697_45822# a_3483_46348# 0.033264f
C26390 a_16855_45546# a_12741_44636# 7.31e-20
C26391 a_15861_45028# a_11415_45002# 0.041647f
C26392 a_2809_45028# a_2609_46660# 5.53e-21
C26393 a_18587_45118# a_19321_45002# 2.02e-19
C26394 a_19778_44110# a_13747_46662# 0.670692f
C26395 a_18184_42460# a_13661_43548# 0.031622f
C26396 a_2903_45348# a_3877_44458# 2.68e-20
C26397 a_413_45260# a_11735_46660# 5.06e-20
C26398 a_7276_45260# a_6755_46942# 4.58e-22
C26399 a_8746_45002# a_10355_46116# 0.002156f
C26400 a_10193_42453# a_9290_44172# 1.23123f
C26401 a_7499_43078# a_10903_43370# 0.888628f
C26402 a_2711_45572# a_10809_44734# 0.037787f
C26403 a_10180_45724# a_11189_46129# 4.36e-20
C26404 a_18443_44721# a_16327_47482# 0.1665f
C26405 a_n2661_43922# a_2063_45854# 0.033229f
C26406 a_10083_42826# a_10533_42308# 0.003061f
C26407 a_5649_42852# a_19647_42308# 1.31e-19
C26408 a_4361_42308# a_20712_42282# 0.013294f
C26409 a_13678_32519# a_13258_32519# 0.055554f
C26410 a_18504_43218# a_18695_43230# 4.61e-19
C26411 a_13467_32519# a_7174_31319# 6e-19
C26412 a_310_45028# DATA[0] 1.08e-20
C26413 a_n881_46662# a_13569_47204# 0.001167f
C26414 a_n1151_42308# a_5257_43370# 0.058425f
C26415 a_n971_45724# a_6969_46634# 0.235123f
C26416 a_2063_45854# a_7927_46660# 0.004156f
C26417 a_n443_46116# a_5072_46660# 3.53e-19
C26418 a_4791_45118# a_5275_47026# 0.004467f
C26419 a_n237_47217# a_10249_46116# 2.78e-20
C26420 a_6491_46660# a_4817_46660# 1.23e-19
C26421 a_5815_47464# a_5907_46634# 0.004583f
C26422 a_4915_47217# a_6540_46812# 1.17e-20
C26423 a_6575_47204# a_3877_44458# 6.28e-20
C26424 a_13507_46334# a_n743_46660# 0.024694f
C26425 a_4883_46098# a_n1925_46634# 0.030451f
C26426 a_11453_44696# a_n2661_46634# 0.032889f
C26427 a_n2312_40392# a_n2840_46634# 3.22e-21
C26428 C0_N_btm VDD 1.02806f
C26429 a_n913_45002# a_7287_43370# 9.35e-21
C26430 a_3232_43370# a_4093_43548# 0.091441f
C26431 a_5147_45002# a_4905_42826# 3.8e-19
C26432 a_2382_45260# a_2982_43646# 0.468592f
C26433 a_n2661_42834# a_11967_42832# 2.11e-20
C26434 a_19778_44110# a_20269_44172# 1.25e-19
C26435 a_9313_44734# a_18579_44172# 3.89e-19
C26436 a_18494_42460# a_19478_44306# 6.46e-21
C26437 a_5883_43914# a_7281_43914# 0.029594f
C26438 a_11827_44484# a_18079_43940# 0.002983f
C26439 a_11691_44458# a_14955_43940# 0.00153f
C26440 a_8103_44636# a_7845_44172# 2.71e-19
C26441 a_18184_42460# a_19862_44208# 0.028217f
C26442 a_16922_45042# a_15493_43940# 0.019907f
C26443 a_17613_45144# a_11341_43940# 7.11e-21
C26444 a_8953_45002# VDD 1.24336f
C26445 a_8191_45002# a_8034_45724# 1.83e-20
C26446 a_7276_45260# a_8049_45260# 5.67e-19
C26447 a_2437_43646# a_n2293_45546# 0.031092f
C26448 a_3357_43084# a_n2661_45546# 0.045914f
C26449 a_n2293_42834# a_2324_44458# 0.168086f
C26450 a_n97_42460# a_584_46384# 0.526796f
C26451 a_n1557_42282# a_n2497_47436# 7.44e-20
C26452 a_18184_42460# a_4185_45028# 0.006813f
C26453 a_9028_43914# a_768_44030# 0.113848f
C26454 a_7542_44172# a_n2293_46634# 5.45e-20
C26455 a_17517_44484# a_6755_46942# 8.4e-20
C26456 a_1209_47178# VDD 0.38145f
C26457 a_n3674_37592# a_n4334_39392# 6.37e-20
C26458 a_6123_31319# a_13258_32519# 0.00105f
C26459 a_14113_42308# a_15959_42545# 0.036113f
C26460 a_15486_42560# a_15764_42576# 0.118759f
C26461 a_15051_42282# a_15803_42450# 0.043619f
C26462 a_4190_30871# a_8530_39574# 1.25e-19
C26463 VREF_GND VCM 2.79113f
C26464 a_13661_43548# a_12741_44636# 0.13948f
C26465 a_19321_45002# a_11415_45002# 0.065361f
C26466 a_2107_46812# a_765_45546# 0.001701f
C26467 a_10554_47026# a_10384_47026# 2.6e-19
C26468 a_10428_46928# a_10768_47026# 0.027606f
C26469 a_6755_46942# a_8189_46660# 0.002345f
C26470 a_10249_46116# a_8270_45546# 1.06e-19
C26471 a_n881_46662# a_2202_46116# 0.051959f
C26472 a_n1613_43370# a_167_45260# 1.05e-19
C26473 a_11453_44696# a_8199_44636# 3.39e-19
C26474 a_4883_46098# a_10355_46116# 0.23167f
C26475 a_11599_46634# a_18985_46122# 0.570252f
C26476 a_16327_47482# a_17583_46090# 1.09e-19
C26477 a_10227_46804# a_14275_46494# 0.18614f
C26478 a_16023_47582# a_15682_46116# 0.001021f
C26479 a_13717_47436# a_20708_46348# 5.9e-22
C26480 a_13381_47204# a_6945_45028# 0.006113f
C26481 a_12861_44030# a_19900_46494# 4.29e-21
C26482 a_4700_47436# a_526_44458# 1.71e-21
C26483 a_4007_47204# a_n1925_42282# 8.11e-20
C26484 a_n237_47217# a_8781_46436# 5.45e-19
C26485 a_n1741_47186# a_10586_45546# 3.67e-20
C26486 a_10729_43914# a_10807_43548# 0.238591f
C26487 a_9313_44734# a_9396_43370# 4.33e-20
C26488 a_18579_44172# a_20974_43370# 2.18e-20
C26489 a_11823_42460# a_12563_42308# 0.039858f
C26490 a_10193_42453# a_15051_42282# 5.96e-19
C26491 a_20193_45348# a_13678_32519# 0.055785f
C26492 a_2127_44172# a_2253_43940# 0.143754f
C26493 a_895_43940# a_1241_43940# 0.054548f
C26494 a_2479_44172# a_1443_43940# 8.09e-20
C26495 a_n2293_42834# a_8387_43230# 4.23e-19
C26496 a_n1059_45260# a_11136_42852# 0.004379f
C26497 a_3537_45260# a_3863_42891# 5.22e-20
C26498 a_2711_45572# a_8120_45572# 7.29e-19
C26499 a_6472_45840# a_8697_45822# 8.93e-21
C26500 a_6598_45938# a_6905_45572# 3.69e-19
C26501 a_6667_45809# a_6977_45572# 0.013793f
C26502 a_10053_45546# a_10180_45724# 0.144403f
C26503 a_9049_44484# a_10193_42453# 6.5e-20
C26504 a_7499_43078# a_8746_45002# 0.153858f
C26505 a_19862_44208# a_12741_44636# 8.5e-21
C26506 a_743_42282# a_12549_44172# 0.119701f
C26507 a_6197_43396# a_5257_43370# 0.001674f
C26508 a_7274_43762# a_4646_46812# 2.49e-19
C26509 a_15743_43084# a_21588_30879# 3.87e-20
C26510 a_n356_44636# a_n357_42282# 0.308599f
C26511 a_n23_44458# a_310_45028# 0.002647f
C26512 a_n4318_38680# a_n2312_39304# 0.0235f
C26513 a_19963_31679# VCM 0.035453f
C26514 en_comp RST_Z 4.34313f
C26515 a_20447_31679# VREF 0.059621f
C26516 a_10768_47026# VDD 0.132317f
C26517 a_1606_42308# VDAC_N 0.010938f
C26518 a_5742_30871# a_2113_38308# 6.13e-20
C26519 a_n2293_46098# a_167_45260# 0.086636f
C26520 a_n1076_46494# a_472_46348# 0.001137f
C26521 a_12741_44636# a_4185_45028# 1.08e-20
C26522 a_948_46660# a_n443_42852# 2.59e-20
C26523 a_3877_44458# a_n2661_45546# 0.026409f
C26524 a_2959_46660# a_n755_45592# 2.79e-21
C26525 a_2443_46660# a_2957_45546# 3.36e-19
C26526 a_1123_46634# a_1609_45822# 8.43e-20
C26527 a_n743_46660# a_603_45572# 1.47e-19
C26528 a_1799_45572# a_3316_45546# 2.21e-21
C26529 a_8189_46660# a_8049_45260# 2.51e-20
C26530 a_8270_45546# a_8781_46436# 2.13e-19
C26531 a_16388_46812# a_18189_46348# 0.0042f
C26532 a_12513_46660# a_10809_44734# 5.68e-19
C26533 a_n2956_37592# a_n2216_38778# 1.2e-19
C26534 a_n97_42460# a_n144_43396# 1.59e-19
C26535 a_3905_42865# a_2905_42968# 2.41e-19
C26536 a_4093_43548# a_4905_42826# 5.66e-20
C26537 a_1568_43370# a_n1557_42282# 3.82e-20
C26538 a_15493_43396# a_17486_43762# 3.67e-19
C26539 a_1049_43396# a_1427_43646# 0.010711f
C26540 a_3422_30871# a_16795_42852# 2.85e-21
C26541 a_3600_43914# a_3681_42891# 2.17e-20
C26542 a_19279_43940# a_19987_42826# 1.18e-19
C26543 a_18579_44172# a_18599_43230# 1.99e-20
C26544 a_2998_44172# a_3935_42891# 3.35e-21
C26545 a_11341_43940# a_19700_43370# 4.45e-20
C26546 a_15493_43940# a_15743_43084# 0.206331f
C26547 a_4235_43370# a_3080_42308# 0.098951f
C26548 a_12429_44172# a_743_42282# 3.38e-21
C26549 a_20679_44626# a_21195_42852# 7.08e-20
C26550 w_11334_34010# EN_VIN_BSTR_N 3.99277f
C26551 SMPL_ON_P a_n1838_35608# 0.399535f
C26552 a_3626_43646# VDD 0.340378f
C26553 a_15037_45618# a_1307_43914# 1.49e-21
C26554 a_15765_45572# a_14537_43396# 3.49e-19
C26555 a_15599_45572# a_15415_45028# 5.19e-19
C26556 a_8696_44636# a_13348_45260# 1.38e-20
C26557 a_11322_45546# a_11361_45348# 9.02e-20
C26558 a_10490_45724# a_n2661_43370# 7.79e-21
C26559 a_19963_31679# a_22959_45572# 0.020087f
C26560 a_2437_43646# a_n2661_45010# 0.15182f
C26561 a_22591_45572# a_20447_31679# 7.75e-19
C26562 a_8147_43396# a_526_44458# 2.13e-19
C26563 a_1443_43940# a_n443_42852# 3.91e-20
C26564 a_n3674_37592# a_n2312_38680# 0.026177f
C26565 a_18249_42858# a_15227_44166# 2.56e-20
C26566 a_11601_46155# VDD 0.001563f
C26567 a_2711_45572# a_n881_46662# 0.170524f
C26568 a_7499_43078# a_4883_46098# 8.38e-19
C26569 a_11823_42460# a_10227_46804# 0.428745f
C26570 a_11682_45822# a_11459_47204# 6.52e-21
C26571 a_14033_45822# a_4915_47217# 0.002034f
C26572 a_n2956_38680# a_n2472_45546# 4.48e-19
C26573 a_n2956_39304# a_n2956_38216# 0.05012f
C26574 a_21487_43396# a_13467_32519# 0.152042f
C26575 a_9885_43646# a_10083_42826# 1.33e-19
C26576 a_8685_43396# a_5534_30871# 4.59e-19
C26577 a_9145_43396# a_12545_42858# 6.25e-19
C26578 a_20512_43084# a_19511_42282# 7.2e-20
C26579 a_3422_30871# a_21335_42336# 0.002526f
C26580 a_4190_30871# a_5649_42852# 0.434284f
C26581 a_4905_42826# a_5457_43172# 2.02e-20
C26582 VDAC_N C1_N_btm 1.7375f
C26583 a_7705_45326# a_5343_44458# 2.71e-19
C26584 a_6431_45366# a_5883_43914# 1.65e-19
C26585 a_5111_44636# a_10057_43914# 0.002052f
C26586 a_3232_43370# a_10157_44484# 0.049345f
C26587 a_7229_43940# a_6298_44484# 0.028942f
C26588 a_15861_45028# a_11967_42832# 6.28e-20
C26589 a_4921_42308# a_1823_45246# 4.85e-19
C26590 a_7227_42852# a_n443_42852# 0.008558f
C26591 a_12379_42858# a_n357_42282# 0.031137f
C26592 a_n784_42308# a_9290_44172# 1.07e-19
C26593 a_327_44734# a_491_47026# 5.88e-21
C26594 a_2382_45260# a_2107_46812# 5.81e-22
C26595 a_5205_44484# a_n2293_46634# 2.48e-19
C26596 a_3357_43084# a_5385_46902# 0.001502f
C26597 a_13490_45394# a_13507_46334# 1.03e-19
C26598 a_16321_45348# a_10227_46804# 9.56e-20
C26599 a_19778_44110# a_11599_46634# 1.94e-19
C26600 a_17613_45144# a_16327_47482# 7.07e-20
C26601 a_21005_45260# a_12861_44030# 1.13e-21
C26602 C10_P_btm VDD 2.40001f
C26603 a_6298_44484# a_n237_47217# 8.52e-20
C26604 a_8701_44490# a_n971_45724# 8.96e-19
C26605 a_742_44458# a_584_46384# 0.031608f
C26606 a_n2267_44484# a_n1151_42308# 2.66e-19
C26607 a_3175_45822# a_n2293_46098# 0.008709f
C26608 a_15599_45572# a_15368_46634# 0.100853f
C26609 a_15765_45572# a_3090_45724# 0.046838f
C26610 a_15903_45785# a_14976_45028# 1.22e-19
C26611 a_9482_43914# a_13747_46662# 1.7e-20
C26612 a_13777_45326# a_5807_45002# 1.7e-21
C26613 a_13556_45296# a_13661_43548# 0.559682f
C26614 a_5342_30871# a_14853_42852# 5e-21
C26615 a_791_42968# a_n784_42308# 1.7e-19
C26616 a_13467_32519# a_5932_42308# 1.17e-19
C26617 a_743_42282# a_7227_42308# 0.008196f
C26618 a_4361_42308# a_6171_42473# 0.008302f
C26619 a_16243_43396# a_14113_42308# 3.98e-19
C26620 a_15781_43660# a_15959_42545# 2.85e-19
C26621 a_2112_39137# VDD 0.284849f
C26622 a_6151_47436# a_12549_44172# 0.214024f
C26623 a_6575_47204# a_8128_46384# 0.105633f
C26624 a_9313_45822# a_n881_46662# 1.00227f
C26625 a_n971_45724# a_n2293_46634# 0.090091f
C26626 a_n1741_47186# a_n743_46660# 0.017496f
C26627 a_n1151_42308# a_5807_45002# 1.52318f
C26628 a_n2109_47186# a_n133_46660# 2.86e-20
C26629 a_n1920_47178# a_n2438_43548# 1.47e-19
C26630 a_n23_47502# a_n2661_46634# 5.47e-19
C26631 a_n2497_47436# a_33_46660# 6.33e-21
C26632 a_19386_47436# a_12465_44636# 2.39e-19
C26633 a_21177_47436# a_13507_46334# 0.329096f
C26634 a_18143_47464# a_11453_44696# 0.001066f
C26635 a_11787_45002# a_11341_43940# 1.39e-22
C26636 a_16751_45260# a_15682_43940# 3.8e-19
C26637 a_13249_42308# a_10341_43396# 0.040208f
C26638 a_14539_43914# a_15433_44458# 2.67e-20
C26639 a_6109_44484# a_5891_43370# 3.31e-20
C26640 a_15004_44636# a_15463_44811# 6.64e-19
C26641 a_8975_43940# a_12553_44484# 1.95e-20
C26642 a_12607_44458# a_12189_44484# 2.07e-20
C26643 a_7640_43914# a_8375_44464# 5.23e-19
C26644 a_11827_44484# a_17730_32519# 0.009382f
C26645 a_18727_42674# a_n357_42282# 4.23e-20
C26646 a_22775_42308# a_20205_31679# 4.58e-21
C26647 a_22165_42308# RST_Z 4.44e-21
C26648 a_14180_45002# a_3483_46348# 2.73e-20
C26649 a_375_42282# a_1138_42852# 7.22e-21
C26650 a_5105_45348# a_n2293_46098# 2.55e-19
C26651 a_18315_45260# a_16388_46812# 5e-21
C26652 a_11967_42832# a_19321_45002# 0.266816f
C26653 a_5891_43370# a_4646_46812# 0.089437f
C26654 a_20159_44458# a_13747_46662# 1.78e-20
C26655 a_20362_44736# a_13661_43548# 5.77e-20
C26656 a_19789_44512# a_12549_44172# 5e-19
C26657 a_15861_45028# a_13259_45724# 0.16873f
C26658 a_16855_45546# a_16375_45002# 2.09e-19
C26659 a_19256_45572# a_8049_45260# 0.007359f
C26660 a_6171_45002# a_9823_46155# 9.16e-22
C26661 a_8191_45002# a_8016_46348# 3.05e-20
C26662 a_413_45260# a_2324_44458# 0.021366f
C26663 a_7229_43940# a_5937_45572# 0.126047f
C26664 a_1606_42308# a_5742_30871# 3.46204f
C26665 a_4921_42308# a_5934_30871# 3.08e-20
C26666 a_6171_42473# a_6761_42308# 3.88e-19
C26667 a_n784_42308# a_15051_42282# 1.37e-19
C26668 a_18707_42852# a_18727_42674# 2.69e-19
C26669 CAL_P a_19120_35138# 0.00106f
C26670 a_n1838_35608# a_n1532_35090# 4.88e-19
C26671 a_n1741_47186# a_11189_46129# 4.54e-19
C26672 a_n971_45724# a_9625_46129# 2.11e-20
C26673 a_2063_45854# a_5164_46348# 0.022664f
C26674 a_n237_47217# a_5937_45572# 0.08715f
C26675 a_2905_45572# a_4419_46090# 1.32e-19
C26676 a_5807_45002# a_14084_46812# 0.006112f
C26677 a_3877_44458# a_5385_46902# 0.021989f
C26678 a_4646_46812# a_4817_46660# 0.588038f
C26679 a_4651_46660# a_4955_46873# 0.140348f
C26680 a_12549_44172# a_19466_46812# 1.6e-19
C26681 a_13747_46662# a_12816_46660# 2.17e-21
C26682 a_n2661_46634# a_10384_47026# 1.14e-19
C26683 a_n1925_46634# a_6682_46660# 1.03e-19
C26684 a_n443_46116# a_2202_46116# 7.93e-21
C26685 a_16327_47482# a_20885_46660# 8.54e-21
C26686 a_13507_46334# a_20841_46902# 0.005806f
C26687 a_4883_46098# a_20411_46873# 0.012008f
C26688 a_11453_44696# a_765_45546# 0.010973f
C26689 a_n2017_45002# a_13113_42826# 1.01e-19
C26690 a_n1059_45260# a_12545_42858# 0.011705f
C26691 a_3537_45260# a_4520_42826# 0.066648f
C26692 a_n913_45002# a_12089_42308# 0.038293f
C26693 a_5343_44458# a_2982_43646# 1.31e-19
C26694 a_n699_43396# a_3626_43646# 2.23e-19
C26695 a_18579_44172# a_17737_43940# 6.7e-20
C26696 a_3905_42865# a_5495_43940# 1.51e-20
C26697 a_11691_44458# a_8685_43396# 5.46e-21
C26698 a_n2661_44458# a_7287_43370# 3.62e-21
C26699 a_11967_42832# a_20623_43914# 7.1e-20
C26700 a_20159_44458# a_20269_44172# 0.001015f
C26701 a_5244_44056# a_5013_44260# 0.094334f
C26702 a_17767_44458# VDD 0.348803f
C26703 a_n4064_39616# C8_P_btm 0.001799f
C26704 a_n3420_39616# C6_P_btm 5.51e-20
C26705 a_7174_31319# VCM 0.076834f
C26706 a_12189_44484# a_10903_43370# 1.63e-19
C26707 a_14621_43646# a_12465_44636# 1.9e-19
C26708 a_19700_43370# a_16327_47482# 1.38e-19
C26709 a_19328_44172# a_3090_45724# 0.153704f
C26710 a_14955_43940# a_15227_44166# 0.134177f
C26711 a_1427_43646# a_n2293_46634# 2.05e-21
C26712 a_288_46660# VDD 0.079457f
C26713 a_n4064_39616# a_n4334_38528# 8.04e-19
C26714 a_1736_39587# comp_n 0.004824f
C26715 a_n4209_39304# a_n4251_39392# 0.00226f
C26716 a_n4209_39590# a_n2302_38778# 7.57e-20
C26717 a_n3565_39304# a_n4064_39072# 0.344587f
C26718 a_5742_30871# C1_N_btm 0.026156f
C26719 a_13059_46348# a_11415_45002# 0.225168f
C26720 a_3090_45724# a_3147_46376# 0.010392f
C26721 a_765_45546# a_17639_46660# 0.094916f
C26722 a_20107_46660# a_22000_46634# 3.29e-20
C26723 a_20841_46902# a_20623_46660# 0.209641f
C26724 a_20273_46660# a_21363_46634# 0.042415f
C26725 a_17339_46660# a_18280_46660# 0.002515f
C26726 a_n743_46660# a_10586_45546# 0.018104f
C26727 a_13661_43548# a_16375_45002# 0.003429f
C26728 a_19321_45002# a_13259_45724# 5.11e-20
C26729 a_5807_45002# a_19240_46482# 0.002625f
C26730 a_n881_46662# a_n1079_45724# 0.002262f
C26731 a_8270_45546# a_5937_45572# 0.29626f
C26732 a_6755_46942# a_13351_46090# 3.38e-19
C26733 a_9863_46634# a_2324_44458# 2.26e-21
C26734 a_n1613_43370# a_n863_45724# 0.027265f
C26735 a_n4318_38216# a_n4064_37984# 0.017009f
C26736 a_n3674_38216# a_n3420_37984# 0.064303f
C26737 a_20835_44721# a_20749_43396# 2e-20
C26738 a_8333_44056# a_8685_43396# 1.53e-20
C26739 a_20512_43084# a_21259_43561# 0.002989f
C26740 a_n2661_43922# a_10083_42826# 6.13e-21
C26741 a_n2293_43922# a_8952_43230# 2.5e-21
C26742 a_9313_44734# a_13635_43156# 0.013436f
C26743 a_18494_42460# a_20256_43172# 0.052522f
C26744 a_n2293_42834# a_1606_42308# 7.69e-19
C26745 a_1307_43914# a_8515_42308# 1.29e-21
C26746 a_19808_44306# a_19319_43548# 1.05e-19
C26747 a_n2661_43370# a_n3674_37592# 2.27e-20
C26748 a_n2017_45002# a_18214_42558# 2.04e-19
C26749 en_comp a_17303_42282# 1.29e-19
C26750 a_n913_45002# a_18907_42674# 1.21e-19
C26751 a_19479_31679# a_22775_42308# 3.61e-21
C26752 a_n1059_45260# a_19332_42282# 8.78e-20
C26753 a_3052_44056# VDD 0.001151f
C26754 a_7499_43078# a_3232_43370# 0.318423f
C26755 a_8568_45546# a_6171_45002# 0.005143f
C26756 a_17786_45822# a_18341_45572# 3.4e-19
C26757 a_2711_45572# a_1307_43914# 0.187968f
C26758 a_16147_45260# a_18479_45785# 0.005418f
C26759 a_6293_42852# a_4185_45028# 1.35e-20
C26760 a_4361_42308# a_19692_46634# 0.004083f
C26761 a_5649_42852# a_15227_44166# 3.43e-20
C26762 a_18429_43548# a_17339_46660# 0.033468f
C26763 a_3499_42826# a_n755_45592# 0.003508f
C26764 a_n2840_42282# a_n2312_39304# 3.28e-20
C26765 a_n3674_38680# a_n2312_40392# 0.025175f
C26766 a_15015_46420# VDD 0.337162f
C26767 a_10053_45546# a_n1741_47186# 8.64e-21
C26768 a_6511_45714# a_n1151_42308# 0.044048f
C26769 a_2711_45572# a_n443_46116# 0.060543f
C26770 a_n4209_38216# a_n3690_37440# 5.18e-19
C26771 a_n3565_38216# a_n4334_37440# 6.61e-19
C26772 a_n2293_46098# a_n863_45724# 0.003336f
C26773 a_n2157_46122# a_n1079_45724# 0.006548f
C26774 a_n1641_46494# a_n2661_45546# 7.41e-20
C26775 a_n1853_46287# a_n2293_45546# 8.68e-20
C26776 a_9823_46155# a_9751_46155# 6.64e-19
C26777 a_11189_46129# a_10586_45546# 0.028266f
C26778 a_13351_46090# a_8049_45260# 0.002917f
C26779 a_n3674_39768# a_n4318_38216# 0.032347f
C26780 a_15095_43370# a_15037_43396# 0.001617f
C26781 a_453_43940# a_961_42354# 2.06e-22
C26782 a_n97_42460# a_8952_43230# 6.13e-21
C26783 a_3905_42865# a_n784_42308# 7.08e-21
C26784 a_10341_43396# a_19700_43370# 0.013451f
C26785 a_15781_43660# a_16243_43396# 7.62e-21
C26786 a_15681_43442# a_16547_43609# 2.74e-20
C26787 a_5807_45002# START 1.22e-19
C26788 a_768_44030# CLK 1.44e-19
C26789 a_13661_43548# RST_Z 1.9e-20
C26790 a_8037_42858# VDD 0.344922f
C26791 a_11823_42460# a_14815_43914# 2.04e-19
C26792 a_2711_45572# a_18579_44172# 0.170319f
C26793 a_13249_42308# a_n2293_43922# 6.65e-19
C26794 a_10216_45572# a_5891_43370# 3.99e-20
C26795 a_6171_45002# a_n2661_43370# 2.37006f
C26796 a_7229_43940# a_7418_45067# 0.006955f
C26797 a_7276_45260# a_7735_45067# 6.64e-19
C26798 a_8191_45002# a_8488_45348# 0.004422f
C26799 a_8685_42308# a_3090_45724# 3.16e-21
C26800 a_n2302_39072# a_n2312_38680# 0.00306f
C26801 a_19862_44208# RST_Z 4.49e-21
C26802 a_n3420_37984# w_1575_34946# 3.98e-19
C26803 a_20273_45572# a_19321_45002# 1.46e-20
C26804 a_3357_43084# a_12891_46348# 6.59e-20
C26805 a_20623_45572# a_13747_46662# 4.02e-19
C26806 a_2437_43646# a_15928_47570# 0.003813f
C26807 a_19479_31679# a_12549_44172# 1.37e-20
C26808 a_n2293_45010# a_n1613_43370# 0.077436f
C26809 a_4558_45348# a_4883_46098# 2.08e-20
C26810 a_9482_43914# a_11599_46634# 8.71e-21
C26811 a_14537_43396# a_12861_44030# 0.015677f
C26812 a_5105_45348# a_4791_45118# 3.48e-19
C26813 a_16414_43172# a_16795_42852# 1.48e-19
C26814 a_3539_42460# a_5742_30871# 2.25e-20
C26815 a_3626_43646# a_11551_42558# 0.005206f
C26816 a_2982_43646# a_12563_42308# 2.07e-19
C26817 a_5649_42852# a_14635_42282# 7.52e-20
C26818 a_19741_43940# a_19647_42308# 5.24e-21
C26819 a_4520_42826# a_4649_43172# 0.010132f
C26820 a_4185_45028# RST_Z 0.005781f
C26821 a_6151_47436# a_6575_47204# 0.047329f
C26822 a_6491_46660# a_7227_47204# 0.001647f
C26823 a_4915_47217# a_11031_47542# 0.125943f
C26824 a_6545_47178# a_7903_47542# 1.49e-19
C26825 a_n1151_42308# a_14311_47204# 0.003307f
C26826 a_4007_47204# a_n1435_47204# 0.001005f
C26827 a_n2017_45002# a_n2661_42282# 0.035164f
C26828 a_3537_45260# a_7281_43914# 1.36e-20
C26829 a_4927_45028# a_5244_44056# 6.1e-21
C26830 a_3232_43370# a_3600_43914# 0.087298f
C26831 a_5147_45002# a_5495_43940# 0.086203f
C26832 a_5111_44636# a_5013_44260# 0.029412f
C26833 a_21363_45546# a_19862_44208# 3.42e-20
C26834 a_16147_45260# a_14021_43940# 2.27e-20
C26835 a_n2267_44484# a_n1821_44484# 2.28e-19
C26836 a_n1699_44726# a_n1190_44850# 2.6e-19
C26837 a_n1917_44484# a_n1809_44850# 0.057222f
C26838 a_13249_42308# a_n97_42460# 0.067568f
C26839 a_20107_45572# a_20935_43940# 1.76e-21
C26840 a_10334_44484# a_10057_43914# 0.002134f
C26841 a_10157_44484# a_8975_43940# 0.045547f
C26842 a_n2661_44458# a_n23_44458# 0.006363f
C26843 a_1576_42282# a_n443_42852# 4.39e-21
C26844 a_3318_42354# a_n755_45592# 0.152654f
C26845 a_3823_42558# a_n357_42282# 1.45e-20
C26846 a_12791_45546# VDD 0.205486f
C26847 a_13467_32519# VREF 1.56e-19
C26848 a_13159_45002# a_13059_46348# 3.4e-19
C26849 a_14180_45002# a_14513_46634# 8.73e-22
C26850 a_18989_43940# a_19321_45002# 2.21e-19
C26851 a_n2293_45010# a_n2293_46098# 5.07e-19
C26852 a_n2661_45010# a_n1853_46287# 1.83e-20
C26853 en_comp a_20820_30879# 3.02e-19
C26854 a_11525_45546# a_8049_45260# 0.002729f
C26855 a_10053_45546# a_10586_45546# 0.024917f
C26856 a_17478_45572# a_17715_44484# 0.017416f
C26857 a_16223_45938# a_15682_46116# 5.37e-19
C26858 a_15861_45028# a_18189_46348# 3.09e-20
C26859 a_12561_45572# a_2324_44458# 4.6e-19
C26860 a_9313_44734# a_n1613_43370# 3.6e-19
C26861 a_15433_44458# a_11453_44696# 9.82e-21
C26862 a_15367_44484# a_10227_46804# 5.42e-20
C26863 a_20835_44721# a_12861_44030# 3.48e-19
C26864 a_n2065_43946# a_n1151_42308# 1.27e-19
C26865 a_n984_44318# a_584_46384# 1.54e-20
C26866 a_895_43940# a_n746_45260# 3.56e-19
C26867 a_n3674_39304# a_n4209_38502# 1.61e-20
C26868 a_n473_42460# a_196_42282# 2.5e-19
C26869 a_n961_42308# a_n784_42308# 0.154417f
C26870 COMP_P a_n3674_37592# 0.054748f
C26871 a_n1736_42282# a_n1630_35242# 0.071684f
C26872 a_22165_42308# a_17303_42282# 0.095988f
C26873 a_n2661_46634# a_948_46660# 0.008972f
C26874 a_n1925_46634# a_n133_46660# 0.053144f
C26875 a_n1021_46688# a_n2438_43548# 0.053225f
C26876 a_n881_46662# a_6540_46812# 3.2e-19
C26877 a_n1613_43370# a_5072_46660# 0.012366f
C26878 a_11599_46634# a_12816_46660# 6.65e-20
C26879 a_14311_47204# a_14084_46812# 2.83e-19
C26880 a_12861_44030# a_3090_45724# 0.496275f
C26881 a_13717_47436# a_14976_45028# 2.92e-20
C26882 a_n23_47502# a_765_45546# 1.93e-20
C26883 a_13777_45326# a_13667_43396# 1.06e-21
C26884 a_11787_45002# a_10341_43396# 1.52e-22
C26885 a_18287_44626# a_11341_43940# 8.01e-21
C26886 a_19279_43940# a_22959_44484# 6.44e-21
C26887 a_5891_43370# a_10405_44172# 0.15894f
C26888 a_13556_45296# a_14579_43548# 1.57e-22
C26889 a_n2293_42834# a_3539_42460# 0.019435f
C26890 a_7499_43078# a_7573_43172# 0.002331f
C26891 a_20193_45348# a_21205_44306# 0.002474f
C26892 a_n2293_43922# a_n1441_43940# 1.93e-20
C26893 a_n699_43396# a_3052_44056# 1.83e-19
C26894 a_n2661_43922# a_261_44278# 3.53e-19
C26895 a_n2661_42834# a_n822_43940# 1.42e-19
C26896 a_n2017_45002# a_16823_43084# 5.82e-19
C26897 a_3357_43084# a_4361_42308# 3.35e-21
C26898 a_n4251_38304# VDD 3.95e-19
C26899 a_5742_30871# C9_P_btm 0.003249f
C26900 a_5932_42308# VCM 0.146001f
C26901 a_11967_42832# a_13059_46348# 2.62e-19
C26902 a_9801_44260# a_2107_46812# 9.76e-19
C26903 a_15037_43940# a_12549_44172# 2.39e-20
C26904 a_626_44172# a_n2661_45546# 0.002437f
C26905 a_2779_44458# a_2324_44458# 0.092751f
C26906 a_10057_43914# a_9290_44172# 0.034053f
C26907 a_2982_43646# a_10227_46804# 6.99e-19
C26908 a_4099_45572# DATA[2] 9.72e-21
C26909 a_13258_32519# a_22775_42308# 6.32e-19
C26910 a_19511_42282# a_21125_42558# 0.01129f
C26911 a_5742_30871# a_n4209_38502# 7.41e-22
C26912 a_n2312_40392# VDD 0.947797f
C26913 a_14097_32519# C6_N_btm 8.47e-20
C26914 a_n971_45724# a_2277_45546# 1.64e-20
C26915 a_n237_47217# a_n443_42852# 5.8e-21
C26916 a_n1151_42308# a_n755_45592# 0.03818f
C26917 a_2063_45854# a_3316_45546# 0.00135f
C26918 a_2905_45572# a_1848_45724# 5.22e-19
C26919 a_2864_46660# a_2698_46116# 4.69e-19
C26920 a_2959_46660# a_3483_46348# 5.18e-19
C26921 a_15009_46634# a_14513_46634# 0.001266f
C26922 a_3090_45724# a_14180_46812# 0.001631f
C26923 a_14084_46812# a_14226_46987# 0.005572f
C26924 a_15368_46634# a_13885_46660# 5.26e-20
C26925 a_14976_45028# a_14035_46660# 7.08e-22
C26926 a_6151_47436# a_n2661_45546# 1.33e-19
C26927 a_10227_46804# a_14371_46494# 1.79e-19
C26928 a_4883_46098# a_10044_46482# 5.79e-19
C26929 a_5534_30871# a_7754_38470# 1.19e-19
C26930 a_13675_47204# a_6945_45028# 6.96e-19
C26931 a_19321_45002# a_18189_46348# 8.52e-20
C26932 a_13661_43548# a_18985_46122# 0.006378f
C26933 a_2107_46812# a_8349_46414# 0.003223f
C26934 a_13747_46662# a_18819_46122# 0.039742f
C26935 a_n743_46660# a_11189_46129# 0.039903f
C26936 a_5807_45002# a_19553_46090# 0.00287f
C26937 a_n881_46662# a_1337_46436# 4.92e-19
C26938 a_n2017_45002# a_3497_42558# 0.0024f
C26939 a_n1059_45260# a_5379_42460# 2.17e-19
C26940 a_n913_45002# a_5267_42460# 0.081794f
C26941 a_13483_43940# a_13565_43940# 0.171361f
C26942 a_18184_42460# a_21671_42860# 0.021213f
C26943 a_11691_44458# a_17333_42852# 2.56e-21
C26944 a_6298_44484# a_5755_42852# 8.19e-21
C26945 a_11967_42832# a_15095_43370# 0.098499f
C26946 a_3905_42865# a_3080_42308# 0.029566f
C26947 a_1414_42308# a_3540_43646# 0.022584f
C26948 a_5343_44458# a_7871_42858# 0.020081f
C26949 a_n1453_44318# VDD 3.29e-19
C26950 a_11823_42460# a_13297_45572# 3.1e-20
C26951 a_8685_43396# a_15227_44166# 0.013522f
C26952 a_9803_43646# a_3090_45724# 0.002871f
C26953 a_9145_43396# a_14976_45028# 4.71e-20
C26954 a_791_42968# a_n2438_43548# 4.47e-21
C26955 a_4520_42826# a_n2293_46634# 4.07e-20
C26956 a_9885_43396# a_8270_45546# 4.58e-19
C26957 a_2982_43646# a_17339_46660# 2.08e-20
C26958 a_7542_44172# a_8049_45260# 1.33e-20
C26959 a_20679_44626# a_n357_42282# 3.64e-21
C26960 a_n2661_42282# a_526_44458# 0.191497f
C26961 a_14021_43940# a_9290_44172# 0.003037f
C26962 a_12603_44260# a_10903_43370# 0.004294f
C26963 a_12991_43230# a_12861_44030# 5.91e-20
C26964 a_n961_42308# SMPL_ON_P 1.43e-19
C26965 a_n1630_35242# w_11334_34010# 3.10971f
C26966 a_n3674_37592# a_n2497_47436# 2.17e-20
C26967 a_8487_44056# a_3483_46348# 5.36e-21
C26968 a_7174_31319# VDAC_Ni 4.91e-19
C26969 a_n1076_46494# a_n967_46494# 0.007416f
C26970 a_n901_46420# a_n722_46482# 0.007399f
C26971 a_n1641_46494# a_n1533_46116# 0.057222f
C26972 a_n1853_46287# a_n914_46116# 3.05e-19
C26973 a_13059_46348# a_13259_45724# 0.812126f
C26974 a_8270_45546# a_n443_42852# 0.063811f
C26975 a_9290_44172# a_11133_46155# 0.051331f
C26976 a_6165_46155# a_2324_44458# 4.51e-19
C26977 a_n97_42460# a_19700_43370# 0.154491f
C26978 a_n2293_43922# a_2123_42473# 3.54e-20
C26979 a_5891_43370# a_6171_42473# 2.02e-20
C26980 a_n356_44636# a_8685_42308# 1.18e-19
C26981 a_20193_45348# a_22775_42308# 1.84e-19
C26982 a_8147_43396# a_8317_43396# 0.001675f
C26983 a_21381_43940# a_21259_43561# 0.013931f
C26984 SMPL_ON_N CAL_P 0.018369f
C26985 a_9067_47204# CLK 1.63e-19
C26986 a_11031_47542# DATA[5] 0.006702f
C26987 a_9313_45822# DATA[4] 0.0373f
C26988 a_14955_47212# RST_Z 1.35e-19
C26989 a_n1435_47204# DATA[1] 0.037154f
C26990 a_18525_43370# VDD 0.263553f
C26991 a_3537_45260# a_6431_45366# 1.48e-19
C26992 a_5147_45002# a_5691_45260# 0.035185f
C26993 a_5111_44636# a_4927_45028# 0.134309f
C26994 a_4558_45348# a_3232_43370# 6.67e-21
C26995 a_n913_45002# a_14537_43396# 0.003001f
C26996 a_8746_45002# a_9838_44484# 6.4e-19
C26997 a_7499_43078# a_8975_43940# 0.519621f
C26998 a_10180_45724# a_10334_44484# 7.3e-20
C26999 a_15861_45028# a_18315_45260# 1.06e-20
C27000 a_17478_45572# a_17719_45144# 3.17e-19
C27001 a_10193_42453# a_10157_44484# 0.001446f
C27002 a_10991_42826# a_4185_45028# 3.72e-20
C27003 a_13258_32519# a_12549_44172# 1.15e-21
C27004 a_17303_42282# a_13661_43548# 9.85e-21
C27005 a_6197_43396# a_n755_45592# 1.2e-20
C27006 a_2813_43396# a_n2661_45546# 2.3e-20
C27007 a_1987_43646# a_n443_42852# 8.61e-20
C27008 a_5755_42852# a_5937_45572# 6.93e-21
C27009 a_n2302_39866# a_n2312_39304# 0.001835f
C27010 a_3422_30871# VREF_GND 0.10463f
C27011 a_11962_45724# a_n2661_46634# 0.020358f
C27012 a_10053_45546# a_n743_46660# 3.51e-20
C27013 a_19431_45546# a_18597_46090# 0.062716f
C27014 a_18787_45572# a_16327_47482# 9.38e-19
C27015 a_16789_45572# a_10227_46804# 1.86e-22
C27016 a_20623_45572# a_11599_46634# 1.32e-21
C27017 a_3357_43084# a_7903_47542# 1.35e-19
C27018 a_2437_43646# a_9863_47436# 0.005338f
C27019 a_5691_45260# a_n2109_47186# 0.113268f
C27020 a_3429_45260# a_n971_45724# 0.171338f
C27021 a_8685_43396# a_14635_42282# 2.12e-19
C27022 a_13678_32519# a_5534_30871# 0.043974f
C27023 a_14021_43940# a_15051_42282# 1.01e-20
C27024 a_9165_43940# a_8685_42308# 3.85e-21
C27025 a_n1557_42282# a_n4318_37592# 0.004047f
C27026 a_19862_44208# a_17303_42282# 4.5e-20
C27027 a_4190_30871# a_17333_42852# 0.001829f
C27028 a_743_42282# a_17701_42308# 0.014357f
C27029 a_4361_42308# a_5342_30871# 0.047616f
C27030 a_5649_42852# a_14543_43071# 8.21e-22
C27031 a_18079_43940# a_18214_42558# 3.88e-21
C27032 a_10933_46660# CLK 0.002047f
C27033 a_7754_38636# VDAC_Ni 1.97e-19
C27034 a_1149_42558# VDD 4.29e-19
C27035 a_n2497_47436# a_n815_47178# 0.003116f
C27036 a_n1920_47178# a_n1741_47186# 0.173125f
C27037 a_n2109_47186# SMPL_ON_P 0.049302f
C27038 a_11963_45334# a_n2661_43922# 4.65e-20
C27039 a_22223_45036# a_18114_32519# 0.15655f
C27040 a_1423_45028# a_8375_44464# 0.032906f
C27041 a_11827_44484# a_19721_31679# 6.72e-20
C27042 a_9482_43914# a_10617_44484# 1.06e-19
C27043 a_6171_45002# a_11909_44484# 3.97e-20
C27044 a_12800_43218# a_n357_42282# 0.002279f
C27045 a_5379_42460# a_n1925_42282# 2.1e-20
C27046 a_6123_31319# a_n2956_39304# 4.63e-21
C27047 a_13657_42558# a_10903_43370# 2.45e-20
C27048 a_17303_42282# a_4185_45028# 0.235259f
C27049 a_16115_45572# a_12741_44636# 2.27e-20
C27050 a_8696_44636# a_11415_45002# 0.10924f
C27051 a_18911_45144# a_13747_46662# 2.43e-19
C27052 a_19778_44110# a_13661_43548# 1.55e-19
C27053 a_11691_44458# a_768_44030# 0.029945f
C27054 a_20193_45348# a_12549_44172# 0.587618f
C27055 a_2809_45348# a_3877_44458# 2.21e-20
C27056 a_18315_45260# a_19321_45002# 5.84e-20
C27057 a_8953_45002# a_10150_46912# 3.4e-19
C27058 a_5205_44484# a_6755_46942# 2.7e-19
C27059 a_n913_45002# a_3090_45724# 0.039732f
C27060 a_20447_31679# a_19692_46634# 2.89e-20
C27061 a_10193_42453# a_10355_46116# 0.058019f
C27062 a_10180_45724# a_9290_44172# 0.037823f
C27063 a_10053_45546# a_11189_46129# 1.92e-19
C27064 a_9838_44484# a_4883_46098# 0.00188f
C27065 a_18287_44626# a_16327_47482# 0.552724f
C27066 a_14539_43914# a_10227_46804# 0.012909f
C27067 a_n356_44636# a_12861_44030# 4.56e-21
C27068 a_n2661_43922# a_584_46384# 0.0255f
C27069 a_9313_44734# a_4791_45118# 5.17e-19
C27070 a_n2661_42834# a_2063_45854# 0.022984f
C27071 a_13467_32519# a_20712_42282# 0.003044f
C27072 a_743_42282# a_21613_42308# 1.39e-19
C27073 a_21487_43396# a_21335_42336# 5.61e-19
C27074 a_21855_43396# a_13258_32519# 2.82e-20
C27075 a_5649_42852# a_19511_42282# 1.09e-19
C27076 a_4361_42308# a_20107_42308# 0.010379f
C27077 a_5534_30871# a_6123_31319# 0.01835f
C27078 a_4190_30871# a_18997_42308# 6.68e-19
C27079 a_n1099_45572# DATA[0] 1.56e-20
C27080 a_n971_45724# a_6755_46942# 0.185154f
C27081 a_2063_45854# a_8145_46902# 0.003229f
C27082 a_n237_47217# a_10554_47026# 3.85e-20
C27083 a_n1151_42308# a_5429_46660# 4.3e-19
C27084 a_4791_45118# a_5072_46660# 7.69e-21
C27085 a_6545_47178# a_4817_46660# 1.23e-20
C27086 a_7227_47204# a_4646_46812# 0.01221f
C27087 a_4915_47217# a_5732_46660# 4.19e-20
C27088 a_10227_46804# a_2107_46812# 0.002063f
C27089 a_12465_44636# a_n2293_46634# 0.012816f
C27090 a_3357_43084# a_7274_43762# 6.44e-21
C27091 a_5111_44636# a_4699_43561# 9.88e-20
C27092 a_n1059_45260# a_7287_43370# 8.2e-20
C27093 a_n913_45002# a_6547_43396# 1.48e-20
C27094 a_5147_45002# a_3080_42308# 1.53e-20
C27095 a_18184_42460# a_19478_44306# 7.63e-21
C27096 a_18494_42460# a_15493_43396# 7.22e-20
C27097 a_11691_44458# a_13483_43940# 7.11e-21
C27098 a_5883_43914# a_6453_43914# 0.051468f
C27099 a_19778_44110# a_19862_44208# 0.213467f
C27100 a_11827_44484# a_17973_43940# 0.004848f
C27101 a_6298_44484# a_7845_44172# 0.007037f
C27102 a_8191_45002# VDD 0.39677f
C27103 COMP_P EN_VIN_BSTR_P 6.4e-19
C27104 a_8333_44056# a_768_44030# 0.006943f
C27105 a_7281_43914# a_n2293_46634# 7.08e-20
C27106 a_n3674_39768# a_n2956_39768# 0.023472f
C27107 a_14539_43914# a_17339_46660# 4.86e-21
C27108 a_20447_31679# a_20692_30879# 9.02991f
C27109 a_15682_43940# a_n881_46662# 8.75e-21
C27110 a_7639_45394# a_2324_44458# 0.001717f
C27111 a_n2661_43370# a_10903_43370# 3.63e-19
C27112 a_n2129_43609# a_n1151_42308# 0.019226f
C27113 a_n447_43370# a_584_46384# 1.6e-19
C27114 a_327_47204# VDD 0.367528f
C27115 a_n3674_37592# a_n4209_39304# 5.44e-20
C27116 a_14113_42308# a_15803_42450# 0.289859f
C27117 a_15051_42282# a_15764_42576# 0.042737f
C27118 a_4190_30871# a_7754_38470# 8.52e-20
C27119 VREF VCM 45.1232f
C27120 a_5807_45002# a_12741_44636# 0.041091f
C27121 a_19321_45002# a_20202_43084# 2.61e-20
C27122 a_948_46660# a_765_45546# 7.87e-19
C27123 a_6755_46942# a_8023_46660# 0.004684f
C27124 a_10554_47026# a_8270_45546# 9.49e-20
C27125 a_n881_46662# a_1823_45246# 0.155149f
C27126 a_4883_46098# a_9823_46155# 0.046689f
C27127 a_11599_46634# a_18819_46122# 0.314824f
C27128 a_10227_46804# a_14493_46090# 0.202633f
C27129 a_16327_47482# a_15682_46116# 0.050548f
C27130 a_11459_47204# a_6945_45028# 0.010682f
C27131 a_2063_45854# a_5066_45546# 0.055269f
C27132 a_4007_47204# a_526_44458# 6.28e-22
C27133 a_n971_45724# a_8049_45260# 0.078318f
C27134 a_n237_47217# a_6633_46155# 0.002406f
C27135 a_18287_44626# a_10341_43396# 2.54e-20
C27136 a_10729_43914# a_10949_43914# 0.418928f
C27137 a_10405_44172# a_10807_43548# 0.004649f
C27138 a_20193_45348# a_21855_43396# 0.001332f
C27139 a_11823_42460# a_11633_42558# 0.039752f
C27140 a_10193_42453# a_14113_42308# 0.007003f
C27141 a_895_43940# a_726_44056# 8.79e-19
C27142 a_1414_42308# a_2455_43940# 1.52e-20
C27143 a_2479_44172# a_1241_43940# 7.25e-20
C27144 a_n2293_42834# a_8605_42826# 1.62e-19
C27145 a_3065_45002# a_4149_42891# 4.76e-19
C27146 a_5111_44636# a_6101_43172# 2.6e-20
C27147 a_9049_44484# a_10180_45724# 3.43e-20
C27148 a_6511_45714# a_6977_45572# 0.001881f
C27149 a_6472_45840# a_8336_45822# 2.77e-20
C27150 a_2711_45572# a_11682_45822# 0.006243f
C27151 a_6667_45809# a_6905_45572# 0.001705f
C27152 a_6598_45938# a_6469_45572# 4.2e-19
C27153 a_8568_45546# a_8746_45002# 1.75e-19
C27154 a_7499_43078# a_10193_42453# 0.298293f
C27155 a_20365_43914# a_11415_45002# 2.15e-20
C27156 a_20623_43914# a_20202_43084# 1.77e-21
C27157 a_6293_42852# a_5257_43370# 0.001148f
C27158 a_20301_43646# a_12549_44172# 0.008227f
C27159 a_n23_44458# a_n1099_45572# 7.95e-21
C27160 a_n356_44636# a_310_45028# 2.32e-19
C27161 a_7845_44172# a_5937_45572# 1.02e-19
C27162 a_n3674_39304# a_n2312_39304# 0.023737f
C27163 a_n4318_38680# a_n2312_40392# 0.025333f
C27164 a_7871_42858# a_10227_46804# 7.12e-22
C27165 a_12379_42858# a_12861_44030# 2.07e-20
C27166 a_19963_31679# VREF_GND 0.001997f
C27167 a_20447_31679# VIN_N 0.028787f
C27168 a_n2293_46098# a_2202_46116# 0.002053f
C27169 a_n901_46420# a_472_46348# 2.86e-20
C27170 a_n1076_46494# a_376_46348# 4.41e-20
C27171 a_20820_30879# a_4185_45028# 2.33e-19
C27172 a_1799_45572# a_3218_45724# 2.5e-21
C27173 a_8023_46660# a_8049_45260# 1.59e-19
C27174 a_5932_42308# VDAC_Ni 5.53e-19
C27175 a_12347_46660# a_10809_44734# 0.001417f
C27176 a_765_45546# a_13925_46122# 4.47e-20
C27177 a_16388_46812# a_17715_44484# 0.032772f
C27178 a_n2956_37592# a_n2860_38778# 3.22e-20
C27179 en_comp a_n2302_38778# 1.86e-19
C27180 a_1209_43370# a_1427_43646# 0.08213f
C27181 a_1049_43396# a_n1557_42282# 0.211757f
C27182 a_n447_43370# a_n144_43396# 0.001377f
C27183 a_742_44458# a_2123_42473# 9.65e-21
C27184 a_2998_44172# a_3681_42891# 6.9e-21
C27185 a_20679_44626# a_21356_42826# 1.01e-20
C27186 a_19279_43940# a_19164_43230# 7.21e-21
C27187 a_11341_43940# a_19268_43646# 5.82e-20
C27188 a_15493_43940# a_18783_43370# 1.32e-19
C27189 a_4093_43548# a_3080_42308# 0.08049f
C27190 a_4235_43370# a_4699_43561# 0.007134f
C27191 a_11750_44172# a_743_42282# 8.68e-22
C27192 a_18079_43940# a_16823_43084# 5.17e-20
C27193 a_20640_44752# a_21195_42852# 2.95e-22
C27194 a_20835_44721# a_20922_43172# 1.53e-20
C27195 a_9313_44734# a_13814_43218# 1.02e-19
C27196 w_11334_34010# a_11530_34132# 37.743603f
C27197 a_3540_43646# VDD 0.209044f
C27198 a_15903_45785# a_14537_43396# 9.9e-21
C27199 a_8746_45002# a_n2661_43370# 0.052623f
C27200 a_8696_44636# a_13159_45002# 7.18e-20
C27201 a_10193_42453# a_11915_45394# 0.001156f
C27202 a_22591_45572# a_22959_45572# 7.52e-19
C27203 a_3357_43084# a_20447_31679# 3.48e-19
C27204 a_17333_42852# a_15227_44166# 0.043277f
C27205 a_n1630_35242# a_n2442_46660# 0.02547f
C27206 a_7112_43396# a_526_44458# 9.09e-20
C27207 a_1241_43940# a_n443_42852# 3.12e-20
C27208 a_13943_43396# a_9290_44172# 0.003427f
C27209 a_8515_42308# a_n1613_43370# 7.89e-20
C27210 a_5742_30871# a_n2312_39304# 6.2e-21
C27211 a_17124_42282# a_16327_47482# 1.39e-20
C27212 a_n3565_39304# SMPL_ON_P 0.001067f
C27213 a_11315_46155# VDD 1.9e-20
C27214 a_2711_45572# a_n1613_43370# 0.028041f
C27215 a_8568_45546# a_4883_46098# 1.93e-19
C27216 a_12427_45724# a_10227_46804# 6.03e-20
C27217 a_n2956_38680# a_n2661_45546# 0.003946f
C27218 a_21259_43561# a_5649_42852# 1.29e-20
C27219 a_8685_43396# a_14543_43071# 4.35e-20
C27220 a_4190_30871# a_13678_32519# 0.032285f
C27221 a_4905_42826# a_5193_43172# 0.00336f
C27222 a_743_42282# a_4361_42308# 7.66647f
C27223 a_3422_30871# a_7174_31319# 2.22059f
C27224 a_10695_43548# a_10341_42308# 1.31e-19
C27225 VDAC_P C0_dummy_P_btm 0.88451f
C27226 VDAC_N C0_N_btm 0.901121f
C27227 a_7309_42852# VDD 0.177437f
C27228 a_n2293_45010# a_n1243_44484# 3.45e-19
C27229 a_3357_43084# a_5891_43370# 0.013053f
C27230 a_3232_43370# a_9838_44484# 0.053106f
C27231 a_n913_45002# a_n356_44636# 0.640597f
C27232 a_7276_45260# a_6298_44484# 0.007535f
C27233 a_6171_45002# a_5883_43914# 0.002503f
C27234 a_8696_44636# a_11967_42832# 9.33e-19
C27235 a_5755_42852# a_n443_42852# 0.008806f
C27236 a_10341_42308# a_n357_42282# 0.057131f
C27237 a_15599_45572# a_14976_45028# 5.65e-21
C27238 a_15903_45785# a_3090_45724# 0.006612f
C27239 a_15143_45578# a_13059_46348# 0.262261f
C27240 a_9482_43914# a_13661_43548# 0.127225f
C27241 a_13556_45296# a_5807_45002# 0.017285f
C27242 a_375_42282# a_768_44030# 3.77e-19
C27243 a_2437_43646# a_5907_46634# 7.11e-20
C27244 a_5111_44636# a_n743_46660# 7.53e-20
C27245 a_7229_43940# a_n2661_46634# 2.93e-22
C27246 a_5691_45260# a_n1925_46634# 1.67e-21
C27247 a_3357_43084# a_4817_46660# 0.005952f
C27248 a_n967_45348# a_n2661_46098# 2.74e-21
C27249 a_2274_45254# a_2107_46812# 2.87e-19
C27250 a_n2661_43370# a_4883_46098# 0.022462f
C27251 a_14309_45028# a_10227_46804# 8.79e-19
C27252 a_17023_45118# a_16327_47482# 0.006152f
C27253 a_18911_45144# a_11599_46634# 1.61e-20
C27254 a_20567_45036# a_12861_44030# 3.84e-21
C27255 a_21589_35634# VDD 0.525446f
C27256 a_8103_44636# a_n971_45724# 0.003603f
C27257 a_n2129_44697# a_n1151_42308# 0.039834f
C27258 a_2711_45572# a_n2293_46098# 0.530463f
C27259 a_4190_30871# a_6123_31319# 0.018095f
C27260 a_16795_42852# a_17141_43172# 0.013377f
C27261 a_10341_43396# a_17124_42282# 9.69e-21
C27262 a_16137_43396# a_14113_42308# 2.26e-19
C27263 a_743_42282# a_6761_42308# 0.01018f
C27264 a_4361_42308# a_5755_42308# 0.010214f
C27265 a_5649_42852# a_4921_42308# 0.133152f
C27266 a_685_42968# a_n784_42308# 9.99e-21
C27267 a_15781_43660# a_15803_42450# 1.76e-20
C27268 a_n2216_39072# VDD 0.00419f
C27269 a_6151_47436# a_12891_46348# 0.169139f
C27270 a_7903_47542# a_8128_46384# 0.109077f
C27271 a_11031_47542# a_n881_46662# 0.183988f
C27272 SMPL_ON_P a_n1925_46634# 1.71e-19
C27273 a_n2109_47186# a_n2438_43548# 5.34e-19
C27274 a_n237_47217# a_n2661_46634# 0.067716f
C27275 a_10227_46804# a_11453_44696# 0.08211f
C27276 a_20990_47178# a_13507_46334# 0.017412f
C27277 a_18597_46090# a_12465_44636# 3.19e-19
C27278 a_19787_47423# a_4883_46098# 8.92e-21
C27279 a_1307_43914# a_15682_43940# 0.028719f
C27280 a_n356_44636# a_556_44484# 0.001314f
C27281 a_14539_43914# a_14815_43914# 0.099149f
C27282 a_10193_42453# a_15781_43660# 5.82e-21
C27283 a_11823_42460# a_12281_43396# 0.049968f
C27284 a_15004_44636# a_15146_44811# 0.005572f
C27285 a_8975_43940# a_12189_44484# 6.54e-20
C27286 a_20193_45348# a_20637_44484# 4.36e-19
C27287 a_11827_44484# a_22591_44484# 0.003361f
C27288 a_2274_45254# a_2253_43940# 2.55e-20
C27289 a_18057_42282# a_n357_42282# 5.64e-20
C27290 a_21671_42860# RST_Z 4.49e-21
C27291 a_1307_43914# a_1823_45246# 0.013371f
C27292 a_13777_45326# a_3483_46348# 0.027519f
C27293 a_4640_45348# a_n2293_46098# 1.74e-19
C27294 a_n2661_44458# a_3090_45724# 0.088502f
C27295 a_17719_45144# a_16388_46812# 5.03e-21
C27296 a_20159_44458# a_13661_43548# 1.06e-19
C27297 a_18545_45144# a_15227_44166# 0.002275f
C27298 a_19006_44850# a_19321_45002# 1.35e-20
C27299 a_20596_44850# a_12549_44172# 2.61e-19
C27300 a_8696_44636# a_13259_45724# 0.259609f
C27301 a_16115_45572# a_16375_45002# 1.66e-19
C27302 a_19431_45546# a_8049_45260# 0.006516f
C27303 a_6171_45002# a_9569_46155# 6.04e-21
C27304 a_413_45260# a_14840_46494# 2.43e-21
C27305 a_7276_45260# a_5937_45572# 0.052629f
C27306 a_7229_43940# a_8199_44636# 1.98e-19
C27307 a_8191_45002# a_7920_46348# 1.55e-20
C27308 a_5755_42308# a_6761_42308# 2.13e-19
C27309 a_1606_42308# a_11323_42473# 1.34e-20
C27310 CAL_P a_18194_35068# 0.010626f
C27311 a_n1838_35608# a_n1386_35608# 0.150796f
C27312 a_n1741_47186# a_9290_44172# 9.99e-21
C27313 a_2063_45854# a_5068_46348# 0.004281f
C27314 a_n237_47217# a_8199_44636# 0.089777f
C27315 a_n971_45724# a_8953_45546# 5.83e-21
C27316 a_n2661_46634# a_8270_45546# 0.037557f
C27317 a_5807_45002# a_13607_46688# 0.002972f
C27318 a_3877_44458# a_4817_46660# 0.017126f
C27319 a_4646_46812# a_4955_46873# 0.047208f
C27320 a_768_44030# a_15227_44166# 3.48e-22
C27321 a_13747_46662# a_12991_46634# 1.32e-20
C27322 a_n1925_46634# a_8035_47026# 2.38e-20
C27323 a_12549_44172# a_19333_46634# 3.59e-19
C27324 a_n1151_42308# a_3483_46348# 8.25e-19
C27325 a_3160_47472# a_3699_46348# 0.109505f
C27326 a_n443_46116# a_1823_45246# 0.217935f
C27327 a_2905_45572# a_4185_45028# 1.92e-21
C27328 a_16327_47482# a_20719_46660# 5.41e-20
C27329 a_18597_46090# a_20528_46660# 8.24e-19
C27330 a_20990_47178# a_20623_46660# 0.004006f
C27331 a_21177_47436# a_20841_46902# 0.001161f
C27332 a_13507_46334# a_20273_46660# 0.026778f
C27333 a_4883_46098# a_20107_46660# 1.93e-19
C27334 a_12465_44636# a_19123_46287# 1.94e-20
C27335 a_11453_44696# a_17339_46660# 0.071641f
C27336 a_n1059_45260# a_12089_42308# 0.022942f
C27337 a_n2017_45002# a_12545_42858# 1.03e-19
C27338 a_n913_45002# a_12379_42858# 0.066604f
C27339 a_3537_45260# a_3935_42891# 0.001584f
C27340 a_n699_43396# a_3540_43646# 7.76e-19
C27341 a_n2661_42834# a_5326_44056# 2.01e-19
C27342 a_9313_44734# a_10651_43940# 2.96e-19
C27343 a_18579_44172# a_15682_43940# 1.06e-20
C27344 a_7499_43078# a_n784_42308# 6.51e-20
C27345 a_11967_42832# a_20365_43914# 7.55e-20
C27346 a_3905_42865# a_5013_44260# 0.182997f
C27347 a_20159_44458# a_19862_44208# 8.53e-20
C27348 a_18287_44626# a_n97_42460# 2.47e-20
C27349 a_16979_44734# VDD 0.256327f
C27350 a_n4064_39616# C9_P_btm 0.215899f
C27351 a_n3420_39616# C7_P_btm 8.17e-19
C27352 a_n3565_39590# C5_P_btm 1.31e-19
C27353 a_n3565_39304# a_n1532_35090# 1.16e-19
C27354 a_18451_43940# a_3090_45724# 0.004024f
C27355 a_13483_43940# a_15227_44166# 1.48e-20
C27356 a_15301_44260# a_6755_46942# 1.12e-19
C27357 a_13076_44458# a_8049_45260# 2.05e-21
C27358 a_18494_42460# a_n357_42282# 0.033084f
C27359 a_7466_43396# a_n1613_43370# 0.001965f
C27360 a_19268_43646# a_16327_47482# 0.024286f
C27361 a_n722_43218# a_n971_45724# 3.38e-19
C27362 a_1983_46706# VDD 0.119964f
C27363 a_n3420_39616# a_n3565_38502# 0.028014f
C27364 a_n4064_39616# a_n4209_38502# 0.02801f
C27365 a_n3565_39590# a_n3420_38528# 0.031237f
C27366 a_n4209_39590# a_n4064_38528# 0.032071f
C27367 a_n4209_39304# a_n2302_39072# 0.407162f
C27368 a_n3565_39304# a_n2946_39072# 0.410957f
C27369 a_n3690_39392# a_n3420_39072# 0.414961f
C27370 a_n4334_39392# a_n4064_39072# 0.410653f
C27371 a_1239_39587# comp_n 0.001233f
C27372 a_1736_39587# a_1736_39043# 1.92825f
C27373 a_5742_30871# C0_N_btm 0.014563f
C27374 a_17339_46660# a_17639_46660# 0.081726f
C27375 a_20273_46660# a_20623_46660# 0.20669f
C27376 a_20107_46660# a_21188_46660# 0.102355f
C27377 a_19123_46287# a_20528_46660# 1.39e-20
C27378 a_2107_46812# a_8034_45724# 0.006608f
C27379 a_5807_45002# a_16375_45002# 0.042941f
C27380 a_2864_46660# a_526_44458# 8.51e-20
C27381 a_n743_46660# a_8379_46155# 1.92e-19
C27382 a_n881_46662# a_n2293_45546# 0.004473f
C27383 a_8270_45546# a_8199_44636# 0.95539f
C27384 a_6755_46942# a_12594_46348# 1.41e-19
C27385 a_8492_46660# a_2324_44458# 1.06e-20
C27386 a_n1613_43370# a_n1079_45724# 0.013012f
C27387 a_n3674_38216# a_n3690_38304# 0.071735f
C27388 a_n4318_38216# a_n2946_37984# 4.19e-20
C27389 a_20679_44626# a_20749_43396# 1.57e-21
C27390 a_3422_30871# a_21487_43396# 0.003721f
C27391 a_n2661_43922# a_8952_43230# 6.16e-22
C27392 a_n2661_42834# a_10083_42826# 2.3e-20
C27393 a_n2293_43922# a_9127_43156# 6.49e-20
C27394 a_9313_44734# a_12895_43230# 0.007885f
C27395 a_18184_42460# a_20256_43172# 0.043416f
C27396 a_375_42282# a_6123_31319# 1.31e-20
C27397 a_1307_43914# a_5934_30871# 3.28e-21
C27398 a_15493_43940# a_3626_43646# 3.83e-20
C27399 a_n2017_45002# a_19332_42282# 1.65e-19
C27400 en_comp a_4958_30871# 0.086457f
C27401 a_n1059_45260# a_18907_42674# 0.001868f
C27402 a_n913_45002# a_18727_42674# 2.28e-19
C27403 a_2455_43940# VDD 0.144352f
C27404 a_6812_45938# a_5205_44484# 4.18e-20
C27405 a_8162_45546# a_6171_45002# 0.008027f
C27406 a_8568_45546# a_3232_43370# 4.2e-21
C27407 a_2711_45572# a_16019_45002# 0.024255f
C27408 a_16147_45260# a_18175_45572# 0.108647f
C27409 a_6197_43396# a_3483_46348# 8.08e-22
C27410 a_6031_43396# a_4185_45028# 4.43e-21
C27411 a_13467_32519# a_19692_46634# 0.015407f
C27412 a_17324_43396# a_17339_46660# 6.45e-20
C27413 a_3499_42826# a_n357_42282# 0.007965f
C27414 a_n2840_42282# a_n2312_40392# 4.5e-20
C27415 a_14275_46494# VDD 0.196859f
C27416 a_3775_45552# a_2063_45854# 1.46e-19
C27417 a_6472_45840# a_n1151_42308# 0.01357f
C27418 a_4099_45572# a_4007_47204# 4.68e-19
C27419 a_2711_45572# a_4791_45118# 0.160646f
C27420 a_1609_45572# a_n443_46116# 2.27e-19
C27421 a_6812_45938# a_n971_45724# 1.09e-19
C27422 a_n4209_38216# a_n3565_37414# 0.031622f
C27423 a_n3565_38216# a_n4209_37414# 5.88577f
C27424 a_n4334_38304# a_n4334_37440# 0.050585f
C27425 a_n2293_46098# a_n1079_45724# 0.003233f
C27426 a_n2157_46122# a_n2293_45546# 6.79e-20
C27427 a_9625_46129# a_10037_46155# 0.006879f
C27428 a_9290_44172# a_10586_45546# 0.264957f
C27429 a_12594_46348# a_8049_45260# 0.069217f
C27430 a_n2956_38680# a_n1533_46116# 9.67e-20
C27431 a_3422_30871# a_5932_42308# 0.022048f
C27432 a_n4318_39768# a_n4318_38216# 0.023318f
C27433 a_n97_42460# a_9127_43156# 1.6e-19
C27434 a_10341_43396# a_19268_43646# 0.010402f
C27435 a_15681_43442# a_16243_43396# 6.39e-21
C27436 a_15781_43660# a_16137_43396# 0.089942f
C27437 a_453_43940# a_1184_42692# 2.56e-21
C27438 a_12549_44172# CLK 3.33e-19
C27439 a_5807_45002# RST_Z 1.85e-19
C27440 a_7765_42852# VDD 0.333322f
C27441 a_3232_43370# a_n2661_43370# 0.077167f
C27442 a_8953_45002# a_n2293_42834# 1.18e-19
C27443 a_7276_45260# a_7418_45067# 0.005572f
C27444 a_6171_45002# a_11361_45348# 8.73e-20
C27445 a_14097_32519# a_20202_43084# 7.09e-21
C27446 a_n4064_39072# a_n2312_38680# 0.002525f
C27447 a_13467_32519# a_20692_30879# 0.051714f
C27448 a_16759_43396# a_n443_42852# 1.02e-20
C27449 a_5907_45546# a_3090_45724# 4.4e-21
C27450 a_20107_45572# a_19321_45002# 0.006336f
C27451 a_16147_45260# a_n743_46660# 0.071228f
C27452 a_2437_43646# a_768_44030# 0.137571f
C27453 a_20841_45814# a_13747_46662# 1.63e-19
C27454 a_3357_43084# a_11309_47204# 8.86e-21
C27455 a_n2661_45010# a_n881_46662# 1.04e-19
C27456 a_5093_45028# a_2063_45854# 1.55e-21
C27457 a_9396_43370# a_5934_30871# 4.98e-19
C27458 a_3626_43646# a_5742_30871# 0.168508f
C27459 a_5649_42852# a_13291_42460# 5.5e-20
C27460 a_n97_42460# a_17124_42282# 5.78e-20
C27461 a_15743_43084# a_20753_42852# 1.06e-19
C27462 a_6491_46660# a_6851_47204# 0.132946f
C27463 a_6151_47436# a_7903_47542# 7.86e-20
C27464 a_4915_47217# a_9863_47436# 0.018512f
C27465 a_5815_47464# a_6575_47204# 0.009009f
C27466 a_6545_47178# a_7227_47204# 0.001559f
C27467 a_3815_47204# a_n1435_47204# 2.24e-19
C27468 a_n1151_42308# a_13487_47204# 1.36e-19
C27469 a_3537_45260# a_6453_43914# 6.46e-19
C27470 a_3232_43370# a_2998_44172# 0.056614f
C27471 a_5147_45002# a_5013_44260# 0.189328f
C27472 a_4927_45028# a_3905_42865# 1.58e-19
C27473 a_5111_44636# a_5244_44056# 0.01138f
C27474 a_20623_45572# a_19862_44208# 7.47e-20
C27475 a_11827_44484# a_9313_44734# 1.07e-19
C27476 a_n2267_44484# a_n1190_44850# 1.46e-19
C27477 a_n1917_44484# a_n2012_44484# 0.049827f
C27478 a_10157_44484# a_10057_43914# 6.36e-19
C27479 a_9838_44484# a_8975_43940# 0.055678f
C27480 a_n2661_44458# a_n356_44636# 0.055568f
C27481 a_n1699_44726# a_n1809_44850# 0.097745f
C27482 a_10334_44484# a_10440_44484# 0.313533f
C27483 a_1067_42314# a_n443_42852# 0.011239f
C27484 a_3318_42354# a_n357_42282# 1.18e-20
C27485 a_2903_42308# a_n755_45592# 0.070479f
C27486 a_11823_42460# VDD 4.44574f
C27487 a_13467_32519# VIN_N 0.078487f
C27488 a_13017_45260# a_13059_46348# 0.022433f
C27489 a_14180_45002# a_14180_46812# 1.22e-20
C27490 a_18374_44850# a_19321_45002# 1.39e-20
C27491 a_n2472_45002# a_n2293_46098# 0.001044f
C27492 a_n2661_45010# a_n2157_46122# 4.29e-20
C27493 a_9049_44484# a_10586_45546# 0.002146f
C27494 a_11322_45546# a_8049_45260# 0.004301f
C27495 a_5891_43370# a_8128_46384# 1.23e-21
C27496 a_15037_45618# a_6945_45028# 3.02e-21
C27497 a_15861_45028# a_17715_44484# 0.184272f
C27498 a_17478_45572# a_17583_46090# 3.05e-19
C27499 a_16020_45572# a_15682_46116# 3.39e-19
C27500 a_14127_45572# a_12594_46348# 6.01e-19
C27501 a_8696_44636# a_18189_46348# 2.18e-21
C27502 a_14815_43914# a_11453_44696# 6.62e-20
C27503 a_17517_44484# a_18479_47436# 0.017833f
C27504 a_15146_44484# a_10227_46804# 2.64e-22
C27505 a_20679_44626# a_12861_44030# 8.93e-19
C27506 a_2127_44172# a_n237_47217# 3.02e-21
C27507 a_n1329_42308# a_n784_42308# 9.6e-19
C27508 a_n3674_38216# a_n1630_35242# 0.333493f
C27509 a_n4318_37592# a_n3674_37592# 3.06402f
C27510 a_19164_43230# a_19332_42282# 0.002067f
C27511 a_21671_42860# a_17303_42282# 3.64e-20
C27512 a_n2661_46634# a_1123_46634# 0.012266f
C27513 a_n2293_46634# a_33_46660# 6.74e-21
C27514 a_n1021_46688# a_n743_46660# 0.11001f
C27515 a_n1925_46634# a_n2438_43548# 0.166008f
C27516 a_n1613_43370# a_6540_46812# 0.05541f
C27517 a_12465_44636# a_6755_46942# 0.021176f
C27518 a_11599_46634# a_12991_46634# 4.06e-20
C27519 a_10227_46804# a_10384_47026# 1.7e-19
C27520 a_13717_47436# a_3090_45724# 2.02e-20
C27521 a_12861_44030# a_15009_46634# 0.058082f
C27522 a_13487_47204# a_14084_46812# 0.012167f
C27523 a_4915_47217# a_12978_47026# 1.2e-19
C27524 a_n1151_42308# a_14513_46634# 0.042579f
C27525 a_n237_47217# a_765_45546# 0.1364f
C27526 a_2063_45854# a_13059_46348# 5.17e-21
C27527 a_22223_45036# a_14401_32519# 3.29e-20
C27528 a_13556_45296# a_13667_43396# 1.26e-20
C27529 a_18248_44752# a_11341_43940# 6.59e-20
C27530 a_19279_43940# a_17730_32519# 1.25e-20
C27531 a_5891_43370# a_9672_43914# 0.009207f
C27532 a_14537_43396# a_9145_43396# 0.129182f
C27533 a_11827_44484# a_20974_43370# 2.22e-20
C27534 a_3363_44484# a_3499_42826# 1.97e-20
C27535 a_21398_44850# a_3422_30871# 2.52e-19
C27536 a_7499_43078# a_7309_43172# 0.001045f
C27537 a_n2293_42834# a_3626_43646# 0.019674f
C27538 a_n2661_42834# a_261_44278# 3.83e-19
C27539 a_18579_44172# a_20512_43084# 3.29e-19
C27540 a_n2302_37984# VDD 0.350854f
C27541 a_5742_30871# C10_P_btm 0.00237f
C27542 a_5932_42308# VREF_GND 0.001404f
C27543 a_9248_44260# a_2107_46812# 1.38e-19
C27544 a_13565_43940# a_12549_44172# 4.78e-21
C27545 a_501_45348# a_n2661_45546# 1.17e-19
C27546 a_949_44458# a_2324_44458# 0.323116f
C27547 a_10440_44484# a_9290_44172# 5.93e-21
C27548 a_13258_32519# a_21613_42308# 0.060546f
C27549 a_22959_47212# VDD 0.245964f
C27550 a_14097_32519# C5_N_btm 0.001712f
C27551 a_3160_47472# a_n755_45592# 0.001373f
C27552 a_n443_46116# a_n2293_45546# 0.004986f
C27553 a_n746_45260# a_n443_42852# 0.136813f
C27554 a_2063_45854# a_3218_45724# 0.004182f
C27555 a_584_46384# a_3316_45546# 1.77e-21
C27556 a_n971_45724# a_1609_45822# 1.47e-19
C27557 a_n1151_42308# a_n357_42282# 0.009369f
C27558 a_3177_46902# a_3483_46348# 2.05e-20
C27559 a_2959_46660# a_3147_46376# 0.010696f
C27560 a_8270_45546# a_765_45546# 5.94e-19
C27561 a_15009_46634# a_14180_46812# 0.123843f
C27562 a_14976_45028# a_13885_46660# 6.33e-20
C27563 a_3090_45724# a_14035_46660# 6.08e-22
C27564 a_10227_46804# a_14180_46482# 0.014179f
C27565 a_4883_46098# a_9823_46482# 2.91e-19
C27566 a_12465_44636# a_8049_45260# 0.027831f
C27567 a_13569_47204# a_6945_45028# 6.5e-19
C27568 a_13661_43548# a_18819_46122# 0.02447f
C27569 a_2107_46812# a_8016_46348# 0.022583f
C27570 a_n743_46660# a_9290_44172# 0.048675f
C27571 a_13747_46662# a_17957_46116# 1.02e-19
C27572 a_5807_45002# a_18985_46122# 0.017912f
C27573 a_n881_46662# a_n914_46116# 1.02e-19
C27574 a_n913_45002# a_3823_42558# 0.029622f
C27575 a_n2017_45002# a_5379_42460# 0.003023f
C27576 a_n1059_45260# a_5267_42460# 6.15e-20
C27577 a_1307_43914# a_16245_42852# 1.03e-20
C27578 a_14673_44172# a_14621_43646# 6.57e-20
C27579 a_18184_42460# a_21195_42852# 0.017258f
C27580 a_11827_44484# a_18599_43230# 5.4e-21
C27581 a_11967_42832# a_14205_43396# 1.68e-19
C27582 a_3905_42865# a_4699_43561# 0.001039f
C27583 a_4223_44672# a_8037_42858# 9.39e-19
C27584 a_5891_43370# a_743_42282# 0.065685f
C27585 a_1414_42308# a_2982_43646# 0.071994f
C27586 a_n1644_44306# VDD 0.082968f
C27587 a_9145_43396# a_3090_45724# 0.189557f
C27588 a_3935_42891# a_n2293_46634# 4.54e-20
C27589 a_5534_30871# a_12549_44172# 2.57e-20
C27590 a_16409_43396# a_6755_46942# 6.64e-20
C27591 a_11341_43940# a_2324_44458# 0.007112f
C27592 a_12495_44260# a_10903_43370# 0.001658f
C27593 a_n1329_42308# SMPL_ON_P 4.56e-20
C27594 a_n1630_35242# w_1575_34946# 3.10971f
C27595 a_18280_46660# VDD 6.19e-19
C27596 a_n1423_46090# a_n1533_46116# 0.097745f
C27597 a_13059_46348# a_14383_46116# 3.09e-20
C27598 a_10355_46116# a_11133_46155# 6.26e-20
C27599 a_9290_44172# a_11189_46129# 0.199578f
C27600 a_12429_44172# a_5534_30871# 3.45e-20
C27601 a_5891_43370# a_5755_42308# 7.45e-19
C27602 a_n97_42460# a_19268_43646# 0.002543f
C27603 a_n2293_43922# a_1755_42282# 1.6e-19
C27604 a_n356_44636# a_8325_42308# 1.57e-19
C27605 a_2982_43646# a_12281_43396# 4.32e-19
C27606 a_20193_45348# a_21613_42308# 0.137559f
C27607 a_8147_43396# a_8229_43396# 0.005781f
C27608 a_14311_47204# RST_Z 0.184572f
C27609 a_n1435_47204# DATA[0] 0.053257f
C27610 a_18429_43548# VDD 0.163446f
C27611 a_4558_45348# a_5691_45260# 1.08e-19
C27612 a_3537_45260# a_6171_45002# 4.04e-19
C27613 a_5147_45002# a_4927_45028# 0.168157f
C27614 a_4574_45260# a_3232_43370# 3.36e-21
C27615 a_n1059_45260# a_14537_43396# 2.86e-21
C27616 a_n2661_45010# a_1307_43914# 0.016415f
C27617 a_8696_44636# a_18315_45260# 4.09e-21
C27618 a_7499_43078# a_10057_43914# 0.262644f
C27619 a_10180_45724# a_10157_44484# 0.001525f
C27620 a_15861_45028# a_17719_45144# 0.002134f
C27621 a_17478_45572# a_17613_45144# 3.37e-20
C27622 a_8746_45002# a_5883_43914# 2.04e-20
C27623 a_15037_45618# a_11827_44484# 3.23e-22
C27624 a_10796_42968# a_4185_45028# 3.58e-20
C27625 a_15597_42852# a_15227_44166# 0.007489f
C27626 a_4958_30871# a_13661_43548# 9.87e-21
C27627 a_14205_43396# a_13259_45724# 1.43e-20
C27628 a_6293_42852# a_n755_45592# 2.52e-20
C27629 a_6197_43396# a_n357_42282# 6.51e-20
C27630 a_1891_43646# a_n443_42852# 1.53e-19
C27631 a_n2302_39866# a_n2312_40392# 8.29e-19
C27632 a_n4064_39616# a_n2312_39304# 2.53e-19
C27633 a_9049_44484# a_n743_46660# 4.38e-19
C27634 a_11652_45724# a_n2661_46634# 1.97e-19
C27635 a_18691_45572# a_18597_46090# 5.99e-19
C27636 a_19256_45572# a_18479_47436# 2.31e-22
C27637 a_19418_45938# a_16327_47482# 1.07e-19
C27638 a_3357_43084# a_7227_47204# 5.7e-19
C27639 a_2437_43646# a_9067_47204# 0.006126f
C27640 a_n2661_45010# a_n443_46116# 0.005128f
C27641 a_3065_45002# a_n971_45724# 0.220337f
C27642 a_n745_45366# a_n1151_42308# 0.004257f
C27643 a_4927_45028# a_n2109_47186# 0.00143f
C27644 a_3232_43370# a_n2497_47436# 0.04813f
C27645 a_413_45260# a_1209_47178# 3.61e-20
C27646 a_8685_43396# a_13291_42460# 2.12e-19
C27647 a_13467_32519# a_5342_30871# 0.028573f
C27648 a_18451_43940# a_18727_42674# 1.72e-21
C27649 a_14021_43940# a_14113_42308# 3.15e-20
C27650 a_n97_42460# a_1755_42282# 0.002698f
C27651 a_n1557_42282# a_n1736_42282# 0.170341f
C27652 a_743_42282# a_17595_43084# 5.58e-20
C27653 a_4190_30871# a_18083_42858# 0.023338f
C27654 a_10861_46660# CLK 9.26e-19
C27655 a_n4064_37984# VDAC_P 2.99e-19
C27656 a_3754_38802# a_3754_38470# 0.02792f
C27657 a_961_42354# VDD 0.091526f
C27658 a_n2497_47436# a_n1605_47204# 0.0417f
C27659 a_n2109_47186# a_n1741_47186# 0.18579f
C27660 a_n2288_47178# SMPL_ON_P 0.002143f
C27661 a_11322_45546# a_11173_44260# 2.01e-20
C27662 a_11787_45002# a_n2661_43922# 2.24e-20
C27663 a_11963_45334# a_n2661_42834# 9.32e-20
C27664 a_11827_44484# a_18114_32519# 0.09907f
C27665 a_1423_45028# a_7640_43914# 0.105665f
C27666 a_21359_45002# a_19721_31679# 2.35e-20
C27667 a_n2661_43370# a_8975_43940# 3.05e-19
C27668 a_3357_43084# a_22315_44484# 1.44e-21
C27669 a_3232_43370# a_11909_44484# 2.99e-20
C27670 a_4958_30871# a_4185_45028# 0.121495f
C27671 a_10752_42852# a_n357_42282# 1.14e-19
C27672 a_5379_42460# a_526_44458# 1.71e-19
C27673 a_22400_42852# a_13259_45724# 0.34531f
C27674 a_13333_42558# a_10903_43370# 0.00168f
C27675 a_16333_45814# a_12741_44636# 1.84e-20
C27676 a_16680_45572# a_11415_45002# 0.003026f
C27677 a_11691_44458# a_12549_44172# 0.025825f
C27678 a_18691_45572# a_19123_46287# 0.009086f
C27679 a_18911_45144# a_13661_43548# 0.03394f
C27680 a_n2661_43370# a_n133_46660# 2.93e-22
C27681 a_19778_44110# a_5807_45002# 0.032504f
C27682 a_2304_45348# a_3877_44458# 6.26e-21
C27683 a_17719_45144# a_19321_45002# 1.57e-20
C27684 a_8953_45002# a_9863_46634# 3.37e-20
C27685 a_6171_45002# a_6969_46634# 1.08e-20
C27686 a_n1059_45260# a_3090_45724# 0.008195f
C27687 a_10193_42453# a_9823_46155# 0.001684f
C27688 a_11652_45724# a_8199_44636# 4.91e-19
C27689 a_7499_43078# a_11133_46155# 1.49e-20
C27690 a_10490_45724# a_9625_46129# 1.99e-19
C27691 a_2711_45572# a_6945_45028# 0.036364f
C27692 a_10053_45546# a_9290_44172# 8.06e-21
C27693 a_5883_43914# a_4883_46098# 0.01188f
C27694 a_16112_44458# a_10227_46804# 0.001281f
C27695 a_18248_44752# a_16327_47482# 0.050926f
C27696 a_9241_44734# a_4791_45118# 6.15e-20
C27697 a_n2661_42834# a_584_46384# 0.079307f
C27698 a_13467_32519# a_20107_42308# 0.001069f
C27699 a_10083_42826# a_9885_42558# 0.001558f
C27700 a_n2293_42282# a_2351_42308# 6.05e-19
C27701 a_4361_42308# a_13258_32519# 0.076336f
C27702 a_20692_30879# VCM 0.035438f
C27703 a_4791_45118# a_6540_46812# 0.001459f
C27704 a_2063_45854# a_7577_46660# 0.032724f
C27705 a_n237_47217# a_10623_46897# 1.75e-20
C27706 a_n1151_42308# a_5263_46660# 0.001012f
C27707 a_6151_47436# a_4817_46660# 1.46e-20
C27708 a_6851_47204# a_4646_46812# 8.39e-20
C27709 a_5129_47502# a_5167_46660# 6.56e-19
C27710 a_n1435_47204# a_3524_46660# 7.47e-21
C27711 a_4915_47217# a_5907_46634# 1.88e-19
C27712 a_6491_46660# a_4651_46660# 1.14e-20
C27713 a_22959_47212# a_22612_30879# 0.156518f
C27714 a_n881_46662# a_15928_47570# 2.48e-20
C27715 a_3232_43370# a_1568_43370# 7.3e-19
C27716 a_n2017_45002# a_7287_43370# 1.12e-20
C27717 a_8696_44636# a_16867_43762# 1.57e-19
C27718 a_14815_43914# a_15146_44484# 2.88e-19
C27719 a_18184_42460# a_15493_43396# 7.78e-20
C27720 a_11691_44458# a_12429_44172# 2.31e-20
C27721 a_5883_43914# a_5663_43940# 0.153361f
C27722 a_19778_44110# a_19478_44306# 0.099524f
C27723 a_11827_44484# a_17737_43940# 0.003402f
C27724 a_n1809_44850# a_n1761_44111# 7.57e-20
C27725 a_6298_44484# a_7542_44172# 0.014735f
C27726 a_16922_45042# a_11341_43940# 0.028038f
C27727 a_7705_45326# VDD 0.211554f
C27728 COMP_P a_n923_35174# 0.003051f
C27729 a_18443_44721# a_16388_46812# 2.06e-20
C27730 a_6453_43914# a_n2293_46634# 6.32e-20
C27731 a_n4318_39768# a_n2956_39768# 0.023595f
C27732 a_8018_44260# a_768_44030# 9.58e-19
C27733 a_22959_45572# a_20692_30879# 4.31e-19
C27734 a_20447_31679# a_20205_31679# 9.01329f
C27735 a_7418_45394# a_2324_44458# 0.00182f
C27736 a_n2661_43370# a_11387_46155# 2.17e-21
C27737 a_n1352_43396# a_584_46384# 1.26e-20
C27738 a_458_43396# a_n971_45724# 1.17e-19
C27739 a_n785_47204# VDD 0.452945f
C27740 a_14113_42308# a_15764_42576# 0.229529f
C27741 a_15051_42282# a_15486_42560# 0.234322f
C27742 a_5932_42308# a_7174_31319# 13.0265f
C27743 VIN_N VCM 1.7189f
C27744 VREF VREF_GND 45.1141f
C27745 a_13747_46662# a_11415_45002# 0.099293f
C27746 a_1123_46634# a_765_45546# 0.025395f
C27747 a_10623_46897# a_8270_45546# 6.27e-20
C27748 a_n881_46662# a_1138_42852# 0.148785f
C27749 a_n1613_43370# a_1823_45246# 1.96e-19
C27750 a_11453_44696# a_8016_46348# 2.61e-20
C27751 a_4883_46098# a_9569_46155# 0.008675f
C27752 a_11599_46634# a_17957_46116# 0.031252f
C27753 a_10227_46804# a_13925_46122# 0.635045f
C27754 a_16241_47178# a_15682_46116# 0.001179f
C27755 a_16327_47482# a_2324_44458# 1.53e-19
C27756 a_13717_47436# a_20075_46420# 3.99e-21
C27757 a_9313_45822# a_6945_45028# 0.035455f
C27758 a_3815_47204# a_526_44458# 4.06e-21
C27759 a_n237_47217# a_6347_46155# 0.001047f
C27760 a_3785_47178# a_n1925_42282# 1.46e-20
C27761 a_n971_45724# a_8781_46436# 2.04e-19
C27762 a_18248_44752# a_10341_43396# 3.47e-20
C27763 a_10405_44172# a_10949_43914# 0.05348f
C27764 a_18579_44172# a_21381_43940# 1.29e-21
C27765 a_20193_45348# a_4361_42308# 7.54e-19
C27766 a_11823_42460# a_11551_42558# 0.138126f
C27767 a_10193_42453# a_13657_42558# 0.009218f
C27768 a_453_43940# a_1443_43940# 0.009173f
C27769 a_n2293_42834# a_8037_42858# 0.009778f
C27770 a_1414_42308# a_2253_43940# 1.35e-19
C27771 a_9672_43914# a_10807_43548# 2.13e-20
C27772 a_n2661_42834# a_n144_43396# 2.02e-19
C27773 a_n913_45002# a_12800_43218# 0.016338f
C27774 a_5111_44636# a_5837_43172# 1.31e-19
C27775 a_3537_45260# a_8292_43218# 1.01e-19
C27776 a_2711_45572# a_11280_45822# 1.69e-19
C27777 a_6472_45840# a_6977_45572# 2.28e-19
C27778 a_9049_44484# a_10053_45546# 0.005221f
C27779 a_15493_43396# a_12741_44636# 1.11e-19
C27780 a_20365_43914# a_20202_43084# 2.68e-21
C27781 a_4190_30871# a_12549_44172# 0.270972f
C27782 a_19319_43548# a_19692_46634# 5.04e-20
C27783 a_6031_43396# a_5257_43370# 0.004037f
C27784 a_n356_44636# a_n1099_45572# 5.17e-21
C27785 a_13720_44458# a_n443_42852# 1.6e-20
C27786 a_7_44811# a_n863_45724# 7.59e-19
C27787 a_7845_44172# a_8199_44636# 7.26e-19
C27788 a_7542_44172# a_5937_45572# 2.83e-19
C27789 a_n3674_39304# a_n2312_40392# 0.025635f
C27790 a_n2293_42282# a_584_46384# 8.38e-19
C27791 a_19963_31679# VREF 0.055795f
C27792 a_12741_44636# a_3483_46348# 0.023452f
C27793 a_n2293_46098# a_1823_45246# 0.107882f
C27794 a_383_46660# a_n443_42852# 1.35e-19
C27795 a_n2661_46098# a_1848_45724# 5.47e-21
C27796 a_2609_46660# a_n755_45592# 4.05e-19
C27797 a_n743_46660# a_n89_45572# 0.003687f
C27798 a_1799_45572# a_2957_45546# 7.87e-21
C27799 a_3090_45724# a_n1925_42282# 0.157861f
C27800 a_12978_47026# a_10809_44734# 1.72e-19
C27801 a_16721_46634# a_15682_46116# 0.010175f
C27802 a_765_45546# a_13759_46122# 9.6e-20
C27803 a_16388_46812# a_17583_46090# 0.033313f
C27804 en_comp a_n4064_38528# 2.01e-21
C27805 a_n2956_37592# a_n2302_38778# 0.006499f
C27806 a_3905_42865# a_1847_42826# 2.52e-20
C27807 a_1049_43396# a_766_43646# 6.4e-21
C27808 a_n699_43396# a_961_42354# 1.36e-21
C27809 a_19279_43940# a_19339_43156# 3.69e-21
C27810 a_3422_30871# a_15567_42826# 5.99e-21
C27811 a_20640_44752# a_21356_42826# 7.48e-22
C27812 a_18579_44172# a_18249_42858# 1.81e-20
C27813 a_2998_44172# a_2905_42968# 3.82e-19
C27814 a_n1441_43940# a_n1641_43230# 5.44e-21
C27815 a_11341_43940# a_15743_43084# 6.7e-19
C27816 a_15493_43940# a_18525_43370# 1.15e-19
C27817 a_14021_43940# a_15781_43660# 0.00563f
C27818 a_4093_43548# a_4699_43561# 7.24e-19
C27819 a_742_44458# a_1755_42282# 0.013027f
C27820 a_1209_43370# a_n1557_42282# 0.113851f
C27821 a_17973_43940# a_16823_43084# 1.54e-20
C27822 a_10807_43548# a_743_42282# 0.011093f
C27823 a_9313_44734# a_13569_43230# 1.23e-19
C27824 a_2982_43646# VDD 1.40372f
C27825 a_10193_42453# a_n2661_43370# 3.69e-19
C27826 a_15599_45572# a_14537_43396# 3.89e-19
C27827 a_8696_44636# a_13017_45260# 1.73e-20
C27828 a_2711_45572# a_11827_44484# 0.033351f
C27829 a_3357_43084# a_22959_45572# 8.46e-19
C27830 a_22591_45572# a_19963_31679# 0.161955f
C27831 a_19479_31679# a_20447_31679# 0.05179f
C27832 a_17364_32525# a_21076_30879# 0.057544f
C27833 a_18083_42858# a_15227_44166# 2.37e-19
C27834 a_7287_43370# a_526_44458# 5.68e-19
C27835 a_8685_43396# a_10809_44734# 1.08e-21
C27836 a_10341_43396# a_2324_44458# 3.06e-19
C27837 a_13837_43396# a_9290_44172# 0.002072f
C27838 a_5934_30871# a_n1613_43370# 9.62e-19
C27839 a_5742_30871# a_n2312_40392# 9.24e-21
C27840 a_14456_42282# a_12465_44636# 1.36e-21
C27841 a_11962_45724# a_10227_46804# 4.98e-21
C27842 a_8696_44636# a_2063_45854# 0.029184f
C27843 a_n2956_39304# a_n2661_45546# 5.38e-20
C27844 a_n2956_38680# a_n2810_45572# 5.73878f
C27845 a_8049_45260# a_10037_46155# 4.8e-19
C27846 a_743_42282# a_13467_32519# 0.003709f
C27847 a_9145_43396# a_12379_42858# 0.001164f
C27848 a_8685_43396# a_13460_43230# 4.34e-20
C27849 a_3422_30871# a_20712_42282# 0.016384f
C27850 a_4905_42826# a_4743_43172# 2.86e-19
C27851 VDAC_P C0_P_btm 0.901219f
C27852 VDAC_N C0_dummy_N_btm 0.885361f
C27853 a_6540_46812# DATA[3] 1.02e-20
C27854 a_5837_42852# VDD 0.1774f
C27855 en_comp a_n2012_44484# 4.42e-20
C27856 a_7229_43940# a_5343_44458# 0.196399f
C27857 a_n1059_45260# a_n356_44636# 0.07487f
C27858 a_8191_45002# a_4223_44672# 1.76e-20
C27859 a_5205_44484# a_6298_44484# 0.085118f
C27860 a_3232_43370# a_5883_43914# 0.337937f
C27861 a_3905_42558# a_1823_45246# 0.010516f
C27862 a_5111_42852# a_n443_42852# 0.005368f
C27863 a_10922_42852# a_n357_42282# 0.006403f
C27864 a_22223_42860# a_13259_45724# 0.007322f
C27865 a_15599_45572# a_3090_45724# 0.022054f
C27866 a_14495_45572# a_13059_46348# 0.004072f
C27867 a_9482_43914# a_5807_45002# 0.018229f
C27868 a_13348_45260# a_13661_43548# 1.86e-19
C27869 a_11652_45724# a_765_45546# 2.49e-20
C27870 a_15297_45822# a_14976_45028# 2.87e-19
C27871 a_5147_45002# a_n743_46660# 9.05e-20
C27872 a_6171_45002# a_n2293_46634# 2.7e-21
C27873 a_13807_45067# a_10227_46804# 4.48e-20
C27874 a_16922_45042# a_16327_47482# 0.060018f
C27875 a_18587_45118# a_11599_46634# 4.52e-20
C27876 a_18494_42460# a_12861_44030# 0.021479f
C27877 a_19864_35138# VDD 0.332629f
C27878 a_n2433_44484# a_n1151_42308# 1.87e-19
C27879 a_5343_44458# a_n237_47217# 0.001668f
C27880 a_n1352_44484# a_584_46384# 7.22e-22
C27881 a_743_42282# a_6773_42558# 0.001159f
C27882 a_421_43172# a_n784_42308# 5.98e-21
C27883 a_16795_42852# a_16877_43172# 0.003935f
C27884 a_15781_43660# a_15764_42576# 3.57e-20
C27885 a_15681_43442# a_15803_42450# 3.32e-19
C27886 a_4361_42308# a_5421_42558# 7.13e-20
C27887 a_n2860_39072# VDD 0.004184f
C27888 a_4915_47217# a_768_44030# 0.187438f
C27889 a_6151_47436# a_11309_47204# 0.065131f
C27890 a_7227_47204# a_8128_46384# 3.24e-20
C27891 a_9863_47436# a_n881_46662# 0.164043f
C27892 a_n2288_47178# a_n2438_43548# 9.47e-19
C27893 a_n746_45260# a_n2661_46634# 0.037885f
C27894 a_n1741_47186# a_n1925_46634# 0.012189f
C27895 SMPL_ON_P a_n2312_38680# 0.041837f
C27896 a_n2109_47186# a_n743_46660# 0.029623f
C27897 a_20894_47436# a_13507_46334# 0.00122f
C27898 a_18780_47178# a_12465_44636# 4.89e-19
C27899 a_20990_47178# a_21177_47436# 0.159555f
C27900 a_18479_47436# a_22223_47212# 7.85e-20
C27901 a_19386_47436# a_4883_46098# 7.49e-21
C27902 a_16019_45002# a_15682_43940# 0.001434f
C27903 a_n2661_43370# a_5495_43940# 2.51e-21
C27904 a_1307_43914# a_14955_43940# 0.00962f
C27905 a_8975_43940# a_11909_44484# 2.14e-19
C27906 a_6109_44484# a_7640_43914# 0.002099f
C27907 a_11827_44484# a_22485_44484# 0.015798f
C27908 a_19929_45028# a_18579_44172# 6.24e-19
C27909 a_413_45260# a_3052_44056# 4.96e-19
C27910 a_n913_45002# a_8487_44056# 1.53e-20
C27911 a_17531_42308# a_n357_42282# 4.24e-20
C27912 a_21195_42852# RST_Z 4.44e-21
C27913 a_5342_30871# VCM 0.325566f
C27914 a_13556_45296# a_3483_46348# 0.375978f
C27915 a_1307_43914# a_1138_42852# 0.123153f
C27916 a_11967_42832# a_13747_46662# 0.021948f
C27917 a_19615_44636# a_13661_43548# 1.88e-21
C27918 a_7640_43914# a_4646_46812# 0.183308f
C27919 a_5343_44458# a_8270_45546# 1.28e-19
C27920 a_14673_44172# a_n2293_46634# 0.100552f
C27921 a_18450_45144# a_15227_44166# 0.002515f
C27922 a_18588_44850# a_19321_45002# 1.03e-20
C27923 a_16333_45814# a_16375_45002# 0.001746f
C27924 a_16680_45572# a_13259_45724# 0.038605f
C27925 a_18691_45572# a_8049_45260# 0.006525f
C27926 a_6171_45002# a_9625_46129# 4.78e-21
C27927 a_7705_45326# a_7920_46348# 1.67e-19
C27928 a_413_45260# a_15015_46420# 5.92e-21
C27929 a_5205_44484# a_5937_45572# 0.481405f
C27930 a_5111_44636# a_9290_44172# 0.031975f
C27931 a_4921_42308# a_6123_31319# 2.25e-19
C27932 a_1606_42308# a_10723_42308# 3.31e-20
C27933 a_6171_42473# a_6481_42558# 6.01e-20
C27934 CAL_P EN_VIN_BSTR_N 0.049856f
C27935 a_4791_45118# a_1823_45246# 0.015359f
C27936 a_3160_47472# a_3483_46348# 0.154179f
C27937 a_n443_46116# a_1138_42852# 0.017807f
C27938 a_n1151_42308# a_3147_46376# 0.001437f
C27939 a_2905_45572# a_3699_46348# 0.004136f
C27940 a_n237_47217# a_8349_46414# 0.047427f
C27941 a_2063_45854# a_4704_46090# 0.004146f
C27942 a_n971_45724# a_5937_45572# 0.027865f
C27943 a_12549_44172# a_15227_44166# 0.354423f
C27944 a_5807_45002# a_12816_46660# 0.004701f
C27945 a_3877_44458# a_4955_46873# 0.029242f
C27946 a_4646_46812# a_4651_46660# 0.844575f
C27947 a_3524_46660# a_3633_46660# 0.007416f
C27948 a_3699_46634# a_3878_46660# 0.007399f
C27949 a_n1925_46634# a_7832_46660# 0.00149f
C27950 a_13717_47436# a_21076_30879# 5.51e-19
C27951 a_18479_47436# a_20731_47026# 0.004016f
C27952 a_17591_47464# a_17639_46660# 1.72e-19
C27953 a_20894_47436# a_20623_46660# 4.85e-19
C27954 a_20990_47178# a_20841_46902# 1.82e-19
C27955 a_21177_47436# a_20273_46660# 0.003694f
C27956 a_11599_46634# a_11415_45002# 0.007504f
C27957 a_13507_46334# a_20411_46873# 0.035522f
C27958 a_12465_44636# a_18285_46348# 2.07e-20
C27959 a_n2017_45002# a_12089_42308# 0.043278f
C27960 a_n1059_45260# a_12379_42858# 0.003827f
C27961 a_n913_45002# a_10341_42308# 0.070067f
C27962 a_3537_45260# a_3681_42891# 3.51e-19
C27963 a_n2661_42834# a_5025_43940# 1.83e-19
C27964 a_9313_44734# a_10555_43940# 0.001497f
C27965 a_n699_43396# a_2982_43646# 0.004394f
C27966 a_n1331_43914# a_n822_43940# 2.6e-19
C27967 a_1307_43914# a_5649_42852# 2.47e-20
C27968 a_3905_42865# a_5244_44056# 0.002415f
C27969 a_19279_43940# a_17973_43940# 5.98e-20
C27970 a_11967_42832# a_20269_44172# 4.03e-20
C27971 a_19615_44636# a_19862_44208# 8.86e-19
C27972 a_18248_44752# a_n97_42460# 1.22e-20
C27973 a_16922_45042# a_10341_43396# 0.048996f
C27974 a_14539_43914# VDD 0.873589f
C27975 a_n4064_39616# C10_P_btm 7.64e-19
C27976 a_n3420_39616# C8_P_btm 0.090298f
C27977 a_n3565_39304# a_n1386_35608# 8.05e-20
C27978 a_19237_31679# a_21076_30879# 0.05495f
C27979 a_18326_43940# a_3090_45724# 5.94e-19
C27980 a_1756_43548# a_n2438_43548# 2.24e-20
C27981 a_n1557_42282# a_n2442_46660# 2.36e-20
C27982 a_15037_44260# a_6755_46942# 2.99e-20
C27983 a_18184_42460# a_n357_42282# 0.106442f
C27984 a_n23_44458# a_526_44458# 3.73e-19
C27985 a_n356_44636# a_n1925_42282# 0.020589f
C27986 a_7221_43396# a_n1613_43370# 2.95e-19
C27987 a_15743_43084# a_16327_47482# 1.21037f
C27988 a_2905_42968# a_n2497_47436# 7.38e-22
C27989 a_n967_43230# a_n971_45724# 4.78e-20
C27990 a_2107_46812# VDD 0.350275f
C27991 a_n3420_39616# a_n4334_38528# 4.91e-19
C27992 a_n3565_39304# a_n3420_39072# 0.241179f
C27993 a_n4209_39304# a_n4064_39072# 0.19711f
C27994 a_1736_39587# a_1239_39043# 0.036194f
C27995 a_5742_30871# C0_dummy_N_btm 2.87e-19
C27996 a_n4318_38216# a_n3420_37984# 0.001387f
C27997 a_13607_46688# a_3483_46348# 2.14e-20
C27998 a_20107_46660# a_21363_46634# 0.043567f
C27999 a_20273_46660# a_20841_46902# 0.17072f
C28000 a_20411_46873# a_20623_46660# 0.007737f
C28001 a_13747_46662# a_13259_45724# 0.093177f
C28002 a_3524_46660# a_526_44458# 4.66e-19
C28003 a_2107_46812# a_8283_46482# 5.51e-19
C28004 a_n743_46660# a_8062_46155# 1.71e-19
C28005 a_8270_45546# a_8349_46414# 0.002654f
C28006 a_6755_46942# a_12005_46116# 1.39e-19
C28007 a_8667_46634# a_2324_44458# 8.29e-21
C28008 a_n1613_43370# a_n2293_45546# 0.020156f
C28009 a_18579_44172# a_5649_42852# 1.35e-22
C28010 a_n2661_43922# a_9127_43156# 2.21e-20
C28011 a_n2661_42834# a_8952_43230# 9.54e-21
C28012 a_n2293_43922# a_8387_43230# 9.06e-21
C28013 a_9313_44734# a_13113_42826# 0.004011f
C28014 a_1307_43914# a_7963_42308# 3.36e-21
C28015 a_18184_42460# a_18707_42852# 3.84e-20
C28016 a_n1059_45260# a_18727_42674# 0.20226f
C28017 a_n2017_45002# a_18907_42674# 6.48e-20
C28018 a_n913_45002# a_18057_42282# 1.34e-19
C28019 a_20447_31679# a_13258_32519# 0.054935f
C28020 a_2253_43940# VDD 0.156797f
C28021 a_7230_45938# a_6171_45002# 0.001502f
C28022 a_8162_45546# a_3232_43370# 8.68e-20
C28023 a_2711_45572# a_15595_45028# 7.51e-20
C28024 a_17499_43370# a_17339_46660# 1.36e-19
C28025 a_7542_44172# a_n443_42852# 1.35e-21
C28026 a_n2661_42282# a_n863_45724# 1.84e-19
C28027 a_15493_43396# a_16375_45002# 1.46e-20
C28028 a_2537_44260# a_n357_42282# 2.9e-20
C28029 a_n97_42460# a_2324_44458# 5.01e-20
C28030 a_5934_30871# a_4791_45118# 2.81e-20
C28031 a_14493_46090# VDD 0.203567f
C28032 a_7227_45028# a_2063_45854# 0.021063f
C28033 a_6194_45824# a_n1151_42308# 4.58e-20
C28034 a_4099_45572# a_3815_47204# 1.36e-21
C28035 a_1260_45572# a_n443_46116# 0.004853f
C28036 a_n1991_46122# a_n2661_45546# 2.49e-20
C28037 a_n2293_46098# a_n2293_45546# 0.04779f
C28038 a_3483_46348# a_16375_45002# 5.28e-20
C28039 a_n4334_38304# a_n4209_37414# 6.38e-20
C28040 a_n4209_38216# a_n4334_37440# 5.82e-19
C28041 a_9625_46129# a_9751_46155# 0.005702f
C28042 a_10355_46116# a_10586_45546# 0.012906f
C28043 a_12005_46116# a_8049_45260# 0.006548f
C28044 a_1568_43370# a_2905_42968# 5.03e-21
C28045 a_15681_43442# a_16137_43396# 2.85e-19
C28046 a_n3674_39768# a_n3674_38680# 0.035445f
C28047 a_n97_42460# a_8387_43230# 2.28e-20
C28048 a_10341_43396# a_15743_43084# 0.464206f
C28049 a_9396_43370# a_5649_42852# 6.62e-21
C28050 a_453_43940# a_1576_42282# 3.54e-21
C28051 a_1414_42308# a_1184_42692# 0.115223f
C28052 a_12891_46348# CLK 8.04e-20
C28053 en_comp a_7754_40130# 0.011333f
C28054 a_7871_42858# VDD 0.395222f
C28055 a_11823_42460# a_13857_44734# 9.1e-21
C28056 a_10193_42453# a_11909_44484# 3.99e-20
C28057 a_8696_44636# a_18374_44850# 9.12e-20
C28058 a_5691_45260# a_n2661_43370# 0.015295f
C28059 a_7229_43940# a_8560_45348# 1.25e-19
C28060 a_8191_45002# a_n2293_42834# 0.084957f
C28061 a_n913_45002# a_18494_42460# 4.44e-19
C28062 a_22400_42852# a_20202_43084# 3.36e-20
C28063 a_13467_32519# a_20205_31679# 0.051513f
C28064 a_20273_45572# a_13747_46662# 0.002644f
C28065 a_2711_45572# a_15559_46634# 2.74e-20
C28066 a_5263_45724# a_3090_45724# 1.96e-19
C28067 a_2437_43646# a_12549_44172# 0.004577f
C28068 a_n2661_45010# a_n1613_43370# 0.223356f
C28069 a_3537_45260# a_4883_46098# 2.75e-19
C28070 a_n2661_43370# SMPL_ON_P 0.002305f
C28071 a_13777_45326# a_12861_44030# 0.00239f
C28072 a_13159_45002# a_11599_46634# 6.88e-21
C28073 a_8147_43396# a_8515_42308# 6.85e-19
C28074 a_8791_43396# a_5934_30871# 5.94e-19
C28075 a_5342_30871# a_16795_42852# 2.89e-20
C28076 a_3626_43646# a_11323_42473# 0.003176f
C28077 a_2982_43646# a_11551_42558# 1.36e-19
C28078 a_19319_43548# a_20107_42308# 1.44e-20
C28079 a_15567_42826# a_16414_43172# 0.001784f
C28080 a_n97_42460# a_16522_42674# 2.08e-19
C28081 a_167_45260# DATA[1] 1.13e-20
C28082 a_6151_47436# a_7227_47204# 3.14e-19
C28083 a_6545_47178# a_6851_47204# 0.134581f
C28084 a_4915_47217# a_9067_47204# 0.061984f
C28085 a_n237_47217# a_10227_46804# 0.00246f
C28086 a_3785_47178# a_n1435_47204# 5.76e-19
C28087 a_n1151_42308# a_12861_44030# 0.029342f
C28088 a_n913_45002# a_3499_42826# 6.51e-19
C28089 a_3537_45260# a_5663_43940# 1.06e-19
C28090 a_5147_45002# a_5244_44056# 0.122327f
C28091 a_5111_44636# a_3905_42865# 0.006261f
C28092 a_4558_45348# a_5013_44260# 3.95e-20
C28093 a_n2433_44484# a_n1821_44484# 0.001881f
C28094 a_n2129_44697# a_n1190_44850# 3.86e-19
C28095 a_n2267_44484# a_n1809_44850# 0.027606f
C28096 a_5883_43914# a_8975_43940# 0.50976f
C28097 a_n1630_35242# a_n443_42852# 6.01e-19
C28098 a_2903_42308# a_n357_42282# 2.49e-20
C28099 a_2713_42308# a_n755_45592# 0.243663f
C28100 a_12427_45724# VDD 0.33808f
C28101 a_14180_45002# a_14035_46660# 3.28e-19
C28102 a_2437_43646# a_1208_46090# 6.09e-20
C28103 a_8560_45348# a_8270_45546# 4.84e-20
C28104 a_18443_44721# a_19321_45002# 6.29e-21
C28105 a_n2661_45010# a_n2293_46098# 1.61e-19
C28106 a_18989_43940# a_13747_46662# 0.002177f
C28107 a_10490_45724# a_8049_45260# 0.006151f
C28108 a_7499_43078# a_10586_45546# 1.07e-19
C28109 a_8375_44464# a_8128_46384# 3.74e-20
C28110 a_15861_45028# a_17583_46090# 1.62e-19
C28111 a_16680_45572# a_18189_46348# 6.45e-21
C28112 a_8696_44636# a_17715_44484# 0.017149f
C28113 a_14033_45572# a_12594_46348# 9.76e-19
C28114 a_11778_45572# a_10809_44734# 2.41e-19
C28115 a_11967_42832# a_11599_46634# 1.61e-22
C28116 a_20640_44752# a_12861_44030# 0.001266f
C28117 COMP_P a_n784_42308# 0.10915f
C28118 a_n1736_42282# a_n3674_37592# 0.006442f
C28119 a_n961_42308# a_n473_42460# 0.011409f
C28120 a_n2104_42282# a_n1630_35242# 0.030917f
C28121 a_21195_42852# a_17303_42282# 3.32e-20
C28122 a_19339_43156# a_19332_42282# 0.004421f
C28123 a_n2312_38680# a_n2438_43548# 0.046935f
C28124 a_n2661_46634# a_383_46660# 0.007768f
C28125 a_n1925_46634# a_n743_46660# 0.193773f
C28126 a_n1613_43370# a_5732_46660# 0.268372f
C28127 a_4883_46098# a_6969_46634# 1.82e-19
C28128 a_11599_46634# a_12251_46660# 7.45e-20
C28129 a_10227_46804# a_8270_45546# 1.67e-19
C28130 a_13717_47436# a_15009_46634# 9.67e-21
C28131 a_12861_44030# a_14084_46812# 0.003999f
C28132 a_13487_47204# a_13607_46688# 2.07e-19
C28133 a_4915_47217# a_10933_46660# 1.75e-19
C28134 a_n1151_42308# a_14180_46812# 0.037471f
C28135 a_n746_45260# a_765_45546# 0.006723f
C28136 a_9482_43914# a_13667_43396# 1.67e-20
C28137 a_21359_45002# a_20974_43370# 5.16e-21
C28138 a_17970_44736# a_11341_43940# 3.63e-21
C28139 a_16979_44734# a_15493_43940# 6.95e-20
C28140 a_19279_43940# a_22591_44484# 1.13e-20
C28141 a_5891_43370# a_9028_43914# 0.001563f
C28142 a_1307_43914# a_8685_43396# 4.34e-20
C28143 a_n2661_42834# a_n1441_43940# 0.004368f
C28144 a_20679_44626# a_19237_31679# 1.41e-20
C28145 a_7499_43078# a_6101_43172# 3.94e-21
C28146 a_n2661_43922# a_n630_44306# 3.27e-19
C28147 a_19479_31679# a_13467_32519# 0.051245f
C28148 a_n4064_37984# VDD 1.70621f
C28149 a_14309_45028# VDD 0.189806f
C28150 a_13565_43940# a_12891_46348# 0.001515f
C28151 a_3422_30871# a_19692_46634# 0.208985f
C28152 a_14761_44260# a_n2293_46634# 0.009374f
C28153 a_18204_44850# a_17339_46660# 1.39e-19
C28154 a_375_42282# a_n2661_45546# 0.001753f
C28155 a_5205_44484# a_n443_42852# 6.5e-20
C28156 a_742_44458# a_2324_44458# 0.00317f
C28157 a_7221_43396# a_4791_45118# 2.22e-20
C28158 a_13258_32519# a_21887_42336# 8.1e-19
C28159 a_20712_42282# a_7174_31319# 3.53e-19
C28160 a_11453_44696# VDD 3.75355f
C28161 a_14097_32519# C4_N_btm 0.030945f
C28162 a_n971_45724# a_n443_42852# 0.329303f
C28163 a_2063_45854# a_2957_45546# 0.002513f
C28164 a_2905_45572# a_n755_45592# 0.168143f
C28165 a_n746_45260# a_509_45822# 4.34e-21
C28166 a_n1151_42308# a_310_45028# 2.08e-20
C28167 a_2959_46660# a_2804_46116# 2.23e-19
C28168 a_2609_46660# a_3483_46348# 0.010427f
C28169 a_3177_46902# a_3147_46376# 0.003463f
C28170 a_14084_46812# a_14180_46812# 0.318161f
C28171 a_3090_45724# a_13885_46660# 1.72e-19
C28172 a_11599_46634# a_13259_45724# 0.249721f
C28173 a_10227_46804# a_12638_46436# 3.98e-20
C28174 a_4883_46098# a_9241_46436# 7.71e-20
C28175 a_n1613_43370# a_n914_46116# 1.68e-19
C28176 a_16119_47582# a_6945_45028# 2.34e-19
C28177 a_768_44030# a_10809_44734# 0.037504f
C28178 a_n2293_46634# a_10903_43370# 0.046902f
C28179 a_2107_46812# a_7920_46348# 0.006995f
C28180 a_n743_46660# a_10355_46116# 0.011802f
C28181 a_13747_46662# a_18189_46348# 0.022348f
C28182 a_5807_45002# a_18819_46122# 0.012467f
C28183 a_n881_46662# a_739_46482# 3.69e-19
C28184 a_n1059_45260# a_3823_42558# 2.04e-20
C28185 a_n913_45002# a_3318_42354# 0.03912f
C28186 a_n2017_45002# a_5267_42460# 0.003851f
C28187 a_2998_44172# a_3080_42308# 6.67e-19
C28188 a_1467_44172# a_2982_43646# 8.78e-21
C28189 a_18184_42460# a_21356_42826# 0.016504f
C28190 a_9313_44734# a_16823_43084# 0.031008f
C28191 a_5343_44458# a_5755_42852# 5.25e-22
C28192 a_5518_44484# a_5111_42852# 2.49e-21
C28193 a_4223_44672# a_7765_42852# 2.94e-20
C28194 a_11967_42832# a_14358_43442# 8.52e-20
C28195 a_3905_42865# a_4235_43370# 0.041971f
C28196 a_1414_42308# a_2896_43646# 0.005191f
C28197 a_n2293_42834# a_7309_42852# 4.09e-20
C28198 a_n3674_39768# VDD 0.398971f
C28199 a_14495_45572# a_8696_44636# 3.04e-20
C28200 a_11682_45822# a_12016_45572# 2.43e-19
C28201 a_12427_45724# a_12749_45572# 0.001367f
C28202 a_11962_45724# a_13297_45572# 0.001004f
C28203 a_11823_42460# a_12649_45572# 5.54e-19
C28204 a_13460_43230# a_768_44030# 6.38e-21
C28205 a_3681_42891# a_n2293_46634# 1.32e-20
C28206 a_16547_43609# a_6755_46942# 7.51e-20
C28207 a_22315_44484# a_20205_31679# 2.01e-21
C28208 a_11816_44260# a_10903_43370# 8.18e-19
C28209 COMP_P SMPL_ON_P 0.03194f
C28210 a_17639_46660# VDD 0.001662f
C28211 a_n1991_46122# a_n1533_46116# 0.034619f
C28212 a_n2293_46098# a_n914_46116# 1.25e-19
C28213 a_19692_46634# a_21167_46155# 0.005265f
C28214 a_13059_46348# a_15194_46482# 6.53e-22
C28215 a_10355_46116# a_11189_46129# 0.001778f
C28216 a_5204_45822# a_2324_44458# 2.51e-21
C28217 a_9625_46129# a_10903_43370# 1.41e-19
C28218 a_9396_43370# a_8685_43396# 0.007917f
C28219 a_n97_42460# a_15743_43084# 0.205305f
C28220 a_13483_43940# a_13460_43230# 2.1e-20
C28221 a_n2293_43922# a_1606_42308# 0.080878f
C28222 a_20193_45348# a_21887_42336# 0.169001f
C28223 a_12861_44030# START 0.006864f
C28224 a_9863_47436# DATA[4] 7.9e-19
C28225 a_13487_47204# RST_Z 0.07884f
C28226 a_13717_47436# SINGLE_ENDED 0.032092f
C28227 a_n1435_47204# CLK_DATA 8.83e-21
C28228 a_17324_43396# VDD 0.274722f
C28229 a_4558_45348# a_4927_45028# 0.123258f
C28230 a_3537_45260# a_3232_43370# 0.530258f
C28231 a_5147_45002# a_5111_44636# 0.562127f
C28232 a_n2017_45002# a_14537_43396# 3.09e-22
C28233 a_7499_43078# a_10440_44484# 3.35e-19
C28234 a_9049_44484# a_10334_44484# 2.09e-20
C28235 a_10053_45546# a_10157_44484# 1.49e-20
C28236 a_8696_44636# a_17719_45144# 3.25e-19
C28237 a_8746_45002# a_8701_44490# 1.65e-19
C28238 a_15861_45028# a_17613_45144# 0.016666f
C28239 a_10835_43094# a_4185_45028# 1.34e-20
C28240 a_19511_42282# a_12549_44172# 5.57e-20
C28241 a_5932_42308# a_4646_46812# 2.43e-19
C28242 a_14358_43442# a_13259_45724# 1.56e-20
C28243 a_6293_42852# a_n357_42282# 0.00795f
C28244 a_6031_43396# a_n755_45592# 2.22e-20
C28245 a_1427_43646# a_n443_42852# 0.002947f
C28246 a_n4064_39616# a_n2312_40392# 9.29e-20
C28247 a_n2946_39866# a_n2312_39304# 2.85e-20
C28248 a_3422_30871# VIN_N 0.057975f
C28249 a_15143_45578# a_13747_46662# 0.040557f
C28250 a_7499_43078# a_n743_46660# 1.36e-19
C28251 a_8746_45002# a_n2293_46634# 3.85e-20
C28252 a_11525_45546# a_n2661_46634# 0.003942f
C28253 a_6469_45572# a_5807_45002# 4.31e-19
C28254 a_20273_45572# a_11599_46634# 0.004992f
C28255 a_18909_45814# a_18597_46090# 8.56e-20
C28256 a_18691_45572# a_18780_47178# 1.83e-20
C28257 a_17668_45572# a_16327_47482# 0.003454f
C28258 a_3357_43084# a_6851_47204# 2.62e-19
C28259 a_2437_43646# a_6575_47204# 0.029543f
C28260 a_2274_45254# a_n237_47217# 3.92e-19
C28261 a_n913_45002# a_n1151_42308# 0.395136f
C28262 a_2680_45002# a_n971_45724# 0.108251f
C28263 a_5111_44636# a_n2109_47186# 0.017519f
C28264 a_n1557_42282# a_n3674_38216# 1.82e-19
C28265 a_3080_42308# COMP_P 4.43551f
C28266 a_4361_42308# a_5534_30871# 0.049795f
C28267 a_15493_43396# a_17303_42282# 1.81e-21
C28268 a_n97_42460# a_1606_42308# 1.2e-19
C28269 a_458_43396# a_564_42282# 1.51e-20
C28270 a_4190_30871# a_17701_42308# 0.008836f
C28271 a_743_42282# a_16795_42852# 1.32e-20
C28272 a_5649_42852# a_13635_43156# 6.61e-20
C28273 a_1568_43370# a_n784_42308# 8.96e-20
C28274 a_14513_46634# RST_Z 1.53e-20
C28275 a_7754_38968# a_3754_38470# 0.209356f
C28276 a_1184_42692# VDD 0.813074f
C28277 a_n2288_47178# a_n1741_47186# 0.001294f
C28278 a_n2109_47186# a_n1920_47178# 0.070142f
C28279 a_n2497_47436# SMPL_ON_P 0.131317f
C28280 a_10951_45334# a_n2661_43922# 4.26e-20
C28281 a_n2661_43370# a_10057_43914# 2.24e-19
C28282 a_1423_45028# a_6109_44484# 0.018788f
C28283 a_21359_45002# a_18114_32519# 2.21e-19
C28284 a_11827_44484# a_20205_45028# 5.4e-19
C28285 a_3232_43370# a_11541_44484# 0.050289f
C28286 a_19479_31679# a_22315_44484# 7.36e-19
C28287 a_3357_43084# a_3422_30871# 1.8e-20
C28288 en_comp a_11967_42832# 5.02e-20
C28289 a_5267_42460# a_526_44458# 3.04e-19
C28290 a_3823_42558# a_n1925_42282# 0.010285f
C28291 a_11554_42852# a_n357_42282# 0.001921f
C28292 a_13249_42558# a_10903_43370# 0.003601f
C28293 a_9885_42308# a_8199_44636# 0.001301f
C28294 a_15765_45572# a_12741_44636# 4.82e-19
C28295 a_16855_45546# a_11415_45002# 0.004485f
C28296 a_1423_45028# a_4646_46812# 0.415897f
C28297 a_18909_45814# a_19123_46287# 5.82e-19
C28298 a_11691_44458# a_12891_46348# 0.141379f
C28299 a_n2661_43370# a_n2438_43548# 0.147387f
C28300 a_18315_45260# a_13747_46662# 1.26e-20
C28301 a_18587_45118# a_13661_43548# 0.087703f
C28302 a_18911_45144# a_5807_45002# 2.35e-20
C28303 a_18596_45572# a_17339_46660# 0.009893f
C28304 a_6171_45002# a_6755_46942# 0.026424f
C28305 a_n2017_45002# a_3090_45724# 2.3e-19
C28306 a_19963_31679# a_19692_46634# 1.27e-19
C28307 a_7499_43078# a_11189_46129# 5.71e-20
C28308 a_10053_45546# a_10355_46116# 1.96e-19
C28309 a_10180_45724# a_9823_46155# 0.002058f
C28310 a_9049_44484# a_9290_44172# 1.37e-20
C28311 a_8746_45002# a_9625_46129# 4.27e-19
C28312 a_556_44484# a_n1151_42308# 9.41e-20
C28313 a_8855_44734# a_4791_45118# 3.24e-21
C28314 a_18989_43940# a_11599_46634# 7.89e-20
C28315 a_17970_44736# a_16327_47482# 0.219775f
C28316 a_15004_44636# a_10227_46804# 0.003988f
C28317 a_20205_31679# VCM 0.035399f
C28318 a_20692_30879# VREF_GND 0.010456f
C28319 a_n357_42282# RST_Z 2.38e-20
C28320 a_743_42282# a_21335_42336# 2.86e-19
C28321 a_n2293_42282# a_2123_42473# 1.62e-19
C28322 a_10341_42308# a_8325_42308# 1.07e-20
C28323 a_4361_42308# a_19647_42308# 0.007305f
C28324 a_13467_32519# a_13258_32519# 11.0084f
C28325 a_14635_42282# a_14853_42852# 0.01129f
C28326 a_n237_47217# a_10467_46802# 2.29e-19
C28327 a_2063_45854# a_7715_46873# 0.178294f
C28328 a_4791_45118# a_5732_46660# 4.55e-19
C28329 a_6851_47204# a_3877_44458# 8.01e-20
C28330 a_5129_47502# a_5385_46902# 0.001505f
C28331 a_n1435_47204# a_3699_46634# 5.5e-20
C28332 a_5815_47464# a_4817_46660# 0.00304f
C28333 a_6491_46660# a_4646_46812# 0.042695f
C28334 a_4883_46098# a_n2293_46634# 0.046481f
C28335 a_11453_44696# a_22612_30879# 0.005655f
C28336 a_22959_47212# a_21588_30879# 0.018188f
C28337 a_9804_47204# a_10037_47542# 5.76e-19
C28338 a_n881_46662# a_768_44030# 0.057002f
C28339 C0_P_btm VDD 1.02806f
C28340 a_3357_43084# a_5565_43396# 0.009914f
C28341 a_n913_45002# a_6197_43396# 2.11e-20
C28342 a_n2017_45002# a_6547_43396# 4.02e-20
C28343 a_4574_45260# a_3080_42308# 5.32e-21
C28344 a_3537_45260# a_4905_42826# 0.339989f
C28345 a_19778_44110# a_15493_43396# 0.015561f
C28346 a_18184_42460# a_19328_44172# 1.54e-19
C28347 a_11827_44484# a_15682_43940# 0.006752f
C28348 a_5343_44458# a_7845_44172# 0.103601f
C28349 a_5883_43914# a_5495_43940# 0.09813f
C28350 a_n1809_44850# a_n2065_43946# 8.2e-20
C28351 a_9313_44734# a_19279_43940# 3.78e-20
C28352 a_11691_44458# a_11750_44172# 5.84e-19
C28353 a_6298_44484# a_7281_43914# 0.010383f
C28354 a_n3565_38216# a_n2956_38216# 0.307285f
C28355 a_6709_45028# VDD 0.390566f
C28356 a_n1630_35242# CAL_P 0.016538f
C28357 COMP_P a_n1532_35090# 4.87e-20
C28358 a_18287_44626# a_16388_46812# 4.61e-22
C28359 a_14673_44172# a_6755_46942# 0.050772f
C28360 a_5663_43940# a_n2293_46634# 5.03e-20
C28361 a_7911_44260# a_768_44030# 0.001075f
C28362 a_22959_45572# a_20205_31679# 0.002292f
C28363 a_6171_45002# a_8049_45260# 0.048422f
C28364 en_comp a_13259_45724# 0.19355f
C28365 a_19963_31679# a_20692_30879# 0.051965f
C28366 a_2437_43646# a_n2661_45546# 0.028152f
C28367 a_6945_45348# a_2324_44458# 4.69e-19
C28368 a_n229_43646# a_n971_45724# 0.059197f
C28369 a_n1177_43370# a_584_46384# 2.93e-20
C28370 a_3080_42308# a_n2497_47436# 2.97e-19
C28371 a_n23_47502# VDD 0.152616f
C28372 a_11551_42558# a_11897_42308# 0.013377f
C28373 a_n4318_37592# a_n4064_39072# 0.019896f
C28374 a_6171_42473# a_7174_31319# 4.88e-21
C28375 a_14113_42308# a_15486_42560# 0.039784f
C28376 VIN_P VCM 1.7189f
C28377 VIN_N VREF_GND 16.4969f
C28378 a_13661_43548# a_11415_45002# 0.107787f
C28379 a_13747_46662# a_20202_43084# 0.308003f
C28380 a_383_46660# a_765_45546# 1.21e-19
C28381 a_10467_46802# a_8270_45546# 3.96e-20
C28382 a_6755_46942# a_6903_46660# 0.003896f
C28383 a_10428_46928# a_10384_47026# 1.46e-19
C28384 a_n881_46662# a_1176_45822# 0.048496f
C28385 a_n1613_43370# a_1138_42852# 1.35e-19
C28386 a_4883_46098# a_9625_46129# 0.164961f
C28387 a_11599_46634# a_18189_46348# 0.101491f
C28388 a_16327_47482# a_14840_46494# 6.83e-21
C28389 a_10227_46804# a_13759_46122# 0.920747f
C28390 a_15673_47210# a_15682_46116# 6.62e-20
C28391 a_13717_47436# a_19335_46494# 1.62e-21
C28392 a_11031_47542# a_6945_45028# 0.007285f
C28393 a_n237_47217# a_8034_45724# 0.0717f
C28394 a_3785_47178# a_526_44458# 2.7e-22
C28395 a_19279_43940# a_20974_43370# 2.3e-20
C28396 a_1414_42308# a_1443_43940# 0.018064f
C28397 a_10405_44172# a_10729_43914# 0.083277f
C28398 a_18579_44172# a_19741_43940# 0.005651f
C28399 a_n2293_42834# a_7765_42852# 0.010796f
C28400 a_n2293_43922# a_3539_42460# 6.26e-20
C28401 a_11823_42460# a_5742_30871# 9.73e-19
C28402 a_20193_45348# a_13467_32519# 0.016015f
C28403 a_453_43940# a_1241_43940# 0.002487f
C28404 a_9672_43914# a_10949_43914# 2.19e-20
C28405 a_5111_44636# a_5457_43172# 0.002744f
C28406 a_n1059_45260# a_12800_43218# 0.002165f
C28407 a_n913_45002# a_10752_42852# 6.19e-19
C28408 a_3537_45260# a_7573_43172# 1e-19
C28409 a_6511_45714# a_6469_45572# 2.56e-19
C28410 a_2711_45572# a_10907_45822# 0.016608f
C28411 a_19862_44208# a_11415_45002# 1.39e-19
C28412 a_20269_44172# a_20202_43084# 9.29e-21
C28413 a_21259_43561# a_12549_44172# 0.001855f
C28414 a_16243_43396# a_n2293_46634# 1.28e-22
C28415 a_n356_44636# a_380_45546# 5.74e-21
C28416 a_14673_44172# a_8049_45260# 8.94e-21
C28417 a_n310_44811# a_n863_45724# 5.09e-19
C28418 a_13076_44458# a_n443_42852# 4.94e-19
C28419 a_7281_43914# a_5937_45572# 9.58e-19
C28420 a_5649_42852# a_n1613_43370# 2.17e-20
C28421 a_19479_31679# VCM 0.03628f
C28422 a_19963_31679# VIN_N 0.029022f
C28423 a_10384_47026# VDD 4.6e-19
C28424 a_n1630_35242# CAL_N 1.66e-19
C28425 a_n1423_46090# a_472_46348# 3.09e-21
C28426 a_n2293_46098# a_1138_42852# 0.029886f
C28427 a_n901_46420# a_n1076_46494# 0.234322f
C28428 a_11415_45002# a_4185_45028# 5.21e-19
C28429 a_16388_46812# a_15682_46116# 0.044769f
C28430 a_765_45546# a_13351_46090# 9.37e-21
C28431 a_1799_45572# a_1848_45724# 0.080562f
C28432 a_2443_46660# a_n755_45592# 5.37e-20
C28433 a_3090_45724# a_526_44458# 0.058033f
C28434 a_n2661_46098# a_997_45618# 4.98e-22
C28435 a_8270_45546# a_8034_45724# 0.031124f
C28436 a_n2956_37592# a_n4064_38528# 0.015398f
C28437 a_n2810_45028# a_n2302_38778# 4.97e-19
C28438 a_n3674_39768# a_n4318_38680# 0.024755f
C28439 a_n97_42460# a_3539_42460# 0.021726f
C28440 a_3422_30871# a_5342_30871# 0.026613f
C28441 a_n699_43396# a_1184_42692# 5.3e-21
C28442 a_11341_43940# a_18783_43370# 3.91e-20
C28443 a_15493_43940# a_18429_43548# 4.75e-20
C28444 a_14021_43940# a_15681_43442# 0.004196f
C28445 a_742_44458# a_1606_42308# 0.001459f
C28446 a_458_43396# a_n1557_42282# 0.027865f
C28447 a_4093_43548# a_4235_43370# 0.515101f
C28448 a_17737_43940# a_16823_43084# 1.26e-20
C28449 a_21115_43940# a_15743_43084# 3.08e-21
C28450 a_2889_44172# a_2905_42968# 5.52e-20
C28451 w_1575_34946# a_n83_35174# 0.001523f
C28452 a_2896_43646# VDD 0.208317f
C28453 a_8696_44636# a_11963_45334# 5.44e-20
C28454 a_10180_45724# a_n2661_43370# 0.038795f
C28455 a_3357_43084# a_19963_31679# 0.009628f
C28456 a_19479_31679# a_22959_45572# 0.004153f
C28457 a_22223_45572# a_20447_31679# 2.46e-19
C28458 a_21513_45002# a_21542_45572# 5.31e-19
C28459 a_19164_43230# a_3090_45724# 4.01e-21
C28460 a_17701_42308# a_15227_44166# 0.172697f
C28461 a_n3674_37592# a_n2442_46660# 0.032368f
C28462 a_7499_43940# a_n357_42282# 8.54e-20
C28463 a_13749_43396# a_9290_44172# 0.00194f
C28464 a_7963_42308# a_n1613_43370# 5.32e-20
C28465 a_n4209_39304# SMPL_ON_P 0.001361f
C28466 a_5891_43370# CLK 8.38e-19
C28467 a_14180_46482# VDD 0.077608f
C28468 a_11652_45724# a_10227_46804# 2.55e-20
C28469 a_15143_45578# a_11599_46634# 0.028879f
C28470 a_n2956_38680# a_n2840_45546# 2.65e-20
C28471 a_n2956_39304# a_n2810_45572# 0.043323f
C28472 a_8049_45260# a_9751_46155# 4.35e-19
C28473 a_2324_44458# a_3503_45724# 9.33e-22
C28474 a_4190_30871# a_4361_42308# 0.06171f
C28475 a_10695_43548# a_10991_42826# 8.2e-19
C28476 a_8685_43396# a_13635_43156# 3.19e-19
C28477 a_3422_30871# a_20107_42308# 3.36e-19
C28478 a_4905_42826# a_4649_43172# 9.93e-20
C28479 VDAC_P C1_P_btm 1.74268f
C28480 a_5193_42852# VDD 0.187605f
C28481 a_n2017_45002# a_n356_44636# 0.036195f
C28482 a_5111_44636# a_10157_44484# 2.31e-20
C28483 a_3537_45260# a_8975_43940# 7.28e-19
C28484 a_5691_45260# a_5883_43914# 3.05e-21
C28485 a_5205_44484# a_5518_44484# 0.135771f
C28486 a_3232_43370# a_8701_44490# 0.062297f
C28487 a_6171_45002# a_8103_44636# 1.07e-20
C28488 a_6431_45366# a_6298_44484# 0.006936f
C28489 a_16855_45546# a_11967_42832# 1.82e-21
C28490 a_4520_42826# a_n443_42852# 5.33e-20
C28491 a_10991_42826# a_n357_42282# 0.005156f
C28492 a_22165_42308# a_13259_45724# 0.001551f
C28493 a_13249_42308# a_13059_46348# 0.306398f
C28494 a_1307_43914# a_768_44030# 1.13357f
C28495 a_13348_45260# a_5807_45002# 9.82e-22
C28496 a_16751_45260# a_12549_44172# 6.99e-22
C28497 a_15225_45822# a_14976_45028# 5.88e-19
C28498 a_15297_45822# a_3090_45724# 8.48e-19
C28499 a_2437_43646# a_5385_46902# 7.1e-20
C28500 a_3357_43084# a_4651_46660# 0.004361f
C28501 a_n37_45144# a_288_46660# 1e-20
C28502 a_5205_44484# a_n2661_46634# 1.71e-21
C28503 a_3232_43370# a_n2293_46634# 0.046281f
C28504 a_5111_44636# a_n1925_46634# 2.77e-20
C28505 a_13490_45067# a_10227_46804# 6.94e-20
C28506 a_18315_45260# a_11599_46634# 2.46e-20
C28507 a_16501_45348# a_16327_47482# 5.1e-19
C28508 a_18184_42460# a_12861_44030# 0.266953f
C28509 a_19120_35138# VDD 0.318963f
C28510 a_n2661_44458# a_n1151_42308# 0.030695f
C28511 a_4743_44484# a_n237_47217# 1.26e-21
C28512 a_743_42282# a_6481_42558# 0.001159f
C28513 a_3080_42308# a_n4209_39304# 4.02e-21
C28514 a_5534_30871# a_13622_42852# 2.49e-19
C28515 a_14543_43071# a_14853_42852# 6.01e-20
C28516 a_15681_43442# a_15764_42576# 4.17e-19
C28517 comp_n VDD 0.504719f
C28518 a_4915_47217# a_12549_44172# 0.316329f
C28519 a_9067_47204# a_n881_46662# 0.073421f
C28520 a_6575_47204# a_7989_47542# 6.62e-20
C28521 a_n443_46116# a_768_44030# 0.177051f
C28522 a_n2497_47436# a_n2438_43548# 0.206216f
C28523 a_n2109_47186# a_n1021_46688# 1.8e-21
C28524 SMPL_ON_P a_n2104_46634# 3.11e-20
C28525 a_n1920_47178# a_n1925_46634# 0.013665f
C28526 a_n971_45724# a_n2661_46634# 0.190714f
C28527 a_18479_47436# a_12465_44636# 7.24e-19
C28528 a_19787_47423# a_13507_46334# 5.57e-21
C28529 a_18597_46090# a_4883_46098# 0.084375f
C28530 a_15004_44636# a_14815_43914# 0.078606f
C28531 a_9482_43914# a_15493_43396# 3.87e-21
C28532 a_18114_32519# a_19279_43940# 3.43e-19
C28533 a_n2661_43370# a_5013_44260# 3.07e-21
C28534 a_1307_43914# a_13483_43940# 0.00928f
C28535 a_11827_44484# a_20512_43084# 0.030456f
C28536 a_8975_43940# a_11541_44484# 0.028558f
C28537 a_2711_45572# a_16823_43084# 1.31e-19
C28538 a_20193_45348# a_22315_44484# 0.002679f
C28539 a_n2293_42834# a_n1644_44306# 5.64e-19
C28540 a_3232_43370# a_11816_44260# 3.27e-19
C28541 a_17303_42282# a_n357_42282# 4.34e-19
C28542 a_18799_45938# VDD 0.132317f
C28543 a_5342_30871# VREF_GND 0.055227f
C28544 a_21356_42826# RST_Z 4.49e-21
C28545 a_9482_43914# a_3483_46348# 0.130172f
C28546 a_11967_42832# a_13661_43548# 0.165876f
C28547 a_19615_44636# a_5807_45002# 0.003455f
C28548 a_6109_44484# a_4646_46812# 0.010238f
C28549 a_17969_45144# a_15227_44166# 5.42e-19
C28550 a_15765_45572# a_16375_45002# 2.15e-19
C28551 a_16855_45546# a_13259_45724# 0.067694f
C28552 a_18909_45814# a_8049_45260# 0.006015f
C28553 a_6171_45002# a_8953_45546# 0.0298f
C28554 a_6431_45366# a_5937_45572# 0.129839f
C28555 a_5205_44484# a_8199_44636# 1.08e-20
C28556 a_961_42354# a_5742_30871# 1.96e-20
C28557 a_4921_42308# a_7227_42308# 1.41e-19
C28558 a_6171_42473# a_5932_42308# 0.224949f
C28559 a_1606_42308# a_10533_42308# 1.94e-20
C28560 a_17364_32525# C10_N_btm 1.08e-19
C28561 CAL_P a_11530_34132# 0.055606f
C28562 a_n443_46116# a_1176_45822# 0.092452f
C28563 a_3160_47472# a_3147_46376# 0.208295f
C28564 a_4700_47436# a_1823_45246# 1.11e-20
C28565 a_2905_45572# a_3483_46348# 0.024106f
C28566 a_n1741_47186# a_9823_46155# 1.05e-20
C28567 a_n971_45724# a_8199_44636# 0.247183f
C28568 a_n237_47217# a_8016_46348# 0.017823f
C28569 a_2063_45854# a_4419_46090# 0.025095f
C28570 a_12861_44030# a_12741_44636# 0.366155f
C28571 a_20894_47436# a_20841_46902# 2.44e-19
C28572 a_20990_47178# a_20273_46660# 1.7e-19
C28573 a_13507_46334# a_20107_46660# 0.031344f
C28574 a_4883_46098# a_19123_46287# 0.022559f
C28575 a_9804_47204# a_10185_46660# 4.55e-19
C28576 a_n1925_46634# a_6086_46660# 2.66e-19
C28577 a_3877_44458# a_4651_46660# 0.032518f
C28578 a_12549_44172# a_18834_46812# 0.01219f
C28579 a_5807_45002# a_12991_46634# 0.006904f
C28580 a_n2017_45002# a_12379_42858# 2.94e-19
C28581 a_n1059_45260# a_10341_42308# 0.032786f
C28582 a_n913_45002# a_10922_42852# 0.01889f
C28583 a_3065_45002# a_3935_42891# 0.01149f
C28584 a_n2661_42834# a_3992_43940# 3.11e-20
C28585 a_n699_43396# a_2896_43646# 0.00787f
C28586 a_2998_44172# a_5013_44260# 0.004647f
C28587 a_n1899_43946# a_n822_43940# 1.46e-19
C28588 a_n1549_44318# a_n1441_43940# 0.057222f
C28589 a_n809_44244# a_n630_44306# 0.007399f
C28590 a_n984_44318# a_n875_44318# 0.007416f
C28591 a_n2661_44458# a_6197_43396# 1.22e-20
C28592 a_11967_42832# a_19862_44208# 3.19e-19
C28593 a_19615_44636# a_19478_44306# 0.004687f
C28594 a_16112_44458# VDD 0.182397f
C28595 a_n3420_39616# C9_P_btm 7.08e-19
C28596 a_n4209_39590# C5_P_btm 5.07e-20
C28597 a_n3565_39590# C7_P_btm 0.00198f
C28598 a_n3565_39304# a_n1838_35608# 1.81e-19
C28599 a_n4209_39304# a_n1532_35090# 1.52e-19
C28600 a_13258_32519# VCM 0.033198f
C28601 a_7174_31319# VIN_N 0.022822f
C28602 a_11967_42832# a_4185_45028# 2.11e-19
C28603 a_5829_43940# a_5257_43370# 0.003839f
C28604 a_9396_43370# a_768_44030# 0.010156f
C28605 a_18079_43940# a_3090_45724# 8.6e-20
C28606 a_1568_43370# a_n2438_43548# 4.4e-21
C28607 a_4905_42826# a_n2293_46634# 0.024749f
C28608 a_14761_44260# a_6755_46942# 2.19e-20
C28609 a_12607_44458# a_8049_45260# 7.47e-21
C28610 a_n356_44636# a_526_44458# 0.142971f
C28611 a_14815_43914# a_13759_46122# 1.02e-21
C28612 a_n2661_43922# a_2324_44458# 0.088002f
C28613 a_8685_43396# a_n1613_43370# 0.016726f
C28614 a_18783_43370# a_16327_47482# 0.026485f
C28615 a_5649_42852# a_4791_45118# 0.075725f
C28616 a_11064_45572# CLK 6.18e-19
C28617 a_948_46660# VDD 0.278482f
C28618 a_n3565_39590# a_n3565_38502# 0.031189f
C28619 a_n3420_39616# a_n4209_38502# 0.028008f
C28620 a_n4209_39590# a_n3420_38528# 0.032196f
C28621 a_n4209_39304# a_n2946_39072# 0.022779f
C28622 a_n4334_39392# a_n3420_39072# 0.004849f
C28623 a_n3565_39304# a_n3690_39392# 0.247167f
C28624 a_1239_39587# a_1239_39043# 0.054961f
C28625 a_5742_30871# C0_dummy_P_btm 2.87e-19
C28626 a_n4318_38216# a_n3690_38304# 7.76e-19
C28627 a_12816_46660# a_3483_46348# 8.76e-22
C28628 a_20107_46660# a_20623_46660# 0.105914f
C28629 a_13661_43548# a_13259_45724# 0.250875f
C28630 a_13747_46662# a_14383_46116# 2.43e-19
C28631 a_3699_46634# a_526_44458# 1.66e-21
C28632 a_n1925_46634# a_8379_46155# 2.63e-19
C28633 a_n2661_46634# a_12005_46436# 8.72e-20
C28634 a_2107_46812# a_8062_46482# 2.73e-19
C28635 a_8270_45546# a_8016_46348# 0.036831f
C28636 a_6755_46942# a_10903_43370# 1.97e-19
C28637 a_5732_46660# a_6945_45028# 1.4e-20
C28638 a_12465_44636# a_n443_42852# 1.42e-19
C28639 a_4743_44484# a_4649_42852# 5.95e-21
C28640 a_15493_43940# a_2982_43646# 6.34e-20
C28641 a_n2661_42834# a_9127_43156# 3.28e-20
C28642 a_n2661_43922# a_8387_43230# 4.36e-21
C28643 a_9313_44734# a_12545_42858# 0.005689f
C28644 a_n2293_43922# a_8605_42826# 7.25e-21
C28645 a_n2293_42834# a_961_42354# 2.18e-20
C28646 a_11341_43940# a_3626_43646# 1.01e-21
C28647 a_3422_30871# a_743_42282# 5.66e-19
C28648 a_n1059_45260# a_18057_42282# 0.141112f
C28649 a_n2017_45002# a_18727_42674# 8.71e-20
C28650 a_n913_45002# a_17531_42308# 2.07e-19
C28651 a_1443_43940# VDD 0.144342f
C28652 a_7499_43078# a_5111_44636# 0.753731f
C28653 a_2711_45572# a_15415_45028# 7.81e-20
C28654 a_6031_43396# a_3483_46348# 5.46e-22
C28655 a_14579_43548# a_11415_45002# 4.66e-21
C28656 a_21487_43396# a_19692_46634# 0.016698f
C28657 a_4361_42308# a_15227_44166# 2.26e-19
C28658 a_16759_43396# a_17339_46660# 7.48e-21
C28659 a_19862_44208# a_13259_45724# 1.06e-20
C28660 a_2253_44260# a_n357_42282# 1.12e-19
C28661 COMP_P a_13507_46334# 2.67e-20
C28662 a_13925_46122# VDD 0.251868f
C28663 a_6598_45938# a_2063_45854# 0.018518f
C28664 a_5907_45546# a_n1151_42308# 6.31e-20
C28665 a_2711_45572# a_4007_47204# 9.84e-20
C28666 a_1176_45572# a_n443_46116# 0.003318f
C28667 a_n4209_38216# a_n4209_37414# 0.041723f
C28668 a_10903_43370# a_8049_45260# 0.114138f
C28669 a_n1853_46287# a_n2661_45546# 0.004849f
C28670 a_n2293_46098# a_n2956_38216# 0.003979f
C28671 a_4185_45028# a_13259_45724# 0.194989f
C28672 a_n2472_46090# a_n2293_45546# 3.06e-19
C28673 a_n4318_39768# a_n3674_38680# 0.027425f
C28674 a_9313_44734# a_19332_42282# 2.91e-20
C28675 a_1414_42308# a_1576_42282# 0.004774f
C28676 a_n97_42460# a_8605_42826# 2.01e-20
C28677 a_1756_43548# a_1847_42826# 4.29e-19
C28678 a_10341_43396# a_18783_43370# 0.010939f
C28679 a_8791_43396# a_5649_42852# 4.06e-22
C28680 a_1568_43370# a_2075_43172# 0.006043f
C28681 a_1115_44172# a_961_42354# 4.94e-20
C28682 a_11309_47204# CLK 0.01087f
C28683 a_12549_44172# DATA[5] 3.42e-20
C28684 a_7227_42852# VDD 0.254613f
C28685 a_10193_42453# a_11541_44484# 6.17e-19
C28686 a_2711_45572# a_19279_43940# 0.001969f
C28687 a_10210_45822# a_9313_44734# 7.56e-21
C28688 a_8696_44636# a_18443_44721# 5.52e-20
C28689 a_4927_45028# a_n2661_43370# 0.007616f
C28690 a_n1059_45260# a_18494_42460# 0.187733f
C28691 a_n913_45002# a_18184_42460# 3.93e-19
C28692 a_7705_45326# a_n2293_42834# 0.071732f
C28693 a_3232_43370# a_8704_45028# 3.4e-20
C28694 a_15959_42545# a_6755_46942# 9.08e-38
C28695 a_n2302_39072# a_n2442_46660# 1.26e-19
C28696 a_16409_43396# a_n443_42852# 2.64e-19
C28697 a_10807_43548# CLK 8.86e-22
C28698 a_11652_45724# a_10467_46802# 4.42e-19
C28699 a_4099_45572# a_3090_45724# 0.004385f
C28700 a_2711_45572# a_15368_46634# 0.0051f
C28701 a_20107_45572# a_13747_46662# 0.012917f
C28702 a_8746_45002# a_6755_46942# 4.26e-20
C28703 a_16377_45572# a_n743_46660# 5.01e-19
C28704 a_2437_43646# a_12891_46348# 0.004901f
C28705 a_21513_45002# a_12549_44172# 0.002562f
C28706 a_1423_45028# a_6545_47178# 4.56e-21
C28707 a_13556_45296# a_12861_44030# 0.028687f
C28708 a_13017_45260# a_11599_46634# 1.1e-20
C28709 a_413_45260# a_22959_47212# 0.024836f
C28710 a_8147_43396# a_5934_30871# 1.84e-20
C28711 a_5342_30871# a_16414_43172# 6.64e-20
C28712 a_n97_42460# a_16104_42674# 0.007062f
C28713 a_3626_43646# a_10723_42308# 0.003809f
C28714 a_2982_43646# a_5742_30871# 0.196805f
C28715 a_4361_42308# a_14635_42282# 0.018479f
C28716 a_16823_43084# a_16877_42852# 0.001502f
C28717 a_19237_31679# C10_N_btm 1.19e-19
C28718 a_6545_47178# a_6491_46660# 0.181574f
C28719 a_6151_47436# a_6851_47204# 0.007871f
C28720 a_4915_47217# a_6575_47204# 0.849579f
C28721 a_2063_45854# a_11599_46634# 0.19861f
C28722 a_3381_47502# a_n1435_47204# 4.12e-19
C28723 a_n1151_42308# a_13717_47436# 2.89e-19
C28724 a_n1059_45260# a_3499_42826# 0.002236f
C28725 a_3232_43370# a_2675_43914# 0.003881f
C28726 a_3537_45260# a_5495_43940# 2.48e-20
C28727 a_5147_45002# a_3905_42865# 0.048808f
C28728 a_5883_43914# a_10057_43914# 2.04e-20
C28729 a_n2129_44697# a_n1809_44850# 0.026556f
C28730 a_8701_44490# a_8975_43940# 9.09e-19
C28731 a_n2267_44484# a_n2012_44484# 0.05936f
C28732 a_10157_44484# a_10334_44484# 0.159555f
C28733 a_564_42282# a_n443_42852# 0.005734f
C28734 a_11962_45724# VDD 0.210594f
C28735 a_13777_45326# a_14035_46660# 4.08e-20
C28736 a_18287_44626# a_19321_45002# 0.00979f
C28737 a_4223_44672# a_2107_46812# 3.28e-20
C28738 a_13076_44458# a_n2661_46634# 7.24e-19
C28739 a_8975_43940# a_n2293_46634# 1.9e-19
C28740 a_18989_43940# a_13661_43548# 0.039099f
C28741 en_comp a_20202_43084# 6.61e-20
C28742 a_8488_45348# a_8270_45546# 3.69e-19
C28743 a_9838_44484# a_n743_46660# 8.79e-21
C28744 a_8746_45002# a_8049_45260# 0.001752f
C28745 a_8696_44636# a_17583_46090# 7.3e-19
C28746 a_15861_45028# a_15682_46116# 0.001207f
C28747 a_16680_45572# a_17715_44484# 0.001431f
C28748 a_14127_45572# a_10903_43370# 0.003658f
C28749 a_n2293_43922# a_n2312_39304# 5.35e-20
C28750 a_20362_44736# a_12861_44030# 0.004923f
C28751 a_1414_42308# a_n237_47217# 8.74e-23
C28752 a_453_43940# a_n746_45260# 0.004985f
C28753 COMP_P a_196_42282# 4.12e-21
C28754 a_5342_30871# a_7174_31319# 0.046616f
C28755 a_n4318_37592# a_n784_42308# 7e-20
C28756 a_n4318_38216# a_n1630_35242# 0.031712f
C28757 a_n3674_38216# a_n3674_37592# 0.048035f
C28758 a_21356_42826# a_17303_42282# 2.46e-20
C28759 a_n2293_46634# a_n133_46660# 1.8e-21
C28760 a_n2661_46634# a_601_46902# 0.009214f
C28761 a_n1925_46634# a_n1021_46688# 0.011448f
C28762 a_n2104_46634# a_n2438_43548# 0.052991f
C28763 a_n2312_38680# a_n743_46660# 0.001509f
C28764 a_n881_46662# a_5167_46660# 7.84e-21
C28765 a_n1613_43370# a_5907_46634# 0.338694f
C28766 a_4883_46098# a_6755_46942# 0.060162f
C28767 a_11599_46634# a_12469_46902# 9.01e-21
C28768 a_12861_44030# a_13607_46688# 0.019182f
C28769 a_n1151_42308# a_14035_46660# 0.026112f
C28770 a_n971_45724# a_765_45546# 0.140618f
C28771 a_13777_45326# a_9145_43396# 1.2e-21
C28772 a_5891_43370# a_8333_44056# 0.070354f
C28773 a_19279_43940# a_22485_44484# 2.14e-20
C28774 a_20679_44626# a_22959_44484# 1.47e-21
C28775 a_n2661_43370# a_4699_43561# 4.75e-21
C28776 a_9482_43914# a_10695_43548# 1.47e-20
C28777 a_14539_43914# a_15493_43940# 0.625897f
C28778 a_20640_44752# a_19237_31679# 7.45e-21
C28779 a_18989_43940# a_19862_44208# 7.01e-21
C28780 a_20193_45348# a_19319_43548# 1.24e-19
C28781 a_n2293_42834# a_2982_43646# 0.019738f
C28782 a_n2661_43922# a_n875_44318# 1.08e-19
C28783 a_11827_44484# a_21381_43940# 0.002761f
C28784 a_n2661_42834# a_n630_44306# 3.44e-19
C28785 a_8953_45002# a_10341_43396# 5.38e-21
C28786 a_n2946_37984# VDD 0.38275f
C28787 a_13807_45067# VDD 2.18e-20
C28788 a_5932_42308# VIN_N 0.023512f
C28789 a_n23_44458# a_167_45260# 7.57e-19
C28790 a_17517_44484# a_17339_46660# 0.020067f
C28791 a_5829_43940# a_5807_45002# 8.28e-21
C28792 a_n2661_43370# a_10586_45546# 0.002741f
C28793 a_8685_43396# a_4791_45118# 4.61e-21
C28794 a_3626_43646# a_16327_47482# 3.96e-19
C28795 a_20107_42308# a_7174_31319# 0.175129f
C28796 a_13258_32519# a_21335_42336# 0.022004f
C28797 a_19511_42282# a_21613_42308# 0.001375f
C28798 a_5934_30871# a_n4209_38216# 1.88e-21
C28799 SMPL_ON_N VDD 0.503419f
C28800 a_n1151_42308# a_n1099_45572# 0.046104f
C28801 a_2063_45854# a_1848_45724# 0.057473f
C28802 a_2609_46660# a_3147_46376# 4.21e-19
C28803 a_2443_46660# a_3483_46348# 1.28e-19
C28804 a_4883_46098# a_8049_45260# 0.469963f
C28805 a_10227_46804# a_12379_46436# 0.001273f
C28806 a_14955_47212# a_13259_45724# 7.31e-21
C28807 a_11599_46634# a_14383_46116# 0.026426f
C28808 a_12861_44030# a_16375_45002# 0.033138f
C28809 a_15928_47570# a_6945_45028# 0.004753f
C28810 a_13661_43548# a_18189_46348# 2.95e-19
C28811 a_12549_44172# a_10809_44734# 2.27272f
C28812 a_2107_46812# a_6419_46155# 0.007575f
C28813 a_n743_46660# a_9823_46155# 0.196587f
C28814 a_n2661_46634# a_12594_46348# 7.33e-20
C28815 a_13747_46662# a_17715_44484# 0.025502f
C28816 a_5807_45002# a_17957_46116# 0.00544f
C28817 a_n881_46662# a_518_46482# 5.79e-19
C28818 a_11813_46116# a_13059_46348# 0.001208f
C28819 a_15009_46634# a_13885_46660# 2.97e-19
C28820 a_12816_46660# a_14513_46634# 1.47e-20
C28821 a_14084_46812# a_14035_46660# 0.086342f
C28822 a_13607_46688# a_14180_46812# 5.9e-19
C28823 a_3357_43084# a_5932_42308# 2.19e-20
C28824 a_n2017_45002# a_3823_42558# 0.005755f
C28825 a_n1059_45260# a_3318_42354# 3.58e-19
C28826 a_n913_45002# a_2903_42308# 0.041908f
C28827 a_3537_45260# a_n784_42308# 5.26e-20
C28828 a_18184_42460# a_20922_43172# 0.018236f
C28829 a_18494_42460# a_19987_42826# 0.098055f
C28830 a_5343_44458# a_5111_42852# 1.38e-21
C28831 a_11827_44484# a_18249_42858# 1.13e-20
C28832 a_11691_44458# a_17595_43084# 7.45e-21
C28833 a_4223_44672# a_7871_42858# 5.46e-20
C28834 a_11967_42832# a_14579_43548# 0.060711f
C28835 a_3905_42865# a_4093_43548# 0.032751f
C28836 a_n1441_43940# a_n1177_43370# 6.39e-20
C28837 a_n4318_39768# VDD 0.469044f
C28838 a_13249_42308# a_8696_44636# 0.021669f
C28839 a_12427_45724# a_12649_45572# 0.001658f
C28840 a_11823_42460# a_12561_45572# 0.004618f
C28841 a_13635_43156# a_768_44030# 5.26e-19
C28842 a_16243_43396# a_6755_46942# 4.46e-20
C28843 a_7845_44172# a_8034_45724# 2.09e-21
C28844 a_20159_44458# a_n357_42282# 5.88e-21
C28845 a_3499_42826# a_n1925_42282# 4.47e-20
C28846 a_11173_44260# a_10903_43370# 0.035423f
C28847 a_12429_44172# a_10809_44734# 2.57e-21
C28848 a_12710_44260# a_9290_44172# 1.37e-19
C28849 a_196_42282# a_n2497_47436# 4.06e-22
C28850 a_n4318_37592# SMPL_ON_P 0.040097f
C28851 a_n1641_46494# a_n1379_46482# 0.001705f
C28852 a_n1423_46090# a_n967_46494# 4.2e-19
C28853 a_n1853_46287# a_n1533_46116# 8.49e-19
C28854 a_19692_46634# a_20850_46155# 0.006879f
C28855 a_13059_46348# a_14949_46494# 6.26e-19
C28856 a_5164_46348# a_2324_44458# 5.59e-20
C28857 a_10355_46116# a_9290_44172# 0.01806f
C28858 a_9823_46155# a_11189_46129# 6.08e-20
C28859 a_13483_43940# a_13635_43156# 4.94e-20
C28860 a_8791_43396# a_8685_43396# 0.086218f
C28861 a_n97_42460# a_18783_43370# 0.00416f
C28862 a_n2661_42834# a_1755_42282# 8.39e-21
C28863 a_3626_43646# a_10341_43396# 5.18e-20
C28864 a_6452_43396# a_6643_43396# 4.61e-19
C28865 a_20193_45348# a_21335_42336# 4.79e-20
C28866 SMPL_ON_N a_22469_39537# 0.017847f
C28867 a_13717_47436# START 0.034426f
C28868 a_9067_47204# DATA[4] 0.354356f
C28869 a_12861_44030# RST_Z 0.290405f
C28870 a_17499_43370# VDD 0.453381f
C28871 a_3429_45260# a_3232_43370# 0.001753f
C28872 a_4558_45348# a_5111_44636# 0.009468f
C28873 a_4574_45260# a_4927_45028# 0.047624f
C28874 a_3537_45260# a_5691_45260# 9.13e-19
C28875 a_2382_45260# a_5205_44484# 1.09e-21
C28876 a_3357_43084# a_1423_45028# 0.02044f
C28877 a_n913_45002# a_13556_45296# 7.49e-21
C28878 a_9049_44484# a_10157_44484# 1.97e-19
C28879 a_7499_43078# a_10334_44484# 1.72e-19
C28880 a_8696_44636# a_17613_45144# 0.09062f
C28881 a_15861_45028# a_17023_45118# 0.076138f
C28882 a_17478_45572# a_16922_45042# 3.77e-20
C28883 a_10518_42984# a_4185_45028# 8.53e-21
C28884 a_22165_42308# a_20202_43084# 0.001287f
C28885 a_6171_42473# a_4646_46812# 2.16e-21
C28886 a_6031_43396# a_n357_42282# 0.012855f
C28887 a_n1557_42282# a_n443_42852# 0.078868f
C28888 a_n2946_39866# a_n2312_40392# 2.19e-20
C28889 a_n3420_39616# a_n2312_39304# 1.17e-19
C28890 a_3422_30871# VIN_P 0.057975f
C28891 a_9049_44484# a_n1925_46634# 2.71e-20
C28892 a_14495_45572# a_13747_46662# 0.288916f
C28893 a_11322_45546# a_n2661_46634# 0.059929f
C28894 a_8568_45546# a_n743_46660# 3.92e-20
C28895 a_4099_45572# a_3699_46634# 4.97e-20
C28896 a_10193_42453# a_n2293_46634# 0.037794f
C28897 a_6229_45572# a_5807_45002# 6.77e-19
C28898 a_18341_45572# a_18597_46090# 0.010006f
C28899 a_18909_45814# a_18780_47178# 1.24e-20
C28900 a_20107_45572# a_11599_46634# 0.246047f
C28901 a_17568_45572# a_16327_47482# 9.92e-19
C28902 a_3357_43084# a_6491_46660# 0.014978f
C28903 a_2437_43646# a_7903_47542# 0.006626f
C28904 a_21363_45546# a_12861_44030# 1.6e-22
C28905 a_2382_45260# a_n971_45724# 0.019144f
C28906 a_n1059_45260# a_n1151_42308# 0.16984f
C28907 a_5147_45002# a_n2109_47186# 0.05864f
C28908 a_1667_45002# a_n237_47217# 0.002992f
C28909 a_20205_31679# a_21167_46155# 4.36e-20
C28910 a_n4318_39768# a_n2860_39866# 4.42e-20
C28911 a_15493_43396# a_4958_30871# 1.31e-20
C28912 a_13467_32519# a_5534_30871# 0.041703f
C28913 a_n1557_42282# a_n2104_42282# 3.45e-19
C28914 a_4190_30871# a_17595_43084# 7.76e-19
C28915 a_743_42282# a_16414_43172# 5.93e-20
C28916 a_5649_42852# a_12895_43230# 9.12e-21
C28917 a_685_42968# a_791_42968# 0.13675f
C28918 a_14180_46812# RST_Z 5.82e-19
C28919 a_n3420_37984# VDAC_P 3.33e-19
C28920 a_3754_38802# VDAC_Ni 0.301032f
C28921 a_7754_39300# a_8530_39574# 3.17e-19
C28922 a_2113_38308# a_4338_37500# 1.76e-20
C28923 a_1576_42282# VDD 0.26017f
C28924 a_n2288_47178# a_n1920_47178# 7.52e-19
C28925 a_n2497_47436# a_n1741_47186# 0.098118f
C28926 a_n2833_47464# SMPL_ON_P 0.002772f
C28927 a_10775_45002# a_n2661_43922# 8.33e-21
C28928 a_10951_45334# a_n2661_42834# 1.25e-20
C28929 a_n2661_43370# a_10440_44484# 9.47e-21
C28930 a_1423_45028# a_5826_44734# 0.003941f
C28931 a_21101_45002# a_18114_32519# 1.7e-19
C28932 a_10193_42453# a_11816_44260# 1.82e-19
C28933 a_19479_31679# a_3422_30871# 2.13e-21
C28934 a_3823_42558# a_526_44458# 0.183187f
C28935 a_3318_42354# a_n1925_42282# 6.66e-20
C28936 a_8483_43230# a_n443_42852# 0.001379f
C28937 a_14113_42308# a_9290_44172# 4.21e-20
C28938 a_14456_42282# a_10903_43370# 3.29e-21
C28939 a_15903_45785# a_12741_44636# 1.65e-19
C28940 a_16115_45572# a_11415_45002# 0.004692f
C28941 a_18341_45572# a_19123_46287# 0.001192f
C28942 a_1423_45028# a_3877_44458# 0.022537f
C28943 a_n2661_43370# a_n743_46660# 7.86e-20
C28944 a_18909_45814# a_18285_46348# 1.07e-21
C28945 a_17719_45144# a_13747_46662# 3.9e-20
C28946 a_18315_45260# a_13661_43548# 0.002575f
C28947 a_18587_45118# a_5807_45002# 5.91e-22
C28948 a_8953_45002# a_8667_46634# 8.44e-19
C28949 a_20447_31679# a_15227_44166# 2.55e-19
C28950 a_10193_42453# a_9625_46129# 0.002796f
C28951 a_10053_45546# a_9823_46155# 8.94e-19
C28952 a_11322_45546# a_8199_44636# 8.36e-19
C28953 a_7499_43078# a_9290_44172# 0.597117f
C28954 a_10490_45724# a_5937_45572# 3.4e-20
C28955 a_8746_45002# a_8953_45546# 0.020026f
C28956 a_484_44484# a_n1151_42308# 2.43e-19
C28957 a_8783_44734# a_4791_45118# 6.39e-21
C28958 a_13720_44458# a_10227_46804# 0.001314f
C28959 a_17767_44458# a_16327_47482# 0.269619f
C28960 a_n2293_42282# a_1755_42282# 0.875855f
C28961 a_743_42282# a_7174_31319# 0.004769f
C28962 a_20556_43646# a_20712_42282# 1.47e-20
C28963 a_4361_42308# a_19511_42282# 0.071032f
C28964 a_5342_30871# a_5932_42308# 0.01856f
C28965 a_20205_31679# VREF_GND 0.001993f
C28966 a_20692_30879# VREF 0.098117f
C28967 a_2063_45854# a_7411_46660# 0.029159f
C28968 a_4791_45118# a_5907_46634# 0.016954f
C28969 a_n237_47217# a_10428_46928# 1.3e-19
C28970 a_n2109_47186# a_5841_46660# 1.94e-19
C28971 a_4915_47217# a_5385_46902# 9.3e-21
C28972 a_5129_47502# a_4817_46660# 0.001806f
C28973 a_6545_47178# a_4646_46812# 0.02302f
C28974 a_6491_46660# a_3877_44458# 0.02519f
C28975 a_22959_47212# a_20916_46384# 9.45e-20
C28976 SMPL_ON_N a_22612_30879# 5.16049f
C28977 a_12465_44636# a_n2661_46634# 1.89e-19
C28978 a_11453_44696# a_21588_30879# 0.075738f
C28979 a_n1613_43370# a_768_44030# 0.028683f
C28980 a_n881_46662# a_12549_44172# 0.225257f
C28981 C1_P_btm VDD 0.264503f
C28982 a_3357_43084# a_4181_43396# 1.16e-20
C28983 a_413_45260# a_2982_43646# 7.3e-22
C28984 a_n1059_45260# a_6197_43396# 4.64e-20
C28985 a_n913_45002# a_6293_42852# 0.001086f
C28986 a_4574_45260# a_4699_43561# 3.74e-21
C28987 a_3537_45260# a_3080_42308# 0.02683f
C28988 a_15463_44811# a_14673_44172# 0.001037f
C28989 a_5883_43914# a_5013_44260# 0.001282f
C28990 a_18494_42460# a_18326_43940# 1.27e-19
C28991 a_16922_45042# a_20935_43940# 1.08e-20
C28992 a_19778_44110# a_19328_44172# 0.064774f
C28993 a_11827_44484# a_14955_43940# 0.005645f
C28994 a_n2012_44484# a_n2065_43946# 7.1e-20
C28995 a_5343_44458# a_7542_44172# 0.014194f
C28996 a_n1177_44458# a_n1441_43940# 7.12e-20
C28997 a_6298_44484# a_6453_43914# 0.002276f
C28998 a_18911_45144# a_15493_43396# 2.88e-21
C28999 a_n4334_38304# a_n2956_38216# 6.77e-20
C29000 a_7229_43940# VDD 0.821851f
C29001 a_n2661_44458# a_12741_44636# 0.004092f
C29002 a_18248_44752# a_16388_46812# 1.08e-21
C29003 a_5495_43940# a_n2293_46634# 8.7e-21
C29004 a_7584_44260# a_768_44030# 6.93e-19
C29005 a_3232_43370# a_8049_45260# 0.003961f
C29006 a_19963_31679# a_20205_31679# 9.023429f
C29007 a_3357_43084# a_20850_46155# 5.34e-19
C29008 a_n2661_43370# a_11189_46129# 7.55e-21
C29009 a_5837_45028# a_2324_44458# 0.003084f
C29010 a_15493_43940# a_11453_44696# 5.75e-20
C29011 a_n1655_43396# a_n971_45724# 2.13e-20
C29012 a_n237_47217# VDD 4.05131f
C29013 a_11551_42558# a_11633_42308# 0.003935f
C29014 a_n784_42308# a_1343_38525# 2.98e-20
C29015 a_5755_42308# a_7174_31319# 9.76e-21
C29016 a_14113_42308# a_15051_42282# 0.077852f
C29017 a_13657_42558# a_15486_42560# 1.21e-20
C29018 VIN_N VREF 0.775904f
C29019 VIN_P VREF_GND 16.4969f
C29020 a_768_44030# a_n2293_46098# 0.039783f
C29021 a_5807_45002# a_11415_45002# 0.05094f
C29022 a_13661_43548# a_20202_43084# 1.29e-19
C29023 a_601_46902# a_765_45546# 1.65e-19
C29024 a_10150_46912# a_10384_47026# 0.006453f
C29025 a_6755_46942# a_6682_46660# 9.82e-21
C29026 a_10428_46928# a_8270_45546# 1.48e-19
C29027 a_n881_46662# a_1208_46090# 0.076994f
C29028 a_n1613_43370# a_1176_45822# 0.004031f
C29029 a_4883_46098# a_8953_45546# 0.078639f
C29030 a_11599_46634# a_17715_44484# 0.031427f
C29031 a_15673_47210# a_2324_44458# 1.57e-19
C29032 a_10227_46804# a_13351_46090# 0.008909f
C29033 a_15811_47375# a_15682_46116# 0.002105f
C29034 a_12861_44030# a_18985_46122# 4.61e-20
C29035 a_13717_47436# a_19553_46090# 3.99e-21
C29036 a_9863_47436# a_6945_45028# 0.0046f
C29037 a_3160_47472# a_3873_46454# 5.76e-19
C29038 a_n237_47217# a_8283_46482# 1.91e-19
C29039 a_n1151_42308# a_n1925_42282# 3.65e-19
C29040 a_n443_46116# a_518_46482# 6.82e-19
C29041 a_3381_47502# a_526_44458# 9.83e-20
C29042 a_1467_44172# a_1443_43940# 0.011516f
C29043 a_1414_42308# a_1241_43940# 0.005139f
C29044 a_20766_44850# a_20974_43370# 4.78e-21
C29045 a_n2293_42834# a_7871_42858# 0.027f
C29046 a_2711_45572# a_19332_42282# 0.004712f
C29047 a_453_43940# a_726_44056# 0.001159f
C29048 a_11823_42460# a_11323_42473# 0.0014f
C29049 a_9672_43914# a_10729_43914# 1.18e-19
C29050 a_n2293_43922# a_3626_43646# 0.03147f
C29051 a_n2661_42834# a_n1243_43396# 9.21e-20
C29052 a_n913_45002# a_11554_42852# 0.016237f
C29053 a_2382_45260# a_3863_42891# 6.79e-20
C29054 a_3537_45260# a_7309_43172# 4.53e-19
C29055 a_n1059_45260# a_10752_42852# 1.72e-19
C29056 a_18204_44850# VDD 4.6e-19
C29057 a_2711_45572# a_10210_45822# 0.007317f
C29058 a_6472_45840# a_6469_45572# 2.36e-20
C29059 a_7499_43078# a_9049_44484# 8.37e-20
C29060 a_19862_44208# a_20202_43084# 0.058613f
C29061 a_n2661_42282# a_1823_45246# 3.88e-19
C29062 a_19268_43646# a_19321_45002# 1.56e-20
C29063 a_16867_43762# a_13661_43548# 6.73e-22
C29064 a_16137_43396# a_n2293_46634# 4.18e-20
C29065 a_n23_44458# a_n863_45724# 0.056041f
C29066 a_n356_44636# a_n452_45724# 7.27e-21
C29067 a_6453_43914# a_5937_45572# 0.144397f
C29068 a_20447_31679# EN_OFFSET_CAL 2.14e-19
C29069 a_19479_31679# VREF_GND 0.00198f
C29070 a_n913_45002# RST_Z 2.65e-19
C29071 a_8270_45546# VDD 1.26092f
C29072 a_5742_30871# a_n4064_37984# 0.004679f
C29073 a_n2293_46098# a_1176_45822# 0.027035f
C29074 a_20202_43084# a_4185_45028# 2.38e-19
C29075 a_n1641_46494# a_n1076_46494# 7.99e-20
C29076 a_765_45546# a_12594_46348# 7.51e-20
C29077 a_n743_46660# a_2307_45899# 2.73e-19
C29078 a_33_46660# a_n443_42852# 1.61e-19
C29079 a_n2661_46098# a_n755_45592# 7.65e-20
C29080 a_n2956_37592# a_n2946_38778# 2.49e-19
C29081 a_14021_43940# a_14621_43646# 0.001689f
C29082 a_458_43396# a_766_43646# 0.017351f
C29083 a_n1177_43370# a_n998_43396# 0.007399f
C29084 a_n1352_43396# a_n1243_43396# 0.007416f
C29085 a_n3674_39768# a_n3674_39304# 0.037712f
C29086 a_n4318_39768# a_n4318_38680# 0.02372f
C29087 a_n699_43396# a_1576_42282# 7.71e-23
C29088 a_18579_44172# a_18083_42858# 2.69e-21
C29089 a_n97_42460# a_3626_43646# 0.394673f
C29090 a_2675_43914# a_2905_42968# 9.88e-21
C29091 a_11341_43940# a_18525_43370# 1.4e-19
C29092 a_15493_43940# a_17324_43396# 1.55e-20
C29093 a_20935_43940# a_15743_43084# 6.65e-21
C29094 a_15682_43940# a_16823_43084# 7.58e-19
C29095 a_11967_42832# a_21671_42860# 1.16e-19
C29096 a_9313_44734# a_13157_43218# 1.2e-19
C29097 w_1575_34946# EN_VIN_BSTR_P 3.99222f
C29098 a_15903_45785# a_13556_45296# 1.89e-19
C29099 a_15037_45618# a_14797_45144# 0.003975f
C29100 a_8696_44636# a_11787_45002# 5.52e-20
C29101 a_3357_43084# a_22591_45572# 0.181818f
C29102 a_19479_31679# a_19963_31679# 0.104687f
C29103 a_2437_43646# a_20447_31679# 1.16e-19
C29104 a_21513_45002# a_21297_45572# 1.2e-19
C29105 a_14209_32519# a_21076_30879# 0.055087f
C29106 a_n4318_37592# a_n2438_43548# 1.35e-19
C29107 a_19339_43156# a_3090_45724# 2.9e-19
C29108 a_17595_43084# a_15227_44166# 0.041195f
C29109 a_n1630_35242# a_n2956_39768# 0.003986f
C29110 a_6123_31319# a_n1613_43370# 0.002625f
C29111 a_12638_46436# VDD 0.002311f
C29112 a_10193_42453# a_18597_46090# 0.001118f
C29113 a_15143_45578# a_14955_47212# 2.5e-21
C29114 a_14495_45572# a_11599_46634# 3.57e-19
C29115 a_n2956_39304# a_n2840_45546# 4.31e-19
C29116 a_2324_44458# a_3316_45546# 1.07e-19
C29117 a_21259_43561# a_4361_42308# 0.005186f
C29118 a_10695_43548# a_10796_42968# 6.99e-20
C29119 a_3422_30871# a_13258_32519# 0.410904f
C29120 a_4190_30871# a_13467_32519# 0.032722f
C29121 a_3626_43646# a_3935_43218# 6.34e-19
C29122 a_n2661_42282# a_5934_30871# 2.9e-20
C29123 a_4649_42852# VDD 0.194775f
C29124 a_n2017_45002# a_n1655_44484# 6.5e-19
C29125 a_3537_45260# a_10057_43914# 0.001231f
C29126 a_3357_43084# a_6109_44484# 0.016236f
C29127 a_5111_44636# a_9838_44484# 1.88e-22
C29128 a_5205_44484# a_5343_44458# 0.129692f
C29129 a_n2293_45010# a_n23_44458# 1.13e-19
C29130 a_3232_43370# a_8103_44636# 0.013825f
C29131 a_6171_45002# a_6298_44484# 0.001994f
C29132 a_8696_44636# a_17325_44484# 5.02e-20
C29133 a_16115_45572# a_11967_42832# 1.12e-20
C29134 a_3497_42558# a_1823_45246# 0.002234f
C29135 a_20712_42282# a_19692_46634# 1.06e-20
C29136 a_3935_42891# a_n443_42852# 5.99e-20
C29137 a_10796_42968# a_n357_42282# 0.048375f
C29138 a_21671_42860# a_13259_45724# 1.9e-20
C29139 a_15037_45618# a_14976_45028# 0.003888f
C29140 a_13904_45546# a_13059_46348# 0.001004f
C29141 a_13159_45002# a_5807_45002# 1.28e-21
C29142 a_1307_43914# a_12549_44172# 1.82879f
C29143 a_13017_45260# a_13661_43548# 6.88e-20
C29144 a_14033_45822# a_15368_46634# 8.96e-21
C29145 a_8696_44636# a_11813_46116# 4.79e-21
C29146 a_15225_45822# a_3090_45724# 7.41e-20
C29147 a_3357_43084# a_4646_46812# 0.024669f
C29148 a_2437_43646# a_4817_46660# 4.02e-20
C29149 a_1667_45002# a_1123_46634# 3.71e-19
C29150 a_4574_45260# a_n743_46660# 5.3e-20
C29151 a_413_45260# a_2107_46812# 0.032665f
C29152 a_5147_45002# a_n1925_46634# 2.49e-20
C29153 a_1423_45028# a_8128_46384# 2.49e-21
C29154 a_17719_45144# a_11599_46634# 1.93e-21
C29155 a_19778_44110# a_12861_44030# 0.113118f
C29156 a_18194_35068# VDD 2.17116f
C29157 a_5343_44458# a_n971_45724# 0.001055f
C29158 a_16414_43172# a_16328_43172# 0.001377f
C29159 a_3080_42308# a_1343_38525# 3.95e-19
C29160 a_4361_42308# a_4921_42308# 0.472085f
C29161 a_743_42282# a_5932_42308# 0.024532f
C29162 a_15681_43442# a_15486_42560# 2.96e-20
C29163 a_1736_39043# VDD 2.8939f
C29164 a_4915_47217# a_12891_46348# 0.156543f
C29165 a_6575_47204# a_n881_46662# 0.708623f
C29166 a_7903_47542# a_7989_47542# 0.006584f
C29167 a_6491_46660# a_8128_46384# 6.19e-21
C29168 a_n2109_47186# a_n1925_46634# 0.033276f
C29169 SMPL_ON_P a_n2293_46634# 9.68e-20
C29170 a_n452_47436# a_n2661_46634# 0.001956f
C29171 a_4791_45118# a_768_44030# 0.03019f
C29172 a_n2497_47436# a_n743_46660# 1.09e-19
C29173 a_n1605_47204# a_n2442_46660# 3.01e-19
C29174 a_18143_47464# a_12465_44636# 0.001005f
C29175 a_20894_47436# a_20990_47178# 0.313533f
C29176 a_19386_47436# a_13507_46334# 6.44e-21
C29177 a_18780_47178# a_4883_46098# 4.43e-20
C29178 a_18479_47436# a_21811_47423# 1.31e-19
C29179 a_21359_45002# a_20512_43084# 7.4e-21
C29180 a_1423_45028# a_9672_43914# 4.02e-19
C29181 a_13249_42308# a_14205_43396# 5.12e-22
C29182 a_20193_45348# a_3422_30871# 0.042753f
C29183 a_n2661_43370# a_5244_44056# 4.22e-21
C29184 a_1307_43914# a_12429_44172# 0.007436f
C29185 a_8975_43940# a_10809_44484# 5.15e-19
C29186 a_20205_45028# a_19279_43940# 6.24e-19
C29187 a_11827_44484# a_21145_44484# 0.001286f
C29188 a_18114_32519# a_20766_44850# 2.21e-19
C29189 a_3232_43370# a_11173_44260# 0.002786f
C29190 a_15890_42674# a_n443_42852# 5.07e-21
C29191 a_4958_30871# a_n357_42282# 0.004392f
C29192 a_18596_45572# VDD 0.077608f
C29193 a_5534_30871# VCM 0.095752f
C29194 a_20922_43172# RST_Z 2.99e-22
C29195 a_13348_45260# a_3483_46348# 0.041217f
C29196 a_16922_45042# a_16388_46812# 4.23e-21
C29197 a_11967_42832# a_5807_45002# 3.26e-19
C29198 a_18579_44172# a_12549_44172# 0.154956f
C29199 a_16115_45572# a_13259_45724# 0.035684f
C29200 a_18341_45572# a_8049_45260# 0.021945f
C29201 a_15903_45785# a_16375_45002# 0.005324f
C29202 a_20447_31679# a_22959_46124# 0.015464f
C29203 a_6171_45002# a_5937_45572# 0.206948f
C29204 a_6709_45028# a_6419_46155# 3.25e-20
C29205 a_3232_43370# a_8953_45546# 0.019509f
C29206 a_1184_42692# a_5742_30871# 1.12e-20
C29207 a_4921_42308# a_6761_42308# 9.41e-19
C29208 a_5755_42308# a_5932_42308# 0.196877f
C29209 a_3823_42558# a_4169_42308# 0.013377f
C29210 a_17364_32525# C9_N_btm 7.29e-20
C29211 a_n443_46116# a_1208_46090# 1.26e-19
C29212 a_2063_45854# a_4185_45028# 0.023928f
C29213 a_n1151_42308# a_2698_46116# 9.22e-21
C29214 a_4007_47204# a_1823_45246# 4.86e-22
C29215 a_2905_45572# a_3147_46376# 0.02017f
C29216 a_3160_47472# a_2804_46116# 4.58e-19
C29217 a_n971_45724# a_8349_46414# 0.01782f
C29218 a_n1741_47186# a_9569_46155# 4.67e-20
C29219 a_n237_47217# a_7920_46348# 0.059304f
C29220 a_584_46384# a_4419_46090# 3.79e-21
C29221 a_10227_46804# a_20731_47026# 0.016434f
C29222 a_13717_47436# a_12741_44636# 5.57e-20
C29223 a_13507_46334# a_19551_46910# 0.002438f
C29224 a_20894_47436# a_20273_46660# 6.02e-20
C29225 a_21177_47436# a_20107_46660# 9.39e-19
C29226 a_4883_46098# a_18285_46348# 0.026239f
C29227 a_12465_44636# a_765_45546# 0.019565f
C29228 a_n1925_46634# a_5841_46660# 1.6e-19
C29229 a_n2661_46634# a_8654_47026# 1.14e-19
C29230 a_3524_46660# a_5072_46660# 5.75e-21
C29231 a_3877_44458# a_4646_46812# 0.056449f
C29232 a_12549_44172# a_17609_46634# 0.487224f
C29233 a_5807_45002# a_12251_46660# 0.003883f
C29234 a_n2017_45002# a_10341_42308# 0.049998f
C29235 a_n1059_45260# a_10922_42852# 0.002568f
C29236 a_n913_45002# a_10991_42826# 0.029878f
C29237 a_3065_45002# a_3681_42891# 1.71e-20
C29238 a_n699_43396# a_1987_43646# 2.2e-19
C29239 a_2998_44172# a_5244_44056# 3.3e-19
C29240 a_n2661_42834# a_3737_43940# 3.81e-20
C29241 a_n1761_44111# a_n822_43940# 2.49e-19
C29242 a_3600_43914# a_3905_42865# 1.98e-20
C29243 a_742_44458# a_3626_43646# 3.38e-20
C29244 a_11827_44484# a_8685_43396# 3.35e-20
C29245 a_n1331_43914# a_n1441_43940# 0.097745f
C29246 a_11967_42832# a_19478_44306# 2.52e-19
C29247 a_8696_44636# a_8495_42852# 8.39e-21
C29248 a_2779_44458# a_2982_43646# 1.05e-20
C29249 a_15004_44636# VDD 0.090175f
C29250 a_n3420_39616# C10_P_btm 2.16e-19
C29251 a_n3565_39590# C8_P_btm 0.384801f
C29252 a_n4064_40160# C2_P_btm 1.17e-19
C29253 a_n4209_39304# a_n1386_35608# 9.16e-20
C29254 a_13258_32519# VREF_GND 0.033872f
C29255 a_7174_31319# VIN_P 0.022822f
C29256 a_17730_32519# a_21076_30879# 0.054832f
C29257 a_5745_43940# a_5257_43370# 0.005229f
C29258 a_17973_43940# a_3090_45724# 0.001042f
C29259 a_1049_43396# a_n2438_43548# 1.79e-20
C29260 a_3080_42308# a_n2293_46634# 0.039273f
C29261 a_8975_43940# a_8049_45260# 6.62e-21
C29262 a_n2661_42834# a_2324_44458# 0.004585f
C29263 a_6809_43396# a_n1613_43370# 0.001918f
C29264 a_18525_43370# a_16327_47482# 0.059008f
C29265 a_1123_46634# VDD 0.469393f
C29266 a_n4334_39392# a_n3690_39392# 8.67e-19
C29267 a_n4209_39304# a_n3420_39072# 0.071714f
C29268 a_5742_30871# C0_P_btm 0.014563f
C29269 a_3090_45724# a_167_45260# 5.35e-19
C29270 a_14035_46660# a_12741_44636# 8.27e-21
C29271 a_20411_46873# a_20273_46660# 0.219954f
C29272 a_20107_46660# a_20841_46902# 0.053479f
C29273 a_5807_45002# a_13259_45724# 0.096565f
C29274 a_2959_46660# a_526_44458# 6.06e-19
C29275 a_12549_44172# a_19443_46116# 3.9e-22
C29276 a_n743_46660# a_9823_46482# 0.004996f
C29277 a_n1925_46634# a_8062_46155# 1.86e-19
C29278 a_n881_46662# a_n2661_45546# 0.02866f
C29279 a_8270_45546# a_7920_46348# 5.66e-19
C29280 a_10249_46116# a_10903_43370# 7.46e-21
C29281 a_n310_47243# a_n755_45592# 3.51e-20
C29282 a_n3674_38680# a_n3420_37984# 2.36e-20
C29283 a_9159_44484# a_8952_43230# 1.71e-20
C29284 a_n2293_43922# a_8037_42858# 1.82e-20
C29285 a_n2661_42834# a_8387_43230# 2.69e-20
C29286 a_9313_44734# a_12089_42308# 0.011899f
C29287 a_n2293_42834# a_1184_42692# 6.11e-20
C29288 a_1307_43914# a_7227_42308# 7.17e-37
C29289 a_n2661_44458# a_11554_42852# 3.79e-20
C29290 a_n1059_45260# a_17531_42308# 0.001278f
C29291 a_n2017_45002# a_18057_42282# 4.4e-19
C29292 a_n913_45002# a_17303_42282# 1.81467f
C29293 a_19963_31679# a_13258_32519# 0.054679f
C29294 a_1241_43940# VDD 0.162129f
C29295 a_2711_45572# a_14797_45144# 4.99e-20
C29296 a_17478_45572# a_17668_45572# 0.045837f
C29297 a_9145_43396# a_12741_44636# 3.38e-20
C29298 a_20556_43646# a_19692_46634# 0.118928f
C29299 a_16977_43638# a_17339_46660# 3.09e-20
C29300 a_6453_43914# a_n443_42852# 4.9e-19
C29301 a_1525_44260# a_n357_42282# 1.47e-19
C29302 a_6123_31319# a_4791_45118# 3.81e-20
C29303 a_n4064_37440# C2_P_btm 0.001797f
C29304 a_13759_46122# VDD 0.399995f
C29305 a_6667_45809# a_2063_45854# 0.029741f
C29306 a_4880_45572# a_n971_45724# 2.82e-20
C29307 a_5263_45724# a_n1151_42308# 0.005089f
C29308 a_2711_45572# a_3815_47204# 3.98e-20
C29309 a_8199_44636# a_10037_46155# 4.91e-19
C29310 a_11387_46155# a_8049_45260# 0.00421f
C29311 a_2324_44458# a_5066_45546# 0.002463f
C29312 a_n1736_46482# a_n1545_46494# 4.61e-19
C29313 a_n2472_46090# a_n2956_38216# 5.66e-19
C29314 a_n2293_46098# a_n2472_45546# 0.015672f
C29315 a_n2157_46122# a_n2661_45546# 5.14e-20
C29316 a_n1761_44111# a_n327_42308# 1.97e-19
C29317 a_9313_44734# a_18907_42674# 4.46e-21
C29318 a_1467_44172# a_1576_42282# 1.16e-20
C29319 a_1414_42308# a_1067_42314# 0.100434f
C29320 a_n97_42460# a_8037_42858# 4.35e-19
C29321 a_10341_43396# a_18525_43370# 0.015853f
C29322 a_1568_43370# a_1847_42826# 0.153113f
C29323 a_1115_44172# a_1184_42692# 1.35e-20
C29324 a_12891_46348# DATA[5] 0.001817f
C29325 a_5755_42852# VDD 0.179985f
C29326 a_17478_45572# a_17970_44736# 3.84e-19
C29327 a_626_44172# a_1423_45028# 0.014461f
C29328 a_8696_44636# a_18287_44626# 8.04e-20
C29329 a_5111_44636# a_n2661_43370# 0.075649f
C29330 a_n1059_45260# a_18184_42460# 0.52106f
C29331 a_n2017_45002# a_18494_42460# 0.002888f
C29332 a_3232_43370# a_7735_45067# 0.001345f
C29333 a_6709_45028# a_n2293_42834# 0.001466f
C29334 a_16547_43609# a_n443_42852# 0.004823f
C29335 a_10949_43914# CLK 1.96e-21
C29336 a_9159_45572# a_4646_46812# 1.29e-20
C29337 a_10193_42453# a_6755_46942# 0.00109f
C29338 a_3175_45822# a_3090_45724# 0.008745f
C29339 a_2711_45572# a_14976_45028# 0.025742f
C29340 a_8746_45002# a_10249_46116# 1.31e-20
C29341 a_16211_45572# a_n743_46660# 8.28e-19
C29342 a_2437_43646# a_11309_47204# 0.003942f
C29343 a_3357_43084# a_9804_47204# 8.68e-20
C29344 a_2903_45348# a_n443_46116# 9.86e-20
C29345 a_8560_45348# a_n971_45724# 0.007243f
C29346 a_1423_45028# a_6151_47436# 2.69e-21
C29347 a_9482_43914# a_12861_44030# 0.021886f
C29348 a_11963_45334# a_11599_46634# 7.4e-22
C29349 a_413_45260# a_11453_44696# 0.032816f
C29350 a_5342_30871# a_15567_42826# 0.024331f
C29351 a_3626_43646# a_10533_42308# 0.002711f
C29352 a_2982_43646# a_11323_42473# 1.02e-19
C29353 a_4361_42308# a_13291_42460# 0.029279f
C29354 a_19319_43548# a_19647_42308# 1.57e-21
C29355 a_2905_42968# a_3059_42968# 0.008678f
C29356 a_n97_42460# a_13921_42308# 0.003369f
C29357 a_4190_30871# a_18695_43230# 1.55e-19
C29358 a_19237_31679# C9_N_btm 3.18e-20
C29359 a_5815_47464# a_6851_47204# 1.23e-20
C29360 a_6151_47436# a_6491_46660# 0.31912f
C29361 a_4915_47217# a_7903_47542# 0.042037f
C29362 a_n1151_42308# a_n1435_47204# 0.002911f
C29363 a_n443_46116# a_6575_47204# 2.21e-20
C29364 a_n2017_45002# a_3499_42826# 4.96e-19
C29365 a_5147_45002# a_3600_43914# 7.58e-20
C29366 a_3537_45260# a_5013_44260# 0.001173f
C29367 a_4558_45348# a_3905_42865# 9.27e-19
C29368 a_n2661_44458# a_n1190_44850# 1.42e-19
C29369 a_8103_44636# a_8975_43940# 1.09e-20
C29370 a_n2433_44484# a_n1809_44850# 9.73e-19
C29371 a_n2129_44697# a_n2012_44484# 0.172424f
C29372 a_20107_45572# a_19862_44208# 4.31e-20
C29373 a_n39_42308# a_n755_45592# 7.86e-19
C29374 a_n3674_37592# a_n443_42852# 6.07e-20
C29375 a_11652_45724# VDD 0.155048f
C29376 a_4190_30871# VCM 1.23535f
C29377 a_17364_32525# RST_Z 0.050609f
C29378 a_13556_45296# a_14035_46660# 1.33e-21
C29379 a_2437_43646# a_472_46348# 1.19e-20
C29380 a_18248_44752# a_19321_45002# 0.004965f
C29381 a_2779_44458# a_2107_46812# 6.26e-21
C29382 a_18374_44850# a_13661_43548# 0.00877f
C29383 a_10057_43914# a_n2293_46634# 0.01757f
C29384 a_18989_43940# a_5807_45002# 5.17e-20
C29385 a_10193_42453# a_8049_45260# 0.082788f
C29386 a_8696_44636# a_15682_46116# 0.00216f
C29387 a_15861_45028# a_2324_44458# 8.69e-19
C29388 a_14033_45572# a_10903_43370# 0.003863f
C29389 a_16855_45546# a_17715_44484# 0.001764f
C29390 a_n2661_43922# a_n2312_39304# 1.13e-20
C29391 a_n2293_43922# a_n2312_40392# 0.002335f
C29392 a_20159_44458# a_12861_44030# 0.014378f
C29393 a_1414_42308# a_n746_45260# 3.24e-20
C29394 a_n1899_43946# a_584_46384# 6.88e-21
C29395 COMP_P a_n473_42460# 1.25e-19
C29396 a_n1736_42282# a_n784_42308# 2.19e-19
C29397 a_n2104_42282# a_n3674_37592# 0.006157f
C29398 a_n1329_42308# a_n961_42308# 0.001982f
C29399 a_n2472_42282# a_n1630_35242# 0.040716f
C29400 a_20922_43172# a_17303_42282# 1.39e-20
C29401 a_18599_43230# a_18907_42674# 0.001393f
C29402 a_18249_42858# a_18214_42558# 2.84e-19
C29403 a_n2661_46634# a_33_46660# 0.050833f
C29404 a_n2293_46634# a_n2438_43548# 0.807205f
C29405 a_n2312_38680# a_n1021_46688# 7.19e-20
C29406 a_n2104_46634# a_n743_46660# 6.41e-20
C29407 a_n881_46662# a_5385_46902# 5.4e-19
C29408 a_8128_46384# a_4646_46812# 5.76e-21
C29409 a_n1613_43370# a_5167_46660# 0.177362f
C29410 a_4883_46098# a_10249_46116# 0.01923f
C29411 a_11599_46634# a_11901_46660# 0.002693f
C29412 a_12861_44030# a_12816_46660# 7.2e-19
C29413 a_13717_47436# a_13607_46688# 6.92e-19
C29414 a_4915_47217# a_12359_47026# 2.51e-19
C29415 a_n1151_42308# a_13885_46660# 0.333314f
C29416 a_21005_45260# a_20974_43370# 3.69e-20
C29417 a_21359_45002# a_21381_43940# 5.38e-20
C29418 a_8375_44464# a_8333_44056# 2.14e-19
C29419 a_9482_43914# a_9803_43646# 9.27e-20
C29420 a_13556_45296# a_9145_43396# 5.5e-21
C29421 a_16979_44734# a_11341_43940# 5.51e-20
C29422 a_19279_43940# a_20512_43084# 1.32e-19
C29423 a_20679_44626# a_17730_32519# 3.62e-21
C29424 a_18989_43940# a_19478_44306# 1.12e-19
C29425 a_11691_44458# a_19319_43548# 4.59e-19
C29426 a_8696_44636# a_9127_43156# 6.2e-21
C29427 a_5891_43370# a_8018_44260# 8.02e-19
C29428 a_16112_44458# a_15493_43940# 4.79e-19
C29429 a_n2661_43922# a_n1287_44306# 5.84e-19
C29430 a_n2661_42834# a_n875_44318# 1.15e-19
C29431 a_8953_45002# a_9885_43646# 1.33e-20
C29432 a_n3420_37984# VDD 0.930532f
C29433 a_13490_45067# VDD 6.34e-20
C29434 a_5932_42308# VIN_P 0.023512f
C29435 a_n356_44636# a_167_45260# 5.64e-19
C29436 a_5745_43940# a_5807_45002# 3.73e-21
C29437 a_14021_43940# a_n2293_46634# 0.202404f
C29438 a_20980_44850# a_19692_46634# 5.34e-20
C29439 a_1307_43914# a_n2661_45546# 0.021108f
C29440 a_6171_45002# a_n443_42852# 2.87e-20
C29441 a_9838_44484# a_9290_44172# 6.21e-19
C29442 a_8975_43940# a_8953_45546# 0.02155f
C29443 a_20107_42308# a_20712_42282# 0.008f
C29444 a_13258_32519# a_7174_31319# 0.02542f
C29445 a_5742_30871# comp_n 1.22e-19
C29446 a_19511_42282# a_21887_42336# 2.03e-19
C29447 a_22731_47423# VDD 0.196667f
C29448 a_n443_46116# a_n2661_45546# 0.136593f
C29449 a_584_46384# a_1848_45724# 3.13e-19
C29450 a_2553_47502# a_n755_45592# 8.3e-22
C29451 a_n971_45724# a_n906_45572# 0.001365f
C29452 a_4883_46098# a_8781_46436# 7.71e-20
C29453 a_14311_47204# a_13259_45724# 4.93e-21
C29454 a_768_44030# a_6945_45028# 0.014703f
C29455 a_2107_46812# a_6165_46155# 0.003422f
C29456 a_n2661_46634# a_12005_46116# 0.038027f
C29457 a_12891_46348# a_10809_44734# 0.102888f
C29458 a_n743_46660# a_9569_46155# 0.104962f
C29459 a_13661_43548# a_17715_44484# 0.003425f
C29460 a_13747_46662# a_17583_46090# 1.47e-19
C29461 a_5807_45002# a_18189_46348# 0.033239f
C29462 a_12816_46660# a_14180_46812# 5.52e-19
C29463 a_13607_46688# a_14035_46660# 0.003044f
C29464 a_14084_46812# a_13885_46660# 0.237373f
C29465 a_1057_46660# a_1176_45822# 1.55e-19
C29466 a_2443_46660# a_3147_46376# 5.77e-19
C29467 a_n913_45002# a_2713_42308# 0.291963f
C29468 a_n1059_45260# a_2903_42308# 0.003187f
C29469 a_n2017_45002# a_3318_42354# 0.01513f
C29470 a_11691_44458# a_16795_42852# 1.42e-19
C29471 a_10807_43548# a_11257_43940# 0.013221f
C29472 a_18494_42460# a_19164_43230# 5.14e-19
C29473 a_11827_44484# a_17333_42852# 3.3e-21
C29474 a_18184_42460# a_19987_42826# 0.208392f
C29475 a_11967_42832# a_13667_43396# 6.68e-20
C29476 a_3600_43914# a_4093_43548# 4.01e-19
C29477 a_2998_44172# a_4235_43370# 2.06e-20
C29478 a_n2293_42834# a_5193_42852# 2.39e-20
C29479 a_7845_44172# VDD 0.11772f
C29480 a_13904_45546# a_8696_44636# 5.54e-21
C29481 a_11823_42460# a_16223_45938# 3.12e-20
C29482 a_12427_45724# a_12561_45572# 0.001089f
C29483 a_10907_45822# a_12016_45572# 3.47e-20
C29484 a_17538_32519# a_21076_30879# 0.054805f
C29485 a_13460_43230# a_12891_46348# 1.83e-20
C29486 a_743_42282# a_4646_46812# 3.55e-19
C29487 a_13635_43156# a_12549_44172# 2.09e-20
C29488 a_16137_43396# a_6755_46942# 1.16e-19
C29489 a_7542_44172# a_8034_45724# 7e-22
C29490 a_14673_44172# a_n443_42852# 1.12e-19
C29491 a_3499_42826# a_526_44458# 0.089844f
C29492 a_11750_44172# a_10809_44734# 6e-21
C29493 a_10555_44260# a_10903_43370# 0.011277f
C29494 a_n1736_42282# SMPL_ON_P 5.11e-20
C29495 a_n784_42308# w_11334_34010# 0.001604f
C29496 a_15890_42674# CAL_N 6.88e-19
C29497 a_n4064_39616# a_n4064_37984# 0.048968f
C29498 a_4958_30871# a_n4064_37440# 0.031235f
C29499 a_n2157_46122# a_n1533_46116# 9.73e-19
C29500 a_n1641_46494# a_n1545_46494# 0.013793f
C29501 a_n1423_46090# a_n1379_46482# 3.69e-19
C29502 a_n1991_46122# a_n967_46494# 2.36e-20
C29503 a_21363_46634# a_8049_45260# 3.11e-20
C29504 a_13059_46348# a_14537_46482# 0.002353f
C29505 a_19692_46634# a_20692_30879# 4.77e-20
C29506 a_9625_46129# a_11133_46155# 4.63e-20
C29507 a_8147_43396# a_8685_43396# 0.077232f
C29508 a_n97_42460# a_18525_43370# 0.005868f
C29509 a_19319_43548# a_4190_30871# 0.188868f
C29510 a_7112_43396# a_7221_43396# 0.007416f
C29511 a_7287_43370# a_7466_43396# 0.007399f
C29512 a_3905_42865# a_5193_43172# 8.11e-19
C29513 a_10949_43914# a_5534_30871# 2.43e-20
C29514 SMPL_ON_N a_22821_38993# 2.28e-19
C29515 a_6575_47204# DATA[4] 0.15718f
C29516 a_13717_47436# RST_Z 4.51263f
C29517 a_16759_43396# VDD 0.191873f
C29518 a_n913_45002# a_9482_43914# 8.96e-20
C29519 a_2437_43646# a_2304_45348# 0.006164f
C29520 a_4558_45348# a_5147_45002# 0.09356f
C29521 a_3537_45260# a_4927_45028# 0.216859f
C29522 a_3065_45002# a_3232_43370# 0.049451f
C29523 a_4574_45260# a_5111_44636# 1.69e-19
C29524 a_9049_44484# a_9838_44484# 8.16e-19
C29525 a_7499_43078# a_10157_44484# 4.34e-20
C29526 a_15861_45028# a_16922_45042# 0.259169f
C29527 a_8696_44636# a_17023_45118# 0.064781f
C29528 a_10083_42826# a_4185_45028# 3.49e-20
C29529 a_21671_42860# a_20202_43084# 0.002893f
C29530 a_13667_43396# a_13259_45724# 0.160676f
C29531 a_766_43646# a_n443_42852# 8.62e-19
C29532 a_n3420_39616# a_n2312_40392# 6.3e-21
C29533 a_19237_31679# RST_Z 0.050685f
C29534 a_15143_45578# a_5807_45002# 3.06e-21
C29535 a_13249_42308# a_13747_46662# 0.134714f
C29536 a_8162_45546# a_n743_46660# 2.28e-21
C29537 a_7499_43078# a_n1925_46634# 9.19e-20
C29538 a_10490_45724# a_n2661_46634# 0.01771f
C29539 a_2211_45572# a_2107_46812# 3.18e-20
C29540 a_18479_45785# a_18597_46090# 0.009071f
C29541 a_18341_45572# a_18780_47178# 1.16e-20
C29542 a_17034_45572# a_16327_47482# 0.002231f
C29543 a_3357_43084# a_6545_47178# 0.005247f
C29544 a_2437_43646# a_7227_47204# 0.006315f
C29545 a_20623_45572# a_12861_44030# 7.98e-22
C29546 a_n2017_45002# a_n1151_42308# 0.058036f
C29547 a_1667_45002# a_n746_45260# 2.7e-22
C29548 a_2274_45254# a_n971_45724# 0.002827f
C29549 a_4558_45348# a_n2109_47186# 5.21e-20
C29550 a_5111_44636# a_n2497_47436# 8.27e-21
C29551 a_20205_31679# a_20850_46155# 4.73e-21
C29552 a_10425_46660# CLK 1.87e-19
C29553 a_n1557_42282# a_n4318_38216# 2.95e-20
C29554 a_n3674_39768# a_n4064_39616# 0.464693f
C29555 a_4190_30871# a_16795_42852# 3.12e-21
C29556 a_743_42282# a_15567_42826# 7.68e-20
C29557 a_5649_42852# a_13113_42826# 3.48e-21
C29558 a_1209_43370# a_n784_42308# 3.67e-21
C29559 a_18079_43940# a_18057_42282# 3.16e-21
C29560 a_14035_46660# RST_Z 1.33e-19
C29561 a_2113_38308# a_3726_37500# 1.83e-19
C29562 a_7754_38968# VDAC_Ni 1.16e-19
C29563 a_1067_42314# VDD 0.128996f
C29564 a_n2833_47464# a_n1741_47186# 3.87e-20
C29565 a_n2497_47436# a_n1920_47178# 0.049461f
C29566 a_n2288_47178# a_n2109_47186# 0.177673f
C29567 a_10775_45002# a_n2661_42834# 1.02e-20
C29568 a_11823_42460# a_11341_43940# 0.087329f
C29569 a_n2661_43370# a_10334_44484# 7.92e-20
C29570 a_14537_43396# a_9313_44734# 1.05e-20
C29571 a_1423_45028# a_5289_44734# 0.002441f
C29572 a_21005_45260# a_18114_32519# 6.8e-20
C29573 a_8953_45002# a_n2661_43922# 5.04e-19
C29574 a_22223_45572# a_3422_30871# 2.45e-20
C29575 a_22465_38105# a_21076_30879# 6.77e-19
C29576 a_3318_42354# a_526_44458# 3.31e-19
C29577 a_2903_42308# a_n1925_42282# 1.31e-19
C29578 a_8292_43218# a_n443_42852# 0.002007f
C29579 a_13657_42558# a_9290_44172# 4.35e-20
C29580 a_13575_42558# a_10903_43370# 8.65e-20
C29581 a_15599_45572# a_12741_44636# 3.13e-19
C29582 a_16333_45814# a_11415_45002# 0.00197f
C29583 a_n2661_43370# a_n1021_46688# 1.67e-22
C29584 a_18341_45572# a_18285_46348# 2.47e-21
C29585 a_17613_45144# a_13747_46662# 1.85e-20
C29586 a_18315_45260# a_5807_45002# 5.54e-21
C29587 a_17719_45144# a_13661_43548# 2.08e-20
C29588 a_16922_45042# a_19321_45002# 0.493823f
C29589 a_11827_44484# a_768_44030# 0.831344f
C29590 a_22223_45036# a_12549_44172# 8.25e-20
C29591 a_18479_45785# a_19123_46287# 3.74e-20
C29592 a_3357_43084# a_19692_46634# 0.046179f
C29593 a_10490_45724# a_8199_44636# 0.019372f
C29594 a_3775_45552# a_2324_44458# 6.98e-21
C29595 a_8746_45002# a_5937_45572# 0.121678f
C29596 a_10180_45724# a_9625_46129# 0.00231f
C29597 a_10193_42453# a_8953_45546# 6e-19
C29598 a_8333_44734# a_4791_45118# 4.95e-19
C29599 a_n89_44484# a_n1151_42308# 0.007033f
C29600 a_6109_44484# a_6151_47436# 1.83e-20
C29601 a_16979_44734# a_16327_47482# 4.27e-19
C29602 a_18443_44721# a_11599_46634# 1.76e-20
C29603 a_13076_44458# a_10227_46804# 1.5e-19
C29604 a_6298_44484# a_4883_46098# 9.77e-21
C29605 a_21487_43396# a_13258_32519# 9.88e-21
C29606 a_10083_42826# a_9803_42558# 0.006054f
C29607 a_n2293_42282# a_1606_42308# 0.192228f
C29608 a_743_42282# a_20712_42282# 0.001163f
C29609 a_13467_32519# a_19511_42282# 0.003538f
C29610 a_4361_42308# a_18548_42308# 5.09e-19
C29611 a_20205_31679# VREF 0.056031f
C29612 a_20692_30879# VIN_N 0.039f
C29613 a_2063_45854# a_5257_43370# 0.426517f
C29614 a_n237_47217# a_10150_46912# 2.7e-19
C29615 a_n1741_47186# a_6969_46634# 7.57e-20
C29616 a_4791_45118# a_5167_46660# 0.008966f
C29617 a_4915_47217# a_4817_46660# 2.69e-19
C29618 a_5815_47464# a_4651_46660# 0.001772f
C29619 a_6151_47436# a_4646_46812# 0.153739f
C29620 a_6545_47178# a_3877_44458# 0.026367f
C29621 a_22731_47423# a_22612_30879# 9.38e-19
C29622 SMPL_ON_N a_21588_30879# 0.119129f
C29623 a_11453_44696# a_20916_46384# 0.021978f
C29624 a_8128_46384# a_9804_47204# 0.001612f
C29625 a_n881_46662# a_12891_46348# 0.026595f
C29626 a_3537_45260# a_4699_43561# 0.024682f
C29627 a_n1059_45260# a_6293_42852# 0.002519f
C29628 a_n913_45002# a_6031_43396# 2.91e-20
C29629 a_n2017_45002# a_6197_43396# 4.71e-20
C29630 a_3065_45002# a_4905_42826# 2.38e-20
C29631 a_n967_45348# a_n998_43396# 4.97e-19
C29632 a_3357_43084# a_3457_43396# 5.15e-19
C29633 a_4558_45348# a_4093_43548# 9.14e-21
C29634 a_15861_45028# a_15743_43084# 1.08e-20
C29635 a_5883_43914# a_5244_44056# 1.47e-19
C29636 a_15146_44811# a_14673_44172# 0.001224f
C29637 a_16922_45042# a_20623_43914# 0.001335f
C29638 a_11827_44484# a_13483_43940# 5.96e-19
C29639 a_5343_44458# a_7281_43914# 8.75e-20
C29640 a_9313_44734# a_20835_44721# 4.17e-21
C29641 a_11691_44458# a_10949_43914# 4.22e-20
C29642 a_n4209_38216# a_n2956_38216# 0.232905f
C29643 a_7276_45260# VDD 0.093163f
C29644 a_19721_31679# a_21076_30879# 0.05488f
C29645 a_9313_44734# a_3090_45724# 2.43867f
C29646 a_5013_44260# a_n2293_46634# 3.03e-20
C29647 a_6756_44260# a_768_44030# 3.81e-19
C29648 a_n1059_45260# a_16375_45002# 0.001787f
C29649 a_n2661_43370# a_9290_44172# 0.185465f
C29650 a_15493_43940# SMPL_ON_N 1.94e-20
C29651 a_15301_44260# a_10227_46804# 2.48e-19
C29652 a_14021_43940# a_18597_46090# 0.0185f
C29653 a_3080_42308# w_11334_34010# 0.001073f
C29654 a_n1821_43396# a_n971_45724# 2.41e-20
C29655 a_n746_45260# VDD 1.41433f
C29656 a_n3674_38216# a_n4064_39072# 0.019725f
C29657 a_5742_30871# a_11633_42308# 0.001223f
C29658 a_5932_42308# a_13258_32519# 5.13e-19
C29659 a_n4318_37592# a_n3420_39072# 0.02033f
C29660 a_14456_42282# a_15803_42450# 5.2e-21
C29661 VIN_P VREF 0.775904f
C29662 a_10150_46912# a_8270_45546# 4.81e-19
C29663 a_33_46660# a_765_45546# 4.44e-20
C29664 a_8492_46660# a_8601_46660# 0.007416f
C29665 a_8667_46634# a_8846_46660# 0.007399f
C29666 a_19594_46812# a_19636_46660# 0.009543f
C29667 a_n881_46662# a_805_46414# 0.011286f
C29668 a_n1613_43370# a_1208_46090# 0.002092f
C29669 a_4883_46098# a_5937_45572# 0.015486f
C29670 a_11599_46634# a_17583_46090# 0.031836f
C29671 a_10227_46804# a_12594_46348# 0.001992f
C29672 a_15811_47375# a_2324_44458# 0.001263f
C29673 a_15507_47210# a_15682_46116# 3.39e-19
C29674 a_12861_44030# a_18819_46122# 0.001599f
C29675 a_13717_47436# a_18985_46122# 1.33e-21
C29676 a_9067_47204# a_6945_45028# 0.014009f
C29677 a_n971_45724# a_8034_45724# 0.027525f
C29678 a_n1151_42308# a_526_44458# 0.003737f
C29679 a_n237_47217# a_8062_46482# 0.001342f
C29680 a_3160_47472# a_n1925_42282# 2.98e-19
C29681 a_2063_45854# a_1337_46116# 4.29e-19
C29682 a_16979_44734# a_10341_43396# 8.24e-21
C29683 a_1467_44172# a_1241_43940# 0.011879f
C29684 a_9672_43914# a_10405_44172# 4.63e-19
C29685 a_20835_44721# a_20974_43370# 5.58e-21
C29686 a_20193_45348# a_21487_43396# 5.6e-20
C29687 a_n2293_42834# a_7227_42852# 0.008564f
C29688 a_10193_42453# a_14456_42282# 0.001037f
C29689 a_1115_44172# a_1443_43940# 0.096132f
C29690 a_18579_44172# a_19478_44056# 2.74e-19
C29691 a_5891_43370# a_6452_43396# 1.68e-20
C29692 a_11823_42460# a_10723_42308# 3.49e-19
C29693 a_2711_45572# a_18907_42674# 2.61e-19
C29694 a_n1059_45260# a_11554_42852# 0.002165f
C29695 a_17517_44484# VDD 2.99662f
C29696 a_2711_45572# a_9241_45822# 1.37e-19
C29697 a_6194_45824# a_6469_45572# 0.007416f
C29698 a_8568_45546# a_9049_44484# 4.21e-19
C29699 a_15493_43396# a_11415_45002# 1.63e-20
C29700 a_n2661_42282# a_1138_42852# 1.46e-20
C29701 a_15743_43084# a_19321_45002# 6.69e-20
C29702 a_3457_43396# a_3877_44458# 3.97e-22
C29703 a_n356_44636# a_n863_45724# 0.301674f
C29704 a_12607_44458# a_n443_42852# 4.46e-20
C29705 a_5663_43940# a_5937_45572# 0.177912f
C29706 a_n901_43156# a_n2312_40392# 1.65e-20
C29707 a_n1059_45260# RST_Z 3.96e-20
C29708 a_19479_31679# VREF 0.056254f
C29709 a_n4064_39616# C0_P_btm 3.27e-20
C29710 a_n1630_35242# VDAC_P 0.00281f
C29711 a_11415_45002# a_3483_46348# 0.057381f
C29712 a_n2293_46098# a_1208_46090# 0.002845f
C29713 a_n1853_46287# a_472_46348# 1.54e-20
C29714 a_n1423_46090# a_n1076_46494# 0.051162f
C29715 a_12359_47026# a_10809_44734# 0.010386f
C29716 a_13059_46348# a_2324_44458# 0.0606f
C29717 a_n743_46660# a_1990_45899# 5.84e-19
C29718 a_n2661_46098# a_n357_42282# 6.61e-20
C29719 a_8035_47026# a_8049_45260# 6.19e-20
C29720 a_171_46873# a_n443_42852# 5.11e-19
C29721 a_1799_45572# a_n755_45592# 0.024036f
C29722 a_n2438_43548# a_2277_45546# 9.99e-20
C29723 a_n2956_37592# a_n3420_38528# 6.26e-20
C29724 a_14021_43940# a_14537_43646# 0.001553f
C29725 a_n2661_42282# a_5649_42852# 0.052118f
C29726 a_2479_44172# a_3681_42891# 1.73e-19
C29727 a_n97_42460# a_3540_43646# 0.027089f
C29728 a_3422_30871# a_5534_30871# 0.023427f
C29729 a_n4318_39768# a_n3674_39304# 0.024426f
C29730 a_19279_43940# a_18249_42858# 5.33e-20
C29731 a_11341_43940# a_18429_43548# 2.54e-20
C29732 a_15493_43940# a_17499_43370# 2.64e-19
C29733 a_20623_43914# a_15743_43084# 1.72e-20
C29734 a_10405_44172# a_743_42282# 1.09e-20
C29735 a_2889_44172# a_1847_42826# 6.94e-19
C29736 a_2675_43914# a_2075_43172# 3.57e-20
C29737 a_9313_44734# a_12991_43230# 2.5e-19
C29738 w_1575_34946# a_n923_35174# 37.7438f
C29739 a_15037_45618# a_14537_43396# 3.1e-20
C29740 a_15599_45572# a_13556_45296# 7.13e-22
C29741 a_8696_44636# a_10951_45334# 0.001322f
C29742 a_9049_44484# a_n2661_43370# 0.030026f
C29743 a_19479_31679# a_22591_45572# 0.011797f
C29744 a_21513_45002# a_20447_31679# 4.16e-20
C29745 a_22223_45572# a_19963_31679# 0.00254f
C29746 a_17364_32525# a_20820_30879# 0.055604f
C29747 a_n784_42308# a_n2442_46660# 3.54e-19
C29748 a_16795_42852# a_15227_44166# 3.87e-19
C29749 a_6197_43396# a_526_44458# 5.62e-19
C29750 a_5829_43940# a_n357_42282# 3.11e-19
C29751 a_15095_43370# a_2324_44458# 5.95e-19
C29752 a_7227_42308# a_n1613_43370# 0.001156f
C29753 a_15720_42674# a_10227_46804# 1.7e-19
C29754 a_n4064_39072# w_1575_34946# 0.016546f
C29755 a_12379_46436# VDD 0.002681f
C29756 a_9241_45822# a_9313_45822# 7.24e-19
C29757 a_11322_45546# a_10227_46804# 6.46e-22
C29758 a_13249_42308# a_11599_46634# 4.64e-20
C29759 a_11823_42460# a_16327_47482# 1.03e-20
C29760 a_2324_44458# a_3218_45724# 1.93e-20
C29761 a_10903_43370# a_n443_42852# 0.176275f
C29762 a_10695_43548# a_10835_43094# 5.89e-20
C29763 a_n97_42460# a_7309_42852# 0.024142f
C29764 a_16823_43084# a_5649_42852# 6.08e-21
C29765 a_3422_30871# a_19647_42308# 6.32e-20
C29766 a_4190_30871# a_19095_43396# 0.046015f
C29767 a_743_42282# a_20556_43646# 0.028541f
C29768 a_3539_42460# a_n2293_42282# 0.010651f
C29769 a_4149_42891# VDD 0.001563f
C29770 a_5111_44636# a_5883_43914# 0.281106f
C29771 a_3232_43370# a_6298_44484# 0.256727f
C29772 a_n2293_45010# a_n356_44636# 0.031375f
C29773 a_5205_44484# a_4743_44484# 8.65e-19
C29774 a_7229_43940# a_4223_44672# 0.014299f
C29775 a_n2017_45002# a_n1821_44484# 0.001578f
C29776 a_3357_43084# a_5826_44734# 2.81e-19
C29777 a_8696_44636# a_17061_44484# 3.53e-19
C29778 a_9482_43914# a_n2661_44458# 0.017706f
C29779 a_16333_45814# a_11967_42832# 2.46e-21
C29780 a_5379_42460# a_1823_45246# 1.01e-20
C29781 a_3681_42891# a_n443_42852# 1.37e-20
C29782 a_10835_43094# a_n357_42282# 0.02434f
C29783 a_21195_42852# a_13259_45724# 1.73e-20
C29784 a_13527_45546# a_13059_46348# 0.017655f
C29785 a_15037_45618# a_3090_45724# 8.98e-19
C29786 a_1307_43914# a_12891_46348# 0.008663f
C29787 a_16019_45002# a_12549_44172# 8.08e-21
C29788 a_13017_45260# a_5807_45002# 4.58e-19
C29789 a_3357_43084# a_3877_44458# 0.02473f
C29790 a_3537_45260# a_n743_46660# 4.3e-20
C29791 a_6171_45002# a_n2661_46634# 0.042529f
C29792 a_2437_43646# a_4955_46873# 1.65e-19
C29793 a_17613_45144# a_11599_46634# 4.99e-21
C29794 a_15060_45348# a_10227_46804# 3.31e-19
C29795 a_18911_45144# a_12861_44030# 0.169f
C29796 EN_VIN_BSTR_N VDD 1.13406f
C29797 a_n699_43396# a_n746_45260# 0.002245f
C29798 a_4223_44672# a_n237_47217# 2.68e-21
C29799 a_15567_42826# a_16328_43172# 1.3e-20
C29800 a_13460_43230# a_13622_42852# 0.006453f
C29801 a_15681_43442# a_15051_42282# 1.21e-19
C29802 a_743_42282# a_6171_42473# 0.007484f
C29803 a_15781_43660# a_14113_42308# 2.97e-21
C29804 a_4361_42308# a_4933_42558# 4.55e-21
C29805 a_1239_39043# VDD 0.507578f
C29806 a_4915_47217# a_11309_47204# 0.045252f
C29807 a_6151_47436# a_9804_47204# 0.095181f
C29808 a_7903_47542# a_n881_46662# 0.178742f
C29809 a_6545_47178# a_8128_46384# 5.48e-21
C29810 a_6575_47204# a_n1613_43370# 0.005913f
C29811 a_n2109_47186# a_n2312_38680# 4.37e-19
C29812 a_n1920_47178# a_n2104_46634# 3.21e-19
C29813 a_n815_47178# a_n2661_46634# 0.003247f
C29814 a_2063_45854# a_5807_45002# 0.074286f
C29815 SMPL_ON_P a_n2442_46660# 0.092029f
C29816 a_n2497_47436# a_n1021_46688# 9.22e-19
C29817 a_10227_46804# a_12465_44636# 0.057431f
C29818 a_19787_47423# a_20990_47178# 4.61e-20
C29819 a_18597_46090# a_13507_46334# 0.093881f
C29820 a_18479_47436# a_4883_46098# 0.038695f
C29821 a_11823_42460# a_10341_43396# 0.088285f
C29822 a_13249_42308# a_14358_43442# 1.53e-20
C29823 a_n2661_43370# a_3905_42865# 6.49e-20
C29824 a_1423_45028# a_9028_43914# 7.39e-20
C29825 a_1307_43914# a_11750_44172# 0.007207f
C29826 a_13720_44458# a_14112_44734# 0.016359f
C29827 a_10057_43914# a_10809_44484# 2.31e-19
C29828 a_n356_44636# a_9313_44734# 2.11e-20
C29829 a_11827_44484# a_21073_44484# 7.17e-19
C29830 a_18114_32519# a_20835_44721# 9.39e-20
C29831 a_15959_42545# a_n443_42852# 1.56e-19
C29832 a_19256_45572# VDD 0.27151f
C29833 a_5534_30871# VREF_GND 0.060532f
C29834 a_19987_42826# RST_Z 8.97e-21
C29835 a_5342_30871# VIN_N 0.00693f
C29836 a_13159_45002# a_3483_46348# 0.017316f
C29837 a_18588_44850# a_13661_43548# 0.005669f
C29838 a_4223_44672# a_8270_45546# 1.84e-19
C29839 a_17801_45144# a_15227_44166# 8.12e-20
C29840 a_16333_45814# a_13259_45724# 0.02201f
C29841 a_15599_45572# a_16375_45002# 1.1e-19
C29842 a_18479_45785# a_8049_45260# 0.0037f
C29843 a_22959_45572# a_22959_46124# 0.025171f
C29844 a_20447_31679# a_10809_44734# 0.005556f
C29845 a_3232_43370# a_5937_45572# 0.662525f
C29846 a_6171_45002# a_8199_44636# 0.163434f
C29847 a_413_45260# a_13925_46122# 9.96e-21
C29848 a_1576_42282# a_5742_30871# 2.87e-20
C29849 a_5755_42308# a_6171_42473# 0.017801f
C29850 a_5379_42460# a_5934_30871# 5.78e-20
C29851 a_n784_42308# a_14456_42282# 3.86e-20
C29852 a_3823_42558# a_3905_42308# 0.003935f
C29853 a_5421_42558# a_5932_42308# 6.5e-19
C29854 a_17364_32525# C8_N_btm 7.96e-19
C29855 a_22717_37285# a_22717_36887# 0.003901f
C29856 a_2063_45854# a_3699_46348# 0.002997f
C29857 a_3160_47472# a_2698_46116# 4.19e-19
C29858 a_2905_45572# a_2804_46116# 3.04e-19
C29859 a_n443_46116# a_805_46414# 9.4e-20
C29860 a_2952_47436# a_3147_46376# 1.09e-19
C29861 a_n1151_42308# a_2521_46116# 2.53e-20
C29862 a_3815_47204# a_1823_45246# 6.25e-21
C29863 a_584_46384# a_4185_45028# 5.71e-19
C29864 a_n237_47217# a_6419_46155# 0.029086f
C29865 a_n1741_47186# a_9625_46129# 6.6e-20
C29866 a_n971_45724# a_8016_46348# 0.029312f
C29867 a_13507_46334# a_19123_46287# 0.034113f
C29868 a_20990_47178# a_20107_46660# 2.98e-20
C29869 a_10227_46804# a_20528_46660# 1.1e-20
C29870 a_12465_44636# a_17339_46660# 6.05e-22
C29871 a_11453_44696# a_16751_46987# 1.13e-21
C29872 a_3177_46902# a_3633_46660# 4.2e-19
C29873 a_n743_46660# a_6969_46634# 1.5e-19
C29874 a_2107_46812# a_8492_46660# 2.24e-20
C29875 a_5807_45002# a_12469_46902# 0.003304f
C29876 a_12549_44172# a_16292_46812# 0.013094f
C29877 a_2382_45260# a_3935_42891# 0.061675f
C29878 a_n913_45002# a_10796_42968# 0.545674f
C29879 a_n1059_45260# a_10991_42826# 0.004257f
C29880 a_n2017_45002# a_10922_42852# 1.02e-20
C29881 a_n699_43396# a_1891_43646# 4.33e-19
C29882 a_1307_43914# a_4361_42308# 7.03e-21
C29883 a_n1899_43946# a_n1441_43940# 0.03441f
C29884 a_2998_44172# a_3905_42865# 3.52e-19
C29885 a_n2661_44458# a_6031_43396# 5.36e-21
C29886 a_742_44458# a_3540_43646# 1.09e-20
C29887 a_16979_44734# a_n97_42460# 1.23e-21
C29888 a_19615_44636# a_19328_44172# 3.27e-21
C29889 a_11967_42832# a_15493_43396# 0.02628f
C29890 a_2779_44458# a_2896_43646# 6.83e-21
C29891 a_13720_44458# VDD 0.202097f
C29892 a_n3565_39590# C9_P_btm 0.001137f
C29893 a_n4064_40160# C3_P_btm 1.27e-19
C29894 a_n4209_39304# a_n1838_35608# 2.06e-19
C29895 a_13258_32519# VREF 9.37e-19
C29896 a_11967_42832# a_3483_46348# 0.264293f
C29897 a_19237_31679# a_20820_30879# 0.053048f
C29898 a_17737_43940# a_3090_45724# 3.24e-20
C29899 a_14021_43940# a_6755_46942# 2.04e-19
C29900 a_1209_43370# a_n2438_43548# 8.21e-21
C29901 a_4699_43561# a_n2293_46634# 0.006722f
C29902 a_8147_43396# a_768_44030# 2.39e-22
C29903 a_n1557_42282# a_n2956_39768# 2.12e-20
C29904 a_3080_42308# a_n2442_46660# 4.94e-21
C29905 a_10057_43914# a_8049_45260# 5.59e-20
C29906 a_13857_44734# a_13759_46122# 2.43e-22
C29907 a_6643_43396# a_n1613_43370# 2.72e-19
C29908 a_16409_43396# a_10227_46804# 6.95e-19
C29909 a_18429_43548# a_16327_47482# 0.057366f
C29910 a_791_42968# a_n2497_47436# 2.18e-21
C29911 a_383_46660# VDD 0.198466f
C29912 a_n4209_39590# a_n3565_38502# 0.031792f
C29913 a_n4334_39392# a_n3565_39304# 0.001004f
C29914 a_n3565_39590# a_n4209_38502# 0.0315f
C29915 a_n4064_40160# a_n4064_38528# 0.055466f
C29916 a_n4209_39304# a_n3690_39392# 0.045342f
C29917 a_5742_30871# C1_P_btm 0.026156f
C29918 a_14513_46634# a_11415_45002# 2.15e-20
C29919 a_20107_46660# a_20273_46660# 0.608339f
C29920 a_19123_46287# a_20623_46660# 1.73e-20
C29921 a_3177_46902# a_526_44458# 0.001189f
C29922 a_5807_45002# a_14383_46116# 0.007691f
C29923 a_6755_46942# a_11133_46155# 1.21e-19
C29924 a_7577_46660# a_2324_44458# 1.05e-20
C29925 a_n1613_43370# a_n2661_45546# 0.029057f
C29926 a_2747_46873# a_n755_45592# 1.74e-20
C29927 a_n3674_38680# a_n3690_38304# 3.4e-19
C29928 a_4883_46098# a_n443_42852# 0.074259f
C29929 a_11341_43940# a_2982_43646# 0.002145f
C29930 a_18579_44172# a_4361_42308# 6.73e-20
C29931 a_3422_30871# a_4190_30871# 12.909901f
C29932 a_9159_44484# a_9127_43156# 7.52e-21
C29933 a_n2661_43922# a_8037_42858# 4.47e-22
C29934 a_n2293_43922# a_7765_42852# 1.03e-20
C29935 a_9313_44734# a_12379_42858# 0.05039f
C29936 a_n2293_42834# a_1576_42282# 5e-20
C29937 a_n1059_45260# a_17303_42282# 0.001091f
C29938 a_n2017_45002# a_17531_42308# 0.00607f
C29939 a_n913_45002# a_4958_30871# 0.058702f
C29940 a_726_44056# VDD 0.001151f
C29941 a_8162_45546# a_5111_44636# 1.13e-21
C29942 a_17478_45572# a_17568_45572# 0.008441f
C29943 a_2711_45572# a_14537_43396# 0.249285f
C29944 a_15861_45028# a_17668_45572# 0.065471f
C29945 a_n4064_37440# C3_P_btm 1.74e-19
C29946 a_743_42282# a_19692_46634# 0.150479f
C29947 a_16409_43396# a_17339_46660# 4.94e-20
C29948 a_5663_43940# a_n443_42852# 3.4e-21
C29949 a_15493_43396# a_13259_45724# 0.021264f
C29950 a_n2661_42282# a_n2956_38216# 3.02e-20
C29951 a_1241_44260# a_n357_42282# 3.97e-19
C29952 a_13351_46090# VDD 0.238036f
C29953 a_6511_45714# a_2063_45854# 0.037319f
C29954 a_4099_45572# a_n1151_42308# 9.09e-21
C29955 a_2711_45572# a_3785_47178# 1.05e-20
C29956 a_3260_45572# a_n237_47217# 6.54e-22
C29957 a_n4064_38528# a_n4064_37440# 0.045121f
C29958 a_8199_44636# a_9751_46155# 7.99e-20
C29959 a_9625_46129# a_10586_45546# 9.22e-19
C29960 a_11133_46155# a_8049_45260# 0.001208f
C29961 a_n2956_39304# a_n1379_46482# 9.59e-21
C29962 a_n2840_46090# a_n2956_38216# 0.004667f
C29963 a_n2293_46098# a_n2661_45546# 3.03243f
C29964 a_n2472_46090# a_n2472_45546# 0.025171f
C29965 a_3483_46348# a_13259_45724# 0.230226f
C29966 a_8685_43396# a_16823_43084# 7.39e-20
C29967 a_1414_42308# a_n1630_35242# 2.24e-20
C29968 a_1568_43370# a_791_42968# 4.67e-20
C29969 a_9145_43396# a_15231_43396# 0.005861f
C29970 a_9313_44734# a_18727_42674# 2.59e-20
C29971 a_1115_44172# a_1576_42282# 2.71e-21
C29972 a_453_43940# a_564_42282# 4.63e-21
C29973 a_15095_43370# a_15743_43084# 0.022008f
C29974 a_n97_42460# a_7765_42852# 0.002083f
C29975 a_10341_43396# a_18429_43548# 0.012565f
C29976 a_9396_43370# a_4361_42308# 3.82e-20
C29977 a_10037_47542# CLK 2.34e-19
C29978 a_11309_47204# DATA[5] 0.080873f
C29979 a_5111_42852# VDD 0.178652f
C29980 a_17478_45572# a_17767_44458# 6.59e-21
C29981 a_8192_45572# a_8375_44464# 1.55e-21
C29982 a_11823_42460# a_n2293_43922# 0.494696f
C29983 a_626_44172# a_1145_45348# 0.009374f
C29984 a_8696_44636# a_18248_44752# 7.61e-21
C29985 a_5147_45002# a_n2661_43370# 0.034793f
C29986 a_7229_43940# a_n2293_42834# 0.148023f
C29987 a_20447_31679# a_22959_45036# 4.88e-19
C29988 a_n2017_45002# a_18184_42460# 0.205351f
C29989 a_6709_45028# a_7639_45394# 0.004982f
C29990 a_3232_43370# a_7418_45067# 0.001221f
C29991 a_6171_45002# a_10903_45394# 5.41e-20
C29992 a_20256_43172# a_20202_43084# 0.006261f
C29993 a_8515_42308# a_3090_45724# 1.5e-21
C29994 a_n3565_39304# a_n2312_38680# 0.418567f
C29995 a_16243_43396# a_n443_42852# 0.001298f
C29996 a_10922_42852# a_526_44458# 2.42e-20
C29997 a_10180_45724# a_6755_46942# 4.84e-20
C29998 a_2711_45572# a_3090_45724# 0.555348f
C29999 a_10193_42453# a_10249_46116# 0.034764f
C30000 a_10490_45724# a_10623_46897# 3.15e-20
C30001 a_20107_45572# a_5807_45002# 4.31e-21
C30002 a_16842_45938# a_n743_46660# 1.64e-19
C30003 a_18953_45572# a_13661_43548# 5.68e-19
C30004 a_2437_43646# a_11117_47542# 5.27e-19
C30005 a_3357_43084# a_8128_46384# 5.77e-20
C30006 a_8488_45348# a_n971_45724# 0.001106f
C30007 a_n2293_42834# a_n237_47217# 0.002403f
C30008 a_2809_45348# a_n443_46116# 0.001393f
C30009 a_n2661_43370# a_n2109_47186# 0.008032f
C30010 a_13348_45260# a_12861_44030# 2.51e-20
C30011 a_11787_45002# a_11599_46634# 1.65e-20
C30012 a_413_45260# SMPL_ON_N 0.199669f
C30013 a_2982_43646# a_10723_42308# 2.53e-19
C30014 a_19319_43548# a_19511_42282# 1.71e-21
C30015 a_2905_42968# a_2987_42968# 0.004999f
C30016 a_15279_43071# a_15567_42826# 7.4e-20
C30017 a_n97_42460# a_13657_42308# 0.005924f
C30018 a_15743_43084# a_14097_32519# 0.001681f
C30019 a_4190_30871# a_18504_43218# 9.82e-19
C30020 a_17730_32519# C10_N_btm 7.64e-19
C30021 a_19237_31679# C8_N_btm 1.71e-20
C30022 a_6151_47436# a_6545_47178# 0.39775f
C30023 a_4915_47217# a_7227_47204# 0.059062f
C30024 a_5815_47464# a_6491_46660# 0.003594f
C30025 a_3160_47472# a_n1435_47204# 5e-19
C30026 a_4791_45118# a_6575_47204# 8.32e-20
C30027 a_n1151_42308# a_13381_47204# 7.76e-20
C30028 a_3537_45260# a_5244_44056# 6.11e-20
C30029 a_5147_45002# a_2998_44172# 7.85e-20
C30030 a_3232_43370# a_2479_44172# 0.003118f
C30031 a_n2661_44458# a_n1809_44850# 0.003338f
C30032 a_11823_42460# a_n97_42460# 0.324041f
C30033 a_n2433_44484# a_n2012_44484# 0.093133f
C30034 a_n39_42308# a_n357_42282# 0.001655f
C30035 a_n327_42308# a_n755_45592# 7.83e-20
C30036 a_7174_31319# a_n2956_39304# 4.27e-21
C30037 a_11525_45546# VDD 0.133093f
C30038 a_4190_30871# VREF_GND 0.105109f
C30039 a_22959_43396# RST_Z 0.001326f
C30040 a_9482_43914# a_14035_46660# 8.69e-20
C30041 a_18443_44721# a_13661_43548# 0.011774f
C30042 a_n2433_44484# a_n2661_46098# 5.13e-22
C30043 a_12607_44458# a_n2661_46634# 1.26e-19
C30044 a_18287_44626# a_13747_46662# 1.75e-20
C30045 a_10440_44484# a_n2293_46634# 3.4e-20
C30046 a_17970_44736# a_19321_45002# 1.04e-21
C30047 a_n2293_42834# a_8270_45546# 1.57e-20
C30048 a_949_44458# a_2107_46812# 8.97e-21
C30049 a_10180_45724# a_8049_45260# 0.002472f
C30050 a_16680_45572# a_15682_46116# 0.006985f
C30051 a_8696_44636# a_2324_44458# 0.033373f
C30052 a_13485_45572# a_10903_43370# 0.001122f
C30053 a_16115_45572# a_17715_44484# 6.11e-20
C30054 a_n2661_43922# a_n2312_40392# 1.45e-20
C30055 a_n2661_42834# a_n2312_39304# 6.52e-20
C30056 a_14815_43914# a_12465_44636# 3.16e-19
C30057 a_16241_44734# a_10227_46804# 4.02e-19
C30058 a_19615_44636# a_12861_44030# 0.094785f
C30059 a_1467_44172# a_n746_45260# 9.96e-21
C30060 a_1414_42308# a_n971_45724# 4.43e-21
C30061 a_n1761_44111# a_584_46384# 1.76e-20
C30062 a_17333_42852# a_18214_42558# 0.00105f
C30063 a_18249_42858# a_19332_42282# 4.14e-19
C30064 a_19987_42826# a_17303_42282# 5.3e-20
C30065 COMP_P a_n961_42308# 0.001912f
C30066 a_18599_43230# a_18727_42674# 1e-19
C30067 a_18817_42826# a_18907_42674# 7.77e-19
C30068 a_n4318_38216# a_n3674_37592# 0.077253f
C30069 a_n3674_38680# a_n1630_35242# 0.020981f
C30070 a_n3674_38216# a_n784_42308# 0.001581f
C30071 a_5534_30871# a_7174_31319# 0.038837f
C30072 a_14097_32519# a_1606_42308# 2.3e-20
C30073 a_n2293_46634# a_n743_46660# 0.001475f
C30074 a_n2661_46634# a_171_46873# 0.007801f
C30075 a_n2312_38680# a_n1925_46634# 0.004049f
C30076 a_n2442_46660# a_n2438_43548# 0.002667f
C30077 a_n881_46662# a_4817_46660# 1.02e-19
C30078 a_8128_46384# a_3877_44458# 1.82e-21
C30079 a_n1613_43370# a_5385_46902# 0.182522f
C30080 a_13507_46334# a_6755_46942# 0.075659f
C30081 a_4883_46098# a_10554_47026# 1.36e-20
C30082 a_11599_46634# a_11813_46116# 0.106062f
C30083 a_12861_44030# a_12991_46634# 0.001474f
C30084 a_4915_47217# a_12156_46660# 7.15e-20
C30085 a_n1435_47204# a_13607_46688# 7.18e-19
C30086 a_n1151_42308# a_13170_46660# 1.42e-19
C30087 a_9482_43914# a_9145_43396# 5.35e-19
C30088 a_8696_44636# a_8387_43230# 7.22e-21
C30089 a_18989_43940# a_15493_43396# 2.4e-19
C30090 a_20679_44626# a_22591_44484# 4.6e-21
C30091 a_n2293_43922# a_n1644_44306# 1.12e-19
C30092 a_14539_43914# a_11341_43940# 0.077754f
C30093 a_n356_44636# a_17737_43940# 3.52e-21
C30094 a_13017_45260# a_13667_43396# 1.23e-20
C30095 a_19279_43940# a_21145_44484# 0.004519f
C30096 a_5891_43370# a_7911_44260# 2.91e-19
C30097 a_n2661_43922# a_n1453_44318# 0.001188f
C30098 a_11827_44484# a_21205_44306# 4.85e-19
C30099 a_n2661_42834# a_n1287_44306# 6.06e-19
C30100 a_n699_43396# a_726_44056# 7.74e-20
C30101 a_3357_43084# a_743_42282# 1.72e-19
C30102 a_n3690_38304# VDD 0.363068f
C30103 a_9313_44734# a_21076_30879# 1.55e-20
C30104 a_3422_30871# a_15227_44166# 2.1e-20
C30105 a_3232_43370# a_n443_42852# 0.02112f
C30106 a_8975_43940# a_5937_45572# 6.52e-19
C30107 a_5883_43914# a_9290_44172# 0.026946f
C30108 a_10057_43914# a_8953_45546# 1.06e-19
C30109 a_2982_43646# a_16327_47482# 0.030062f
C30110 a_19647_42308# a_7174_31319# 0.006018f
C30111 a_13258_32519# a_20712_42282# 0.016015f
C30112 a_5742_30871# a_1736_39043# 4.53e-20
C30113 a_19511_42282# a_21335_42336# 0.011904f
C30114 a_22223_47212# VDD 0.236555f
C30115 a_14097_32519# C1_N_btm 5.88e-20
C30116 a_13487_47204# a_13259_45724# 1.12e-20
C30117 a_584_46384# a_997_45618# 2.73e-20
C30118 a_2124_47436# a_1848_45724# 6.36e-22
C30119 a_2063_45854# a_n755_45592# 0.074611f
C30120 a_4791_45118# a_n2661_45546# 0.012117f
C30121 a_n971_45724# a_n1013_45572# 0.004752f
C30122 a_13507_46334# a_8049_45260# 0.086137f
C30123 a_14311_47204# a_14383_46116# 9.92e-21
C30124 a_11309_47204# a_10809_44734# 5.65e-20
C30125 a_n1613_43370# a_n1533_46116# 0.012221f
C30126 a_12549_44172# a_6945_45028# 0.028827f
C30127 a_2107_46812# a_5497_46414# 0.003373f
C30128 a_n743_46660# a_9625_46129# 0.206271f
C30129 a_n2661_46634# a_10903_43370# 0.663878f
C30130 a_13747_46662# a_15682_46116# 0.001312f
C30131 a_5807_45002# a_17715_44484# 0.045558f
C30132 a_n881_46662# a_n722_46482# 6.07e-19
C30133 a_12816_46660# a_14035_46660# 5.75e-20
C30134 a_13607_46688# a_13885_46660# 0.11044f
C30135 a_12991_46634# a_14180_46812# 2e-20
C30136 a_19466_46812# a_19692_46634# 0.001654f
C30137 a_2443_46660# a_2804_46116# 0.006742f
C30138 a_3524_46660# a_1823_45246# 2.12e-19
C30139 a_2609_46660# a_2698_46116# 4.2e-21
C30140 a_4743_44484# a_4520_42826# 6.49e-21
C30141 a_1414_42308# a_1427_43646# 0.006859f
C30142 a_2998_44172# a_4093_43548# 2.37e-19
C30143 a_4223_44672# a_5755_42852# 5.06e-21
C30144 a_11827_44484# a_18083_42858# 3.77e-21
C30145 a_18494_42460# a_19339_43156# 4.88e-20
C30146 a_18184_42460# a_19164_43230# 0.001269f
C30147 a_10807_43548# a_11173_43940# 0.013678f
C30148 a_n2293_42834# a_4649_42852# 4.54e-19
C30149 a_10949_43914# a_11257_43940# 0.001366f
C30150 a_n1059_45260# a_2713_42308# 0.002489f
C30151 a_n2017_45002# a_2903_42308# 0.013263f
C30152 a_3357_43084# a_5755_42308# 2.11e-20
C30153 a_3065_45002# a_n784_42308# 1.67e-20
C30154 a_n913_45002# a_2725_42558# 0.005368f
C30155 a_7542_44172# VDD 0.412456f
C30156 a_13527_45546# a_8696_44636# 2.77e-21
C30157 a_11823_42460# a_16020_45572# 5.14e-20
C30158 a_11962_45724# a_12561_45572# 1.59e-19
C30159 a_7466_43396# a_3090_45724# 9.39e-20
C30160 a_11967_42832# a_n357_42282# 0.153035f
C30161 a_10807_43548# a_10809_44734# 1.71e-19
C30162 a_15493_43396# a_18189_46348# 4.56e-21
C30163 a_n2293_42282# a_n2312_39304# 4.65e-20
C30164 a_n961_42308# a_n2497_47436# 1.14e-20
C30165 a_n784_42308# w_1575_34946# 0.001423f
C30166 a_n3674_38216# SMPL_ON_P 0.044338f
C30167 a_20731_47026# VDD 0.132317f
C30168 a_15959_42545# CAL_N 3.77e-19
C30169 a_n1641_46494# a_n1736_46482# 0.049827f
C30170 a_n1423_46090# a_n1545_46494# 3.16e-19
C30171 a_n2293_46098# a_n1533_46116# 0.002776f
C30172 a_19692_46634# a_20205_31679# 0.001591f
C30173 a_13059_46348# a_12839_46116# 0.098052f
C30174 a_14513_46634# a_13259_45724# 2.83e-21
C30175 a_9625_46129# a_11189_46129# 0.003371f
C30176 a_9823_46155# a_10355_46116# 0.001471f
C30177 a_8199_44636# a_10903_43370# 8.9e-20
C30178 a_3626_43646# a_14955_43396# 4.11e-21
C30179 a_n97_42460# a_18429_43548# 0.003367f
C30180 a_2982_43646# a_10341_43396# 0.029008f
C30181 a_20193_45348# a_20712_42282# 0.010791f
C30182 a_n2293_43922# a_961_42354# 5.68e-20
C30183 a_n356_44636# a_8515_42308# 1.17e-19
C30184 a_2813_43396# a_3457_43396# 0.026697f
C30185 a_7112_43396# a_8685_43396# 2.65e-19
C30186 SMPL_ON_N a_22545_38993# 1.95e-21
C30187 a_7903_47542# DATA[4] 2.01e-19
C30188 a_6575_47204# DATA[3] 0.055018f
C30189 a_n1435_47204# RST_Z 0.179508f
C30190 a_16977_43638# VDD 0.206333f
C30191 a_16680_45572# a_17023_45118# 0.002499f
C30192 a_8696_44636# a_16922_45042# 0.10244f
C30193 a_9049_44484# a_5883_43914# 0.025986f
C30194 a_7499_43078# a_9838_44484# 2.03e-20
C30195 a_2437_43646# a_2232_45348# 0.001172f
C30196 a_3537_45260# a_5111_44636# 1.36722f
C30197 a_4574_45260# a_5147_45002# 0.001891f
C30198 a_21195_42852# a_20202_43084# 0.018373f
C30199 a_8952_43230# a_4185_45028# 3.54e-21
C30200 a_4905_42826# a_n443_42852# 0.037419f
C30201 a_648_43396# a_n357_42282# 0.003365f
C30202 a_n3565_39590# a_n2312_39304# 0.491833f
C30203 a_22959_44484# RST_Z 0.001339f
C30204 a_13249_42308# a_13661_43548# 0.486588f
C30205 a_14495_45572# a_5807_45002# 0.012666f
C30206 a_13904_45546# a_13747_46662# 0.031534f
C30207 a_2711_45572# a_3699_46634# 0.001403f
C30208 a_10907_45822# a_768_44030# 7.18e-20
C30209 a_8746_45002# a_n2661_46634# 3.38e-20
C30210 a_7230_45938# a_n743_46660# 8.13e-19
C30211 a_18175_45572# a_18597_46090# 0.002203f
C30212 a_18479_45785# a_18780_47178# 1.02e-21
C30213 a_18341_45572# a_18479_47436# 3.11e-21
C30214 a_16789_45572# a_16327_47482# 4.55e-19
C30215 a_3357_43084# a_6151_47436# 0.025786f
C30216 a_2437_43646# a_6851_47204# 0.003764f
C30217 a_413_45260# a_n237_47217# 0.030002f
C30218 a_327_44734# a_n746_45260# 0.256943f
C30219 a_1667_45002# a_n971_45724# 1.51e-19
C30220 a_20205_31679# a_20692_30879# 0.055565f
C30221 a_13259_45724# a_n357_42282# 0.056511f
C30222 a_458_43396# a_n784_42308# 1.67e-20
C30223 a_5649_42852# a_12545_42858# 3.24e-20
C30224 a_4361_42308# a_13635_43156# 2.7e-19
C30225 a_743_42282# a_5342_30871# 0.035916f
C30226 a_16823_43084# a_17333_42852# 5.93e-19
C30227 a_n97_42460# a_961_42354# 5.71e-22
C30228 a_14021_43940# a_14456_42282# 3.19e-21
C30229 a_n4318_39768# a_n4064_39616# 0.047349f
C30230 a_n1557_42282# a_n2472_42282# 3.44e-20
C30231 a_n3674_39768# a_n2946_39866# 4.03e-21
C30232 a_17678_43396# a_17701_42308# 1.14e-19
C30233 a_15743_43084# a_22959_42860# 0.001327f
C30234 a_13885_46660# RST_Z 2.35e-19
C30235 a_7754_38968# a_7754_38636# 0.296258f
C30236 a_3754_39134# a_3754_38470# 2.48e-19
C30237 a_n1630_35242# VDD 3.16282f
C30238 a_n2497_47436# a_n2109_47186# 0.197671f
C30239 a_n2661_43370# a_10157_44484# 7.91e-20
C30240 a_1307_43914# a_5891_43370# 0.084799f
C30241 a_1423_45028# a_5205_44734# 0.001252f
C30242 a_20567_45036# a_18114_32519# 1.7e-20
C30243 a_11691_44458# a_16981_45144# 1.91e-19
C30244 a_8191_45002# a_n2661_43922# 8.71e-21
C30245 a_8953_45002# a_n2661_42834# 2.09e-19
C30246 a_6171_45002# a_15433_44458# 2.27e-20
C30247 a_2437_43646# a_3422_30871# 4.22e-21
C30248 a_9114_42852# a_n357_42282# 1.14e-19
C30249 a_18707_42852# a_13259_45724# 1.69e-20
C30250 a_2713_42308# a_n1925_42282# 7.52e-20
C30251 a_2903_42308# a_526_44458# 5.08e-21
C30252 a_5932_42308# a_n2956_39304# 3.95e-21
C30253 a_7573_43172# a_n443_42852# 4.79e-19
C30254 a_13070_42354# a_10903_43370# 0.04369f
C30255 a_22469_40625# a_13507_46334# 7e-21
C30256 a_15765_45572# a_11415_45002# 0.003223f
C30257 a_15143_45578# a_3483_46348# 1.45e-21
C30258 a_13249_42308# a_4185_45028# 3.74e-20
C30259 a_11827_44484# a_12549_44172# 1.40268f
C30260 a_18175_45572# a_19123_46287# 7.15e-20
C30261 a_18479_45785# a_18285_46348# 2.17e-20
C30262 a_17719_45144# a_5807_45002# 4.18e-21
C30263 a_17613_45144# a_13661_43548# 1.21e-20
C30264 a_n2661_43370# a_n1925_46634# 1.37e-20
C30265 a_3357_43084# a_19466_46812# 0.006916f
C30266 a_6171_45002# a_10623_46897# 1.49e-20
C30267 a_19479_31679# a_19692_46634# 5.21e-19
C30268 a_7227_45028# a_2324_44458# 0.035814f
C30269 a_10053_45546# a_9625_46129# 0.086776f
C30270 a_8746_45002# a_8199_44636# 0.680077f
C30271 a_10193_42453# a_5937_45572# 4.34e-20
C30272 a_8238_44734# a_4791_45118# 0.001045f
C30273 a_n310_44484# a_n1151_42308# 0.00221f
C30274 a_14539_43914# a_16327_47482# 0.031714f
C30275 a_18287_44626# a_11599_46634# 3.51e-19
C30276 a_743_42282# a_20107_42308# 0.00961f
C30277 a_5649_42852# a_19332_42282# 1.31e-19
C30278 a_4190_30871# a_7174_31319# 0.153555f
C30279 a_5534_30871# a_5932_42308# 0.025879f
C30280 a_4361_42308# a_18310_42308# 9.35e-19
C30281 a_20205_31679# VIN_N 0.028894f
C30282 a_17538_32519# C10_N_btm 2.16e-19
C30283 a_n1435_47204# a_2609_46660# 5.42e-20
C30284 a_4915_47217# a_4955_46873# 0.00958f
C30285 a_5129_47502# a_4651_46660# 0.002499f
C30286 a_5815_47464# a_4646_46812# 2.49e-19
C30287 a_6151_47436# a_3877_44458# 0.034088f
C30288 a_n1151_42308# a_5275_47026# 0.002003f
C30289 a_n1741_47186# a_6755_46942# 0.017537f
C30290 a_n237_47217# a_9863_46634# 0.008748f
C30291 a_4791_45118# a_5385_46902# 0.007028f
C30292 a_n443_46116# a_4817_46660# 0.020386f
C30293 a_2905_45572# a_3878_46660# 2.98e-19
C30294 a_22731_47423# a_21588_30879# 0.014331f
C30295 SMPL_ON_N a_20916_46384# 4.07e-20
C30296 a_4883_46098# a_n2661_46634# 0.030655f
C30297 a_n881_46662# a_11309_47204# 0.028783f
C30298 a_8696_44636# a_15743_43084# 3.96e-21
C30299 a_5518_44484# a_5663_43940# 3.51e-19
C30300 a_11691_44458# a_10729_43914# 0.001834f
C30301 a_15433_44458# a_14673_44172# 0.027789f
C30302 a_9313_44734# a_20679_44626# 1.18e-20
C30303 a_5343_44458# a_6453_43914# 1.64e-20
C30304 a_11827_44484# a_12429_44172# 6.51e-20
C30305 a_16922_45042# a_20365_43914# 0.021687f
C30306 a_4223_44672# a_7845_44172# 0.004668f
C30307 a_18184_42460# a_18079_43940# 2.26e-21
C30308 a_5883_43914# a_3905_42865# 5.97e-20
C30309 a_3065_45002# a_3080_42308# 0.171466f
C30310 a_3537_45260# a_4235_43370# 0.010714f
C30311 a_n2017_45002# a_6293_42852# 2.51e-19
C30312 a_n1059_45260# a_6031_43396# 5.04e-20
C30313 a_3357_43084# a_2813_43396# 3.3e-19
C30314 a_n967_45348# a_n1243_43396# 1.73e-19
C30315 a_n3565_38216# a_n2810_45572# 0.104999f
C30316 a_5205_44484# VDD 0.508148f
C30317 COMP_P a_22717_36887# 0.001989f
C30318 a_18114_32519# a_21076_30879# 0.054909f
C30319 a_n2661_42282# a_768_44030# 0.002669f
C30320 a_5244_44056# a_n2293_46634# 1.54e-20
C30321 a_8953_45002# a_5066_45546# 0.013782f
C30322 a_3357_43084# a_20205_31679# 3.97e-19
C30323 a_19479_31679# a_20692_30879# 0.051569f
C30324 a_11361_45348# a_9290_44172# 4.93e-19
C30325 a_11341_43940# a_11453_44696# 0.006646f
C30326 a_15037_44260# a_10227_46804# 2.81e-19
C30327 a_3080_42308# w_1575_34946# 0.001676f
C30328 a_n1190_43762# a_n971_45724# 3.04e-20
C30329 a_n971_45724# VDD 4.911799f
C30330 a_11323_42473# a_11633_42308# 7.95e-20
C30331 a_13657_42558# a_14113_42308# 0.001685f
C30332 a_5742_30871# a_10149_42308# 3.62e-19
C30333 a_14456_42282# a_15764_42576# 4.16e-21
C30334 a_6755_46942# a_7832_46660# 0.025487f
C30335 a_9863_46634# a_8270_45546# 7.01e-19
C30336 a_19321_45002# a_19636_46660# 6.42e-19
C30337 a_n881_46662# a_472_46348# 0.022658f
C30338 a_n1613_43370# a_805_46414# 2.86e-19
C30339 a_4883_46098# a_8199_44636# 0.242f
C30340 a_11599_46634# a_15682_46116# 1.8289f
C30341 a_15507_47210# a_2324_44458# 4e-21
C30342 a_10227_46804# a_12005_46116# 8.43e-19
C30343 a_13717_47436# a_18819_46122# 8.56e-21
C30344 a_12861_44030# a_17957_46116# 0.01013f
C30345 a_6575_47204# a_6945_45028# 0.06375f
C30346 a_3160_47472# a_526_44458# 0.026069f
C30347 a_584_46384# a_1337_46116# 0.044678f
C30348 a_n237_47217# a_5527_46155# 0.001111f
C30349 a_2905_45572# a_n1925_42282# 1.51e-21
C30350 a_n1741_47186# a_8049_45260# 0.003545f
C30351 a_2063_45854# a_835_46155# 1.26e-20
C30352 a_20679_44626# a_20974_43370# 1.79e-20
C30353 a_14539_43914# a_10341_43396# 0.041922f
C30354 a_18579_44172# a_18533_43940# 0.011624f
C30355 a_5891_43370# a_9396_43370# 0.004592f
C30356 a_11827_44484# a_21855_43396# 1e-20
C30357 a_n2293_42834# a_5755_42852# 0.007961f
C30358 a_11823_42460# a_10533_42308# 0.002582f
C30359 a_10193_42453# a_13575_42558# 0.175489f
C30360 a_2711_45572# a_18727_42674# 1.2e-21
C30361 a_1115_44172# a_1241_43940# 0.143754f
C30362 a_19279_43940# a_19741_43940# 6.62e-20
C30363 a_20193_45348# a_20556_43646# 0.009643f
C30364 a_n2661_42834# a_3626_43646# 2.47e-20
C30365 a_n2293_43922# a_2982_43646# 0.094429f
C30366 a_18184_42460# a_14209_32519# 0.006261f
C30367 a_3537_45260# a_5837_43172# 0.001f
C30368 a_17061_44734# VDD 0.17647f
C30369 a_8568_45546# a_7499_43078# 0.070368f
C30370 a_8162_45546# a_9049_44484# 6.68e-20
C30371 a_2711_45572# a_8697_45822# 0.003205f
C30372 a_5841_44260# a_1823_45246# 1.17e-20
C30373 a_19700_43370# a_13661_43548# 0.042923f
C30374 a_8975_43940# a_n443_42852# 0.001317f
C30375 a_18989_43940# a_n357_42282# 6.13e-20
C30376 a_5495_43940# a_5937_45572# 3.03e-19
C30377 a_4361_42308# a_n1613_43370# 1.74e-19
C30378 a_19963_31679# EN_OFFSET_CAL 4.91e-20
C30379 a_n2017_45002# RST_Z 1.48e-20
C30380 a_19479_31679# VIN_N 0.029355f
C30381 a_n4064_39616# C1_P_btm 3.84e-20
C30382 a_5742_30871# a_n3420_37984# 0.004679f
C30383 a_12156_46660# a_10809_44734# 9.31e-19
C30384 a_13059_46348# a_14840_46494# 0.031849f
C30385 a_765_45546# a_10903_43370# 1.58e-19
C30386 a_n2293_46634# a_509_45572# 3.2e-19
C30387 a_n2438_43548# a_1609_45822# 0.002001f
C30388 a_n133_46660# a_n443_42852# 0.001534f
C30389 a_n2661_46098# a_310_45028# 5.46e-20
C30390 a_n743_46660# a_2277_45546# 8.23e-21
C30391 a_6755_46942# a_10586_45546# 1.39e-19
C30392 a_n1991_46122# a_n1076_46494# 0.124988f
C30393 a_n2293_46098# a_805_46414# 0.00328f
C30394 a_20159_44458# a_19987_42826# 4.85e-21
C30395 a_895_43940# a_2075_43172# 1.77e-19
C30396 a_2675_43914# a_1847_42826# 2.13e-20
C30397 a_19862_44208# a_19700_43370# 3.23e-19
C30398 a_20365_43914# a_15743_43084# 1.24e-20
C30399 a_n699_43396# a_n1630_35242# 1.22e-20
C30400 a_2479_44172# a_2905_42968# 0.163227f
C30401 a_15493_43940# a_16759_43396# 8.32e-19
C30402 a_11341_43940# a_17324_43396# 1.91e-20
C30403 a_11967_42832# a_21356_42826# 4.18e-21
C30404 a_n97_42460# a_2982_43646# 0.180648f
C30405 a_375_42282# a_7174_31319# 1.7e-20
C30406 a_15493_43396# a_16867_43762# 0.02646f
C30407 a_9313_44734# a_12800_43218# 0.001591f
C30408 a_n2956_37592# a_n3690_38528# 1.91e-20
C30409 a_n2810_45028# a_n3420_38528# 3.16e-21
C30410 w_1575_34946# a_n1532_35090# 0.796778f
C30411 a_1427_43646# VDD 0.19291f
C30412 a_8696_44636# a_10775_45002# 0.00249f
C30413 a_7499_43078# a_n2661_43370# 0.027764f
C30414 a_22223_45572# a_22591_45572# 7.52e-19
C30415 a_19479_31679# a_3357_43084# 0.058337f
C30416 a_2437_43646# a_19963_31679# 5.48e-19
C30417 a_19700_43370# a_4185_45028# 1.48e-22
C30418 a_13887_32519# a_21076_30879# 0.055154f
C30419 a_n3674_38216# a_n2438_43548# 5.26e-20
C30420 a_n3674_37592# a_n2956_39768# 0.031375f
C30421 a_6293_42852# a_526_44458# 0.029694f
C30422 a_6761_42308# a_n1613_43370# 4.15e-20
C30423 a_15890_42674# a_10227_46804# 0.159412f
C30424 a_10193_42453# a_18479_47436# 8.24e-21
C30425 a_10490_45724# a_10227_46804# 0.031f
C30426 a_13904_45546# a_11599_46634# 6.03e-20
C30427 a_8049_45260# a_10586_45546# 0.038262f
C30428 a_4190_30871# a_21487_43396# 0.001675f
C30429 a_n97_42460# a_5837_42852# 0.011979f
C30430 a_8685_43396# a_12545_42858# 5.31e-20
C30431 a_3422_30871# a_19511_42282# 0.025144f
C30432 a_20301_43646# a_20556_43646# 0.114664f
C30433 a_4093_43548# a_4743_43172# 8.1e-19
C30434 a_3626_43646# a_n2293_42282# 3.32e-19
C30435 a_n2661_42282# a_6123_31319# 0.017717f
C30436 a_19721_31679# C10_N_btm 2.25e-20
C30437 a_3863_42891# VDD 8.63e-19
C30438 a_15765_45572# a_11967_42832# 8.39e-21
C30439 a_3232_43370# a_5518_44484# 0.01014f
C30440 a_6171_45002# a_5343_44458# 2.23e-19
C30441 a_n2661_45010# a_n23_44458# 0.049334f
C30442 a_5147_45002# a_5883_43914# 0.008506f
C30443 a_13258_32519# a_19692_46634# 1.9e-20
C30444 a_7174_31319# a_15227_44166# 5.34e-21
C30445 a_2905_42968# a_n443_42852# 3.32e-21
C30446 a_10518_42984# a_n357_42282# 0.010947f
C30447 a_21356_42826# a_13259_45724# 1.24e-20
C30448 a_15037_45618# a_15009_46634# 1.9e-20
C30449 a_13163_45724# a_13059_46348# 0.00596f
C30450 a_15595_45028# a_12549_44172# 6.29e-22
C30451 a_8746_45002# a_765_45546# 2.27e-20
C30452 a_2437_43646# a_4651_46660# 7.1e-21
C30453 a_327_44734# a_383_46660# 1.22e-20
C30454 a_3429_45260# a_n743_46660# 1.28e-20
C30455 a_4574_45260# a_n1925_46634# 2.53e-20
C30456 a_3232_43370# a_n2661_46634# 3e-21
C30457 a_5111_44636# a_n2293_46634# 0.130609f
C30458 a_14976_45348# a_10227_46804# 7.06e-20
C30459 a_17023_45118# a_11599_46634# 3.91e-20
C30460 a_18587_45118# a_12861_44030# 0.011009f
C30461 a_11530_34132# VDD 0.362839f
C30462 a_n699_43396# a_n971_45724# 0.139047f
C30463 a_2779_44458# a_n237_47217# 8.08e-21
C30464 a_743_42282# a_5755_42308# 0.00936f
C30465 a_15567_42826# a_15785_43172# 0.007234f
C30466 a_4361_42308# a_3905_42558# 0.001685f
C30467 a_5649_42852# a_5379_42460# 0.35554f
C30468 a_4190_30871# a_5932_42308# 0.018227f
C30469 a_n4318_38680# a_n1630_35242# 7.78e-20
C30470 a_n3607_39392# VDD 2.79e-20
C30471 a_4915_47217# a_11117_47542# 0.003021f
C30472 a_6151_47436# a_8128_46384# 0.052868f
C30473 a_7227_47204# a_n881_46662# 0.001451f
C30474 a_n2497_47436# a_n1925_46634# 0.052533f
C30475 SMPL_ON_P a_n2472_46634# 2.91e-19
C30476 a_n2288_47178# a_n2312_38680# 4.65e-20
C30477 a_n2109_47186# a_n2104_46634# 0.009799f
C30478 a_n1741_47186# a_n2442_46660# 0.014004f
C30479 a_n1605_47204# a_n2661_46634# 0.006062f
C30480 a_16327_47482# a_11453_44696# 0.038815f
C30481 a_17591_47464# a_12465_44636# 0.001005f
C30482 a_19386_47436# a_20990_47178# 1.56e-20
C30483 a_18780_47178# a_13507_46334# 3.23e-20
C30484 a_18479_47436# a_21496_47436# 4.29e-19
C30485 a_14797_45144# a_14955_43940# 4.38e-20
C30486 a_10334_44484# a_11541_44484# 4.15e-20
C30487 a_14537_43396# a_15682_43940# 0.01288f
C30488 a_n2293_42834# a_7845_44172# 0.008819f
C30489 a_1423_45028# a_8333_44056# 1.17e-19
C30490 a_1307_43914# a_10807_43548# 0.016974f
C30491 a_13720_44458# a_13857_44734# 0.126609f
C30492 a_11827_44484# a_20637_44484# 9.54e-20
C30493 a_18114_32519# a_20679_44626# 6.99e-19
C30494 a_15803_42450# a_n443_42852# 6.37e-21
C30495 a_13258_32519# a_20692_30879# 0.055049f
C30496 a_19431_45546# VDD 0.342308f
C30497 a_19164_43230# RST_Z 1.35e-21
C30498 a_5342_30871# VIN_P 0.00693f
C30499 a_13017_45260# a_3483_46348# 0.51131f
C30500 a_20193_45348# a_19692_46634# 0.060606f
C30501 a_15765_45572# a_13259_45724# 0.025388f
C30502 a_18175_45572# a_8049_45260# 0.014402f
C30503 a_10193_42453# a_n443_42852# 0.026599f
C30504 a_19963_31679# a_22959_46124# 3.42e-20
C30505 a_22959_45572# a_10809_44734# 3.06e-19
C30506 a_3232_43370# a_8199_44636# 0.32342f
C30507 a_6171_45002# a_8349_46414# 1.52e-21
C30508 a_413_45260# a_13759_46122# 1.21e-20
C30509 a_5691_45260# a_5937_45572# 0.061637f
C30510 a_3537_45260# a_9290_44172# 2.24e-20
C30511 a_20447_31679# a_22223_46124# 9.73e-19
C30512 a_1067_42314# a_5742_30871# 1.17e-20
C30513 a_5267_42460# a_5934_30871# 1.28e-20
C30514 a_n784_42308# a_13575_42558# 2.06e-20
C30515 a_14635_42282# a_7174_31319# 4.88e-21
C30516 a_17364_32525# C7_N_btm 0.072179f
C30517 a_2063_45854# a_3483_46348# 0.164542f
C30518 a_2905_45572# a_2698_46116# 2.3e-20
C30519 a_n1151_42308# a_167_45260# 8.02e-20
C30520 a_n443_46116# a_472_46348# 0.025699f
C30521 a_3785_47178# a_1823_45246# 4.37e-19
C30522 a_3160_47472# a_2521_46116# 1.93e-19
C30523 a_n1741_47186# a_8953_45546# 2.11e-19
C30524 a_n237_47217# a_6165_46155# 0.021223f
C30525 a_13507_46334# a_18285_46348# 0.041986f
C30526 a_4883_46098# a_765_45546# 0.055532f
C30527 a_20894_47436# a_20107_46660# 3.26e-20
C30528 a_13717_47436# a_22591_46660# 4.57e-19
C30529 a_12861_44030# a_11415_45002# 0.081894f
C30530 a_10227_46804# a_22000_46634# 5.39e-19
C30531 a_768_44030# a_15368_46634# 6.08e-22
C30532 a_3221_46660# a_3877_44458# 1.36e-19
C30533 a_2609_46660# a_3633_46660# 2.36e-20
C30534 a_n743_46660# a_6755_46942# 0.044888f
C30535 a_2107_46812# a_8667_46634# 1.72e-19
C30536 a_5807_45002# a_11901_46660# 0.003131f
C30537 a_13747_46662# a_11735_46660# 2.58e-21
C30538 a_12549_44172# a_15559_46634# 0.012304f
C30539 a_11967_42832# a_19328_44172# 1.02e-19
C30540 a_17517_44484# a_15493_43940# 7.18e-20
C30541 a_2998_44172# a_3600_43914# 0.012242f
C30542 a_n699_43396# a_1427_43646# 0.00477f
C30543 a_5518_44484# a_4905_42826# 7.14e-20
C30544 a_742_44458# a_2982_43646# 9.65e-20
C30545 a_626_44172# a_743_42282# 6.2e-19
C30546 a_14539_43914# a_n97_42460# 0.05616f
C30547 a_n1549_44318# a_n1287_44306# 0.001705f
C30548 a_n1331_43914# a_n875_44318# 4.2e-19
C30549 a_n1761_44111# a_n1441_43940# 8.49e-19
C30550 a_n2661_42834# a_3052_44056# 1.84e-19
C30551 a_2382_45260# a_3681_42891# 0.067836f
C30552 a_n1059_45260# a_10796_42968# 0.01348f
C30553 a_n913_45002# a_10835_43094# 0.053818f
C30554 a_n2017_45002# a_10991_42826# 1.61e-19
C30555 a_13076_44458# VDD 0.180665f
C30556 a_n3565_39590# C10_P_btm 9.75e-19
C30557 a_n4064_40160# C4_P_btm 1.47e-19
C30558 a_n4209_39590# C8_P_btm 0.002806f
C30559 a_13258_32519# VIN_N 0.143165f
C30560 a_15682_43940# a_3090_45724# 0.001971f
C30561 a_458_43396# a_n2438_43548# 8.26e-20
C30562 a_4235_43370# a_n2293_46634# 0.012147f
C30563 a_7112_43396# a_768_44030# 4.37e-21
C30564 a_14955_43940# a_14976_45028# 2.22e-19
C30565 a_9159_44484# a_2324_44458# 1.37e-20
C30566 a_11541_44484# a_9290_44172# 0.001162f
C30567 a_7274_43762# a_n1613_43370# 2.77e-19
C30568 a_10341_43396# a_11453_44696# 1.84e-21
C30569 a_17324_43396# a_16327_47482# 0.216094f
C30570 a_16547_43609# a_10227_46804# 8.56e-19
C30571 a_685_42968# a_n2497_47436# 9.26e-22
C30572 a_4361_42308# a_4791_45118# 0.111224f
C30573 a_601_46902# VDD 0.204253f
C30574 a_n4209_39304# a_n3565_39304# 6.82668f
C30575 a_n4315_30879# a_n2302_38778# 6.48e-20
C30576 a_n4064_40160# a_n2946_38778# 1.87e-20
C30577 a_n3607_39616# a_n3420_39072# 3.77e-20
C30578 a_3090_45724# a_1823_45246# 0.038665f
C30579 a_14180_46812# a_11415_45002# 8.77e-22
C30580 a_20107_46660# a_20411_46873# 0.316529f
C30581 a_19551_46910# a_20273_46660# 2.93e-19
C30582 a_19123_46287# a_20841_46902# 3.69e-21
C30583 a_n743_46660# a_8049_45260# 2.07544f
C30584 a_2609_46660# a_526_44458# 2.13e-19
C30585 a_2107_46812# a_6640_46482# 8.98e-19
C30586 a_10623_46897# a_10903_43370# 1.59e-19
C30587 a_6755_46942# a_11189_46129# 6.12e-20
C30588 a_10249_46116# a_11133_46155# 0.007085f
C30589 a_7715_46873# a_2324_44458# 2.47e-20
C30590 a_5343_44458# a_8292_43218# 0.01105f
C30591 a_21115_43940# a_2982_43646# 5.25e-20
C30592 a_3422_30871# a_21259_43561# 1.69e-19
C30593 a_21398_44850# a_4190_30871# 8.73e-21
C30594 a_n2661_43922# a_7765_42852# 2.66e-21
C30595 a_n2293_43922# a_7871_42858# 1.21e-20
C30596 a_n2661_42834# a_8037_42858# 7.33e-22
C30597 a_9313_44734# a_10341_42308# 0.019286f
C30598 a_10807_43548# a_9396_43370# 2.23e-20
C30599 a_n1059_45260# a_4958_30871# 0.005345f
C30600 a_n2017_45002# a_17303_42282# 0.006515f
C30601 en_comp a_17124_42282# 4.59e-20
C30602 a_2711_45572# a_14180_45002# 0.147337f
C30603 a_15861_45028# a_17568_45572# 0.004094f
C30604 a_8696_44636# a_17668_45572# 2.03e-19
C30605 a_9049_44484# a_3537_45260# 1.31e-19
C30606 a_n4064_37440# C4_P_btm 1.74e-19
C30607 a_n3420_37440# C2_P_btm 2.75e-19
C30608 VDAC_N EN_VIN_BSTR_N 0.341739f
C30609 a_20301_43646# a_19692_46634# 0.110092f
C30610 a_5495_43940# a_n443_42852# 1.65e-21
C30611 a_3499_42826# a_n863_45724# 9.47e-19
C30612 a_6761_42308# a_4791_45118# 0.001495f
C30613 a_12594_46348# VDD 1.03351f
C30614 a_6472_45840# a_2063_45854# 0.545607f
C30615 a_2211_45572# a_n237_47217# 0.005215f
C30616 a_3175_45822# a_n1151_42308# 2.87e-20
C30617 a_8953_45546# a_10586_45546# 2.02e-20
C30618 a_8016_46348# a_10037_46155# 0.002633f
C30619 a_9823_46155# a_10044_46482# 0.007833f
C30620 a_11189_46129# a_8049_45260# 0.03932f
C30621 a_n2956_38680# a_n1736_46482# 1.43e-19
C30622 a_n2956_39304# a_n1545_46494# 1.4e-20
C30623 a_n2472_46090# a_n2661_45546# 0.00558f
C30624 a_n2293_46098# a_n2810_45572# 0.013787f
C30625 a_20202_43084# a_n357_42282# 0.062522f
C30626 a_1115_44172# a_1067_42314# 2.43e-21
C30627 a_15681_43442# a_15781_43660# 0.167615f
C30628 a_7287_43370# a_5649_42852# 1.08e-21
C30629 a_8791_43396# a_4361_42308# 2.28e-21
C30630 a_10341_43396# a_17324_43396# 0.010417f
C30631 a_1049_43396# a_791_42968# 5.89e-19
C30632 a_n97_42460# a_7871_42858# 0.001218f
C30633 a_9313_44734# a_18057_42282# 2.51e-20
C30634 a_9145_43396# a_15125_43396# 0.001605f
C30635 a_1568_43370# a_685_42968# 1.82e-20
C30636 a_1414_42308# a_564_42282# 1.31e-20
C30637 a_15037_43940# a_5342_30871# 6.83e-20
C30638 a_9804_47204# CLK 5.1e-19
C30639 a_11117_47542# DATA[5] 3.92e-19
C30640 a_13759_47204# RST_Z 9.49e-19
C30641 a_4520_42826# VDD 0.142755f
C30642 a_n2956_37592# a_n2216_37984# 1.2e-19
C30643 a_11823_42460# a_n2661_43922# 0.005005f
C30644 a_17478_45572# a_16979_44734# 9.61e-20
C30645 a_7499_43078# a_11909_44484# 7.77e-22
C30646 a_8696_44636# a_17970_44736# 4.11e-19
C30647 a_22959_45572# a_22959_45036# 0.026152f
C30648 a_4558_45348# a_n2661_43370# 0.018142f
C30649 a_7276_45260# a_n2293_42834# 1.85e-19
C30650 a_6171_45002# a_8560_45348# 0.004926f
C30651 a_3357_43084# a_20193_45348# 1.08e-20
C30652 a_21188_45572# a_19721_31679# 3.94e-20
C30653 a_5934_30871# a_3090_45724# 2.22e-20
C30654 a_16137_43396# a_n443_42852# 0.020044f
C30655 a_10991_42826# a_526_44458# 2.56e-21
C30656 a_16867_43762# a_n357_42282# 8.18e-21
C30657 a_10405_44172# CLK 6.38e-19
C30658 a_10053_45546# a_6755_46942# 1.29e-20
C30659 a_10490_45724# a_10467_46802# 2.95e-19
C30660 a_19418_45938# a_13747_46662# 6.02e-19
C30661 a_18787_45572# a_13661_43548# 0.001493f
C30662 a_1609_45572# a_3090_45724# 1.86e-20
C30663 a_2437_43646# a_10037_47542# 9.04e-19
C30664 a_n2293_42834# a_n746_45260# 1.39e-21
C30665 a_2304_45348# a_n443_46116# 0.008048f
C30666 a_8137_45348# a_n971_45724# 7.49e-20
C30667 a_13159_45002# a_12861_44030# 0.008506f
C30668 a_6171_45002# a_10227_46804# 0.087616f
C30669 a_413_45260# a_22731_47423# 0.005286f
C30670 a_15279_43071# a_5342_30871# 0.214197f
C30671 a_15743_43084# a_22400_42852# 0.010325f
C30672 a_2982_43646# a_10533_42308# 1.49e-19
C30673 a_n97_42460# a_11897_42308# 7.16e-19
C30674 a_7112_43396# a_6123_31319# 1.32e-19
C30675 a_17730_32519# C9_N_btm 0.215899f
C30676 a_19237_31679# C7_N_btm 1.43e-20
C30677 a_15720_42674# VDD 4.6e-19
C30678 a_5815_47464# a_6545_47178# 0.001457f
C30679 a_4915_47217# a_6851_47204# 0.172567f
C30680 a_5129_47502# a_6491_46660# 1.6e-20
C30681 a_2905_45572# a_n1435_47204# 5.63e-19
C30682 a_n1151_42308# a_11459_47204# 3.65e-19
C30683 a_n2661_44458# a_n2012_44484# 0.003432f
C30684 a_18494_42460# a_9313_44734# 0.028817f
C30685 a_n4318_40392# a_n1809_44850# 5.8e-21
C30686 a_3537_45260# a_3905_42865# 0.258917f
C30687 a_n967_45348# a_n875_44318# 4.26e-20
C30688 a_4558_45348# a_2998_44172# 2.03e-19
C30689 a_n784_42308# a_n443_42852# 0.005038f
C30690 a_2351_42308# a_n755_45592# 0.057532f
C30691 a_n327_42308# a_n357_42282# 0.00216f
C30692 a_3318_42354# a_n863_45724# 9.94e-19
C30693 a_11322_45546# VDD 0.370908f
C30694 a_14209_32519# RST_Z 0.049869f
C30695 a_9482_43914# a_13885_46660# 3.2e-20
C30696 a_18287_44626# a_13661_43548# 0.021421f
C30697 a_8975_43940# a_n2661_46634# 1.39e-19
C30698 a_18248_44752# a_13747_46662# 2.31e-20
C30699 a_10334_44484# a_n2293_46634# 2.78e-20
C30700 a_n913_45002# a_11415_45002# 4.59e-20
C30701 a_17767_44458# a_19321_45002# 1.52e-37
C30702 a_4185_45348# a_3090_45724# 1.98e-19
C30703 a_10053_45546# a_8049_45260# 0.002369f
C30704 a_8696_44636# a_14840_46494# 1.02e-21
C30705 a_16855_45546# a_15682_46116# 0.011741f
C30706 a_13385_45572# a_10903_43370# 0.006432f
C30707 a_15765_45572# a_18189_46348# 7.83e-21
C30708 a_16333_45814# a_17715_44484# 2.81e-19
C30709 a_5891_43370# a_n1613_43370# 0.064769f
C30710 a_n2661_42834# a_n2312_40392# 8.33e-20
C30711 a_n2293_43922# a_11453_44696# 1.93e-20
C30712 a_15433_44458# a_4883_46098# 2.94e-21
C30713 a_14673_44172# a_10227_46804# 0.012944f
C30714 a_11967_42832# a_12861_44030# 0.209245f
C30715 a_n2065_43946# a_584_46384# 2.03e-21
C30716 a_1115_44172# a_n746_45260# 2.04e-19
C30717 a_18083_42858# a_18214_42558# 0.001378f
C30718 a_18249_42858# a_18907_42674# 0.001692f
C30719 a_18817_42826# a_18727_42674# 0.001214f
C30720 a_19164_43230# a_17303_42282# 9.77e-21
C30721 a_n2840_42282# a_n1630_35242# 0.040623f
C30722 COMP_P a_n1329_42308# 0.232443f
C30723 a_n2472_42282# a_n3674_37592# 0.007439f
C30724 a_5342_30871# a_13258_32519# 0.030303f
C30725 a_n2104_42282# a_n784_42308# 8.09e-20
C30726 a_n2293_46634# a_n1021_46688# 2.69e-22
C30727 a_n2661_46634# a_n133_46660# 0.022138f
C30728 a_n2104_46634# a_n1925_46634# 0.167849f
C30729 a_n2472_46634# a_n2438_43548# 0.008762f
C30730 a_768_44030# a_2864_46660# 1.39e-19
C30731 a_n881_46662# a_4955_46873# 0.066882f
C30732 a_n1613_43370# a_4817_46660# 0.330391f
C30733 a_4883_46098# a_10623_46897# 1.58e-19
C30734 a_11599_46634# a_11735_46660# 0.268769f
C30735 a_n1435_47204# a_12816_46660# 7.47e-21
C30736 a_n1151_42308# a_12925_46660# 5.47e-20
C30737 a_949_44458# a_1443_43940# 2.54e-19
C30738 a_8696_44636# a_8605_42826# 4.39e-21
C30739 a_10057_43914# a_10555_44260# 0.041594f
C30740 a_18374_44850# a_15493_43396# 3.95e-21
C30741 a_20835_44721# a_20512_43084# 1.67e-21
C30742 a_20679_44626# a_22485_44484# 8.1e-21
C30743 a_n2293_43922# a_n3674_39768# 0.018871f
C30744 a_18989_43940# a_19328_44172# 4.08e-19
C30745 a_n356_44636# a_15682_43940# 3.38e-21
C30746 a_20766_44850# a_21145_44484# 3.16e-19
C30747 a_19279_43940# a_21073_44484# 0.002178f
C30748 a_20640_44752# a_22591_44484# 8.79e-21
C30749 a_5891_43370# a_7584_44260# 2.54e-20
C30750 a_7640_43914# a_8018_44260# 9.16e-20
C30751 a_13348_45260# a_9145_43396# 9.73e-20
C30752 a_n2661_43922# a_n1644_44306# 0.002488f
C30753 a_n2661_42834# a_n1453_44318# 0.001232f
C30754 a_5742_30871# EN_VIN_BSTR_N 0.643089f
C30755 a_n356_44636# a_1823_45246# 4.79e-19
C30756 a_18374_44850# a_3483_46348# 1.41e-21
C30757 a_8975_43940# a_8199_44636# 0.028334f
C30758 a_10695_43548# a_2063_45854# 3.18e-19
C30759 a_19511_42282# a_7174_31319# 0.240861f
C30760 a_13258_32519# a_20107_42308# 0.021019f
C30761 a_5742_30871# a_1239_39043# 5.42e-20
C30762 a_17303_42282# a_21973_42336# 5.22e-19
C30763 a_12465_44636# VDD 0.773277f
C30764 a_12861_44030# a_13259_45724# 0.435853f
C30765 a_n1151_42308# a_n863_45724# 0.081395f
C30766 a_584_46384# a_n755_45592# 0.020619f
C30767 a_1431_47204# a_1848_45724# 2.87e-19
C30768 a_2063_45854# a_n357_42282# 1.15e-20
C30769 a_n971_45724# a_7_45899# 3.69e-19
C30770 a_n1613_43370# a_n722_46482# 0.002104f
C30771 a_n2661_46634# a_11387_46155# 0.0013f
C30772 a_n2293_46634# a_9290_44172# 0.102393f
C30773 a_2107_46812# a_5204_45822# 0.002125f
C30774 a_12891_46348# a_6945_45028# 0.013255f
C30775 a_n743_46660# a_8953_45546# 0.062066f
C30776 a_13747_46662# a_2324_44458# 0.025909f
C30777 a_13661_43548# a_15682_46116# 1.42e-19
C30778 a_5807_45002# a_17583_46090# 0.008151f
C30779 a_n881_46662# a_n967_46494# 8.68e-20
C30780 a_19333_46634# a_19692_46634# 0.005582f
C30781 a_12816_46660# a_13885_46660# 8.55e-20
C30782 a_n2661_46098# a_2804_46116# 1.71e-20
C30783 a_3699_46634# a_1823_45246# 1.1e-20
C30784 a_2609_46660# a_2521_46116# 1.95e-19
C30785 a_2443_46660# a_2698_46116# 9.84e-20
C30786 a_9313_44734# a_15940_43402# 4.1e-19
C30787 a_n699_43396# a_4520_42826# 8.42e-22
C30788 a_1467_44172# a_1427_43646# 0.104539f
C30789 a_n1441_43940# a_n2267_43396# 4.29e-19
C30790 a_11691_44458# a_15567_42826# 4.44e-21
C30791 a_11827_44484# a_17701_42308# 5.54e-22
C30792 a_4223_44672# a_5111_42852# 3.04e-21
C30793 a_18184_42460# a_19339_43156# 0.004558f
C30794 a_10729_43914# a_11257_43940# 0.007166f
C30795 a_10949_43914# a_11173_43940# 4.93e-19
C30796 a_10807_43548# a_10867_43940# 9.12e-19
C30797 a_2479_44172# a_3080_42308# 0.001674f
C30798 a_1414_42308# a_n1557_42282# 2.99e-21
C30799 a_n2661_44458# a_10835_43094# 8.47e-20
C30800 a_n1059_45260# a_2725_42558# 2.97e-19
C30801 a_n2017_45002# a_2713_42308# 0.011694f
C30802 en_comp a_1755_42282# 9.98e-21
C30803 a_7281_43914# VDD 0.198809f
C30804 a_11280_45822# a_11136_45572# 6.84e-19
C30805 a_15143_45578# a_15765_45572# 1.5e-19
C30806 a_14401_32519# a_21076_30879# 0.057698f
C30807 a_12545_42858# a_768_44030# 2.24e-19
C30808 a_10949_43914# a_10809_44734# 0.002017f
C30809 a_15493_43396# a_17715_44484# 3.2e-19
C30810 a_n2293_42282# a_n2312_40392# 0.001844f
C30811 a_n2104_42282# SMPL_ON_P 5.11e-20
C30812 a_20528_46660# VDD 0.077608f
C30813 a_15803_42450# CAL_N 0.002185f
C30814 a_n1991_46122# a_n1545_46494# 2.28e-19
C30815 a_n2157_46122# a_n967_46494# 2.56e-19
C30816 a_n1641_46494# a_n2956_38680# 2.13e-19
C30817 a_20841_46902# a_8049_45260# 8.01e-21
C30818 a_14513_46634# a_14383_46116# 4.21e-20
C30819 a_14180_46812# a_13259_45724# 1.49e-21
C30820 a_15227_44166# a_20850_46155# 8.44e-19
C30821 a_3483_46348# a_17715_44484# 0.059106f
C30822 a_9625_46129# a_9290_44172# 4.14e-20
C30823 a_n4064_39616# a_n3420_37984# 0.050009f
C30824 a_n3420_39616# a_n4064_37984# 0.046151f
C30825 a_4958_30871# a_n3420_37440# 0.033151f
C30826 a_4419_46090# a_2324_44458# 2.42e-20
C30827 SMPL_ON_N a_22521_39511# 1.24e-19
C30828 a_7227_47204# DATA[4] 1.74e-19
C30829 a_n97_42460# a_17324_43396# 0.003115f
C30830 a_13483_43940# a_12545_42858# 6.25e-20
C30831 a_n2293_43922# a_1184_42692# 3.75e-20
C30832 a_n356_44636# a_5934_30871# 0.095373f
C30833 a_3626_43646# a_15095_43370# 1.07e-19
C30834 a_7287_43370# a_8685_43396# 7.31e-19
C30835 a_7903_47542# DATA[3] 0.01066f
C30836 a_13381_47204# RST_Z 2.25e-20
C30837 a_16409_43396# VDD 0.250832f
C30838 a_10193_42453# CAL_N 0.00219f
C30839 a_4574_45260# a_4558_45348# 0.19344f
C30840 a_3537_45260# a_5147_45002# 0.092965f
C30841 a_2382_45260# a_3232_43370# 0.239776f
C30842 a_3065_45002# a_4927_45028# 1.12e-20
C30843 a_3429_45260# a_5111_44636# 3.89e-22
C30844 a_16680_45572# a_16922_45042# 5.89e-20
C30845 a_16855_45546# a_17023_45118# 4.36e-19
C30846 a_9049_44484# a_8701_44490# 0.100038f
C30847 a_7499_43078# a_5883_43914# 0.100372f
C30848 a_n2017_45002# a_9482_43914# 2.97e-21
C30849 a_2437_43646# a_1423_45028# 0.023818f
C30850 a_9127_43156# a_4185_45028# 9.18e-20
C30851 a_21356_42826# a_20202_43084# 0.011854f
C30852 a_17141_43172# a_15227_44166# 4.12e-20
C30853 a_3080_42308# a_n443_42852# 0.029846f
C30854 a_548_43396# a_n357_42282# 0.001387f
C30855 a_17730_32519# RST_Z 0.049818f
C30856 a_8162_45546# a_n1925_46634# 0.104508f
C30857 a_13249_42308# a_5807_45002# 0.725941f
C30858 a_10193_42453# a_n2661_46634# 0.351509f
C30859 a_13527_45546# a_13747_46662# 5.21e-20
C30860 a_2711_45572# a_2959_46660# 2.89e-21
C30861 a_13904_45546# a_13661_43548# 9.04e-21
C30862 a_10907_45822# a_12549_44172# 9.26e-20
C30863 a_6812_45938# a_n743_46660# 0.002228f
C30864 a_18175_45572# a_18780_47178# 2.7e-19
C30865 a_18479_45785# a_18479_47436# 2.68e-19
C30866 a_18799_45938# a_16327_47482# 0.013823f
C30867 a_19418_45938# a_11599_46634# 1.59e-19
C30868 a_3357_43084# a_5815_47464# 0.029103f
C30869 a_2437_43646# a_6491_46660# 0.002468f
C30870 a_n2293_45010# a_n1151_42308# 0.020357f
C30871 a_413_45260# a_n746_45260# 0.031693f
C30872 a_3537_45260# a_n2109_47186# 5.89e-19
C30873 a_16823_43084# a_18083_42858# 4.78e-20
C30874 a_15743_43084# a_22223_42860# 0.021215f
C30875 a_5649_42852# a_12089_42308# 3.26e-20
C30876 a_4361_42308# a_12895_43230# 5.63e-20
C30877 a_743_42282# a_15279_43071# 4.98e-21
C30878 a_4190_30871# a_15567_42826# 6.55e-21
C30879 a_n97_42460# a_1184_42692# 8.23e-20
C30880 a_n3674_39768# a_n3420_39616# 0.073948f
C30881 a_n4318_39768# a_n2946_39866# 7.88e-20
C30882 a_7754_39300# a_3754_38470# 0.082848f
C30883 a_564_42282# VDD 0.293756f
C30884 a_n2497_47436# a_n2288_47178# 0.067981f
C30885 a_n2833_47464# a_n2109_47186# 0.002667f
C30886 a_5907_45546# a_5829_43940# 5.47e-21
C30887 a_n2661_43370# a_9838_44484# 1.69e-20
C30888 a_1307_43914# a_8375_44464# 3.91e-20
C30889 a_20567_45036# a_20205_45028# 2.35e-20
C30890 a_1423_45028# a_4181_44734# 0.002332f
C30891 a_413_45260# a_17517_44484# 0.013023f
C30892 a_6171_45002# a_14815_43914# 2.54e-21
C30893 a_n913_45002# a_11967_42832# 0.156551f
C30894 a_21513_45002# a_3422_30871# 9.94e-20
C30895 a_17124_42282# a_4185_45028# 1.64e-19
C30896 a_2713_42308# a_526_44458# 6.21e-21
C30897 a_7309_43172# a_n443_42852# 0.00116f
C30898 a_12563_42308# a_10903_43370# 0.002814f
C30899 a_22521_40599# a_13507_46334# 2.03e-20
C30900 a_15903_45785# a_11415_45002# 0.02962f
C30901 a_14495_45572# a_3483_46348# 9.37e-21
C30902 a_18175_45572# a_18285_46348# 0.010439f
C30903 a_11827_44484# a_12891_46348# 0.020579f
C30904 a_17023_45118# a_13661_43548# 1.73e-20
C30905 a_16922_45042# a_13747_46662# 0.00477f
C30906 a_17613_45144# a_5807_45002# 8.23e-21
C30907 a_21359_45002# a_12549_44172# 9.07e-19
C30908 a_n2661_43370# a_n2312_38680# 1.32e-20
C30909 a_6171_45002# a_10467_46802# 4.36e-22
C30910 a_3357_43084# a_19333_46634# 2.08e-20
C30911 a_22223_45572# a_19692_46634# 1.03e-19
C30912 a_10193_42453# a_8199_44636# 0.236934f
C30913 a_6598_45938# a_2324_44458# 2.88e-20
C30914 a_9049_44484# a_9625_46129# 0.00226f
C30915 a_10180_45724# a_5937_45572# 8.62e-20
C30916 a_10490_45724# a_8016_46348# 2.74e-21
C30917 a_5891_43370# a_4791_45118# 0.066388f
C30918 a_18989_43940# a_12861_44030# 0.047422f
C30919 a_12607_44458# a_10227_46804# 3.68e-19
C30920 a_16112_44458# a_16327_47482# 3.69e-19
C30921 a_18248_44752# a_11599_46634# 2.26e-19
C30922 a_5343_44458# a_4883_46098# 6.41e-22
C30923 a_9127_43156# a_9803_42558# 0.001572f
C30924 a_8952_43230# a_9223_42460# 2.08e-19
C30925 a_5649_42852# a_18907_42674# 5.66e-20
C30926 a_4190_30871# a_20712_42282# 1.12e-20
C30927 a_20301_43646# a_20107_42308# 5.1e-21
C30928 a_743_42282# a_13258_32519# 0.030886f
C30929 a_4361_42308# a_18220_42308# 6.69e-19
C30930 a_17538_32519# C9_N_btm 7.08e-19
C30931 a_n1435_47204# a_2443_46660# 5.41e-20
C30932 a_4915_47217# a_4651_46660# 1.15e-19
C30933 a_5129_47502# a_4646_46812# 1.7e-20
C30934 a_5815_47464# a_3877_44458# 2.22e-20
C30935 a_n237_47217# a_8492_46660# 0.002629f
C30936 a_n1741_47186# a_10249_46116# 5.18e-19
C30937 a_n443_46116# a_4955_46873# 0.126551f
C30938 a_4791_45118# a_4817_46660# 0.020367f
C30939 a_n1151_42308# a_5072_46660# 0.009494f
C30940 a_2905_45572# a_3633_46660# 3.11e-19
C30941 a_2063_45854# a_5263_46660# 1.33e-19
C30942 a_22223_47212# a_21588_30879# 0.164932f
C30943 a_12465_44636# a_22612_30879# 7.45e-19
C30944 a_22731_47423# a_20916_46384# 1.06e-19
C30945 a_18587_45118# a_18451_43940# 1.13e-20
C30946 a_n2267_44484# a_n1441_43940# 1.52e-19
C30947 a_5518_44484# a_5495_43940# 3.48e-20
C30948 a_14815_43914# a_14673_44172# 0.173231f
C30949 a_16922_45042# a_20269_44172# 0.010825f
C30950 a_4223_44672# a_7542_44172# 0.052366f
C30951 a_11827_44484# a_11750_44172# 8.34e-20
C30952 a_3537_45260# a_4093_43548# 0.001642f
C30953 a_3065_45002# a_4699_43561# 1.24e-20
C30954 a_n2017_45002# a_6031_43396# 5.49e-20
C30955 a_2382_45260# a_4905_42826# 7.37e-21
C30956 a_n4334_38304# a_n2810_45572# 3.54e-20
C30957 a_6431_45366# VDD 0.203167f
C30958 a_n784_42308# CAL_P 0.006719f
C30959 a_n2661_44458# a_11415_45002# 2.26e-19
C30960 a_3905_42865# a_n2293_46634# 0.039006f
C30961 a_6101_44260# a_768_44030# 4.28e-19
C30962 a_9482_43914# a_526_44458# 0.001072f
C30963 a_6171_45002# a_8034_45724# 0.002969f
C30964 a_5111_44636# a_8049_45260# 0.00103f
C30965 a_8191_45002# a_5066_45546# 7.35e-19
C30966 a_n913_45002# a_13259_45724# 0.142601f
C30967 a_19479_31679# a_20205_31679# 0.06173f
C30968 a_9801_44260# a_4883_46098# 1.5e-19
C30969 a_14761_44260# a_10227_46804# 6.06e-20
C30970 a_14021_43940# a_18479_47436# 1.76e-19
C30971 a_n2129_43609# a_584_46384# 6.92e-20
C30972 a_n1809_43762# a_n971_45724# 8.16e-19
C30973 a_n452_47436# VDD 0.092189f
C30974 a_14456_42282# a_15486_42560# 6.85e-20
C30975 a_4921_42308# a_7174_31319# 1.72e-20
C30976 a_n1630_35242# a_n2302_39866# 5.02e-20
C30977 a_n784_42308# a_1736_39587# 3.17e-20
C30978 a_n4318_38216# a_n4064_39072# 0.023072f
C30979 a_5742_30871# a_9885_42308# 1.65e-19
C30980 a_n3674_38216# a_n3420_39072# 0.020386f
C30981 a_16137_43396# CAL_N 7.09e-19
C30982 a_8492_46660# a_8270_45546# 0.007406f
C30983 a_n133_46660# a_765_45546# 7.71e-20
C30984 a_n881_46662# a_376_46348# 0.016146f
C30985 a_n1613_43370# a_472_46348# 3.32e-19
C30986 a_4883_46098# a_8349_46414# 0.007204f
C30987 a_10227_46804# a_10903_43370# 0.041882f
C30988 a_11599_46634# a_2324_44458# 0.428445f
C30989 a_12861_44030# a_18189_46348# 0.004513f
C30990 a_7903_47542# a_6945_45028# 0.005336f
C30991 a_2905_45572# a_526_44458# 0.142766f
C30992 a_584_46384# a_835_46155# 0.001103f
C30993 a_n237_47217# a_5210_46155# 0.002744f
C30994 a_3160_47472# a_2981_46116# 4.76e-19
C30995 a_20640_44752# a_20974_43370# 2.23e-21
C30996 a_5891_43370# a_8791_43396# 0.194389f
C30997 a_18579_44172# a_19319_43548# 0.031277f
C30998 a_11827_44484# a_4361_42308# 1.05e-20
C30999 a_18184_42460# a_22591_43396# 8.5e-19
C31000 a_20193_45348# a_743_42282# 0.007306f
C31001 a_n2293_42834# a_5111_42852# 0.009675f
C31002 a_10193_42453# a_13070_42354# 1.07e-19
C31003 a_9028_43914# a_9672_43914# 2.65e-19
C31004 a_11823_42460# a_10545_42558# 1.52e-20
C31005 a_3537_45260# a_5457_43172# 0.001869f
C31006 a_n913_45002# a_9114_42852# 4.02e-19
C31007 a_16241_44734# VDD 0.189894f
C31008 a_n3565_38216# VCM 0.03544f
C31009 a_5907_45546# a_6229_45572# 0.007399f
C31010 a_8162_45546# a_7499_43078# 0.021916f
C31011 a_2711_45572# a_8336_45822# 2.46e-19
C31012 a_17973_43940# a_12741_44636# 1.04e-20
C31013 a_3820_44260# a_1823_45246# 7.74e-19
C31014 a_15743_43084# a_13747_46662# 6.22e-21
C31015 a_19268_43646# a_13661_43548# 0.136251f
C31016 a_6655_43762# a_4646_46812# 8.82e-19
C31017 a_16823_43084# a_12549_44172# 8.9e-20
C31018 a_n356_44636# a_n2293_45546# 1.65e-19
C31019 a_10057_43914# a_n443_42852# 0.06562f
C31020 a_5013_44260# a_5937_45572# 4.74e-20
C31021 a_n1423_42826# a_n2312_40392# 4.82e-21
C31022 a_3357_43084# CLK 2.63944f
C31023 a_8654_47026# VDD 4.6e-19
C31024 a_n3420_39616# C0_P_btm 1.63e-20
C31025 a_n784_42308# CAL_N 0.00432f
C31026 a_n1630_35242# VDAC_N 0.003372f
C31027 a_13059_46348# a_15015_46420# 0.002269f
C31028 a_15227_46910# a_14840_46494# 2e-19
C31029 a_n2293_46634# a_n89_45572# 4.13e-19
C31030 a_10249_46116# a_10586_45546# 1.88e-19
C31031 a_n743_46660# a_1609_45822# 5.99e-19
C31032 a_n2438_43548# a_n443_42852# 3.03e-19
C31033 a_n2661_46098# a_n1099_45572# 7.03e-20
C31034 a_2107_46812# a_3503_45724# 7.75e-22
C31035 a_n1423_46090# a_n1641_46494# 0.209641f
C31036 a_n2157_46122# a_376_46348# 2.25e-21
C31037 a_n1991_46122# a_n901_46420# 0.041816f
C31038 a_n1853_46287# a_n1076_46494# 0.056078f
C31039 a_n2293_46098# a_472_46348# 0.009446f
C31040 a_895_43940# a_1847_42826# 2.53e-19
C31041 a_20269_44172# a_15743_43084# 8.8e-21
C31042 a_19478_44306# a_19700_43370# 0.008781f
C31043 a_1568_43370# a_1756_43548# 0.094732f
C31044 a_742_44458# a_1184_42692# 1.39e-19
C31045 a_15493_43940# a_16977_43638# 5.19e-19
C31046 a_11341_43940# a_17499_43370# 2.28e-19
C31047 a_19279_43940# a_18083_42858# 9.26e-20
C31048 a_n699_43396# a_564_42282# 1.29e-22
C31049 a_n1699_43638# a_n1243_43396# 4.2e-19
C31050 a_n97_42460# a_2896_43646# 0.027089f
C31051 a_15493_43396# a_16664_43396# 0.016417f
C31052 a_2479_44172# a_2075_43172# 0.034186f
C31053 a_n2129_43609# a_n144_43396# 7.58e-20
C31054 a_n2956_37592# a_n3565_38502# 0.024508f
C31055 w_1575_34946# a_n1386_35608# 0.005843f
C31056 a_n1557_42282# VDD 0.355513f
C31057 a_8568_45546# a_n2661_43370# 6.03e-21
C31058 a_14033_45822# a_14180_45002# 2.17e-20
C31059 a_8746_45002# a_8560_45348# 0.044092f
C31060 a_2711_45572# a_18494_42460# 0.1183f
C31061 a_8696_44636# a_8953_45002# 0.018854f
C31062 a_2437_43646# a_22591_45572# 2.94e-19
C31063 a_22223_45572# a_3357_43084# 0.07533f
C31064 a_21513_45002# a_19963_31679# 3.07e-19
C31065 a_14209_32519# a_20820_30879# 0.053104f
C31066 a_n2104_42282# a_n2438_43548# 0.009764f
C31067 a_15567_42826# a_15227_44166# 0.075768f
C31068 a_18249_42858# a_3090_45724# 1.21e-20
C31069 COMP_P a_n2312_38680# 4.95e-19
C31070 a_6031_43396# a_526_44458# 0.002054f
C31071 a_14021_43940# a_n443_42852# 0.05804f
C31072 a_6773_42558# a_n1613_43370# 1.71e-19
C31073 a_15959_42545# a_10227_46804# 0.152289f
C31074 a_n3420_39072# w_1575_34946# 0.023412f
C31075 a_10037_46155# VDD 0.001395f
C31076 a_15143_45578# a_12861_44030# 4.39e-20
C31077 a_13249_42308# a_14311_47204# 1.62e-21
C31078 a_8746_45002# a_10227_46804# 0.117547f
C31079 a_13527_45546# a_11599_46634# 5.7e-19
C31080 a_4880_45572# a_4883_46098# 7.06e-20
C31081 a_8049_45260# a_8379_46155# 1.85e-19
C31082 a_17715_44484# a_n357_42282# 1.41e-20
C31083 a_10695_43548# a_10083_42826# 0.005272f
C31084 a_9145_43396# a_10835_43094# 4.2e-20
C31085 a_20301_43646# a_743_42282# 0.09203f
C31086 a_19177_43646# a_19095_43396# 8.13e-19
C31087 a_21259_43561# a_21487_43396# 0.08444f
C31088 a_4190_30871# a_20556_43646# 0.021112f
C31089 a_4093_43548# a_4649_43172# 0.001356f
C31090 a_n1557_42282# a_873_42968# 8.49e-21
C31091 a_n2661_42282# a_7227_42308# 3.35e-19
C31092 a_8685_43396# a_12089_42308# 3.95e-19
C31093 a_18114_32519# C10_N_btm 0.460005f
C31094 a_19721_31679# C9_N_btm 1.91e-20
C31095 a_16751_45260# a_16981_45144# 0.004937f
C31096 a_5691_45260# a_5518_44484# 8.35e-19
C31097 a_3232_43370# a_5343_44458# 0.654021f
C31098 a_n2661_45010# a_n356_44636# 0.091266f
C31099 a_5205_44484# a_4223_44672# 0.235572f
C31100 a_5111_44636# a_8103_44636# 0.001535f
C31101 a_n2017_45002# a_n1809_44850# 0.001936f
C31102 a_3823_42558# a_1823_45246# 0.137565f
C31103 a_1755_42282# a_4185_45028# 0.023564f
C31104 a_2075_43172# a_n443_42852# 1.18e-20
C31105 a_10083_42826# a_n357_42282# 0.017324f
C31106 a_20922_43172# a_13259_45724# 7.71e-21
C31107 a_n784_42308# a_8199_44636# 3.13e-20
C31108 a_17538_32519# RST_Z 0.050782f
C31109 a_10193_42453# a_765_45546# 1.36e-19
C31110 a_14495_45572# a_14513_46634# 1.75e-20
C31111 a_11787_45002# a_5807_45002# 1.03e-21
C31112 a_15415_45028# a_12549_44172# 1.12e-20
C31113 a_16147_45260# a_6755_46942# 0.001071f
C31114 a_2437_43646# a_4646_46812# 9.69e-20
C31115 a_3065_45002# a_n743_46660# 4.32e-20
C31116 a_3537_45260# a_n1925_46634# 4.08e-19
C31117 a_413_45260# a_383_46660# 1.7e-20
C31118 a_5147_45002# a_n2293_46634# 0.009806f
C31119 a_327_44734# a_601_46902# 6.92e-20
C31120 a_14403_45348# a_10227_46804# 1.32e-19
C31121 a_16922_45042# a_11599_46634# 1.05e-19
C31122 a_18315_45260# a_12861_44030# 0.009909f
C31123 a_n83_35174# VDD 0.313947f
C31124 a_949_44458# a_n237_47217# 0.002359f
C31125 a_4223_44672# a_n971_45724# 0.006952f
C31126 a_n2129_44697# a_584_46384# 1.52e-20
C31127 a_3080_42308# a_1736_39587# 1.8e-19
C31128 a_5649_42852# a_5267_42460# 0.016079f
C31129 a_n3674_39304# a_n1630_35242# 2.14e-19
C31130 a_743_42282# a_5421_42558# 0.001222f
C31131 a_n4251_39392# VDD 3.95e-19
C31132 a_4915_47217# a_10037_47542# 1.22e-19
C31133 a_6851_47204# a_n881_46662# 0.002875f
C31134 a_7227_47204# a_n1613_43370# 2.15e-20
C31135 a_n2288_47178# a_n2104_46634# 3.21e-19
C31136 SMPL_ON_P a_n2661_46634# 0.0112f
C31137 a_n2497_47436# a_n2312_38680# 3.06e-19
C31138 a_n2109_47186# a_n2293_46634# 3.45e-19
C31139 a_n1920_47178# a_n2442_46660# 0.00281f
C31140 a_n1605_47204# a_n2956_39768# 2.5e-19
C31141 a_16588_47582# a_12465_44636# 1.91e-19
C31142 a_10227_46804# a_4883_46098# 0.200137f
C31143 a_18479_47436# a_13507_46334# 0.033523f
C31144 a_22223_45036# a_22315_44484# 0.011923f
C31145 a_n2661_43370# a_2998_44172# 9.42e-20
C31146 a_14537_43396# a_14955_43940# 0.104291f
C31147 a_n2293_42834# a_7542_44172# 0.010138f
C31148 a_1307_43914# a_10949_43914# 0.062121f
C31149 a_13249_42308# a_13667_43396# 0.004219f
C31150 a_11823_42460# a_14955_43396# 5.12e-19
C31151 a_12607_44458# a_14815_43914# 6.91e-21
C31152 a_18114_32519# a_20640_44752# 9.12e-19
C31153 a_11322_45546# a_12293_43646# 9.9e-20
C31154 a_11827_44484# a_20397_44484# 3.81e-19
C31155 a_15764_42576# a_n443_42852# 1.17e-20
C31156 a_13258_32519# a_20205_31679# 0.054848f
C31157 a_18691_45572# VDD 0.191893f
C31158 a_5534_30871# VIN_N 0.00357f
C31159 a_11963_45334# a_3483_46348# 0.016005f
C31160 a_17517_44484# a_20916_46384# 4.81e-21
C31161 a_20193_45348# a_19466_46812# 0.00748f
C31162 a_19279_43940# a_12549_44172# 0.062614f
C31163 a_n2661_43922# a_2107_46812# 0.027806f
C31164 a_15903_45785# a_13259_45724# 0.064252f
C31165 a_16147_45260# a_8049_45260# 0.005281f
C31166 a_19963_31679# a_10809_44734# 1.75e-20
C31167 a_413_45260# a_13351_46090# 3.41e-21
C31168 a_6171_45002# a_8016_46348# 0.022961f
C31169 a_5205_44484# a_6419_46155# 1.38e-21
C31170 a_4927_45028# a_5937_45572# 2.22e-19
C31171 a_5111_44636# a_8953_45546# 0.181796f
C31172 a_20447_31679# a_6945_45028# 5.49e-19
C31173 a_4921_42308# a_5932_42308# 0.194195f
C31174 a_3823_42558# a_5934_30871# 1.35e-20
C31175 a_5379_42460# a_6123_31319# 0.011994f
C31176 a_n784_42308# a_13070_42354# 1.96e-20
C31177 a_13291_42460# a_7174_31319# 4.88e-21
C31178 a_5421_42558# a_5755_42308# 1.68e-19
C31179 a_n1630_35242# a_5742_30871# 1.85829f
C31180 a_17364_32525# C6_N_btm 2.76e-20
C31181 a_22609_37990# a_22717_36887# 0.08947f
C31182 a_22705_37990# a_22717_37285# 9.87e-19
C31183 a_18479_47436# a_20623_46660# 0.005343f
C31184 a_13717_47436# a_11415_45002# 4.62e-20
C31185 a_10227_46804# a_21188_46660# 0.22222f
C31186 a_12861_44030# a_20202_43084# 0.020377f
C31187 a_18597_46090# a_20273_46660# 3.9e-19
C31188 a_2063_45854# a_3147_46376# 0.005517f
C31189 a_n443_46116# a_376_46348# 0.025241f
C31190 a_n1151_42308# a_2202_46116# 1.13e-21
C31191 a_584_46384# a_3483_46348# 0.00258f
C31192 a_3160_47472# a_167_45260# 2.66e-19
C31193 a_3381_47502# a_1823_45246# 1.03e-19
C31194 a_n237_47217# a_5497_46414# 0.021428f
C31195 a_n971_45724# a_6419_46155# 0.001374f
C31196 a_n1741_47186# a_5937_45572# 4.26e-20
C31197 a_11453_44696# a_16721_46634# 4.18e-21
C31198 a_12465_44636# a_14447_46660# 1.13e-19
C31199 a_4883_46098# a_17339_46660# 0.071433f
C31200 a_13507_46334# a_17829_46910# 8.95e-19
C31201 a_3055_46660# a_3877_44458# 2.12e-19
C31202 a_n2661_46634# a_8035_47026# 0.002111f
C31203 a_2443_46660# a_3633_46660# 2.56e-19
C31204 a_n1925_46634# a_6969_46634# 0.007338f
C31205 a_2107_46812# a_7927_46660# 5.88e-20
C31206 a_n743_46660# a_10249_46116# 0.004613f
C31207 a_5807_45002# a_11813_46116# 0.037525f
C31208 a_12549_44172# a_15368_46634# 0.012256f
C31209 a_5343_44458# a_4905_42826# 7.39e-21
C31210 a_n2065_43946# a_n1441_43940# 9.73e-19
C31211 a_n699_43396# a_n1557_42282# 0.02911f
C31212 a_742_44458# a_2896_43646# 8.3e-20
C31213 a_n1549_44318# a_n1453_44318# 0.013793f
C31214 a_n1331_43914# a_n1287_44306# 3.69e-19
C31215 a_n1899_43946# a_n875_44318# 2.36e-20
C31216 a_n2661_42834# a_2455_43940# 0.002019f
C31217 a_11967_42832# a_18451_43940# 0.01235f
C31218 a_14815_43914# a_14761_44260# 1.48e-19
C31219 a_16112_44458# a_n97_42460# 1.17e-19
C31220 a_n984_44318# a_n3674_39768# 4.73e-20
C31221 a_n913_45002# a_10518_42984# 0.058603f
C31222 a_n2017_45002# a_10796_42968# 1.01e-19
C31223 a_n1059_45260# a_10835_43094# 0.004669f
C31224 a_2382_45260# a_2905_42968# 7.68e-19
C31225 a_3065_45002# a_1847_42826# 2.79e-20
C31226 a_12883_44458# VDD 0.263743f
C31227 a_n4209_39590# C9_P_btm 0.786375f
C31228 a_n4064_40160# C5_P_btm 1.78e-19
C31229 a_22465_38105# RST_Z 0.034434f
C31230 a_17730_32519# a_20820_30879# 0.052913f
C31231 a_4093_43548# a_n2293_46634# 0.007782f
C31232 a_7287_43370# a_768_44030# 6.62e-20
C31233 a_14955_43940# a_3090_45724# 0.018423f
C31234 a_10341_43396# SMPL_ON_N 4.16e-20
C31235 a_17499_43370# a_16327_47482# 0.34052f
C31236 a_16243_43396# a_10227_46804# 0.001446f
C31237 a_n13_43084# a_n746_45260# 7.03e-21
C31238 a_33_46660# VDD 0.272723f
C31239 a_n4209_39304# a_n4334_39392# 0.253307f
C31240 a_n4315_30879# a_n4064_38528# 0.034153f
C31241 a_n4064_40160# a_n3420_38528# 0.057096f
C31242 a_n4209_39590# a_n4209_38502# 0.031979f
C31243 a_14035_46660# a_11415_45002# 3.1e-21
C31244 a_11901_46660# a_3483_46348# 4.96e-21
C31245 a_19551_46910# a_20411_46873# 6.03e-20
C31246 a_16388_46812# a_18280_46660# 3.41e-20
C31247 a_19123_46287# a_20273_46660# 7.53e-20
C31248 a_2443_46660# a_526_44458# 3.42e-19
C31249 a_2609_46660# a_2981_46116# 0.001665f
C31250 a_2107_46812# a_6419_46482# 5.65e-19
C31251 a_6755_46942# a_9290_44172# 3.62e-19
C31252 a_10467_46802# a_10903_43370# 8.89e-21
C31253 a_10249_46116# a_11189_46129# 1.33e-19
C31254 a_7411_46660# a_2324_44458# 1.67e-21
C31255 a_4817_46660# a_6945_45028# 8.99e-21
C31256 a_18579_44172# a_19095_43396# 1.8e-19
C31257 a_n2293_42834# a_n1630_35242# 0.007885f
C31258 a_n2661_43922# a_7871_42858# 7.71e-21
C31259 a_n2661_42834# a_7765_42852# 2.1e-21
C31260 a_9313_44734# a_10922_42852# 0.002978f
C31261 a_n2661_42282# a_6643_43396# 1.74e-19
C31262 a_n2017_45002# a_4958_30871# 0.053522f
C31263 a_19479_31679# a_13258_32519# 0.054577f
C31264 a_n1059_45260# a_16269_42308# 1.17e-19
C31265 a_16680_45572# a_17668_45572# 1.69e-19
C31266 a_2711_45572# a_13777_45326# 0.008866f
C31267 a_8696_44636# a_17568_45572# 2.55e-19
C31268 a_7499_43078# a_3537_45260# 0.586701f
C31269 VDAC_P EN_VIN_BSTR_P 0.340512f
C31270 a_n3420_37440# C3_P_btm 2.18e-19
C31271 a_n4064_37440# C5_P_btm 1.49e-19
C31272 VDAC_N a_11530_34132# 0.022899f
C31273 a_9145_43396# a_11415_45002# 8.88e-21
C31274 a_4190_30871# a_19692_46634# 0.013919f
C31275 a_5649_42852# a_3090_45724# 4.39e-22
C31276 a_5013_44260# a_n443_42852# 6.73e-20
C31277 a_10555_44260# a_10586_45546# 3.3e-20
C31278 a_17973_43940# a_16375_45002# 8.39e-19
C31279 a_261_44278# a_n357_42282# 1.78e-19
C31280 a_19721_31679# RST_Z 0.050546f
C31281 a_12005_46116# VDD 0.518463f
C31282 a_6194_45824# a_2063_45854# 0.041827f
C31283 a_2711_45572# a_n1151_42308# 0.039506f
C31284 a_4099_45572# a_2905_45572# 1.64e-20
C31285 a_1990_45572# a_n237_47217# 2.46e-19
C31286 a_3175_45822# a_3160_47472# 7.95e-19
C31287 a_n4064_38528# a_n3420_37440# 0.050813f
C31288 a_n3420_38528# a_n4064_37440# 0.045626f
C31289 a_5937_45572# a_10586_45546# 1.5e-19
C31290 a_8016_46348# a_9751_46155# 0.001112f
C31291 a_9290_44172# a_8049_45260# 0.041148f
C31292 a_n2956_39304# a_n1736_46482# 1.91e-20
C31293 a_n2293_46098# a_n2840_45546# 0.004047f
C31294 a_n2840_46090# a_n2661_45546# 0.003502f
C31295 a_8147_43396# a_4361_42308# 2.94e-21
C31296 a_10341_43396# a_17499_43370# 0.022768f
C31297 a_n97_42460# a_7227_42852# 0.117893f
C31298 a_9313_44734# a_17531_42308# 4.72e-20
C31299 a_9145_43396# a_15037_43396# 5.99e-20
C31300 a_1414_42308# a_n3674_37592# 2.19e-21
C31301 a_8685_43396# a_16855_43396# 8.49e-20
C31302 a_3935_42891# VDD 0.096403f
C31303 a_n2956_37592# a_n2860_37984# 9.05e-19
C31304 a_n2810_45028# a_n2216_37984# 3.1e-19
C31305 a_12427_45724# a_n2661_43922# 1.65e-19
C31306 a_11823_42460# a_n2661_42834# 4.26e-20
C31307 a_15861_45028# a_16979_44734# 4.51e-19
C31308 a_7499_43078# a_11541_44484# 0.048175f
C31309 a_8696_44636# a_17767_44458# 3.64e-19
C31310 a_4574_45260# a_n2661_43370# 0.007993f
C31311 a_5205_44484# a_n2293_42834# 4.84e-20
C31312 a_6171_45002# a_8488_45348# 8.23e-19
C31313 a_19963_31679# a_22959_45036# 0.002114f
C31314 a_21363_45546# a_19721_31679# 2.83e-19
C31315 a_7963_42308# a_3090_45724# 4e-21
C31316 a_n4209_39304# a_n2312_38680# 0.062228f
C31317 a_10796_42968# a_526_44458# 1.9e-20
C31318 a_8192_45572# a_4646_46812# 1.94e-19
C31319 a_9049_44484# a_6755_46942# 5.93e-20
C31320 a_10193_42453# a_10623_46897# 5.98e-20
C31321 a_10490_45724# a_10428_46928# 1.87e-20
C31322 a_17668_45572# a_13747_46662# 2.27e-19
C31323 a_2711_45572# a_14084_46812# 1.95e-20
C31324 a_2437_43646# a_9804_47204# 0.005678f
C31325 a_n2661_43370# a_n2497_47436# 0.031125f
C31326 a_n2293_42834# a_n971_45724# 0.088674f
C31327 a_2232_45348# a_n443_46116# 8.27e-19
C31328 a_3232_43370# a_10227_46804# 0.028168f
C31329 a_13017_45260# a_12861_44030# 0.032265f
C31330 a_413_45260# a_22223_47212# 0.001872f
C31331 a_7287_43370# a_6123_31319# 2.73e-19
C31332 a_5534_30871# a_5342_30871# 11.128201f
C31333 a_7112_43396# a_7227_42308# 4.93e-21
C31334 a_n97_42460# a_11633_42308# 0.00291f
C31335 a_15743_43084# a_20836_43172# 3.08e-19
C31336 a_17730_32519# C8_N_btm 0.001799f
C31337 a_19237_31679# C6_N_btm 1.26e-20
C31338 a_15890_42674# VDD 0.203548f
C31339 a_5815_47464# a_6151_47436# 0.235454f
C31340 a_4915_47217# a_6491_46660# 0.19739f
C31341 a_5129_47502# a_6545_47178# 1.1e-19
C31342 a_2952_47436# a_n1435_47204# 2.1e-19
C31343 a_n1151_42308# a_9313_45822# 0.024431f
C31344 a_4791_45118# a_7227_47204# 6.26e-19
C31345 a_18184_42460# a_9313_44734# 0.069472f
C31346 a_n4318_40392# a_n2012_44484# 7.25e-20
C31347 a_5343_44458# a_8975_43940# 1.49e-20
C31348 a_4574_45260# a_2998_44172# 1.08e-19
C31349 a_3537_45260# a_3600_43914# 0.157156f
C31350 a_n913_45002# a_n822_43940# 1.95e-19
C31351 a_2903_42308# a_n863_45724# 0.007352f
C31352 a_196_42282# a_n443_42852# 3.14e-19
C31353 a_2123_42473# a_n755_45592# 0.022891f
C31354 a_10490_45724# VDD 0.162001f
C31355 a_4190_30871# VIN_N 0.049977f
C31356 a_22591_43396# RST_Z 3.24e-19
C31357 a_18248_44752# a_13661_43548# 0.019034f
C31358 a_6298_44484# a_n743_46660# 1.32e-20
C31359 a_10157_44484# a_n2293_46634# 5.67e-21
C31360 a_n913_45002# a_20202_43084# 0.322116f
C31361 a_n2661_44458# a_1799_45572# 3.78e-20
C31362 a_3602_45348# a_3090_45724# 4.94e-19
C31363 a_9049_44484# a_8049_45260# 0.002717f
C31364 a_8746_45002# a_8034_45724# 2.6e-20
C31365 a_16115_45572# a_15682_46116# 0.008647f
C31366 a_8696_44636# a_15015_46420# 5.75e-21
C31367 a_13297_45572# a_10903_43370# 0.00546f
C31368 a_15765_45572# a_17715_44484# 4.5e-19
C31369 a_12649_45572# a_12594_46348# 2.33e-19
C31370 a_n2661_43922# a_11453_44696# 0.009016f
C31371 a_14581_44484# a_10227_46804# 1.42e-20
C31372 a_18204_44850# a_16327_47482# 1.7e-19
C31373 a_19006_44850# a_12861_44030# 0.008813f
C31374 a_2998_44172# a_n2497_47436# 1.03e-19
C31375 a_644_44056# a_n746_45260# 9.68e-19
C31376 a_n4318_37592# a_n1329_42308# 7.71e-21
C31377 a_19339_43156# a_17303_42282# 4.17e-21
C31378 a_18249_42858# a_18727_42674# 6.54e-20
C31379 a_n3674_38680# a_n3674_37592# 0.028019f
C31380 a_n4318_38216# a_n784_42308# 3.7e-22
C31381 a_n2661_46634# a_n2438_43548# 0.493975f
C31382 a_n2104_46634# a_n2312_38680# 0.154937f
C31383 a_n2293_46634# a_n1925_46634# 0.051324f
C31384 a_n2442_46660# a_n1021_46688# 2.1e-20
C31385 a_n881_46662# a_4651_46660# 1.63e-19
C31386 a_n1613_43370# a_4955_46873# 0.051259f
C31387 a_4883_46098# a_10467_46802# 7.03e-19
C31388 a_11599_46634# a_11186_47026# 1.68e-20
C31389 a_n1435_47204# a_12991_46634# 6.91e-20
C31390 a_n1151_42308# a_12513_46660# 1.2e-19
C31391 a_949_44458# a_1241_43940# 3.56e-19
C31392 a_10440_44484# a_10555_44260# 0.001321f
C31393 a_8696_44636# a_8037_42858# 2.6e-21
C31394 a_15004_44636# a_11341_43940# 2.28e-20
C31395 a_18443_44721# a_15493_43396# 1.69e-21
C31396 a_20679_44626# a_20512_43084# 0.003019f
C31397 a_11967_42832# a_19237_31679# 2.2e-20
C31398 a_n2661_43922# a_n3674_39768# 0.152656f
C31399 a_18989_43940# a_18451_43940# 0.114286f
C31400 a_14537_43396# a_8685_43396# 0.007467f
C31401 a_18184_42460# a_20974_43370# 3.83e-20
C31402 a_20835_44721# a_21145_44484# 0.013793f
C31403 a_20766_44850# a_21073_44484# 3.69e-19
C31404 a_n2661_42834# a_n1644_44306# 0.006513f
C31405 a_19279_43940# a_20637_44484# 9.22e-19
C31406 a_20640_44752# a_22485_44484# 8.77e-20
C31407 a_n2293_43922# a_n4318_39768# 3.58e-19
C31408 a_5891_43370# a_6756_44260# 4.32e-21
C31409 a_7640_43914# a_7911_44260# 1.97e-19
C31410 a_21513_45002# a_21487_43396# 9.71e-22
C31411 en_comp a_15743_43084# 5.37e-21
C31412 a_5111_44636# a_10149_43396# 0.001625f
C31413 a_5742_30871# a_11530_34132# 7.08e-19
C31414 a_n356_44636# a_1138_42852# 0.29814f
C31415 a_18443_44721# a_3483_46348# 1.15e-20
C31416 a_9313_44734# a_12741_44636# 1.82e-21
C31417 a_20980_44850# a_15227_44166# 7.56e-21
C31418 a_9420_43940# a_768_44030# 0.001442f
C31419 a_10057_43914# a_8199_44636# 0.113262f
C31420 a_19647_42308# a_20107_42308# 4.99e-19
C31421 a_19511_42282# a_20712_42282# 0.05034f
C31422 a_18907_42674# a_18997_42308# 0.004764f
C31423 a_5934_30871# a_1177_38525# 1.19e-19
C31424 a_17303_42282# a_22465_38105# 3.32e-19
C31425 a_21811_47423# VDD 0.201359f
C31426 a_4883_46098# a_8034_45724# 0.004608f
C31427 a_11599_46634# a_12839_46116# 0.042002f
C31428 a_13717_47436# a_13259_45724# 2.52e-20
C31429 a_12861_44030# a_14383_46116# 1.08e-19
C31430 a_n2109_47186# a_2277_45546# 3e-21
C31431 a_n746_45260# a_n23_45546# 0.004336f
C31432 a_n1151_42308# a_n1079_45724# 0.012662f
C31433 a_584_46384# a_n357_42282# 0.107436f
C31434 a_n237_47217# a_n356_45724# 1.25e-20
C31435 a_4007_47204# a_n2661_45546# 2.2e-21
C31436 a_n971_45724# a_n310_45899# 0.002723f
C31437 a_11309_47204# a_6945_45028# 0.010402f
C31438 a_n1613_43370# a_n967_46494# 2.95e-19
C31439 a_5807_45002# a_15682_46116# 0.062679f
C31440 a_2107_46812# a_5164_46348# 0.002137f
C31441 a_n743_46660# a_5937_45572# 0.02494f
C31442 a_13661_43548# a_2324_44458# 0.307974f
C31443 a_12549_44172# a_20708_46348# 1.12e-20
C31444 a_19333_46634# a_19466_46812# 0.167526f
C31445 a_12469_46902# a_14180_46812# 4.58e-22
C31446 a_15227_44166# a_19692_46634# 0.116169f
C31447 a_n2661_46098# a_2698_46116# 3.89e-20
C31448 a_2443_46660# a_2521_46116# 5.25e-19
C31449 a_4955_46873# a_n2293_46098# 0.002285f
C31450 a_9313_44734# a_15868_43402# 6.39e-20
C31451 a_11967_42832# a_9145_43396# 8.37e-19
C31452 a_n699_43396# a_3935_42891# 9.41e-22
C31453 a_4223_44672# a_4520_42826# 6.71e-22
C31454 a_11827_44484# a_17595_43084# 1.44e-20
C31455 a_11691_44458# a_5342_30871# 1.35e-19
C31456 a_18494_42460# a_18817_42826# 5.74e-19
C31457 a_18184_42460# a_18599_43230# 1.68e-19
C31458 a_15493_43940# a_15301_44260# 1.97e-19
C31459 a_10729_43914# a_11173_43940# 0.00134f
C31460 a_10949_43914# a_10867_43940# 3.29e-19
C31461 a_10807_43548# a_10651_43940# 3.34e-19
C31462 a_1467_44172# a_n1557_42282# 7.5e-21
C31463 a_n356_44636# a_5649_42852# 0.023625f
C31464 a_2382_45260# a_n784_42308# 1.58e-20
C31465 en_comp a_1606_42308# 0.022666f
C31466 a_n2017_45002# a_2725_42558# 6.21e-19
C31467 a_6453_43914# VDD 0.194953f
C31468 a_15143_45578# a_15903_45785# 8.61e-19
C31469 a_10907_45822# a_11136_45572# 0.080042f
C31470 a_10490_45724# a_12749_45572# 4.85e-22
C31471 a_14495_45572# a_15765_45572# 1.19e-20
C31472 a_17538_32519# a_20820_30879# 0.052874f
C31473 a_8685_43396# a_3090_45724# 2.11639f
C31474 a_12545_42858# a_12549_44172# 3.73e-20
C31475 a_10341_43396# a_8270_45546# 5.91e-19
C31476 a_10729_43914# a_10809_44734# 6.71e-21
C31477 a_11173_44260# a_9290_44172# 0.0082f
C31478 a_n4318_38216# SMPL_ON_P 0.037528f
C31479 COMP_P a_n2497_47436# 1.63e-20
C31480 a_22000_46634# VDD 0.257047f
C31481 a_15764_42576# CAL_N 9.17e-19
C31482 a_n3565_39590# a_n2302_37984# 8.95e-20
C31483 a_n1991_46122# a_n1736_46482# 0.06121f
C31484 a_n1641_46494# a_n2956_39304# 2.7e-20
C31485 a_n1423_46090# a_n2956_38680# 7.5e-20
C31486 a_n2293_46098# a_n967_46494# 4.35e-20
C31487 a_14035_46660# a_13259_45724# 1.96e-19
C31488 a_20273_46660# a_8049_45260# 2.63e-21
C31489 a_14180_46812# a_14383_46116# 1.22e-20
C31490 a_15227_44166# a_20692_30879# 1.69e-19
C31491 a_4185_45028# a_2324_44458# 0.015434f
C31492 a_9625_46129# a_10355_46116# 0.001354f
C31493 a_8199_44636# a_11133_46155# 2.47e-20
C31494 a_8016_46348# a_10903_43370# 6.55e-20
C31495 a_8953_45546# a_9290_44172# 0.373944f
C31496 a_3626_43646# a_14205_43396# 3.91e-21
C31497 a_2982_43646# a_14955_43396# 1.35e-20
C31498 a_n97_42460# a_17499_43370# 0.005876f
C31499 a_20193_45348# a_13258_32519# 0.001033f
C31500 a_n2661_42834# a_961_42354# 1.54e-21
C31501 a_n2293_43922# a_1576_42282# 8.6e-20
C31502 a_n356_44636# a_7963_42308# 1.17e-19
C31503 a_6765_43638# a_7221_43396# 4.2e-19
C31504 a_3905_42865# a_3059_42968# 4.87e-20
C31505 a_6151_47436# CLK 0.036587f
C31506 a_7227_47204# DATA[3] 0.357377f
C31507 a_16547_43609# VDD 0.31275f
C31508 a_3537_45260# a_4558_45348# 0.236111f
C31509 a_3065_45002# a_5111_44636# 9.21e-21
C31510 a_16855_45546# a_16922_45042# 0.002263f
C31511 a_7499_43078# a_8701_44490# 0.011795f
C31512 a_8387_43230# a_4185_45028# 1.29e-20
C31513 a_20922_43172# a_20202_43084# 2.39e-19
C31514 a_1755_42282# a_5257_43370# 2.9e-20
C31515 a_14113_42308# a_n2293_46634# 1.19e-21
C31516 a_16877_43172# a_15227_44166# 1.05e-20
C31517 a_9145_43396# a_13259_45724# 0.155949f
C31518 a_4699_43561# a_n443_42852# 0.004673f
C31519 a_n144_43396# a_n357_42282# 5.4e-19
C31520 a_n4209_39590# a_n2312_39304# 0.065703f
C31521 a_22591_44484# RST_Z 5.01e-19
C31522 a_13904_45546# a_5807_45002# 0.009766f
C31523 a_7499_43078# a_n2293_46634# 0.14773f
C31524 a_13163_45724# a_13747_46662# 8.69e-21
C31525 a_10180_45724# a_n2661_46634# 3.78e-20
C31526 a_13527_45546# a_13661_43548# 5.13e-20
C31527 a_17478_45572# a_11453_44696# 5.17e-21
C31528 a_13485_45572# a_13507_46334# 1.11e-19
C31529 a_18175_45572# a_18479_47436# 1.22e-21
C31530 a_18479_45785# a_18143_47464# 2.32e-21
C31531 a_17668_45572# a_11599_46634# 5.66e-19
C31532 a_18596_45572# a_16327_47482# 0.00301f
C31533 a_20107_45572# a_12861_44030# 2.65e-22
C31534 a_2437_43646# a_6545_47178# 0.010642f
C31535 a_3357_43084# a_5129_47502# 0.001711f
C31536 a_413_45260# a_n971_45724# 0.937818f
C31537 a_n37_45144# a_n746_45260# 0.031257f
C31538 a_n913_45002# a_2063_45854# 2.32e-21
C31539 a_16823_43084# a_17701_42308# 2.64e-19
C31540 a_15743_43084# a_22165_42308# 0.008223f
C31541 a_5649_42852# a_12379_42858# 5.88e-20
C31542 a_4361_42308# a_13113_42826# 1.92e-20
C31543 a_743_42282# a_5534_30871# 0.030281f
C31544 a_n4318_39768# a_n3420_39616# 0.002167f
C31545 a_n3674_39768# a_n3690_39616# 0.07198f
C31546 a_4190_30871# a_5342_30871# 0.0276f
C31547 a_7754_39632# a_8530_39574# 1.05e-19
C31548 a_3754_39134# VDAC_Ni 0.00194f
C31549 a_n3674_37592# VDD 0.357168f
C31550 a_n2833_47464# a_n2288_47178# 0.003549f
C31551 a_11652_45724# a_11341_43940# 8.54e-21
C31552 a_n2661_43370# a_5883_43914# 1.78e-19
C31553 a_1307_43914# a_7640_43914# 0.006778f
C31554 a_7499_43078# a_11816_44260# 0.002269f
C31555 a_18494_42460# a_20205_45028# 0.001453f
C31556 a_8953_45002# a_9159_44484# 1.62e-19
C31557 a_n1059_45260# a_11967_42832# 0.627158f
C31558 a_22465_38105# a_20820_30879# 5.82e-19
C31559 a_8495_42852# a_n755_45592# 0.001078f
C31560 a_6101_43172# a_n443_42852# 7.15e-19
C31561 a_14456_42282# a_9290_44172# 1.41e-20
C31562 a_11633_42558# a_10903_43370# 9.37e-21
C31563 CAL_N a_13507_46334# 0.004017f
C31564 a_15037_45618# a_12741_44636# 1.47e-21
C31565 a_15599_45572# a_11415_45002# 0.007945f
C31566 a_13249_42308# a_3483_46348# 0.338396f
C31567 a_17478_45572# a_17639_46660# 2.83e-21
C31568 a_16922_45042# a_13661_43548# 0.080391f
C31569 a_17023_45118# a_5807_45002# 1.36e-21
C31570 a_21101_45002# a_12549_44172# 0.00335f
C31571 a_18341_45572# a_17339_46660# 0.015732f
C31572 a_2437_43646# a_19692_46634# 0.293918f
C31573 a_3357_43084# a_15227_44166# 0.026794f
C31574 a_8191_45002# a_7577_46660# 7.23e-22
C31575 a_10180_45724# a_8199_44636# 0.216999f
C31576 a_6667_45809# a_2324_44458# 4.9e-20
C31577 a_9049_44484# a_8953_45546# 0.03092f
C31578 a_8746_45002# a_8016_46348# 0.078716f
C31579 a_10053_45546# a_5937_45572# 1.28e-19
C31580 a_8375_44464# a_4791_45118# 0.010645f
C31581 a_3363_44484# a_584_46384# 2.51e-20
C31582 a_18374_44850# a_12861_44030# 0.004423f
C31583 a_8975_43940# a_10227_46804# 0.037352f
C31584 a_17970_44736# a_11599_46634# 1.08e-19
C31585 a_4743_44484# a_4883_46098# 5.83e-20
C31586 a_9127_43156# a_9223_42460# 0.001251f
C31587 a_n2293_42282# a_961_42354# 2.32e-19
C31588 a_8952_43230# a_8791_42308# 6.34e-19
C31589 a_5649_42852# a_18727_42674# 1.1e-19
C31590 a_4190_30871# a_20107_42308# 2.08e-20
C31591 a_743_42282# a_19647_42308# 0.005892f
C31592 a_14209_32519# a_4958_30871# 0.030901f
C31593 a_4361_42308# a_18214_42558# 9.81e-20
C31594 a_10341_42308# a_5934_30871# 3.73e-20
C31595 a_20692_30879# EN_OFFSET_CAL 0.004501f
C31596 a_17538_32519# C8_N_btm 0.090298f
C31597 a_14401_32519# C10_N_btm 3.37e-20
C31598 a_13507_46334# a_n2661_46634# 2.61e-20
C31599 a_4915_47217# a_4646_46812# 1.43e-19
C31600 a_n1435_47204# a_n2661_46098# 6.55e-20
C31601 a_n1151_42308# a_6540_46812# 4.39e-20
C31602 a_n1741_47186# a_10554_47026# 1.58e-20
C31603 a_n237_47217# a_8667_46634# 0.171086f
C31604 a_4791_45118# a_4955_46873# 0.001577f
C31605 a_n443_46116# a_4651_46660# 0.060179f
C31606 a_11453_44696# a_19594_46812# 0.041136f
C31607 a_12465_44636# a_21588_30879# 0.053175f
C31608 a_22223_47212# a_20916_46384# 4.95e-19
C31609 a_n1059_45260# a_648_43396# 1.51e-19
C31610 a_2382_45260# a_3080_42308# 0.006891f
C31611 a_7229_43940# a_n97_42460# 6.25e-19
C31612 a_3065_45002# a_4235_43370# 2.44e-20
C31613 a_3357_43084# a_6655_43762# 3.75e-19
C31614 a_17613_45144# a_15493_43396# 1.5e-21
C31615 a_5518_44484# a_5013_44260# 1.4e-19
C31616 a_5343_44458# a_5495_43940# 7.49e-21
C31617 a_4223_44672# a_7281_43914# 0.01814f
C31618 a_16922_45042# a_19862_44208# 0.038132f
C31619 a_14112_44734# a_14673_44172# 5.17e-20
C31620 a_5883_43914# a_2998_44172# 7.17e-21
C31621 a_n4209_38216# a_n2810_45572# 0.195791f
C31622 a_6171_45002# VDD 0.441339f
C31623 a_19721_31679# a_20820_30879# 0.052985f
C31624 a_16922_45042# a_4185_45028# 9.87e-21
C31625 a_2127_44172# a_n2438_43548# 1.46e-19
C31626 a_3600_43914# a_n2293_46634# 2.97e-20
C31627 a_5841_44260# a_768_44030# 1.86e-19
C31628 a_3232_43370# a_8034_45724# 7.93e-21
C31629 a_22223_45572# a_20205_31679# 9.5e-19
C31630 a_7705_45326# a_5066_45546# 3.84e-20
C31631 a_n1059_45260# a_13259_45724# 0.390886f
C31632 a_2437_43646# a_20692_30879# 4.72e-20
C31633 a_1423_45028# a_10809_44734# 3.48e-20
C31634 a_14485_44260# a_10227_46804# 1.37e-20
C31635 a_104_43370# a_n746_45260# 9.55e-19
C31636 a_n2012_43396# a_n971_45724# 1.54e-19
C31637 a_n815_47178# VDD 0.380339f
C31638 a_14456_42282# a_15051_42282# 2.66e-19
C31639 a_n784_42308# a_1239_39587# 6.81e-20
C31640 a_n1630_35242# a_n4064_39616# 7.67e-20
C31641 a_n4318_37592# a_n4334_39392# 7.52e-20
C31642 COMP_P a_n4209_39304# 1.25e-21
C31643 a_20916_46384# a_20731_47026# 6.18e-20
C31644 a_8667_46634# a_8270_45546# 0.046604f
C31645 a_n2438_43548# a_765_45546# 0.081258f
C31646 a_8145_46902# a_8601_46660# 4.2e-19
C31647 a_n743_46660# a_17829_46910# 1.56e-20
C31648 a_n881_46662# a_n1076_46494# 0.018649f
C31649 a_n1613_43370# a_376_46348# 4.03e-19
C31650 a_2747_46873# a_2804_46116# 0.001759f
C31651 a_4883_46098# a_8016_46348# 0.289691f
C31652 a_11599_46634# a_14840_46494# 0.051732f
C31653 a_16327_47482# a_13759_46122# 1.11e-21
C31654 a_12861_44030# a_17715_44484# 3.76e-19
C31655 a_7227_47204# a_6945_45028# 0.01947f
C31656 a_584_46384# a_518_46155# 0.002222f
C31657 a_5891_43370# a_8147_43396# 0.029069f
C31658 a_20679_44626# a_21381_43940# 0.001413f
C31659 a_n356_44636# a_8685_43396# 2.93e-20
C31660 a_14539_43914# a_14955_43396# 0.00238f
C31661 a_n2293_42834# a_4520_42826# 0.01065f
C31662 a_10193_42453# a_12563_42308# 2.67e-19
C31663 a_2711_45572# a_17531_42308# 2.41e-21
C31664 a_644_44056# a_726_44056# 0.004767f
C31665 a_20193_45348# a_20301_43646# 0.005382f
C31666 a_18184_42460# a_13887_32519# 0.03303f
C31667 a_18579_44172# a_19808_44306# 3.69e-19
C31668 a_11827_44484# a_13467_32519# 1.16e-20
C31669 a_3537_45260# a_5193_43172# 0.003266f
C31670 a_n1059_45260# a_9114_42852# 1.72e-19
C31671 a_14673_44172# VDD 0.381917f
C31672 a_n3565_38216# VREF_GND 0.001975f
C31673 a_8162_45546# a_8568_45546# 0.078784f
C31674 a_7230_45938# a_7499_43078# 2.81e-21
C31675 a_2711_45572# a_6977_45572# 0.001232f
C31676 a_3499_42826# a_1823_45246# 0.003055f
C31677 a_17737_43940# a_12741_44636# 2.79e-21
C31678 a_15743_43084# a_13661_43548# 0.092364f
C31679 a_6452_43396# a_4646_46812# 0.013786f
C31680 a_15781_43660# a_n2293_46634# 3.39e-19
C31681 a_10440_44484# a_n443_42852# 1.3e-20
C31682 a_3422_30871# a_22223_46124# 3.23e-21
C31683 a_5244_44056# a_5937_45572# 2.04e-20
C31684 a_3357_43084# EN_OFFSET_CAL 6.03e-21
C31685 a_n3420_39616# C1_P_btm 1.92e-20
C31686 a_n784_42308# a_11206_38545# 3.18e-20
C31687 a_n1630_35242# a_6886_37412# 2.07e-19
C31688 a_13059_46348# a_14275_46494# 0.036863f
C31689 a_15227_46910# a_15015_46420# 3.17e-20
C31690 a_n2293_46634# a_n310_45572# 1.08e-19
C31691 a_19692_46634# a_22959_46124# 1.54e-19
C31692 a_n743_46660# a_n443_42852# 0.378464f
C31693 a_n1925_46634# a_2277_45546# 1.47e-20
C31694 a_10554_47026# a_10586_45546# 8.4e-19
C31695 a_n1991_46122# a_n1641_46494# 0.219633f
C31696 a_n2157_46122# a_n1076_46494# 0.102355f
C31697 a_n1853_46287# a_n901_46420# 0.049679f
C31698 a_n2293_46098# a_376_46348# 0.004986f
C31699 a_n2810_45028# a_n3565_38502# 0.031875f
C31700 en_comp a_n4209_38502# 0.006885f
C31701 a_2127_44172# a_2075_43172# 8.71e-21
C31702 a_8333_44056# a_743_42282# 9.61e-22
C31703 a_19862_44208# a_15743_43084# 0.022478f
C31704 a_2479_44172# a_1847_42826# 0.141223f
C31705 a_1414_42308# a_3681_42891# 0.001924f
C31706 a_15493_43940# a_16409_43396# 0.004011f
C31707 a_11341_43940# a_16759_43396# 1.49e-20
C31708 a_19478_44306# a_19268_43646# 9.35e-20
C31709 a_15493_43396# a_19700_43370# 0.001674f
C31710 a_895_43940# a_791_42968# 5.63e-21
C31711 a_11967_42832# a_19987_42826# 9.2e-21
C31712 a_742_44458# a_1576_42282# 8.56e-19
C31713 a_n1809_43762# a_n1557_42282# 3.46e-21
C31714 a_n2267_43396# a_n1243_43396# 2.36e-20
C31715 a_9313_44734# a_11554_42852# 0.001434f
C31716 a_n2129_43609# a_n998_43396# 0.002155f
C31717 a_n97_42460# a_1987_43646# 5.54e-19
C31718 a_n699_43396# a_n3674_37592# 3.66e-22
C31719 a_n2661_42282# a_4361_42308# 0.034761f
C31720 a_5343_44458# a_n784_42308# 1.26e-20
C31721 a_766_43646# VDD 0.009527f
C31722 a_15037_45618# a_13556_45296# 1.52e-19
C31723 a_2711_45572# a_18184_42460# 0.367034f
C31724 a_10180_45724# a_10903_45394# 8.17e-20
C31725 a_7499_43078# a_8704_45028# 0.001053f
C31726 a_2437_43646# a_3357_43084# 0.424652f
C31727 a_22223_45572# a_19479_31679# 0.155323f
C31728 a_15743_43084# a_4185_45028# 0.061074f
C31729 a_5342_30871# a_15227_44166# 0.01169f
C31730 a_n4318_37592# a_n2312_38680# 0.02327f
C31731 a_n4318_38216# a_n2438_43548# 0.00199f
C31732 a_n784_42308# a_n2956_39768# 8.06e-21
C31733 a_1512_43396# a_526_44458# 3.44e-19
C31734 a_12281_43396# a_10903_43370# 1.87e-19
C31735 a_10149_43396# a_9290_44172# 4.47e-19
C31736 a_15803_42450# a_10227_46804# 0.296174f
C31737 a_15761_42308# a_12861_44030# 2.44e-20
C31738 a_9313_44734# RST_Z 0.002698f
C31739 a_9751_46155# VDD 7.28e-19
C31740 a_14495_45572# a_12861_44030# 2.03e-19
C31741 a_10193_42453# a_10227_46804# 0.039217f
C31742 a_13163_45724# a_11599_46634# 3.12e-20
C31743 a_22959_46124# a_20692_30879# 0.155635f
C31744 a_8049_45260# a_8062_46155# 1.21e-20
C31745 a_9803_43646# a_10083_42826# 0.008857f
C31746 a_18579_44172# a_7174_31319# 0.002404f
C31747 a_21259_43561# a_20556_43646# 9.91e-19
C31748 a_9145_43396# a_10518_42984# 6.43e-20
C31749 a_8685_43396# a_12379_42858# 1.07e-19
C31750 a_16823_43084# a_4361_42308# 1.45e-19
C31751 a_n2661_42282# a_6761_42308# 0.001468f
C31752 a_4190_30871# a_743_42282# 0.18536f
C31753 a_2982_43646# a_n2293_42282# 0.010686f
C31754 a_n1557_42282# a_133_42852# 4.96e-19
C31755 a_18114_32519# C9_N_btm 0.003109f
C31756 a_19721_31679# C8_N_btm 1.65e-20
C31757 a_8292_43218# VDD 0.08228f
C31758 a_n2017_45002# a_n2012_44484# 0.013231f
C31759 a_4927_45028# a_5518_44484# 0.00158f
C31760 a_5691_45260# a_5343_44458# 4.08e-20
C31761 a_3232_43370# a_4743_44484# 1.9e-19
C31762 a_5111_44636# a_6298_44484# 8.64e-20
C31763 a_n2293_45010# a_n1190_44850# 2.46e-19
C31764 a_15599_45572# a_11967_42832# 1.11e-21
C31765 a_11361_45348# a_n2661_43370# 0.009376f
C31766 a_16751_45260# a_16886_45144# 0.008535f
C31767 a_1307_43914# a_16981_45144# 8.73e-21
C31768 a_3318_42354# a_1823_45246# 0.055532f
C31769 a_1606_42308# a_4185_45028# 5.4e-20
C31770 a_19511_42282# a_19692_46634# 1.1e-20
C31771 a_1847_42826# a_n443_42852# 9.74e-19
C31772 a_8952_43230# a_n357_42282# 0.011989f
C31773 a_19987_42826# a_13259_45724# 2.7e-20
C31774 a_20974_43370# RST_Z 0.001986f
C31775 a_2711_45572# a_12741_44636# 0.044854f
C31776 a_11823_42460# a_13059_46348# 0.256727f
C31777 a_14495_45572# a_14180_46812# 3.41e-19
C31778 a_10951_45334# a_5807_45002# 1.45e-20
C31779 a_14797_45144# a_12549_44172# 1.61e-20
C31780 a_10193_42453# a_17339_46660# 0.023481f
C31781 a_14537_43396# a_768_44030# 9.19e-20
C31782 a_10180_45724# a_765_45546# 2.49e-20
C31783 a_2437_43646# a_3877_44458# 9.39e-20
C31784 a_2382_45260# a_n2438_43548# 4.79e-21
C31785 a_327_44734# a_33_46660# 1.67e-20
C31786 a_3429_45260# a_n1925_46634# 2.79e-22
C31787 a_n2017_45002# a_n2661_46098# 1.63e-20
C31788 a_1423_45028# a_n881_46662# 1.63e-19
C31789 a_14309_45348# a_10227_46804# 1.15e-19
C31790 a_17719_45144# a_12861_44030# 2.48e-19
C31791 EN_VIN_BSTR_P VDD 0.917313f
C31792 a_n2661_44458# a_2063_45854# 0.029811f
C31793 a_2779_44458# a_n971_45724# 0.009966f
C31794 a_949_44458# a_n746_45260# 0.00147f
C31795 a_742_44458# a_n237_47217# 0.002559f
C31796 a_n13_43084# a_n1630_35242# 3.65e-20
C31797 a_5342_30871# a_14635_42282# 0.012123f
C31798 a_3080_42308# a_1239_39587# 3.4e-19
C31799 a_n4318_38680# a_n3674_37592# 0.02489f
C31800 a_13113_42826# a_13622_42852# 2.6e-19
C31801 a_743_42282# a_5337_42558# 0.001061f
C31802 a_n2302_39072# VDD 0.355374f
C31803 a_4915_47217# a_9804_47204# 0.072476f
C31804 a_6491_46660# a_n881_46662# 1.53e-19
C31805 a_6851_47204# a_n1613_43370# 2.26e-20
C31806 a_n2497_47436# a_n2104_46634# 0.002384f
C31807 a_n2109_47186# a_n2442_46660# 0.004864f
C31808 a_n2833_47464# a_n2312_38680# 6.08e-20
C31809 a_n2288_47178# a_n2293_46634# 0.011283f
C31810 a_n1741_47186# a_n2661_46634# 0.22396f
C31811 SMPL_ON_P a_n2956_39768# 0.039986f
C31812 a_16763_47508# a_12465_44636# 8.56e-19
C31813 a_18597_46090# a_20894_47436# 2.7e-21
C31814 a_10227_46804# a_21496_47436# 0.007515f
C31815 a_17591_47464# a_4883_46098# 4.46e-20
C31816 a_18479_47436# a_21177_47436# 0.001742f
C31817 a_19386_47436# a_19787_47423# 0.002814f
C31818 a_22223_45036# a_3422_30871# 0.011196f
C31819 a_1307_43914# a_10729_43914# 0.051086f
C31820 a_18184_42460# a_22485_44484# 1.09e-21
C31821 a_11823_42460# a_15095_43370# 0.003619f
C31822 a_18494_42460# a_20512_43084# 0.115057f
C31823 a_13076_44458# a_13468_44734# 0.016359f
C31824 a_12607_44458# a_14112_44734# 2.6e-19
C31825 a_11827_44484# a_22315_44484# 0.013f
C31826 a_20193_45348# a_20596_44850# 1.95e-19
C31827 a_15486_42560# a_n443_42852# 3.9e-21
C31828 a_18909_45814# VDD 0.205795f
C31829 a_18599_43230# RST_Z 8.97e-22
C31830 a_5534_30871# VIN_P 0.00357f
C31831 a_11787_45002# a_3483_46348# 0.019413f
C31832 a_11691_44458# a_19466_46812# 0.008122f
C31833 a_16237_45028# a_15227_44166# 8.33e-19
C31834 a_20766_44850# a_12549_44172# 1.16e-19
C31835 a_n2661_42834# a_2107_46812# 0.028012f
C31836 a_18545_45144# a_3090_45724# 2.17e-19
C31837 a_15599_45572# a_13259_45724# 0.205417f
C31838 a_13249_42308# a_n357_42282# 0.024753f
C31839 a_17786_45822# a_8049_45260# 0.001566f
C31840 a_n1059_45260# a_18189_46348# 7.59e-21
C31841 a_413_45260# a_12594_46348# 4.56e-21
C31842 a_5111_44636# a_5937_45572# 0.06133f
C31843 a_5205_44484# a_6165_46155# 3.92e-22
C31844 a_6171_45002# a_7920_46348# 8.34e-21
C31845 a_3232_43370# a_8016_46348# 0.025981f
C31846 a_564_42282# a_5742_30871# 2.87e-20
C31847 a_4921_42308# a_6171_42473# 0.004176f
C31848 a_3318_42354# a_5934_30871# 1.28e-20
C31849 a_5267_42460# a_6123_31319# 1.13e-20
C31850 a_1606_42308# a_9803_42558# 1.77e-20
C31851 a_n784_42308# a_12563_42308# 3.86e-20
C31852 a_5337_42558# a_5755_42308# 1.15e-19
C31853 a_17364_32525# C5_N_btm 2.13e-20
C31854 a_14209_32519# C7_N_btm 1.64e-19
C31855 a_13507_46334# a_765_45546# 0.045587f
C31856 a_18597_46090# a_20411_46873# 0.070431f
C31857 a_10227_46804# a_21363_46634# 0.273017f
C31858 a_18479_47436# a_20841_46902# 0.006861f
C31859 a_16327_47482# a_16434_46660# 7.88e-19
C31860 a_13717_47436# a_20202_43084# 1.46e-20
C31861 a_2905_45572# a_167_45260# 0.001572f
C31862 a_2063_45854# a_2804_46116# 0.007304f
C31863 a_n443_46116# a_n1076_46494# 0.002776f
C31864 a_n1151_42308# a_1823_45246# 1.93e-19
C31865 a_3160_47472# a_2202_46116# 1.2e-19
C31866 a_584_46384# a_3147_46376# 6.53e-20
C31867 a_n237_47217# a_5204_45822# 0.019965f
C31868 a_n971_45724# a_6165_46155# 1.18e-20
C31869 a_n1741_47186# a_8199_44636# 4.26e-20
C31870 a_11453_44696# a_16388_46812# 0.019353f
C31871 a_n2661_46634# a_7832_46660# 0.001683f
C31872 a_768_44030# a_3090_45724# 0.115303f
C31873 a_n1925_46634# a_6755_46942# 0.12389f
C31874 a_2107_46812# a_8145_46902# 5.47e-21
C31875 a_5807_45002# a_11735_46660# 0.005164f
C31876 a_12549_44172# a_14976_45028# 0.005173f
C31877 a_n913_45002# a_10083_42826# 0.052028f
C31878 a_n1059_45260# a_10518_42984# 0.004826f
C31879 a_n2017_45002# a_10835_43094# 1e-19
C31880 a_2382_45260# a_2075_43172# 3.99e-21
C31881 a_4743_44484# a_4905_42826# 2.27e-19
C31882 a_15433_44458# a_14021_43940# 4.46e-21
C31883 a_2889_44172# a_2998_44172# 0.179664f
C31884 a_11967_42832# a_18326_43940# 0.058879f
C31885 a_17517_44484# a_11341_43940# 7.52e-20
C31886 a_375_42282# a_743_42282# 0.006396f
C31887 a_n1549_44318# a_n1644_44306# 0.049827f
C31888 a_n1331_43914# a_n1453_44318# 3.16e-19
C31889 a_n2661_42834# a_2253_43940# 0.004238f
C31890 a_5891_43370# a_10555_43940# 2.09e-19
C31891 a_n699_43396# a_766_43646# 0.001138f
C31892 a_742_44458# a_1987_43646# 2.71e-19
C31893 a_n809_44244# a_n3674_39768# 1.06e-21
C31894 a_12607_44458# VDD 0.188171f
C31895 a_n4209_39590# C10_P_btm 0.002325f
C31896 a_n4064_40160# C6_P_btm 2.2e-19
C31897 a_17325_44484# a_3483_46348# 0.001497f
C31898 a_19237_31679# a_20202_43084# 2.47e-20
C31899 a_13483_43940# a_3090_45724# 2.45e-20
C31900 a_6547_43396# a_768_44030# 8.31e-20
C31901 a_3080_42308# a_n2956_39768# 4.45e-21
C31902 a_1756_43548# a_n2293_46634# 3.05e-19
C31903 a_13213_44734# a_13351_46090# 1.41e-20
C31904 a_5708_44484# a_2324_44458# 7.43e-19
C31905 a_14955_43396# a_11453_44696# 3.7e-22
C31906 a_16759_43396# a_16327_47482# 0.152273f
C31907 a_16137_43396# a_10227_46804# 0.001438f
C31908 a_16664_43396# a_12861_44030# 2.54e-20
C31909 a_n13_43084# a_n971_45724# 1.75e-19
C31910 a_n1076_43230# a_n746_45260# 8.81e-21
C31911 a_171_46873# VDD 0.539781f
C31912 a_n4064_40160# a_n3690_38528# 2.54e-19
C31913 a_5934_30871# C10_N_btm 1.89e-19
C31914 a_11813_46116# a_3483_46348# 8.59e-21
C31915 a_3090_45724# a_1176_45822# 5.71e-21
C31916 a_19123_46287# a_20411_46873# 1.69e-20
C31917 a_16388_46812# a_17639_46660# 1.85e-19
C31918 a_18285_46348# a_20273_46660# 8.45e-20
C31919 a_2107_46812# a_5066_45546# 0.004218f
C31920 a_2443_46660# a_2981_46116# 1.22e-19
C31921 a_n1925_46634# a_8049_45260# 0.088663f
C31922 a_n2661_46634# a_10586_45546# 0.001458f
C31923 a_5807_45002# a_14537_46482# 6.7e-19
C31924 a_12549_44172# a_18051_46116# 2.41e-20
C31925 a_n743_46660# a_6633_46155# 1.23e-19
C31926 a_5257_43370# a_2324_44458# 0.067403f
C31927 a_6755_46942# a_10355_46116# 3.41e-20
C31928 a_10467_46802# a_11387_46155# 5.52e-19
C31929 a_10428_46928# a_10903_43370# 1.9e-19
C31930 a_10249_46116# a_9290_44172# 2.05e-19
C31931 a_19279_43940# a_4361_42308# 4.21e-21
C31932 a_18579_44172# a_21487_43396# 2.15e-21
C31933 a_n2661_42834# a_7871_42858# 1.63e-20
C31934 a_742_44458# a_4649_42852# 5.01e-21
C31935 a_n2293_43922# a_5755_42852# 3.26e-21
C31936 a_9313_44734# a_10991_42826# 0.007504f
C31937 a_n2293_42834# a_564_42282# 5.42e-20
C31938 a_1307_43914# a_5932_42308# 0.00164f
C31939 a_n2661_43370# a_n4318_37592# 2.73e-20
C31940 a_n2661_42282# a_7274_43762# 9.24e-21
C31941 a_7227_45028# a_8191_45002# 8.51e-20
C31942 a_5437_45600# a_5111_44636# 3.47e-19
C31943 a_2711_45572# a_13556_45296# 0.00137f
C31944 a_8696_44636# a_17034_45572# 4.18e-19
C31945 a_3539_42460# a_4185_45028# 0.065262f
C31946 a_6197_43396# a_1823_45246# 5.44e-21
C31947 a_743_42282# a_15227_44166# 3.95e-19
C31948 a_21259_43561# a_19692_46634# 0.014184f
C31949 a_16137_43396# a_17339_46660# 1.34e-19
C31950 a_17737_43940# a_16375_45002# 0.001093f
C31951 a_5244_44056# a_n443_42852# 5.78e-21
C31952 a_n2661_42282# a_n2810_45572# 3.31e-20
C31953 a_18326_43940# a_13259_45724# 8.21e-19
C31954 a_261_44278# a_310_45028# 6.05e-20
C31955 a_n784_42308# a_10227_46804# 8.64e-21
C31956 a_22469_40625# a_22717_36887# 0.011861f
C31957 VDAC_P a_n923_35174# 0.015621f
C31958 a_n3420_37440# C4_P_btm 2.18e-19
C31959 a_n4064_37440# C6_P_btm 1.49e-19
C31960 a_18114_32519# RST_Z 0.049686f
C31961 a_10903_43370# VDD 2.60588f
C31962 a_5907_45546# a_2063_45854# 0.023999f
C31963 a_3175_45822# a_2905_45572# 0.046585f
C31964 a_n4064_39072# VDAC_P 0.002951f
C31965 a_n3565_38502# a_n2302_37690# 6.13e-19
C31966 a_10355_46116# a_8049_45260# 0.003592f
C31967 a_8199_44636# a_10586_45546# 0.057648f
C31968 a_n2956_39304# a_n2956_38680# 0.163045f
C31969 a_n2840_46090# a_n2810_45572# 4.48e-19
C31970 a_458_43396# a_791_42968# 3.18e-19
C31971 a_10341_43396# a_16759_43396# 0.010617f
C31972 a_n97_42460# a_5755_42852# 0.149651f
C31973 a_9313_44734# a_17303_42282# 9.64e-19
C31974 a_14579_43548# a_15743_43084# 1.21e-19
C31975 a_1414_42308# a_n327_42558# 2.72e-21
C31976 a_n356_44636# a_18997_42308# 1.66e-20
C31977 a_10037_47542# DATA[4] 1.79e-19
C31978 a_3681_42891# VDD 0.223661f
C31979 a_8696_44636# a_16979_44734# 0.005402f
C31980 a_15861_45028# a_14539_43914# 2.35e-19
C31981 a_1307_43914# a_1423_45028# 0.054616f
C31982 a_375_42282# a_626_44172# 0.017957f
C31983 a_7499_43078# a_10809_44484# 3.94e-19
C31984 a_11962_45724# a_n2661_43922# 2.11e-20
C31985 a_3537_45260# a_n2661_43370# 0.087747f
C31986 a_7276_45260# a_7418_45394# 0.007833f
C31987 a_22223_45572# a_20193_45348# 1.1e-19
C31988 a_6171_45002# a_8137_45348# 1.04e-19
C31989 a_6123_31319# a_3090_45724# 3.25e-20
C31990 a_n2946_39072# a_n2956_39768# 0.004795f
C31991 a_19700_43370# a_n357_42282# 6.27e-20
C31992 a_10835_43094# a_526_44458# 1.38e-20
C31993 a_10490_45724# a_10150_46912# 5.77e-22
C31994 a_7499_43078# a_6755_46942# 4.83e-20
C31995 a_10180_45724# a_10623_46897# 5.76e-20
C31996 a_10193_42453# a_10467_46802# 5.21e-20
C31997 a_1423_45028# a_n443_46116# 0.022652f
C31998 a_413_45260# a_12465_44636# 0.28925f
C31999 en_comp a_n2312_39304# 0.001599f
C32000 a_n967_45348# a_n2312_40392# 4.63e-20
C32001 a_2437_43646# a_8128_46384# 0.005098f
C32002 a_509_45822# a_603_45572# 1.26e-19
C32003 a_6547_43396# a_6123_31319# 1.98e-19
C32004 a_7287_43370# a_7227_42308# 1.42e-19
C32005 a_20974_43370# a_17303_42282# 5.91e-22
C32006 a_5534_30871# a_15279_43071# 0.00177f
C32007 a_14543_43071# a_5342_30871# 5.56e-19
C32008 a_7112_43396# a_6761_42308# 1.62e-20
C32009 a_743_42282# a_14635_42282# 0.02914f
C32010 a_15743_43084# a_20573_43172# 3.04e-20
C32011 a_n97_42460# a_10149_42308# 8.69e-19
C32012 a_1847_42826# a_1793_42852# 2.52e-20
C32013 a_17730_32519# C7_N_btm 1.47e-19
C32014 a_19237_31679# C5_N_btm 1.11e-20
C32015 a_15959_42545# VDD 0.19373f
C32016 a_4915_47217# a_6545_47178# 0.033555f
C32017 a_5129_47502# a_6151_47436# 1.77e-19
C32018 a_2553_47502# a_n1435_47204# 4.12e-19
C32019 a_4791_45118# a_6851_47204# 4.68e-20
C32020 a_3537_45260# a_2998_44172# 0.059736f
C32021 a_3232_43370# a_1414_42308# 0.248035f
C32022 a_3065_45002# a_3905_42865# 0.034773f
C32023 a_n473_42460# a_n443_42852# 0.001248f
C32024 a_2713_42308# a_n863_45724# 0.044499f
C32025 a_1755_42282# a_n755_45592# 1.52791f
C32026 a_2123_42473# a_n357_42282# 1.65e-20
C32027 a_8746_45002# VDD 0.970181f
C32028 a_4190_30871# VIN_P 0.049977f
C32029 a_13887_32519# RST_Z 0.048332f
C32030 a_13017_45260# a_14035_46660# 1.07e-19
C32031 a_n2661_43370# a_6969_46634# 5.75e-22
C32032 a_8103_44636# a_n1925_46634# 5.79e-21
C32033 a_18248_44752# a_5807_45002# 4.21e-21
C32034 a_9838_44484# a_n2293_46634# 2.45e-22
C32035 a_17970_44736# a_13661_43548# 2.76e-21
C32036 a_17767_44458# a_13747_46662# 5.22e-21
C32037 a_n356_44636# a_768_44030# 0.098499f
C32038 a_3495_45348# a_3090_45724# 6.6e-19
C32039 a_7499_43078# a_8049_45260# 0.00119f
C32040 a_2711_45572# a_16375_45002# 0.00407f
C32041 a_6109_44484# a_n881_46662# 0.001229f
C32042 a_16333_45814# a_15682_46116# 0.011944f
C32043 a_8696_44636# a_14275_46494# 9.68e-21
C32044 a_15599_45572# a_18189_46348# 2.91e-37
C32045 a_12749_45572# a_10903_43370# 1.89e-20
C32046 a_7640_43914# a_n1613_43370# 2.1e-20
C32047 a_n2661_42834# a_11453_44696# 4.17e-19
C32048 a_13468_44734# a_12465_44636# 1.06e-20
C32049 a_13940_44484# a_10227_46804# 1.36e-20
C32050 a_17517_44484# a_16327_47482# 0.090308f
C32051 a_18588_44850# a_12861_44030# 0.006708f
C32052 a_175_44278# a_n746_45260# 0.159759f
C32053 a_18249_42858# a_18057_42282# 1.52e-19
C32054 a_18599_43230# a_17303_42282# 1.61e-20
C32055 a_n2840_42282# a_n3674_37592# 0.007977f
C32056 a_18083_42858# a_18907_42674# 1.44e-20
C32057 a_5534_30871# a_13258_32519# 0.04166f
C32058 a_n1736_42282# a_n1329_42308# 0.050456f
C32059 a_n4318_37592# COMP_P 0.001501f
C32060 a_n3674_38216# a_n961_42308# 7.46e-20
C32061 a_n3674_39304# a_n4251_39392# 8.42e-19
C32062 a_n2661_46634# a_n743_46660# 0.037388f
C32063 a_n2293_46634# a_n2312_38680# 0.131017f
C32064 a_n2956_39768# a_n2438_43548# 8.21e-19
C32065 a_n2442_46660# a_n1925_46634# 6.55e-19
C32066 a_n881_46662# a_4646_46812# 0.024758f
C32067 a_n1613_43370# a_4651_46660# 0.686447f
C32068 a_4883_46098# a_10428_46928# 0.001889f
C32069 a_13381_47204# a_12991_46634# 4.07e-19
C32070 a_n1741_47186# a_765_45546# 0.536367f
C32071 a_n1151_42308# a_12347_46660# 2.21e-19
C32072 a_13720_44458# a_11341_43940# 2.52e-20
C32073 a_18287_44626# a_15493_43396# 1.74e-20
C32074 a_18374_44850# a_18451_43940# 6.12e-19
C32075 a_11967_42832# a_22959_44484# 4.39e-22
C32076 a_20640_44752# a_20512_43084# 4.38e-19
C32077 a_11691_44458# a_15037_43940# 2.9e-20
C32078 a_n2661_43922# a_n4318_39768# 0.010131f
C32079 a_5891_43370# a_n2661_42282# 0.032052f
C32080 a_1423_45028# a_9396_43370# 5.93e-21
C32081 a_11827_44484# a_19319_43548# 0.00137f
C32082 a_18494_42460# a_21381_43940# 2.36e-20
C32083 a_n2293_42834# a_n1557_42282# 0.034384f
C32084 a_20766_44850# a_20637_44484# 4.2e-19
C32085 a_20835_44721# a_21073_44484# 0.001705f
C32086 a_n2661_42834# a_n3674_39768# 0.150968f
C32087 a_8975_43940# a_9248_44260# 0.001408f
C32088 a_18989_43940# a_18326_43940# 3.26e-20
C32089 a_19279_43940# a_20397_44484# 0.002084f
C32090 a_20679_44626# a_21145_44484# 3.82e-19
C32091 a_7640_43914# a_7584_44260# 5.72e-19
C32092 a_18184_42460# a_14401_32519# 4.69e-20
C32093 a_n1059_45260# a_16867_43762# 1.11e-19
C32094 a_5111_44636# a_9885_43396# 0.004113f
C32095 a_18287_44626# a_3483_46348# 2.49e-19
C32096 a_9313_44734# a_20820_30879# 1.42e-20
C32097 a_9165_43940# a_768_44030# 0.00651f
C32098 a_7911_44260# a_4646_46812# 2.43e-21
C32099 a_5111_44636# a_n443_42852# 0.584506f
C32100 a_9145_43396# a_2063_45854# 1.47e-19
C32101 a_8975_43940# a_8016_46348# 0.01976f
C32102 a_10440_44484# a_8199_44636# 8.12e-19
C32103 a_2711_45572# RST_Z 4.2e-20
C32104 a_19647_42308# a_13258_32519# 0.153411f
C32105 a_19511_42282# a_20107_42308# 0.043647f
C32106 a_17303_42282# a_22397_42558# 0.012536f
C32107 a_4883_46098# VDD 1.12729f
C32108 a_4883_46098# a_8283_46482# 7.98e-20
C32109 a_n746_45260# a_n356_45724# 0.030083f
C32110 a_n237_47217# a_3503_45724# 6.04e-21
C32111 a_n1151_42308# a_n2293_45546# 0.01733f
C32112 a_584_46384# a_310_45028# 0.024195f
C32113 a_1431_47204# a_n755_45592# 1.62e-21
C32114 a_3815_47204# a_n2661_45546# 1.03e-20
C32115 a_n971_45724# a_n23_45546# 4.37e-19
C32116 a_n1613_43370# a_n1379_46482# 0.001903f
C32117 a_2107_46812# a_5068_46348# 0.007279f
C32118 a_n2661_46634# a_11189_46129# 1.44e-19
C32119 a_5807_45002# a_2324_44458# 0.232399f
C32120 a_16131_47204# a_15682_46116# 6.99e-20
C32121 a_n743_46660# a_8199_44636# 0.046048f
C32122 a_13747_46662# a_15015_46420# 1.31e-19
C32123 a_13661_43548# a_14840_46494# 4.52e-20
C32124 a_18834_46812# a_19692_46634# 1.69e-19
C32125 a_12991_46634# a_13170_46660# 0.007399f
C32126 a_12816_46660# a_12925_46660# 0.007416f
C32127 a_15227_44166# a_19466_46812# 0.310201f
C32128 a_n2661_46098# a_2521_46116# 7.45e-20
C32129 a_2443_46660# a_167_45260# 0.012819f
C32130 a_n2017_45002# a_n39_42308# 6.45e-19
C32131 a_n913_45002# a_2351_42308# 0.023646f
C32132 a_3357_43084# a_4921_42308# 2.67e-20
C32133 a_17517_44484# a_10341_43396# 0.001868f
C32134 a_1115_44172# a_n1557_42282# 3.9e-19
C32135 a_n1441_43940# a_n2433_43396# 2.36e-19
C32136 a_4223_44672# a_3935_42891# 8.13e-21
C32137 a_n2661_44458# a_10083_42826# 9.84e-22
C32138 a_18494_42460# a_18249_42858# 8.63e-19
C32139 a_18184_42460# a_18817_42826# 6.72e-20
C32140 a_10405_44172# a_11173_43940# 7.97e-21
C32141 a_10729_43914# a_10867_43940# 0.00501f
C32142 a_10807_43548# a_10555_43940# 1.21e-19
C32143 a_2479_44172# a_4235_43370# 1.29e-20
C32144 a_11691_44458# a_15279_43071# 1.05e-19
C32145 a_5663_43940# VDD 0.133666f
C32146 a_15143_45578# a_15599_45572# 2.96e-19
C32147 a_14495_45572# a_15903_45785# 3.7e-21
C32148 a_11823_42460# a_8696_44636# 0.026654f
C32149 a_10907_45822# a_11064_45572# 0.007306f
C32150 a_10490_45724# a_12649_45572# 4.67e-19
C32151 a_15781_43660# a_6755_46942# 1.89e-20
C32152 a_12379_42858# a_768_44030# 1.38e-20
C32153 a_12545_42858# a_12891_46348# 1.12e-20
C32154 a_9885_43646# a_8270_45546# 0.002107f
C32155 a_12089_42308# a_12549_44172# 1.47e-19
C32156 a_10555_44260# a_9290_44172# 3.43e-21
C32157 a_n2472_42282# SMPL_ON_P 2.48e-19
C32158 a_21188_46660# VDD 0.284105f
C32159 a_n3565_39590# a_n4064_37984# 0.031327f
C32160 a_n3420_39616# a_n3420_37984# 0.047086f
C32161 a_n1853_46287# a_n1736_46482# 0.170096f
C32162 a_n1423_46090# a_n2956_39304# 7.61e-21
C32163 a_n2157_46122# a_n1545_46494# 3.82e-19
C32164 a_n1991_46122# a_n2956_38680# 0.004896f
C32165 a_n2293_46098# a_n1379_46482# 2.44e-19
C32166 a_20411_46873# a_8049_45260# 0.003303f
C32167 a_13885_46660# a_13259_45724# 1.34e-21
C32168 a_13059_46348# a_14371_46494# 0.004662f
C32169 a_15227_44166# a_20205_31679# 3.84e-19
C32170 a_765_45546# a_10586_45546# 4.93e-20
C32171 a_8199_44636# a_11189_46129# 8.81e-19
C32172 a_9625_46129# a_9823_46155# 0.321686f
C32173 a_8953_45546# a_10355_46116# 3.1e-20
C32174 a_12429_44172# a_12089_42308# 1.7e-21
C32175 a_3626_43646# a_14358_43442# 1.37e-20
C32176 a_n97_42460# a_16759_43396# 0.003171f
C32177 a_13483_43940# a_12379_42858# 5.33e-20
C32178 a_n2661_42834# a_1184_42692# 6.05e-21
C32179 a_n2293_43922# a_1067_42314# 3.58e-20
C32180 a_n356_44636# a_6123_31319# 0.169259f
C32181 a_7112_43396# a_7274_43762# 0.006453f
C32182 a_6547_43396# a_6809_43396# 0.001705f
C32183 a_6197_43396# a_7221_43396# 2.36e-20
C32184 a_3905_42865# a_2987_42968# 4.66e-20
C32185 a_2982_43646# a_15095_43370# 4.05e-20
C32186 SMPL_ON_N a_22459_39145# 0.00803f
C32187 a_6851_47204# DATA[3] 0.146601f
C32188 a_16243_43396# VDD 0.39865f
C32189 a_8162_45546# a_5883_43914# 1.03e-21
C32190 a_7499_43078# a_8103_44636# 3.16e-19
C32191 a_9049_44484# a_6298_44484# 2.08e-21
C32192 a_2437_43646# a_626_44172# 2.83e-21
C32193 a_3537_45260# a_4574_45260# 0.234297f
C32194 a_3065_45002# a_5147_45002# 4.34e-21
C32195 a_9127_43156# a_3483_46348# 0.001097f
C32196 a_19987_42826# a_20202_43084# 0.177726f
C32197 a_8605_42826# a_4185_45028# 1.07e-20
C32198 a_4235_43370# a_n443_42852# 0.026532f
C32199 a_n4209_39590# a_n2312_40392# 1.62e-19
C32200 a_22485_44484# RST_Z 4.8e-19
C32201 a_13527_45546# a_5807_45002# 2.96e-20
C32202 a_10053_45546# a_n2661_46634# 2.08e-20
C32203 a_2711_45572# a_2609_46660# 7.29e-21
C32204 a_6428_45938# a_n743_46660# 1.23e-19
C32205 a_8192_45572# a_8128_46384# 2.19e-19
C32206 a_15861_45028# a_11453_44696# 0.044605f
C32207 a_19256_45572# a_16327_47482# 0.235006f
C32208 a_18479_45785# a_10227_46804# 6.39e-22
C32209 a_2437_43646# a_6151_47436# 0.017593f
C32210 a_3357_43084# a_4915_47217# 0.028255f
C32211 a_n143_45144# a_n746_45260# 0.043399f
C32212 a_3537_45260# a_n2497_47436# 7.77e-19
C32213 a_n2661_45010# a_n1151_42308# 0.155007f
C32214 a_n913_45002# a_584_46384# 7.62e-20
C32215 a_n1059_45260# a_2063_45854# 1.14e-20
C32216 a_17737_43940# a_17303_42282# 7.23e-21
C32217 a_104_43370# a_n1630_35242# 5.25e-21
C32218 a_16823_43084# a_17595_43084# 8.04e-20
C32219 a_15743_43084# a_21671_42860# 0.004756f
C32220 a_5649_42852# a_10341_42308# 1.31e-20
C32221 a_4361_42308# a_12545_42858# 1.78e-19
C32222 a_743_42282# a_14543_43071# 2.19e-20
C32223 a_15493_43396# a_17124_42282# 2.88e-21
C32224 a_n3674_39768# a_n3565_39590# 0.128683f
C32225 a_n4318_39768# a_n3690_39616# 3.79e-19
C32226 a_n327_42558# VDD 0.198414f
C32227 a_n2833_47464# a_n2497_47436# 0.217831f
C32228 a_11525_45546# a_11341_43940# 2.62e-20
C32229 a_10907_45822# a_10807_43548# 0.002089f
C32230 a_n2661_43370# a_8701_44490# 2.05e-19
C32231 a_9482_43914# a_9313_44734# 0.060868f
C32232 a_7499_43078# a_11173_44260# 5.58e-19
C32233 a_1307_43914# a_6109_44484# 0.00821f
C32234 a_19778_44110# a_18114_32519# 5.95e-20
C32235 a_11691_44458# a_20193_45348# 0.003224f
C32236 a_18184_42460# a_20205_45028# 0.001438f
C32237 a_n2017_45002# a_11967_42832# 0.086561f
C32238 a_7229_43940# a_n2661_43922# 0.030151f
C32239 a_8495_42852# a_n357_42282# 0.002316f
C32240 a_5837_43172# a_n443_42852# 2.77e-19
C32241 a_13575_42558# a_9290_44172# 0.001995f
C32242 a_11551_42558# a_10903_43370# 9.18e-20
C32243 a_13904_45546# a_3483_46348# 0.125708f
C32244 a_18479_45785# a_17339_46660# 0.027772f
C32245 a_15861_45028# a_17639_46660# 4.98e-21
C32246 a_16922_45042# a_5807_45002# 0.030945f
C32247 a_21005_45260# a_12549_44172# 0.002789f
C32248 a_1307_43914# a_4646_46812# 0.031289f
C32249 a_n2661_43370# a_n2293_46634# 2.59564f
C32250 a_2437_43646# a_19466_46812# 1.21e-19
C32251 a_7705_45326# a_7577_46660# 3.37e-20
C32252 a_21513_45002# a_19692_46634# 0.098725f
C32253 a_n2661_43922# a_n237_47217# 1.49e-20
C32254 a_556_44484# a_584_46384# 0.004299f
C32255 a_7640_43914# a_4791_45118# 0.027432f
C32256 a_18443_44721# a_12861_44030# 0.007707f
C32257 a_10057_43914# a_10227_46804# 0.054198f
C32258 a_17767_44458# a_11599_46634# 0.001378f
C32259 a_7499_43078# a_8953_45546# 0.108436f
C32260 a_9049_44484# a_5937_45572# 0.311862f
C32261 a_6511_45714# a_2324_44458# 0.001394f
C32262 a_10053_45546# a_8199_44636# 0.014322f
C32263 a_10193_42453# a_8016_46348# 0.125497f
C32264 a_4190_30871# a_13258_32519# 0.039476f
C32265 a_8952_43230# a_8685_42308# 0.008199f
C32266 a_n2293_42282# a_1184_42692# 1.61e-19
C32267 a_5649_42852# a_18057_42282# 6.29e-20
C32268 a_743_42282# a_19511_42282# 0.00872f
C32269 a_4361_42308# a_19332_42282# 0.009695f
C32270 a_945_42968# a_n784_42308# 7.59e-20
C32271 a_13887_32519# a_17303_42282# 0.0067f
C32272 a_20205_31679# EN_OFFSET_CAL 0.002855f
C32273 a_14401_32519# C9_N_btm 5.77e-20
C32274 a_17538_32519# C7_N_btm 8.17e-19
C32275 a_12465_44636# a_20916_46384# 3.77e-19
C32276 a_11453_44696# a_19321_45002# 0.023175f
C32277 a_4883_46098# a_22612_30879# 9.37e-21
C32278 a_21811_47423# a_21588_30879# 8.73e-19
C32279 a_n1435_47204# a_1799_45572# 3.59e-20
C32280 a_4915_47217# a_3877_44458# 8.8e-20
C32281 a_n971_45724# a_8492_46660# 0.016456f
C32282 a_n1151_42308# a_5732_46660# 9.82e-22
C32283 a_4700_47436# a_4955_46873# 0.001297f
C32284 a_n443_46116# a_4646_46812# 0.077958f
C32285 a_4791_45118# a_4651_46660# 0.020454f
C32286 a_n237_47217# a_7927_46660# 0.008694f
C32287 a_7989_47542# a_8128_46384# 5.76e-19
C32288 a_n881_46662# a_9804_47204# 0.061323f
C32289 a_n2433_44484# a_n1441_43940# 4.71e-20
C32290 a_5343_44458# a_5013_44260# 1.37e-19
C32291 a_9313_44734# a_20159_44458# 1.77e-20
C32292 a_5518_44484# a_5244_44056# 2.08e-19
C32293 a_4223_44672# a_6453_43914# 0.019918f
C32294 a_13857_44734# a_14673_44172# 2.8e-20
C32295 a_11827_44484# a_10949_43914# 5.25e-20
C32296 a_15861_45028# a_17324_43396# 1.36e-19
C32297 a_3065_45002# a_4093_43548# 0.003025f
C32298 a_2382_45260# a_4699_43561# 6.05e-21
C32299 en_comp a_3626_43646# 5.78e-20
C32300 a_2437_43646# a_2813_43396# 0.012852f
C32301 a_3357_43084# a_6452_43396# 5.12e-19
C32302 a_3232_43370# VDD 2.96597f
C32303 COMP_P a_22609_37990# 0.010152f
C32304 a_18114_32519# a_20820_30879# 0.053f
C32305 a_20205_45028# a_12741_44636# 0.001258f
C32306 a_14539_43914# a_13059_46348# 0.05997f
C32307 a_453_43940# a_n2438_43548# 0.001215f
C32308 a_2998_44172# a_n2293_46634# 0.06774f
C32309 a_n2661_43922# a_8270_45546# 0.025118f
C32310 a_3820_44260# a_768_44030# 3.84e-19
C32311 a_n2017_45002# a_13259_45724# 0.065062f
C32312 a_2437_43646# a_20205_31679# 3.32e-19
C32313 a_3357_43084# a_20850_46482# 7.81e-19
C32314 a_14021_43940# a_10227_46804# 0.062062f
C32315 a_n97_42460# a_n746_45260# 2.64e-19
C32316 a_1049_43396# a_n2497_47436# 3.45e-20
C32317 a_104_43370# a_n971_45724# 0.156156f
C32318 a_14456_42282# a_14113_42308# 0.038993f
C32319 a_n1630_35242# a_n2946_39866# 6.3e-21
C32320 COMP_P a_1343_38525# 0.004705f
C32321 a_n3674_38680# a_n4064_39072# 0.020036f
C32322 a_n4318_38216# a_n3420_39072# 0.032825f
C32323 a_n1605_47204# VDD 0.20224f
C32324 a_7927_46660# a_8270_45546# 8.4e-21
C32325 a_n743_46660# a_765_45546# 0.148721f
C32326 a_7577_46660# a_8601_46660# 2.36e-20
C32327 a_13661_43548# a_19636_46660# 3.05e-20
C32328 a_n881_46662# a_n901_46420# 0.053662f
C32329 a_n1613_43370# a_n1076_46494# 0.232314f
C32330 a_2747_46873# a_2698_46116# 0.006795f
C32331 a_4883_46098# a_7920_46348# 0.006584f
C32332 a_11599_46634# a_15015_46420# 0.040858f
C32333 a_10227_46804# a_11133_46155# 0.019137f
C32334 a_14955_47212# a_14840_46494# 7.46e-21
C32335 a_12861_44030# a_17583_46090# 2.84e-20
C32336 a_6851_47204# a_6945_45028# 0.013916f
C32337 a_1239_47204# a_1337_46116# 6.31e-21
C32338 a_2063_45854# a_n1925_42282# 0.025501f
C32339 a_n1151_42308# a_n914_46116# 2.87e-19
C32340 a_8375_44464# a_8147_43396# 3.2e-20
C32341 a_8333_44056# a_9028_43914# 0.007993f
C32342 a_5891_43370# a_7112_43396# 5.95e-19
C32343 a_14539_43914# a_15095_43370# 4.59e-20
C32344 a_20193_45348# a_4190_30871# 0.02125f
C32345 a_1307_43914# a_15567_42826# 2.68e-20
C32346 a_n2293_42834# a_3935_42891# 0.008823f
C32347 a_18494_42460# a_5649_42852# 1.97e-19
C32348 a_10193_42453# a_11633_42558# 0.017236f
C32349 a_2711_45572# a_17303_42282# 3.67e-19
C32350 a_18579_44172# a_18797_44260# 4.08e-20
C32351 a_17517_44484# a_n97_42460# 7.31e-22
C32352 a_3537_45260# a_4743_43172# 0.002397f
C32353 a_n4209_38216# VCM 0.035453f
C32354 a_n3565_38216# VREF 0.057702f
C32355 a_2711_45572# a_6905_45572# 6.06e-19
C32356 a_15682_43940# a_12741_44636# 0.003137f
C32357 a_18783_43370# a_13661_43548# 0.057336f
C32358 a_15037_43940# a_15227_44166# 0.010516f
C32359 a_15681_43442# a_n2293_46634# 1.89e-19
C32360 a_14021_43940# a_17339_46660# 0.037923f
C32361 a_3539_42460# a_5257_43370# 5.78e-20
C32362 a_10334_44484# a_n443_42852# 1.29e-20
C32363 a_18287_44626# a_n357_42282# 1.16e-21
C32364 a_n1853_43023# a_n2312_40392# 2.89e-21
C32365 a_3905_42865# a_5937_45572# 6.25e-21
C32366 a_19479_31679# EN_OFFSET_CAL 3.97e-20
C32367 a_3357_43084# DATA[5] 0.032568f
C32368 a_5934_30871# VDAC_Pi 1.75e-19
C32369 a_n784_42308# VDAC_P 0.005848f
C32370 a_19692_46634# a_10809_44734# 0.014397f
C32371 a_765_45546# a_11189_46129# 2.79e-21
C32372 a_13059_46348# a_14493_46090# 0.029059f
C32373 a_2443_46660# a_n863_45724# 5.17e-22
C32374 a_10623_46897# a_10586_45546# 5.93e-19
C32375 a_n743_46660# a_509_45822# 0.039863f
C32376 a_8035_47026# a_8034_45724# 1.67e-20
C32377 a_n1991_46122# a_n1423_46090# 0.175891f
C32378 a_n2157_46122# a_n901_46420# 0.043559f
C32379 a_n2293_46098# a_n1076_46494# 0.006462f
C32380 a_n1853_46287# a_n1641_46494# 0.033696f
C32381 a_9313_44734# a_11301_43218# 2.3e-19
C32382 a_19615_44636# a_19339_43156# 1.43e-21
C32383 a_2127_44172# a_1847_42826# 8.79e-22
C32384 a_1414_42308# a_2905_42968# 0.00136f
C32385 a_19478_44306# a_15743_43084# 7.05e-21
C32386 a_15493_43396# a_19268_43646# 0.024436f
C32387 a_15493_43940# a_16547_43609# 0.002713f
C32388 a_11341_43940# a_16977_43638# 6.41e-21
C32389 a_19328_44172# a_19700_43370# 1.6e-19
C32390 a_11967_42832# a_19164_43230# 1.58e-20
C32391 a_n2129_43609# a_n1243_43396# 9.68e-19
C32392 a_n97_42460# a_1891_43646# 0.001075f
C32393 a_1049_43396# a_1568_43370# 2.09e-20
C32394 a_n2956_37592# a_n4209_38502# 0.090878f
C32395 en_comp a_2112_39137# 1.51e-20
C32396 a_4905_42826# VDD 0.439034f
C32397 a_15037_45618# a_9482_43914# 2.11e-19
C32398 a_2711_45572# a_19778_44110# 0.003443f
C32399 a_2437_43646# a_19479_31679# 0.004873f
C32400 a_21513_45002# a_3357_43084# 0.04265f
C32401 a_18783_43370# a_4185_45028# 1.92e-21
C32402 a_13887_32519# a_20820_30879# 0.053104f
C32403 a_13678_32519# a_21076_30879# 0.05537f
C32404 a_15279_43071# a_15227_44166# 0.002075f
C32405 a_18083_42858# a_3090_45724# 9.89e-21
C32406 a_n1736_42282# a_n2312_38680# 2.73e-20
C32407 a_n1329_42308# a_n2442_46660# 3.57e-20
C32408 a_648_43396# a_526_44458# 0.04105f
C32409 a_15764_42576# a_10227_46804# 0.024352f
C32410 a_7174_31319# a_4791_45118# 9.47e-21
C32411 a_13904_45546# a_13487_47204# 3e-19
C32412 a_13249_42308# a_12861_44030# 4.25e-19
C32413 a_10180_45724# a_10227_46804# 0.03118f
C32414 a_12791_45546# a_11599_46634# 5.33e-20
C32415 a_22959_46124# a_20205_31679# 0.012679f
C32416 a_2324_44458# a_n755_45592# 1.99e-20
C32417 a_10809_44734# a_20692_30879# 0.006707f
C32418 a_9290_44172# a_n443_42852# 0.483812f
C32419 a_6945_45028# a_21167_46155# 7.16e-19
C32420 a_21259_43561# a_743_42282# 2.87e-19
C32421 a_9145_43396# a_10083_42826# 6.91e-20
C32422 a_4190_30871# a_20301_43646# 0.00107f
C32423 a_8685_43396# a_10341_42308# 3.51e-19
C32424 a_18114_32519# C8_N_btm 4.06e-19
C32425 a_19721_31679# C7_N_btm 1.43e-20
C32426 a_1307_43914# a_16886_45144# 9.14e-21
C32427 a_8704_45028# a_n2661_43370# 3.79e-19
C32428 a_6171_45002# a_4223_44672# 1.27e-20
C32429 a_5111_44636# a_5518_44484# 0.124556f
C32430 a_4927_45028# a_5343_44458# 1.54e-19
C32431 a_3537_45260# a_5883_43914# 0.018824f
C32432 a_3232_43370# a_n699_43396# 0.074855f
C32433 a_n2017_45002# a_18989_43940# 1.19e-20
C32434 a_2903_42308# a_1823_45246# 0.002746f
C32435 a_5932_42308# a_n2293_46098# 1.61e-20
C32436 a_791_42968# a_n443_42852# 0.04806f
C32437 a_9127_43156# a_n357_42282# 0.021342f
C32438 a_19164_43230# a_13259_45724# 4.12e-20
C32439 a_8387_43230# a_n755_45592# 0.010497f
C32440 a_14401_32519# RST_Z 0.048069f
C32441 a_11823_42460# a_15227_46910# 9.32e-22
C32442 a_10053_45546# a_765_45546# 1.49e-20
C32443 a_14180_45002# a_768_44030# 0.003277f
C32444 a_14537_43396# a_12549_44172# 0.037266f
C32445 a_2274_45254# a_n2438_43548# 1.51e-21
C32446 a_413_45260# a_33_46660# 4.39e-19
C32447 a_3065_45002# a_n1925_46634# 1.56e-20
C32448 a_4574_45260# a_n2293_46634# 1.72e-21
C32449 a_1423_45028# a_n1613_43370# 0.023846f
C32450 a_13711_45394# a_10227_46804# 2.22e-20
C32451 a_n923_35174# VDD 0.340432f
C32452 a_742_44458# a_n746_45260# 0.0971f
C32453 a_n2661_44458# a_584_46384# 0.031143f
C32454 a_n1076_43230# a_n1630_35242# 2.32e-20
C32455 a_15279_43071# a_14635_42282# 2.87e-19
C32456 a_n1533_42852# COMP_P 0.001038f
C32457 a_743_42282# a_4921_42308# 0.015669f
C32458 a_4361_42308# a_5379_42460# 0.045451f
C32459 a_12545_42858# a_13622_42852# 1.46e-19
C32460 a_5342_30871# a_13291_42460# 0.031084f
C32461 a_n3674_39304# a_n3674_37592# 0.024803f
C32462 a_n4064_39072# VDD 1.74897f
C32463 a_4915_47217# a_8128_46384# 0.070866f
C32464 a_6545_47178# a_n881_46662# 0.020203f
C32465 a_6491_46660# a_n1613_43370# 0.071408f
C32466 a_n1435_47204# a_2747_46873# 1.47e-19
C32467 a_n2497_47436# a_n2293_46634# 0.174929f
C32468 SMPL_ON_P a_n2840_46634# 8.18e-19
C32469 a_n2288_47178# a_n2442_46660# 0.009097f
C32470 a_n1920_47178# a_n2661_46634# 1.7e-19
C32471 a_n1741_47186# a_n2956_39768# 1.86e-19
C32472 a_16023_47582# a_12465_44636# 4.1e-19
C32473 a_10227_46804# a_13507_46334# 0.120657f
C32474 a_18479_47436# a_20990_47178# 0.003332f
C32475 a_16588_47582# a_4883_46098# 6.92e-21
C32476 a_18597_46090# a_19787_47423# 0.001396f
C32477 a_11827_44484# a_3422_30871# 0.076229f
C32478 a_n2661_43370# a_2675_43914# 6.77e-21
C32479 a_1307_43914# a_10405_44172# 0.010378f
C32480 a_11823_42460# a_14205_43396# 0.176571f
C32481 a_18184_42460# a_20512_43084# 0.00468f
C32482 a_10193_42453# a_12281_43396# 0.006314f
C32483 a_13076_44458# a_13213_44734# 0.126609f
C32484 a_12883_44458# a_13468_44734# 2.6e-19
C32485 a_12607_44458# a_13857_44734# 0.002706f
C32486 a_6171_45002# a_15493_43940# 5.86e-20
C32487 a_17124_42282# a_n357_42282# 0.011823f
C32488 a_15051_42282# a_n443_42852# 9.06e-21
C32489 a_21973_42336# a_13259_45724# 5.32e-20
C32490 a_18341_45572# VDD 0.2432f
C32491 a_18817_42826# RST_Z 4.49e-21
C32492 a_10951_45334# a_3483_46348# 0.027449f
C32493 a_1423_45028# a_n2293_46098# 0.017396f
C32494 a_14309_45028# a_13059_46348# 0.050896f
C32495 a_15433_44458# a_n743_46660# 1.16e-21
C32496 a_20835_44721# a_12549_44172# 0.002438f
C32497 a_16335_44484# a_13661_43548# 0.002382f
C32498 a_19113_45348# a_19466_46812# 6.36e-19
C32499 a_20193_45348# a_15227_44166# 1.63e-20
C32500 a_15297_45822# a_13259_45724# 1.06e-19
C32501 a_3357_43084# a_10809_44734# 0.035293f
C32502 a_n1059_45260# a_17715_44484# 2.97e-20
C32503 a_5111_44636# a_8199_44636# 0.024227f
C32504 a_5147_45002# a_5937_45572# 8.8e-19
C32505 a_5205_44484# a_5497_46414# 6.8e-22
C32506 a_6171_45002# a_6419_46155# 1.62e-19
C32507 a_413_45260# a_12005_46116# 5.61e-21
C32508 a_4921_42308# a_5755_42308# 0.175841f
C32509 a_2903_42308# a_5934_30871# 2.52e-20
C32510 a_3823_42558# a_6123_31319# 1.19e-20
C32511 a_5379_42460# a_6761_42308# 1.12e-19
C32512 a_1606_42308# a_9223_42460# 1.69e-20
C32513 a_17364_32525# C4_N_btm 1.7e-20
C32514 a_14209_32519# C6_N_btm 0.001467f
C32515 a_3080_42308# VDAC_P 0.009713f
C32516 a_22609_37990# a_22705_37990# 0.087835f
C32517 a_11453_44696# a_13059_46348# 0.039573f
C32518 a_13507_46334# a_17339_46660# 0.05814f
C32519 a_18479_47436# a_20273_46660# 0.018124f
C32520 a_18597_46090# a_20107_46660# 0.001674f
C32521 a_10227_46804# a_20623_46660# 0.156341f
C32522 a_3160_47472# a_1823_45246# 0.002764f
C32523 a_2063_45854# a_2698_46116# 0.006352f
C32524 a_n443_46116# a_n901_46420# 0.367344f
C32525 a_n1151_42308# a_1138_42852# 1.84e-20
C32526 a_2553_47502# a_2521_46116# 7.08e-19
C32527 a_584_46384# a_2804_46116# 1.93e-19
C32528 a_n237_47217# a_5164_46348# 0.081549f
C32529 a_n2109_47186# a_5937_45572# 0.00225f
C32530 a_5807_45002# a_11186_47026# 0.003092f
C32531 a_2443_46660# a_5072_46660# 1.72e-21
C32532 a_2107_46812# a_7577_46660# 1.05e-19
C32533 a_n743_46660# a_10623_46897# 7.67e-20
C32534 a_12549_44172# a_3090_45724# 0.082348f
C32535 a_949_44458# a_1427_43646# 2.11e-19
C32536 a_2675_43914# a_2998_44172# 0.173844f
C32537 a_11967_42832# a_18079_43940# 0.052453f
C32538 a_14815_43914# a_14021_43940# 6.02e-20
C32539 a_4743_44484# a_3080_42308# 5.3e-21
C32540 a_n1899_43946# a_n1453_44318# 2.28e-19
C32541 a_n2065_43946# a_n875_44318# 2.56e-19
C32542 a_n2661_42834# a_1443_43940# 0.001546f
C32543 a_14673_44172# a_15493_43940# 4.52e-20
C32544 a_2479_44172# a_3905_42865# 1.7e-19
C32545 a_742_44458# a_1891_43646# 8.56e-19
C32546 a_5891_43370# a_9801_43940# 8.91e-19
C32547 a_n1549_44318# a_n3674_39768# 1.64e-19
C32548 a_n1059_45260# a_10083_42826# 0.006796f
C32549 a_n913_45002# a_8952_43230# 0.04786f
C32550 a_n2017_45002# a_10518_42984# 4.7e-20
C32551 a_2382_45260# a_1847_42826# 8.82e-20
C32552 a_8975_43940# VDD 0.257588f
C32553 a_n4064_40160# C7_P_btm 2.94e-19
C32554 a_12429_44172# a_3090_45724# 1.23e-21
C32555 a_6765_43638# a_768_44030# 1.04e-20
C32556 a_3626_43646# a_13661_43548# 2.98e-20
C32557 a_1568_43370# a_n2293_46634# 2.04e-19
C32558 a_n2661_43370# a_2277_45546# 5.63e-21
C32559 a_13105_45348# a_n443_42852# 1.05e-20
C32560 a_13943_43396# a_10227_46804# 2.15e-20
C32561 a_16977_43638# a_16327_47482# 0.15941f
C32562 a_19700_43370# a_12861_44030# 1.67e-20
C32563 a_n1076_43230# a_n971_45724# 0.003103f
C32564 a_n1533_42852# a_n2497_47436# 2.22e-19
C32565 a_n2302_39866# a_n2302_39072# 0.052227f
C32566 a_n4315_30879# a_n3420_38528# 0.034192f
C32567 a_n4064_40160# a_n3565_38502# 0.028121f
C32568 a_n133_46660# VDD 0.483405f
C32569 a_5934_30871# C9_N_btm 1.37e-19
C32570 a_11735_46660# a_3483_46348# 6.06e-21
C32571 a_19123_46287# a_20107_46660# 4.05e-20
C32572 a_18285_46348# a_20411_46873# 3.41e-21
C32573 a_2107_46812# a_5431_46482# 8.38e-19
C32574 a_n743_46660# a_6347_46155# 1.92e-19
C32575 a_10249_46116# a_10355_46116# 0.182836f
C32576 a_10467_46802# a_11133_46155# 0.001412f
C32577 a_10554_47026# a_9290_44172# 0.003141f
C32578 a_4651_46660# a_6945_45028# 2.58e-21
C32579 a_18989_43940# a_19164_43230# 1.22e-19
C32580 a_18579_44172# a_20556_43646# 2.61e-19
C32581 a_n2293_43922# a_5111_42852# 9.71e-21
C32582 a_9313_44734# a_10796_42968# 0.009402f
C32583 a_1307_43914# a_6171_42473# 5.75e-21
C32584 a_742_44458# a_4149_42891# 2.67e-20
C32585 a_n2293_42834# a_n3674_37592# 0.025586f
C32586 a_16922_45042# a_20256_43172# 0.001682f
C32587 a_2711_45572# a_9482_43914# 0.01017f
C32588 a_8696_44636# a_16789_45572# 3.81e-20
C32589 a_8162_45546# a_3537_45260# 2.11e-19
C32590 a_13249_42308# a_n913_45002# 0.019571f
C32591 a_7227_45028# a_7705_45326# 1.68e-19
C32592 a_5932_42308# a_4791_45118# 0.212275f
C32593 a_3626_43646# a_4185_45028# 0.035503f
C32594 a_19177_43646# a_19692_46634# 8.77e-21
C32595 a_15682_43940# a_16375_45002# 5.84e-19
C32596 a_3905_42865# a_n443_42852# 0.043488f
C32597 a_1525_44260# a_n863_45724# 2.55e-19
C32598 a_18079_43940# a_13259_45724# 0.007888f
C32599 a_22469_40625# a_22717_37285# 0.002464f
C32600 a_22521_40599# a_22717_36887# 1.4e-19
C32601 a_n3420_37440# C5_P_btm 1.87e-19
C32602 a_n4064_37440# C7_P_btm 1.83e-20
C32603 a_11387_46155# VDD 0.099732f
C32604 a_5263_45724# a_2063_45854# 0.030969f
C32605 a_2711_45572# a_2905_45572# 0.041827f
C32606 a_n3565_38502# a_n4064_37440# 0.028296f
C32607 a_n4064_38528# a_n3565_37414# 0.029213f
C32608 a_n3420_38528# a_n3420_37440# 0.051118f
C32609 a_9823_46155# a_8049_45260# 0.004922f
C32610 a_n2840_46090# a_n2840_45546# 0.025171f
C32611 a_10807_43548# a_11136_42852# 0.006177f
C32612 a_7287_43370# a_4361_42308# 2.93e-20
C32613 a_10341_43396# a_16977_43638# 0.008076f
C32614 a_6197_43396# a_5649_42852# 4.06e-21
C32615 a_458_43396# a_685_42968# 5.82e-20
C32616 a_n1557_42282# a_n13_43084# 0.006682f
C32617 a_n97_42460# a_5111_42852# 5.6e-19
C32618 a_644_44056# a_564_42282# 9.77e-22
C32619 a_9313_44734# a_4958_30871# 5.59e-19
C32620 a_1414_42308# a_n784_42308# 0.017857f
C32621 a_8685_43396# a_15940_43402# 3.06e-19
C32622 a_9804_47204# DATA[4] 0.015379f
C32623 a_2905_42968# VDD 0.142081f
C32624 a_11652_45724# a_n2661_43922# 3.34e-21
C32625 a_8696_44636# a_14539_43914# 0.005592f
C32626 a_15861_45028# a_16112_44458# 2.52e-20
C32627 a_375_42282# a_501_45348# 0.009374f
C32628 a_11962_45724# a_n2661_42834# 3.66e-22
C32629 a_3429_45260# a_n2661_43370# 0.004377f
C32630 a_7229_43940# a_5837_45028# 5.34e-21
C32631 a_6171_45002# a_n2293_42834# 0.035829f
C32632 a_2437_43646# a_20193_45348# 2.74e-21
C32633 a_7227_42308# a_3090_45724# 4.26e-20
C32634 a_n3420_39072# a_n2956_39768# 8.07e-19
C32635 a_19268_43646# a_n357_42282# 1.71e-20
C32636 a_10518_42984# a_526_44458# 1.06e-19
C32637 a_1423_45028# a_4791_45118# 0.721318f
C32638 a_2711_45572# a_12816_46660# 2.6e-20
C32639 a_10193_42453# a_10428_46928# 3.41e-20
C32640 a_8696_44636# a_2107_46812# 0.025973f
C32641 a_8746_45002# a_10150_46912# 1.91e-19
C32642 a_413_45260# a_21811_47423# 8.86e-20
C32643 a_n2956_37592# a_n2312_39304# 0.047801f
C32644 en_comp a_n2312_40392# 0.036842f
C32645 a_3357_43084# a_n881_46662# 0.028875f
C32646 a_509_45822# a_509_45572# 6.96e-20
C32647 a_n443_42852# a_n89_45572# 5.42e-19
C32648 a_14543_43071# a_15279_43071# 4.07e-20
C32649 a_3626_43646# a_9803_42558# 0.006512f
C32650 a_12281_43396# a_n784_42308# 2.26e-20
C32651 a_743_42282# a_13291_42460# 0.068071f
C32652 a_15743_43084# a_20256_43172# 0.006046f
C32653 a_n97_42460# a_9885_42308# 0.003237f
C32654 a_1847_42826# a_1709_42852# 7.79e-21
C32655 a_6765_43638# a_6123_31319# 1.83e-19
C32656 a_17730_32519# C6_N_btm 1.1e-19
C32657 a_19237_31679# C4_N_btm 9.91e-21
C32658 a_15803_42450# VDD 0.448709f
C32659 a_5129_47502# a_5815_47464# 4.88e-20
C32660 a_4915_47217# a_6151_47436# 0.783303f
C32661 a_n1741_47186# a_10227_46804# 0.020904f
C32662 a_2063_45854# a_n1435_47204# 0.001106f
C32663 a_4791_45118# a_6491_46660# 0.002326f
C32664 a_n443_46116# a_6545_47178# 0.001077f
C32665 a_8701_44490# a_5883_43914# 1.13e-20
C32666 a_3065_45002# a_3600_43914# 0.011102f
C32667 a_n2661_45010# a_2537_44260# 6.6e-20
C32668 a_1755_42282# a_n357_42282# 2.68e-19
C32669 a_1606_42308# a_n755_45592# 0.104938f
C32670 a_2725_42558# a_n863_45724# 0.003172f
C32671 a_10193_42453# VDD 2.18892f
C32672 a_22223_43396# RST_Z 5.55e-20
C32673 a_5343_44458# a_n743_46660# 5.3e-23
C32674 a_5883_43914# a_n2293_46634# 0.00136f
C32675 a_17767_44458# a_13661_43548# 5.86e-21
C32676 a_n2017_45002# a_20202_43084# 0.005245f
C32677 a_8568_45546# a_8049_45260# 0.003997f
C32678 a_413_45260# a_22000_46634# 4.39e-20
C32679 a_15765_45572# a_15682_46116# 0.015911f
C32680 a_15599_45572# a_17715_44484# 1.85e-19
C32681 a_12649_45572# a_10903_43370# 0.006357f
C32682 a_6109_44484# a_n1613_43370# 0.099934f
C32683 a_11649_44734# a_11453_44696# 3.12e-19
C32684 a_13213_44734# a_12465_44636# 1.97e-20
C32685 a_n984_44318# a_n746_45260# 4.22e-20
C32686 a_2675_43914# a_n2497_47436# 6.16e-20
C32687 a_17333_42852# a_18057_42282# 3.02e-19
C32688 a_18817_42826# a_17303_42282# 2.65e-20
C32689 a_n1736_42282# COMP_P 0.005447f
C32690 a_18083_42858# a_18727_42674# 3.76e-20
C32691 a_n4318_38680# a_n4064_39072# 0.050323f
C32692 a_n3674_38216# a_n1329_42308# 2.22e-19
C32693 a_n2661_46634# a_n1021_46688# 0.009022f
C32694 a_n2472_46634# a_n1925_46634# 0.001266f
C32695 a_n2293_46634# a_n2104_46634# 0.042499f
C32696 a_n2442_46660# a_n2312_38680# 0.068683f
C32697 a_n2840_46634# a_n2438_43548# 0.002664f
C32698 a_n881_46662# a_3877_44458# 0.142507f
C32699 a_n1613_43370# a_4646_46812# 1.38979f
C32700 a_4883_46098# a_10150_46912# 0.001971f
C32701 a_n1151_42308# a_12978_47026# 1.07e-19
C32702 a_10951_45334# a_10695_43548# 1.93e-21
C32703 a_8696_44636# a_7871_42858# 3.01e-21
C32704 a_18248_44752# a_15493_43396# 1.52e-20
C32705 a_18443_44721# a_18451_43940# 5.21e-19
C32706 a_18287_44626# a_19328_44172# 0.011011f
C32707 a_19279_43940# a_22315_44484# 1.97e-20
C32708 a_11967_42832# a_17730_32519# 9.29e-22
C32709 a_1307_43914# a_3457_43396# 0.005402f
C32710 a_18374_44850# a_18326_43940# 9.6e-19
C32711 a_1423_45028# a_8791_43396# 1.85e-20
C32712 a_18184_42460# a_21381_43940# 0.003589f
C32713 a_20640_44752# a_21145_44484# 2.28e-19
C32714 a_n2661_42834# a_n4318_39768# 0.031793f
C32715 a_11827_44484# a_19808_44306# 2.85e-19
C32716 a_n913_45002# a_19700_43370# 4.09e-21
C32717 a_n1059_45260# a_16664_43396# 9.44e-22
C32718 a_5934_30871# RST_Z 0.003901f
C32719 a_5742_30871# EN_VIN_BSTR_P 0.645417f
C32720 a_3457_43396# a_n443_46116# 3.38e-20
C32721 a_18248_44752# a_3483_46348# 2.73e-21
C32722 a_6109_44484# a_n2293_46098# 2.32e-19
C32723 a_18579_44172# a_19692_46634# 3.19e-19
C32724 a_7584_44260# a_4646_46812# 5.27e-19
C32725 a_n2661_43370# a_8049_45260# 0.013528f
C32726 a_10057_43914# a_8016_46348# 0.09388f
C32727 a_10334_44484# a_8199_44636# 6.58e-19
C32728 a_9838_44484# a_8953_45546# 9.26e-20
C32729 a_5147_45002# a_n443_42852# 0.004185f
C32730 a_19511_42282# a_13258_32519# 0.072135f
C32731 a_6123_31319# a_1177_38525# 1.36e-19
C32732 a_17303_42282# a_21421_42336# 1.17e-19
C32733 a_21496_47436# VDD 0.198362f
C32734 a_4883_46098# a_8062_46482# 6.26e-20
C32735 a_10227_46804# a_10586_45546# 0.306536f
C32736 a_13381_47204# a_13259_45724# 4.87e-21
C32737 a_n2497_47436# a_2277_45546# 8.01e-22
C32738 a_n971_45724# a_n356_45724# 0.030873f
C32739 a_n237_47217# a_3316_45546# 1.38e-19
C32740 a_584_46384# a_n1099_45572# 0.021537f
C32741 a_1239_47204# a_n755_45592# 4.63e-21
C32742 a_3785_47178# a_n2661_45546# 8.89e-21
C32743 a_n1151_42308# a_n2956_38216# 4.1e-20
C32744 a_n881_46662# a_n1736_46482# 1.29e-19
C32745 a_13747_46662# a_14275_46494# 0.002369f
C32746 a_13661_43548# a_15015_46420# 0.001123f
C32747 a_n743_46660# a_8349_46414# 0.004029f
C32748 a_5807_45002# a_14840_46494# 8.3e-21
C32749 a_n2661_46634# a_9290_44172# 2.69e-19
C32750 a_2107_46812# a_4704_46090# 0.008508f
C32751 a_n1925_46634# a_5937_45572# 6.05e-20
C32752 a_n1613_43370# a_n1545_46494# 1.79e-19
C32753 a_2747_46873# a_526_44458# 5.38e-20
C32754 a_17609_46634# a_19692_46634# 3.12e-20
C32755 a_15227_44166# a_19333_46634# 0.065741f
C32756 a_2609_46660# a_1823_45246# 3.24e-19
C32757 a_4646_46812# a_n2293_46098# 1.72e-21
C32758 a_n2661_46098# a_167_45260# 1.31e-19
C32759 a_644_44056# a_n1557_42282# 5.83e-21
C32760 a_1414_42308# a_3080_42308# 1.53e-19
C32761 a_895_43940# a_1756_43548# 1.47e-19
C32762 a_n699_43396# a_2905_42968# 2.16e-19
C32763 a_18184_42460# a_18249_42858# 0.003882f
C32764 a_18494_42460# a_17333_42852# 0.00528f
C32765 a_10729_43914# a_10651_43940# 0.004213f
C32766 a_10405_44172# a_10867_43940# 0.022925f
C32767 a_n2293_42834# a_8292_43218# 1.73e-19
C32768 a_2479_44172# a_4093_43548# 1.25e-20
C32769 a_n1441_43940# a_n4318_39304# 1.27e-19
C32770 a_n2017_45002# a_n327_42308# 2.31e-19
C32771 a_n913_45002# a_2123_42473# 0.029944f
C32772 a_n1059_45260# a_2351_42308# 0.001198f
C32773 a_5495_43940# VDD 0.173477f
C32774 a_14495_45572# a_15599_45572# 5.49e-21
C32775 a_11823_42460# a_16680_45572# 3.71e-20
C32776 a_12427_45724# a_8696_44636# 4.63e-21
C32777 a_15143_45578# a_15297_45822# 0.008535f
C32778 a_10907_45822# a_10544_45572# 4.32e-19
C32779 a_10490_45724# a_12561_45572# 0.001961f
C32780 a_14401_32519# a_20820_30879# 0.055735f
C32781 a_12379_42858# a_12549_44172# 3.65e-20
C32782 a_n1736_43218# a_n2438_43548# 2.63e-20
C32783 a_15493_43396# a_2324_44458# 4.05e-19
C32784 a_9895_44260# a_9290_44172# 3.38e-19
C32785 a_18326_43940# a_17715_44484# 0.003424f
C32786 a_18079_43940# a_18189_46348# 1.25e-19
C32787 COMP_P w_11334_34010# 0.004781f
C32788 a_n3674_38680# SMPL_ON_P 0.038963f
C32789 a_n1736_42282# a_n2497_47436# 3.98e-19
C32790 a_21363_46634# VDD 0.357368f
C32791 a_n4209_39590# a_n2302_37984# 7.57e-20
C32792 a_n1853_46287# a_n2956_38680# 6.64e-19
C32793 a_n2157_46122# a_n1736_46482# 0.086708f
C32794 a_n1991_46122# a_n2956_39304# 2.14e-20
C32795 a_n2293_46098# a_n1545_46494# 4.26e-19
C32796 a_3090_45724# a_n2661_45546# 0.561435f
C32797 a_20107_46660# a_8049_45260# 5.25e-21
C32798 a_19692_46634# a_19443_46116# 1.33e-19
C32799 a_13885_46660# a_14383_46116# 2.54e-21
C32800 a_13059_46348# a_14180_46482# 0.025233f
C32801 a_15227_44166# a_20062_46116# 1.82e-19
C32802 a_3483_46348# a_2324_44458# 0.668551f
C32803 a_8953_45546# a_9823_46155# 6.18e-19
C32804 a_8199_44636# a_9290_44172# 0.516297f
C32805 a_9625_46129# a_9569_46155# 0.204034f
C32806 a_12429_44172# a_12379_42858# 5.92e-19
C32807 a_3626_43646# a_14579_43548# 1.34e-19
C32808 a_2982_43646# a_14205_43396# 1.37e-20
C32809 a_n97_42460# a_16977_43638# 0.002871f
C32810 a_5891_43370# a_5379_42460# 1.75e-20
C32811 a_n356_44636# a_7227_42308# 2.77e-19
C32812 a_6547_43396# a_6643_43396# 0.013793f
C32813 a_6765_43638# a_6809_43396# 3.69e-19
C32814 a_18494_42460# a_18997_42308# 0.002891f
C32815 a_n2293_43922# a_n1630_35242# 0.019388f
C32816 a_20193_45348# a_19511_42282# 1.04e-19
C32817 a_2998_44172# a_3059_42968# 5.55e-20
C32818 a_6197_43396# a_8685_43396# 6.89e-20
C32819 SMPL_ON_N a_22521_40055# 5.57e-20
C32820 a_6151_47436# DATA[5] 0.19492f
C32821 a_6491_46660# DATA[3] 0.011549f
C32822 a_16137_43396# VDD 0.483673f
C32823 a_7499_43078# a_6298_44484# 1.09e-19
C32824 a_3357_43084# a_1307_43914# 0.197864f
C32825 a_3065_45002# a_4558_45348# 0.001793f
C32826 a_2382_45260# a_5111_44636# 1.01e-20
C32827 a_8037_42858# a_4185_45028# 2.64e-20
C32828 a_19164_43230# a_20202_43084# 1.12e-19
C32829 a_8387_43230# a_3483_46348# 7.21e-22
C32830 a_18727_42674# a_12549_44172# 1.47e-21
C32831 a_14853_42852# a_3090_45724# 4.1e-19
C32832 a_15785_43172# a_15227_44166# 9.28e-19
C32833 a_4093_43548# a_n443_42852# 0.028988f
C32834 a_3539_42460# a_n755_45592# 0.008691f
C32835 a_1512_43396# a_n863_45724# 1.35e-19
C32836 a_n2216_40160# a_n2312_40392# 0.001083f
C32837 a_20512_43084# RST_Z 4.49e-21
C32838 a_13163_45724# a_5807_45002# 7.62e-21
C32839 a_11823_42460# a_13747_46662# 0.521845f
C32840 a_2711_45572# a_2443_46660# 5.4e-21
C32841 a_7227_45028# a_2107_46812# 7.51e-20
C32842 a_9049_44484# a_n2661_46634# 4.26e-20
C32843 a_8696_44636# a_11453_44696# 2.67247f
C32844 a_19431_45546# a_16327_47482# 0.344862f
C32845 a_18175_45572# a_10227_46804# 1.6e-21
C32846 a_18787_45572# a_12861_44030# 1.98e-19
C32847 a_2437_43646# a_5815_47464# 0.00818f
C32848 a_n467_45028# a_n746_45260# 0.054826f
C32849 a_n1059_45260# a_584_46384# 6.25e-20
C32850 a_n2017_45002# a_2063_45854# 1.9e-20
C32851 a_3357_43084# a_n443_46116# 0.006081f
C32852 a_n97_42460# a_n1630_35242# 0.035802f
C32853 a_16823_43084# a_16795_42852# 0.065873f
C32854 a_15743_43084# a_21195_42852# 0.004294f
C32855 a_5649_42852# a_10922_42852# 1.52e-20
C32856 a_4361_42308# a_12089_42308# 0.006552f
C32857 a_743_42282# a_13460_43230# 1.8e-20
C32858 a_15493_43940# a_15959_42545# 1.59e-20
C32859 a_n3674_39768# a_n4334_39616# 0.05081f
C32860 a_4190_30871# a_5534_30871# 0.020828f
C32861 a_2982_43646# a_22400_42852# 3.1e-21
C32862 a_n4318_39768# a_n3565_39590# 9.85e-20
C32863 a_3754_39466# a_3754_38470# 7.8e-20
C32864 VDAC_Pi a_8530_39574# 1.79e-20
C32865 a_n784_42308# VDD 0.597561f
C32866 a_11322_45546# a_11341_43940# 2.88e-20
C32867 a_10907_45822# a_10949_43914# 2.73e-20
C32868 a_n2661_43370# a_8103_44636# 5.82e-21
C32869 a_7499_43078# a_10555_44260# 0.03816f
C32870 a_626_44172# a_700_44734# 1.02e-19
C32871 a_18184_42460# a_19929_45028# 0.001333f
C32872 a_7229_43940# a_n2661_42834# 0.023622f
C32873 a_22775_42308# a_21076_30879# 6.58e-21
C32874 a_9306_43218# a_n357_42282# 1.74e-19
C32875 a_2351_42308# a_n1925_42282# 5.44e-20
C32876 a_17749_42852# a_13259_45724# 0.001312f
C32877 a_5457_43172# a_n443_42852# 2.37e-19
C32878 a_5742_30871# a_10903_43370# 5.9e-20
C32879 a_13070_42354# a_9290_44172# 0.140007f
C32880 a_n2661_43922# a_n746_45260# 0.037244f
C32881 a_n2293_43922# a_n971_45724# 2.81e-19
C32882 a_6109_44484# a_4791_45118# 3.61e-20
C32883 a_484_44484# a_584_46384# 0.001797f
C32884 a_13527_45546# a_3483_46348# 4.96e-19
C32885 a_18175_45572# a_17339_46660# 0.019286f
C32886 a_20567_45036# a_12549_44172# 0.176249f
C32887 a_1307_43914# a_3877_44458# 4.73e-20
C32888 a_n2661_43370# a_n2442_46660# 1.23e-19
C32889 a_13105_45348# a_n2661_46634# 0.009374f
C32890 a_6171_45002# a_9863_46634# 1.59e-22
C32891 a_2437_43646# a_19333_46634# 3.78e-21
C32892 a_8191_45002# a_7411_46660# 2.65e-23
C32893 a_7705_45326# a_7715_46873# 0.001207f
C32894 a_18287_44626# a_12861_44030# 0.029719f
C32895 a_10440_44484# a_10227_46804# 0.025362f
C32896 a_7499_43078# a_5937_45572# 0.033831f
C32897 a_6472_45840# a_2324_44458# 2.1e-19
C32898 a_10180_45724# a_8016_46348# 0.259851f
C32899 a_9049_44484# a_8199_44636# 0.029722f
C32900 a_8568_45546# a_8953_45546# 0.136365f
C32901 a_21259_43561# a_13258_32519# 3.03e-20
C32902 a_9127_43156# a_8685_42308# 2.44e-19
C32903 a_8387_43230# a_8791_42308# 0.001415f
C32904 a_n2293_42282# a_1576_42282# 3.68e-19
C32905 a_5649_42852# a_17531_42308# 5.44e-20
C32906 a_4190_30871# a_19647_42308# 0.001077f
C32907 a_4361_42308# a_18907_42674# 0.010379f
C32908 a_13887_32519# a_4958_30871# 0.030919f
C32909 a_n2661_45546# CLK_DATA 1.81e-19
C32910 a_14401_32519# C8_N_btm 8.3e-20
C32911 a_17538_32519# C6_N_btm 5.51e-20
C32912 a_4883_46098# a_21588_30879# 4.72e-19
C32913 a_21811_47423# a_20916_46384# 0.109084f
C32914 a_10227_46804# a_n743_46660# 0.134234f
C32915 a_n1741_47186# a_10467_46802# 9.36e-19
C32916 a_n971_45724# a_8667_46634# 0.006462f
C32917 a_n237_47217# a_8145_46902# 3.42e-20
C32918 a_4700_47436# a_4651_46660# 4.72e-19
C32919 a_n443_46116# a_3877_44458# 0.06318f
C32920 a_4791_45118# a_4646_46812# 0.485113f
C32921 a_n881_46662# a_8128_46384# 0.206292f
C32922 a_8696_44636# a_17324_43396# 5.68e-21
C32923 a_16922_45042# a_15493_43396# 5.34e-20
C32924 a_5343_44458# a_5244_44056# 8.23e-19
C32925 a_9313_44734# a_19615_44636# 1.67e-21
C32926 a_4223_44672# a_5663_43940# 0.01368f
C32927 a_15861_45028# a_17499_43370# 6.09e-20
C32928 a_n2661_43370# a_11173_44260# 2.7e-19
C32929 a_n1352_44484# a_n4318_39768# 3e-19
C32930 a_2437_43646# a_2437_43396# 0.009374f
C32931 a_2382_45260# a_4235_43370# 0.006145f
C32932 a_n1059_45260# a_n144_43396# 8.85e-20
C32933 a_5205_44484# a_n97_42460# 1.83e-20
C32934 a_5691_45260# VDD 0.205518f
C32935 a_16922_45042# a_3483_46348# 3.56e-19
C32936 a_19721_31679# a_11415_45002# 0.001159f
C32937 a_19929_45028# a_12741_44636# 0.001258f
C32938 a_1414_42308# a_n2438_43548# 0.001019f
C32939 a_n2661_42834# a_8270_45546# 0.034362f
C32940 a_2889_44172# a_n2293_46634# 1.86e-19
C32941 a_3499_42826# a_768_44030# 0.034429f
C32942 a_7229_43940# a_5066_45546# 4.19e-21
C32943 a_n2661_43370# a_8953_45546# 0.02624f
C32944 a_1423_45028# a_6945_45028# 1.15e-19
C32945 a_11341_43940# a_12465_44636# 0.002963f
C32946 a_13829_44260# a_10227_46804# 1.01e-19
C32947 a_n97_42460# a_n971_45724# 0.581616f
C32948 a_1209_43370# a_n2497_47436# 1.74e-20
C32949 SMPL_ON_P VDD 0.614138f
C32950 a_13575_42558# a_14113_42308# 0.11418f
C32951 a_n1630_35242# a_n3420_39616# 0.001297f
C32952 a_n3674_38216# a_n4334_39392# 9.02e-20
C32953 a_n3674_37592# a_n4064_39616# 0.019733f
C32954 a_8145_46902# a_8270_45546# 4.35e-20
C32955 a_8492_46660# a_8654_47026# 0.006453f
C32956 a_7927_46660# a_8189_46660# 0.001705f
C32957 a_n743_46660# a_17339_46660# 2.36e-19
C32958 a_13661_43548# a_18900_46660# 0.003751f
C32959 a_n881_46662# a_n1641_46494# 4.9e-19
C32960 a_n1613_43370# a_n901_46420# 0.406381f
C32961 a_2747_46873# a_2521_46116# 7.97e-20
C32962 a_4883_46098# a_6419_46155# 0.007342f
C32963 a_11599_46634# a_14275_46494# 0.029786f
C32964 a_10227_46804# a_11189_46129# 0.001224f
C32965 a_14955_47212# a_15015_46420# 4.84e-19
C32966 a_13717_47436# a_17583_46090# 1.18e-21
C32967 a_12861_44030# a_15682_46116# 0.030474f
C32968 a_6151_47436# a_10809_44734# 5.72e-19
C32969 a_6491_46660# a_6945_45028# 0.0023f
C32970 a_n1741_47186# a_8034_45724# 3.32e-21
C32971 a_2063_45854# a_526_44458# 0.039908f
C32972 a_n237_47217# a_5066_45546# 1.48406f
C32973 a_584_46384# a_n1925_42282# 0.194054f
C32974 a_15004_44636# a_14955_43396# 6.17e-20
C32975 a_14539_43914# a_14205_43396# 0.001533f
C32976 a_5891_43370# a_7287_43370# 0.008619f
C32977 a_20193_45348# a_21259_43561# 6.39e-21
C32978 a_11827_44484# a_21487_43396# 3.48e-20
C32979 a_19279_43940# a_19319_43548# 0.023499f
C32980 a_n2293_42834# a_3681_42891# 0.006112f
C32981 a_1307_43914# a_5342_30871# 5.9e-20
C32982 a_10193_42453# a_11551_42558# 0.228057f
C32983 a_18184_42460# a_5649_42852# 0.028842f
C32984 a_18579_44172# a_18533_44260# 0.001461f
C32985 a_10057_43914# a_12281_43396# 5.88e-20
C32986 a_2711_45572# a_4958_30871# 1.35e-20
C32987 a_11691_44458# a_4190_30871# 0.002426f
C32988 a_n913_45002# a_8495_42852# 0.030544f
C32989 a_3537_45260# a_4649_43172# 5.06e-19
C32990 a_n4209_38216# VREF_GND 0.001997f
C32991 a_7230_45938# a_8162_45546# 1.68e-19
C32992 a_2711_45572# a_6469_45572# 2.38e-19
C32993 a_18525_43370# a_13661_43548# 0.031188f
C32994 a_3626_43646# a_5257_43370# 5.37e-20
C32995 a_19478_44056# a_3090_45724# 0.002976f
C32996 a_14621_43646# a_n2293_46634# 0.002737f
C32997 a_n356_44636# a_n2661_45546# 3.08e-21
C32998 a_10157_44484# a_n443_42852# 1.48e-20
C32999 a_18248_44752# a_n357_42282# 9.12e-22
C33000 a_n2157_42858# a_n2312_40392# 5.78e-21
C33001 a_2437_43646# CLK 0.101524f
C33002 a_3357_43084# DATA[4] 0.035981f
C33003 a_8035_47026# VDD 0.132317f
C33004 COMP_P a_22469_40625# 0.120018f
C33005 a_19692_46634# a_22223_46124# 0.001994f
C33006 a_765_45546# a_9290_44172# 4.14e-20
C33007 a_13059_46348# a_13925_46122# 0.056739f
C33008 a_14513_46634# a_2324_44458# 1.3e-19
C33009 a_19466_46812# a_10809_44734# 0.007455f
C33010 a_10249_46116# a_10044_46482# 0.00124f
C33011 a_3699_46634# a_n2661_45546# 5.3e-21
C33012 a_10467_46802# a_10586_45546# 5.92e-20
C33013 a_2107_46812# a_2957_45546# 1.23e-20
C33014 a_n2661_46098# a_n863_45724# 4.3e-20
C33015 a_n1925_46634# a_n443_42852# 5.96e-20
C33016 a_8270_45546# a_5066_45546# 0.189476f
C33017 a_n2157_46122# a_n1641_46494# 0.105995f
C33018 a_n2293_46098# a_n901_46420# 0.007523f
C33019 a_n1853_46287# a_n1423_46090# 0.043126f
C33020 a_9313_44734# a_11229_43218# 1.2e-19
C33021 a_18248_44752# a_18707_42852# 7.68e-22
C33022 a_11967_42832# a_19339_43156# 9.23e-20
C33023 a_19328_44172# a_19268_43646# 9.49e-19
C33024 a_15493_43396# a_15743_43084# 0.517624f
C33025 a_104_43370# a_n1557_42282# 6.03e-21
C33026 a_15493_43940# a_16243_43396# 0.006124f
C33027 a_11341_43940# a_16409_43396# 4.02e-20
C33028 a_n2433_43396# a_n1243_43396# 2.56e-19
C33029 a_n97_42460# a_1427_43646# 0.047018f
C33030 a_1209_43370# a_1568_43370# 9.57e-19
C33031 a_n2810_45028# a_n4209_38502# 0.022376f
C33032 a_3080_42308# VDD 0.849483f
C33033 a_2711_45572# a_18911_45144# 3.83e-20
C33034 a_14033_45822# a_9482_43914# 8.97e-21
C33035 a_2437_43646# a_22223_45572# 0.165664f
C33036 a_21513_45002# a_19479_31679# 0.005077f
C33037 a_15743_43084# a_3483_46348# 8.98e-20
C33038 a_22591_43396# a_11415_45002# 1.64e-20
C33039 a_n3674_38680# a_n2438_43548# 8.18e-20
C33040 COMP_P a_n2442_46660# 0.024155f
C33041 a_n3674_38216# a_n2312_38680# 0.023419f
C33042 a_548_43396# a_526_44458# 0.002535f
C33043 a_10849_43646# a_10903_43370# 0.003042f
C33044 a_15486_42560# a_10227_46804# 0.227612f
C33045 a_13904_45546# a_12861_44030# 0.027907f
C33046 a_10053_45546# a_10227_46804# 0.009863f
C33047 a_11823_42460# a_11599_46634# 5.18e-19
C33048 a_10809_44734# a_20205_31679# 0.039075f
C33049 a_2324_44458# a_n357_42282# 1.23e-19
C33050 a_22223_46124# a_20692_30879# 2.55e-19
C33051 a_9145_43396# a_8952_43230# 1.61e-20
C33052 a_9803_43646# a_9127_43156# 3.02e-19
C33053 a_20512_43084# a_17303_42282# 4.29e-20
C33054 a_n2661_42282# a_6481_42558# 0.001754f
C33055 a_4646_46812# DATA[3] 0.001949f
C33056 a_18114_32519# C7_N_btm 2.94e-19
C33057 a_19721_31679# C6_N_btm 1.26e-20
C33058 a_17478_45572# a_17517_44484# 7.16e-22
C33059 a_1307_43914# a_16237_45028# 0.056593f
C33060 a_7735_45067# a_n2661_43370# 2.56e-19
C33061 a_3232_43370# a_4223_44672# 0.033907f
C33062 a_5111_44636# a_5343_44458# 0.477401f
C33063 a_4927_45028# a_4743_44484# 3.54e-19
C33064 a_5147_45002# a_5518_44484# 0.064422f
C33065 a_3537_45260# a_8701_44490# 5.76e-20
C33066 a_n2661_45010# a_n1190_44850# 2.49e-19
C33067 a_2713_42308# a_1823_45246# 2.25e-19
C33068 a_6171_42473# a_n2293_46098# 1.9e-21
C33069 a_685_42968# a_n443_42852# 0.104532f
C33070 a_8387_43230# a_n357_42282# 0.009479f
C33071 a_19339_43156# a_13259_45724# 7.95e-21
C33072 a_8605_42826# a_n755_45592# 0.003535f
C33073 a_21381_43940# RST_Z 3.55e-21
C33074 a_11962_45724# a_13059_46348# 0.001121f
C33075 a_13904_45546# a_14180_46812# 2.21e-22
C33076 a_14495_45572# a_13885_46660# 1.27e-20
C33077 a_13777_45326# a_768_44030# 0.011242f
C33078 a_14537_43396# a_12891_46348# 5.09e-20
C33079 a_9049_44484# a_765_45546# 2.74e-20
C33080 a_n37_45144# a_33_46660# 3.74e-22
C33081 a_327_44734# a_n133_46660# 9.06e-21
C33082 a_8953_45002# a_5807_45002# 7.32e-20
C33083 a_1667_45002# a_n2438_43548# 0.001763f
C33084 a_3537_45260# a_n2293_46634# 0.155982f
C33085 a_n2293_45010# a_n2661_46098# 1.46e-20
C33086 a_5147_45002# a_n2661_46634# 2.08e-20
C33087 a_n2293_42834# a_4883_46098# 2.72e-20
C33088 a_13490_45394# a_10227_46804# 1.9e-20
C33089 a_n1532_35090# VDD 2.19114f
C33090 a_n452_44636# a_n746_45260# 0.042999f
C33091 a_n901_43156# a_n1630_35242# 3e-19
C33092 a_n13_43084# a_n3674_37592# 1.17e-20
C33093 a_5534_30871# a_14635_42282# 0.020227f
C33094 a_4361_42308# a_5267_42460# 0.005989f
C33095 a_n2293_42282# a_4649_42852# 5.38e-20
C33096 a_743_42282# a_4933_42558# 0.001023f
C33097 a_n2946_39072# VDD 0.383374f
C33098 a_6151_47436# a_n881_46662# 1.58776f
C33099 a_4915_47217# a_5159_47243# 7.22e-19
C33100 a_6545_47178# a_n1613_43370# 0.006198f
C33101 a_n1151_42308# a_768_44030# 0.019901f
C33102 a_n2497_47436# a_n2442_46660# 0.045496f
C33103 a_n2288_47178# a_n2472_46634# 3.21e-19
C33104 a_n2109_47186# a_n2661_46634# 0.038259f
C33105 a_n1920_47178# a_n2956_39768# 6.13e-19
C33106 a_16327_47482# a_12465_44636# 6.07e-19
C33107 a_18597_46090# a_19386_47436# 0.007892f
C33108 a_18780_47178# a_19787_47423# 2.54e-20
C33109 a_17591_47464# a_13507_46334# 3.36e-20
C33110 a_16763_47508# a_4883_46098# 8.86e-22
C33111 a_18479_47436# a_20894_47436# 0.032517f
C33112 a_10227_46804# a_21177_47436# 9.07e-19
C33113 a_13777_45326# a_13483_43940# 5.57e-20
C33114 a_13249_42308# a_9145_43396# 0.072489f
C33115 a_13556_45296# a_14955_43940# 0.059957f
C33116 a_n2293_42834# a_5663_43940# 4.43e-21
C33117 a_1307_43914# a_9672_43914# 0.007152f
C33118 a_11823_42460# a_14358_43442# 0.122636f
C33119 a_12883_44458# a_13213_44734# 0.002706f
C33120 a_12607_44458# a_13468_44734# 1.09e-19
C33121 a_11827_44484# a_21398_44850# 0.003647f
C33122 a_11691_44458# a_18753_44484# 0.005052f
C33123 a_13076_44458# a_n2293_43922# 5.37e-19
C33124 a_10193_42453# a_12293_43646# 9.47e-19
C33125 a_19610_45572# a_19319_43548# 1.39e-20
C33126 a_22465_38105# a_13259_45724# 1.69e-19
C33127 a_14113_42308# a_n443_42852# 3.7e-20
C33128 a_18479_45785# VDD 0.536075f
C33129 a_18249_42858# RST_Z 6.28e-21
C33130 a_10775_45002# a_3483_46348# 0.025931f
C33131 a_11691_44458# a_15227_44166# 0.443265f
C33132 a_20679_44626# a_12549_44172# 0.006058f
C33133 a_22223_45036# a_19692_46634# 8.92e-20
C33134 a_9159_44484# a_2107_46812# 5.96e-19
C33135 a_16241_44484# a_13661_43548# 5.03e-19
C33136 a_7499_43078# a_n443_42852# 0.375366f
C33137 a_15225_45822# a_13259_45724# 7.2e-20
C33138 a_413_45260# a_10903_43370# 4.56e-21
C33139 a_n2017_45002# a_17715_44484# 7.39e-21
C33140 a_4558_45348# a_5937_45572# 1.53e-20
C33141 a_5205_44484# a_5204_45822# 2.74e-21
C33142 a_6171_45002# a_6165_46155# 9.99e-20
C33143 a_3357_43084# a_22223_46124# 2.09e-20
C33144 a_2713_42308# a_5934_30871# 1.48e-20
C33145 a_3318_42354# a_6123_31319# 1.13e-20
C33146 a_1606_42308# a_8791_42308# 3.31e-20
C33147 a_n784_42308# a_11551_42558# 2.06e-20
C33148 a_5267_42460# a_6761_42308# 6.68e-20
C33149 a_16877_42852# a_4958_30871# 6.91e-19
C33150 a_14209_32519# C5_N_btm 0.042017f
C33151 a_17364_32525# C3_N_btm 1.38e-20
C33152 a_13887_32519# C7_N_btm 4.26e-20
C33153 CAL_P a_22717_36887# 9.62e-21
C33154 a_22705_38406# a_22705_37990# 0.003483f
C33155 a_22609_38406# a_22717_37285# 0.08753f
C33156 a_13507_46334# a_15312_46660# 5.88e-21
C33157 a_10227_46804# a_20841_46902# 0.164019f
C33158 a_18479_47436# a_20411_46873# 0.192791f
C33159 a_2905_45572# a_1823_45246# 1.3e-19
C33160 a_2063_45854# a_2521_46116# 0.011365f
C33161 a_n1151_42308# a_1176_45822# 1.53e-19
C33162 a_584_46384# a_2698_46116# 1.53e-19
C33163 a_n237_47217# a_5068_46348# 0.033474f
C33164 a_n971_45724# a_5204_45822# 4.32e-20
C33165 a_n1741_47186# a_8016_46348# 3.91e-20
C33166 a_12891_46348# a_3090_45724# 1.19e-21
C33167 a_3524_46660# a_4817_46660# 1.33e-19
C33168 a_2107_46812# a_7715_46873# 0.032178f
C33169 a_768_44030# a_14084_46812# 0.013767f
C33170 a_n743_46660# a_10467_46802# 9.14e-20
C33171 a_12549_44172# a_15009_46634# 0.009008f
C33172 a_949_44458# a_n1557_42282# 1.2e-19
C33173 a_n699_43396# a_3080_42308# 0.001343f
C33174 a_2675_43914# a_2889_44172# 0.083573f
C33175 a_n1899_43946# a_n1644_44306# 0.06121f
C33176 a_17517_44484# a_20935_43940# 1.78e-20
C33177 a_895_43940# a_2998_44172# 2.2e-19
C33178 a_11967_42832# a_17973_43940# 0.070514f
C33179 a_1307_43914# a_743_42282# 5.15e-19
C33180 a_4223_44672# a_4905_42826# 3.85e-20
C33181 a_742_44458# a_1427_43646# 5.41e-19
C33182 a_4743_44484# a_4699_43561# 6.57e-20
C33183 a_n2661_42834# a_1241_43940# 0.003456f
C33184 a_5891_43370# a_9420_43940# 4.11e-19
C33185 a_n1331_43914# a_n3674_39768# 6.83e-20
C33186 a_n1059_45260# a_8952_43230# 0.010945f
C33187 a_n913_45002# a_9127_43156# 0.038139f
C33188 a_n2017_45002# a_10083_42826# 1.71e-19
C33189 a_10057_43914# VDD 0.399284f
C33190 a_n4064_40160# C8_P_btm 4.06e-19
C33191 a_n4064_39616# EN_VIN_BSTR_P 0.072552f
C33192 a_22591_44484# a_11415_45002# 6.11e-19
C33193 a_2982_43646# a_13747_46662# 0.010585f
C33194 a_11750_44172# a_3090_45724# 3.43e-21
C33195 a_3626_43646# a_5807_45002# 2.2e-22
C33196 a_6197_43396# a_768_44030# 4.37e-20
C33197 a_n2661_43370# a_1609_45822# 0.008983f
C33198 a_5883_43914# a_8049_45260# 3.03e-20
C33199 a_16922_45042# a_n357_42282# 9.6e-19
C33200 a_3363_44484# a_2324_44458# 0.004792f
C33201 a_10341_43396# a_12465_44636# 8.52e-20
C33202 a_14205_43396# a_11453_44696# 1.6e-22
C33203 a_13837_43396# a_10227_46804# 1.96e-20
C33204 a_16409_43396# a_16327_47482# 0.022593f
C33205 a_19268_43646# a_12861_44030# 9.01e-21
C33206 a_743_42282# a_n443_46116# 1.1e-19
C33207 a_n901_43156# a_n971_45724# 0.019025f
C33208 a_n4318_38680# SMPL_ON_P 0.039103f
C33209 a_n4064_40160# a_n4334_38528# 0.007725f
C33210 a_n3420_39616# a_n3607_39392# 6.01e-19
C33211 a_n2438_43548# VDD 3.40589f
C33212 a_6123_31319# C10_N_btm 1.34e-19
C33213 a_5934_30871# C8_N_btm 1.41e-19
C33214 a_n743_46660# a_8034_45724# 0.021079f
C33215 a_n2661_46098# a_1431_46436# 2.82e-19
C33216 a_2107_46812# a_5210_46482# 8.98e-19
C33217 a_10623_46897# a_9290_44172# 0.00174f
C33218 a_10249_46116# a_9823_46155# 0.082191f
C33219 a_6755_46942# a_9569_46155# 1.96e-19
C33220 a_10467_46802# a_11189_46129# 0.005012f
C33221 a_10428_46928# a_11133_46155# 6.41e-19
C33222 a_4646_46812# a_6945_45028# 0.090679f
C33223 a_n2293_42834# a_n327_42558# 0.001338f
C33224 a_19478_44306# a_3626_43646# 6.67e-20
C33225 a_18579_44172# a_743_42282# 9.34e-19
C33226 a_n2293_43922# a_4520_42826# 1.13e-20
C33227 a_n2661_43922# a_5111_42852# 3.12e-21
C33228 a_n2661_42834# a_5755_42852# 1.12e-20
C33229 a_9313_44734# a_10835_43094# 0.050385f
C33230 a_3422_30871# a_16823_43084# 4.23e-21
C33231 a_n356_44636# a_17701_42308# 0.065679f
C33232 a_1307_43914# a_5755_42308# 1.01e-20
C33233 a_742_44458# a_3863_42891# 4.92e-20
C33234 a_n2661_43370# a_n3674_38216# 1.63e-20
C33235 a_n913_45002# a_17124_42282# 4.89e-19
C33236 a_3232_43370# a_5742_30871# 6.51e-20
C33237 a_14021_43940# VDD 1.60583f
C33238 a_2711_45572# a_13348_45260# 7.14e-20
C33239 a_16680_45572# a_16789_45572# 0.007416f
C33240 a_16855_45546# a_17034_45572# 0.007399f
C33241 a_7227_45028# a_6709_45028# 0.115677f
C33242 a_4880_45572# a_5111_44636# 3.99e-20
C33243 a_13249_42308# a_n1059_45260# 0.026496f
C33244 a_11823_42460# en_comp 8.68e-21
C33245 a_6171_42473# a_4791_45118# 5.34e-19
C33246 a_22469_40625# a_22705_37990# 0.010408f
C33247 a_22521_40599# a_22717_37285# 0.010048f
C33248 a_n3420_37440# C6_P_btm 1.87e-19
C33249 a_n4209_37414# C2_P_btm 0.001057f
C33250 a_n3565_37414# C4_P_btm 9.91e-21
C33251 a_8685_43396# a_12741_44636# 5.43e-21
C33252 a_6031_43396# a_1823_45246# 3.31e-19
C33253 a_4361_42308# a_3090_45724# 1.2e-19
C33254 a_4190_30871# a_15227_44166# 2.91e-20
C33255 a_17973_43940# a_13259_45724# 0.025372f
C33256 a_1241_44260# a_n863_45724# 1.7e-19
C33257 a_14097_32519# SMPL_ON_N 0.029158f
C33258 a_8530_39574# RST_Z 0.431385f
C33259 a_11133_46155# VDD 0.176249f
C33260 a_3775_45552# a_n237_47217# 1.02e-19
C33261 a_4099_45572# a_2063_45854# 1.09e-19
C33262 a_3733_45822# a_n971_45724# 3.4e-19
C33263 a_n4209_38502# a_n2302_37690# 4.92e-19
C33264 a_n3565_38502# a_n2946_37690# 4.07e-19
C33265 a_2684_37794# a_3754_38470# 5.6e-20
C33266 a_n4064_38528# a_n4334_37440# 1.78e-19
C33267 a_n3420_39072# VDAC_P 2.6e-19
C33268 a_9569_46155# a_8049_45260# 0.009377f
C33269 a_8016_46348# a_10586_45546# 2.29e-19
C33270 a_n984_44318# a_n1630_35242# 1.73e-21
C33271 a_6547_43396# a_4361_42308# 2.77e-20
C33272 a_9396_43370# a_743_42282# 5.17e-20
C33273 a_10341_43396# a_16409_43396# 0.028466f
C33274 a_n1557_42282# a_n1076_43230# 3.53e-20
C33275 a_n97_42460# a_4520_42826# 4.68e-20
C33276 a_12281_43396# a_13943_43396# 6.37e-21
C33277 a_8685_43396# a_15868_43402# 4.99e-20
C33278 a_6293_42852# a_5649_42852# 2.33e-19
C33279 a_1414_42308# a_196_42282# 6.32e-21
C33280 a_8128_46384# DATA[4] 6.38e-19
C33281 a_2075_43172# VDD 0.001106f
C33282 a_11525_45546# a_n2661_43922# 1.39e-20
C33283 a_16680_45572# a_14539_43914# 2.31e-19
C33284 a_16855_45546# a_16979_44734# 2.49e-21
C33285 a_8696_44636# a_16112_44458# 0.004409f
C33286 a_2711_45572# a_19615_44636# 2.24e-21
C33287 a_1307_43914# a_626_44172# 6.24e-19
C33288 a_3065_45002# a_n2661_43370# 0.356646f
C33289 a_19479_31679# a_22959_45036# 0.018372f
C33290 a_3232_43370# a_n2293_42834# 0.041207f
C33291 a_21513_45002# a_20193_45348# 3.14e-20
C33292 a_6171_45002# a_7639_45394# 3.69e-19
C33293 a_n4209_39304# a_n2442_46660# 2.66e-20
C33294 a_10083_42826# a_526_44458# 0.012145f
C33295 a_15781_43660# a_n443_42852# 0.22553f
C33296 a_15743_43084# a_n357_42282# 0.055032f
C33297 a_626_44172# a_n443_46116# 2.44e-20
C33298 a_10193_42453# a_10150_46912# 1.25e-20
C33299 a_19256_45572# a_19594_46812# 2.98e-19
C33300 a_8746_45002# a_9863_46634# 5.88e-19
C33301 a_10053_45546# a_10467_46802# 1.61e-20
C33302 a_5111_44636# a_10227_46804# 7.06e-20
C33303 a_413_45260# a_4883_46098# 2.47e-19
C33304 a_n2810_45028# a_n2312_39304# 0.043636f
C33305 a_n2956_37592# a_n2312_40392# 0.060336f
C33306 a_3357_43084# a_n1613_43370# 0.228593f
C33307 a_20528_45572# a_12549_44172# 1.17e-19
C33308 a_6547_43396# a_6761_42308# 1.18e-20
C33309 a_6197_43396# a_6123_31319# 1.52e-19
C33310 a_15743_43084# a_18707_42852# 8.78e-20
C33311 a_19319_43548# a_19332_42282# 8.34e-20
C33312 a_14543_43071# a_5534_30871# 0.196814f
C33313 a_13460_43230# a_15279_43071# 2.03e-20
C33314 a_13635_43156# a_5342_30871# 0.001254f
C33315 a_21381_43940# a_17303_42282# 4.27e-20
C33316 a_3626_43646# a_9223_42460# 0.002263f
C33317 a_14401_32519# a_4958_30871# 0.079459f
C33318 a_3935_42891# a_4156_43218# 0.007833f
C33319 a_n97_42460# a_15720_42674# 5.52e-19
C33320 a_472_46348# DATA[0] 3.54e-20
C33321 a_17730_32519# C5_N_btm 8.54e-20
C33322 a_15764_42576# VDD 0.258303f
C33323 a_4915_47217# a_5815_47464# 0.064955f
C33324 a_584_46384# a_n1435_47204# 5e-19
C33325 a_4791_45118# a_6545_47178# 0.112353f
C33326 a_n1151_42308# a_9067_47204# 6.01e-21
C33327 a_n443_46116# a_6151_47436# 1.3e-19
C33328 a_4223_44672# a_8975_43940# 1.67e-19
C33329 a_3065_45002# a_2998_44172# 0.024536f
C33330 a_2382_45260# a_3905_42865# 0.291572f
C33331 a_n2293_45010# a_1241_44260# 1.56e-19
C33332 a_n2661_45010# a_2253_44260# 5.46e-19
C33333 a_3537_45260# a_2675_43914# 2.19e-19
C33334 a_n967_45348# a_n3674_39768# 2.29e-20
C33335 a_1606_42308# a_n357_42282# 0.001349f
C33336 a_3823_42558# a_n2661_45546# 7.7e-21
C33337 a_10180_45724# VDD 0.336512f
C33338 a_5649_42852# RST_Z 6.96e-19
C33339 a_4743_44484# a_n743_46660# 1.08e-21
C33340 a_14539_43914# a_13747_46662# 1.14e-20
C33341 a_16979_44734# a_13661_43548# 5.5e-20
C33342 a_17767_44458# a_5807_45002# 1.7e-21
C33343 a_3357_43084# a_n2293_46098# 0.16657f
C33344 a_8162_45546# a_8049_45260# 0.057007f
C33345 a_413_45260# a_21188_46660# 4.93e-21
C33346 a_15903_45785# a_15682_46116# 0.011633f
C33347 a_15765_45572# a_2324_44458# 0.005634f
C33348 a_8696_44636# a_13925_46122# 7.96e-21
C33349 a_12561_45572# a_10903_43370# 0.002063f
C33350 a_n2293_43922# a_12465_44636# 0.025736f
C33351 a_16241_44734# a_16327_47482# 4.54e-20
C33352 a_n809_44244# a_n746_45260# 1.75e-19
C33353 a_n984_44318# a_n971_45724# 0.003098f
C33354 a_895_43940# a_n2497_47436# 0.0309f
C33355 a_18083_42858# a_18057_42282# 9.91e-19
C33356 a_18249_42858# a_17303_42282# 4.65e-20
C33357 a_n1736_42282# a_n4318_37592# 0.153911f
C33358 a_n3674_39304# a_n4064_39072# 0.539144f
C33359 a_n4318_38216# a_n961_42308# 1.13e-20
C33360 a_n3674_38216# COMP_P 2.04e-19
C33361 a_n2472_46634# a_n2312_38680# 0.039578f
C33362 a_n2661_46634# a_n1925_46634# 4.75867f
C33363 a_n2442_46660# a_n2104_46634# 0.001169f
C33364 a_n1613_43370# a_3877_44458# 1.43013f
C33365 a_5063_47570# a_4955_46873# 3.3e-22
C33366 a_4883_46098# a_9863_46634# 0.007473f
C33367 a_12861_44030# a_11735_46660# 4.6e-21
C33368 a_n1435_47204# a_11901_46660# 7.78e-20
C33369 a_n2109_47186# a_765_45546# 0.126431f
C33370 a_10775_45002# a_10695_43548# 1.22e-21
C33371 a_12883_44458# a_11341_43940# 9.36e-21
C33372 a_13556_45296# a_8685_43396# 6.99e-19
C33373 a_18443_44721# a_18326_43940# 0.007036f
C33374 a_18287_44626# a_18451_43940# 0.005619f
C33375 a_11967_42832# a_22591_44484# 2.53e-20
C33376 a_n2661_43922# a_7542_44172# 5.03e-21
C33377 a_18248_44752# a_19328_44172# 1.49e-20
C33378 a_n2661_42834# a_7845_44172# 0.009718f
C33379 a_18989_43940# a_17973_43940# 8.65e-20
C33380 a_1307_43914# a_2813_43396# 6.65e-19
C33381 a_n2293_42834# a_4905_42826# 0.046599f
C33382 a_1423_45028# a_8147_43396# 2e-21
C33383 a_20159_44458# a_20512_43084# 9.66e-22
C33384 a_18579_44172# a_19789_44512# 0.003679f
C33385 a_20679_44626# a_20637_44484# 2.56e-19
C33386 a_18184_42460# a_19741_43940# 4.62e-19
C33387 a_19279_43940# a_3422_30871# 0.02352f
C33388 a_6109_44484# a_6756_44260# 2.02e-19
C33389 a_11827_44484# a_18797_44260# 5.32e-19
C33390 a_n913_45002# a_19268_43646# 1.96e-21
C33391 a_5742_30871# a_n923_35174# 0.099784f
C33392 a_5934_30871# C2_P_btm 0.011047f
C33393 a_2813_43396# a_n443_46116# 0.124521f
C33394 a_9885_43646# a_n971_45724# 9.07e-21
C33395 a_17970_44736# a_3483_46348# 1.12e-19
C33396 a_18579_44172# a_19466_46812# 0.003312f
C33397 a_14021_43940# a_22612_30879# 1.68e-20
C33398 a_10440_44484# a_8016_46348# 0.001273f
C33399 a_5883_43914# a_8953_45546# 0.262126f
C33400 a_10157_44484# a_8199_44636# 5.53e-20
C33401 a_13507_46334# VDD 1.4135f
C33402 a_19511_42282# a_19647_42308# 0.038787f
C33403 a_19386_47436# a_8049_45260# 2.52e-22
C33404 a_n971_45724# a_3503_45724# 0.011412f
C33405 a_n237_47217# a_3218_45724# 1.35e-20
C33406 a_584_46384# a_380_45546# 0.0075f
C33407 a_n2497_47436# a_1609_45822# 1.24e-19
C33408 a_2107_46812# a_4419_46090# 0.007223f
C33409 a_n881_46662# a_n2956_38680# 5.42e-20
C33410 a_12549_44172# a_19335_46494# 3.43e-19
C33411 a_n1925_46634# a_8199_44636# 0.007627f
C33412 a_13747_46662# a_14493_46090# 5.42e-19
C33413 a_n2661_46634# a_10355_46116# 6.98e-21
C33414 a_n743_46660# a_8016_46348# 0.155955f
C33415 a_5807_45002# a_15015_46420# 1.7e-19
C33416 a_n1613_43370# a_n1736_46482# 2.61e-19
C33417 a_9804_47204# a_6945_45028# 0.028722f
C33418 a_18834_46812# a_19333_46634# 3.48e-20
C33419 a_1799_45572# a_167_45260# 0.061186f
C33420 a_2443_46660# a_1823_45246# 0.001195f
C33421 a_n2661_46098# a_2202_46116# 0.002327f
C33422 a_3877_44458# a_n2293_46098# 0.030683f
C33423 a_n1644_44306# a_n1699_43638# 2.06e-19
C33424 a_895_43940# a_1568_43370# 3.85e-20
C33425 a_1414_42308# a_4699_43561# 4.09e-21
C33426 a_22959_43948# a_14021_43940# 3.06e-19
C33427 a_n2661_44458# a_9127_43156# 6.51e-21
C33428 a_11827_44484# a_15567_42826# 8.21e-22
C33429 a_7281_43914# a_n97_42460# 4.63e-19
C33430 a_18494_42460# a_18083_42858# 0.002227f
C33431 a_18184_42460# a_17333_42852# 1.09e-19
C33432 a_10405_44172# a_10651_43940# 0.014272f
C33433 a_n356_44636# a_4361_42308# 0.030056f
C33434 a_10729_43914# a_10555_43940# 6.54e-19
C33435 a_2479_44172# a_1756_43548# 1.44e-20
C33436 a_742_44458# a_4520_42826# 9.98e-21
C33437 a_n2293_42834# a_7573_43172# 1.55e-19
C33438 a_n913_45002# a_1755_42282# 0.169955f
C33439 a_n1059_45260# a_2123_42473# 0.002629f
C33440 a_n2017_45002# a_2351_42308# 0.0062f
C33441 a_3357_43084# a_3905_42558# 2.81e-19
C33442 a_5013_44260# VDD 0.198233f
C33443 a_13249_42308# a_15599_45572# 6.02e-22
C33444 a_13904_45546# a_15903_45785# 8.4e-22
C33445 a_15143_45578# a_15225_45822# 0.004937f
C33446 a_10210_45822# a_10544_45572# 2.43e-19
C33447 a_10907_45822# a_10306_45572# 2.2e-19
C33448 a_17538_32519# a_20202_43084# 2.29e-20
C33449 a_12379_42858# a_12891_46348# 0.001173f
C33450 a_n4318_38680# a_n2438_43548# 0.001622f
C33451 a_7274_43762# a_3090_45724# 1.37e-19
C33452 a_18079_43940# a_17715_44484# 4.31e-19
C33453 a_17973_43940# a_18189_46348# 4.22e-19
C33454 a_n2840_42282# SMPL_ON_P 6.32e-19
C33455 COMP_P w_1575_34946# 2.48e-19
C33456 a_20623_46660# VDD 0.194217f
C33457 a_14113_42308# CAL_N 0.001678f
C33458 a_n1853_46287# a_n2956_39304# 8.18e-20
C33459 a_n2293_46098# a_n1736_46482# 0.002983f
C33460 a_n2157_46122# a_n2956_38680# 0.001648f
C33461 a_13059_46348# a_12638_46436# 0.053952f
C33462 a_19466_46812# a_19443_46116# 0.004595f
C33463 a_15227_44166# a_21071_46482# 0.004602f
C33464 a_3147_46376# a_2324_44458# 2.35e-21
C33465 a_8199_44636# a_10355_46116# 0.176325f
C33466 a_8953_45546# a_9569_46155# 0.014447f
C33467 a_8016_46348# a_11189_46129# 1.23e-20
C33468 a_n4209_39590# a_n4064_37984# 0.032388f
C33469 a_n3565_39590# a_n3420_37984# 0.031465f
C33470 a_2982_43646# a_14358_43442# 8.47e-21
C33471 a_n97_42460# a_16409_43396# 0.002137f
C33472 a_n2293_43922# a_564_42282# 8.6e-20
C33473 a_n356_44636# a_6761_42308# 1.57e-19
C33474 a_6765_43638# a_6643_43396# 3.16e-19
C33475 a_6031_43396# a_7221_43396# 2.56e-19
C33476 a_10807_43548# a_12089_42308# 0.002697f
C33477 a_18184_42460# a_18997_42308# 2.46e-19
C33478 a_11967_42832# a_17665_42852# 4.85e-19
C33479 a_4915_47217# CLK 0.198293f
C33480 a_6151_47436# DATA[4] 2.92e-19
C33481 a_6545_47178# DATA[3] 0.178561f
C33482 a_8162_45546# a_8103_44636# 5.17e-20
C33483 a_15903_45785# a_17023_45118# 6.24e-21
C33484 a_9049_44484# a_5343_44458# 1.3e-20
C33485 a_3429_45260# a_3537_45260# 0.138977f
C33486 a_3065_45002# a_4574_45260# 4.96e-19
C33487 a_413_45260# a_3232_43370# 0.004402f
C33488 a_7765_42852# a_4185_45028# 1.44e-20
C33489 a_19339_43156# a_20202_43084# 2.42e-20
C33490 a_n2302_40160# a_n2312_39304# 3.32e-19
C33491 a_648_43396# a_n863_45724# 6.1e-19
C33492 a_3626_43646# a_n755_45592# 0.095572f
C33493 a_3539_42460# a_n357_42282# 0.019382f
C33494 a_1756_43548# a_n443_42852# 0.006388f
C33495 a_11823_42460# a_13661_43548# 0.116839f
C33496 a_12791_45546# a_5807_45002# 7.66e-21
C33497 a_7499_43078# a_n2661_46634# 3.96e-20
C33498 a_6598_45938# a_2107_46812# 1.55e-20
C33499 a_3175_45822# a_1799_45572# 6.77e-21
C33500 a_16680_45572# a_11453_44696# 2.06e-21
C33501 a_18691_45572# a_16327_47482# 0.162157f
C33502 a_16147_45260# a_10227_46804# 0.001138f
C33503 a_2437_43646# a_5129_47502# 0.004f
C33504 a_3357_43084# a_4791_45118# 0.144996f
C33505 a_3065_45002# a_n2497_47436# 0.022803f
C33506 a_n467_45028# a_n971_45724# 2.65e-20
C33507 a_n2017_45002# a_584_46384# 4e-20
C33508 a_n955_45028# a_n746_45260# 2.13e-20
C33509 a_15682_43940# a_4958_30871# 2.92e-20
C33510 a_104_43370# a_n3674_37592# 2.95e-21
C33511 a_16823_43084# a_16414_43172# 0.024882f
C33512 a_15743_43084# a_21356_42826# 0.004418f
C33513 a_5649_42852# a_10991_42826# 3.31e-20
C33514 a_4361_42308# a_12379_42858# 2.98e-19
C33515 a_743_42282# a_13635_43156# 4.32e-19
C33516 a_n97_42460# a_564_42282# 4.81e-20
C33517 a_11341_43940# a_15890_42674# 3.39e-22
C33518 a_15493_43940# a_15803_42450# 1.43e-21
C33519 a_n4318_39768# a_n4334_39616# 0.084616f
C33520 a_n3674_39768# a_n4209_39590# 0.044895f
C33521 a_n2661_42282# a_7174_31319# 2.04e-20
C33522 a_15227_44166# EN_OFFSET_CAL 2.2e-20
C33523 a_7754_39964# a_8530_39574# 9.77e-19
C33524 VDAC_Pi a_7754_38470# 0.008396f
C33525 a_7754_39632# a_3754_38470# 0.002634f
C33526 a_196_42282# VDD 0.291844f
C33527 a_10907_45822# a_10729_43914# 0.00119f
C33528 a_n2661_43370# a_6298_44484# 6.23e-19
C33529 a_10193_42453# a_15493_43940# 0.597095f
C33530 a_19778_44110# a_19929_45028# 0.001438f
C33531 a_5205_44484# a_n2661_43922# 0.032439f
C33532 a_22465_38105# a_20202_43084# 1.3e-19
C33533 a_9061_43230# a_n357_42282# 7.05e-20
C33534 a_2351_42308# a_526_44458# 8.58e-19
C33535 a_2123_42473# a_n1925_42282# 5.44e-20
C33536 a_8649_43218# a_n755_45592# 1.17e-19
C33537 a_5193_43172# a_n443_42852# 4.01e-19
C33538 a_12563_42308# a_9290_44172# 0.052279f
C33539 a_n2661_42834# a_n746_45260# 0.01463f
C33540 a_n2661_43922# a_n971_45724# 0.052944f
C33541 a_5826_44734# a_4791_45118# 3.51e-20
C33542 a_15037_45618# a_11415_45002# 5.65e-19
C33543 a_13163_45724# a_3483_46348# 5.34e-20
C33544 a_11823_42460# a_4185_45028# 3.07e-19
C33545 a_14309_45028# a_13747_46662# 1.11e-19
C33546 a_16147_45260# a_17339_46660# 0.006901f
C33547 a_18494_42460# a_12549_44172# 0.331306f
C33548 a_16321_45348# a_13661_43548# 3.11e-19
C33549 a_18248_44752# a_12861_44030# 0.072535f
C33550 a_14539_43914# a_11599_46634# 5.29e-21
C33551 a_10334_44484# a_10227_46804# 0.020432f
C33552 a_7499_43078# a_8199_44636# 0.859274f
C33553 a_8568_45546# a_5937_45572# 0.028968f
C33554 a_6194_45824# a_2324_44458# 0.001699f
C33555 a_10053_45546# a_8016_46348# 0.017312f
C33556 a_6709_45028# a_7715_46873# 3.14e-19
C33557 a_7229_43940# a_7577_46660# 1.48e-22
C33558 a_3357_43084# a_16292_46812# 1.44e-20
C33559 a_2437_43646# a_15227_44166# 0.167451f
C33560 a_7705_45326# a_7411_46660# 2.02e-20
C33561 a_8387_43230# a_8685_42308# 1.16e-19
C33562 a_16823_43084# a_7174_31319# 7.12e-22
C33563 a_n2293_42282# a_1067_42314# 1.58e-19
C33564 a_8605_42826# a_8791_42308# 0.001071f
C33565 a_5649_42852# a_17303_42282# 0.060649f
C33566 a_4361_42308# a_18727_42674# 0.006318f
C33567 a_4190_30871# a_19511_42282# 0.005903f
C33568 a_133_42852# a_n784_42308# 1.2e-19
C33569 a_14401_32519# C7_N_btm 9.48e-19
C33570 a_17538_32519# C5_N_btm 4.27e-20
C33571 a_11453_44696# a_13747_46662# 0.046437f
C33572 a_12465_44636# a_20843_47204# 8.77e-22
C33573 a_4883_46098# a_20916_46384# 0.471396f
C33574 a_21496_47436# a_21588_30879# 6.1e-19
C33575 a_n971_45724# a_7927_46660# 0.035261f
C33576 a_n1741_47186# a_10428_46928# 3.82e-19
C33577 a_n1151_42308# a_5167_46660# 0.011285f
C33578 a_4700_47436# a_4646_46812# 0.010115f
C33579 a_4791_45118# a_3877_44458# 0.024145f
C33580 a_n237_47217# a_7577_46660# 0.032223f
C33581 a_584_46384# a_3633_46660# 1.85e-22
C33582 a_2063_45854# a_5275_47026# 1.75e-19
C33583 a_8696_44636# a_17499_43370# 5.21e-19
C33584 a_17719_45144# a_18079_43940# 2.13e-20
C33585 a_n1699_44726# a_n1644_44306# 3.98e-19
C33586 a_9313_44734# a_11967_42832# 0.216837f
C33587 a_4223_44672# a_5495_43940# 0.06577f
C33588 a_1307_43914# a_15037_43940# 0.004228f
C33589 a_n1177_44458# a_n4318_39768# 1.8e-20
C33590 en_comp a_2982_43646# 0.021697f
C33591 a_4927_45028# VDD 0.159822f
C33592 COMP_P a_22609_38406# 0.00369f
C33593 a_18114_32519# a_11415_45002# 0.002006f
C33594 a_19721_31679# a_20202_43084# 3.09e-20
C33595 a_18545_45144# a_12741_44636# 2.26e-19
C33596 a_15004_44636# a_13059_46348# 2.9e-20
C33597 a_5891_43370# a_3090_45724# 0.166094f
C33598 a_1467_44172# a_n2438_43548# 9.81e-19
C33599 a_2675_43914# a_n2293_46634# 0.026226f
C33600 a_2537_44260# a_768_44030# 1.56e-20
C33601 a_5111_44636# a_8034_45724# 9.19e-22
C33602 a_3537_45260# a_8049_45260# 7.55e-20
C33603 a_n2661_43370# a_5937_45572# 0.202031f
C33604 a_6517_45366# a_2324_44458# 0.002583f
C33605 a_13565_44260# a_10227_46804# 8.58e-20
C33606 a_n447_43370# a_n971_45724# 0.113797f
C33607 a_458_43396# a_n2497_47436# 4.17e-20
C33608 a_n3674_38680# a_n3420_39072# 0.172947f
C33609 a_13575_42558# a_13657_42558# 0.171361f
C33610 a_13070_42354# a_14113_42308# 1.66e-20
C33611 a_5934_30871# a_4958_30871# 0.018095f
C33612 a_n1630_35242# a_n3690_39616# 9.65e-20
C33613 a_n1741_47186# VDD 0.912651f
C33614 DATA[5] CLK 0.059607f
C33615 a_768_44030# a_12741_44636# 0.03898f
C33616 a_n1925_46634# a_765_45546# 0.029508f
C33617 a_13661_43548# a_18280_46660# 4.34e-19
C33618 a_20916_46384# a_21188_46660# 0.003748f
C33619 a_7577_46660# a_8270_45546# 1.63e-19
C33620 a_6755_46942# a_6969_46634# 0.085936f
C33621 a_7927_46660# a_8023_46660# 0.013793f
C33622 a_8145_46902# a_8189_46660# 3.69e-19
C33623 a_7411_46660# a_8601_46660# 2.56e-19
C33624 a_n743_46660# a_15312_46660# 1.45e-21
C33625 a_n881_46662# a_n1423_46090# 4.07e-19
C33626 a_n1613_43370# a_n1641_46494# 0.152421f
C33627 a_4883_46098# a_6165_46155# 0.006098f
C33628 a_11599_46634# a_14493_46090# 0.018622f
C33629 a_10227_46804# a_9290_44172# 0.918064f
C33630 a_13717_47436# a_15682_46116# 9.15e-21
C33631 a_12861_44030# a_2324_44458# 0.95556f
C33632 a_6545_47178# a_6945_45028# 0.09952f
C33633 a_584_46384# a_526_44458# 0.458472f
C33634 a_2063_45854# a_2981_46116# 0.001617f
C33635 a_11967_42832# a_20974_43370# 2.01e-20
C33636 a_14539_43914# a_14358_43442# 2.26e-19
C33637 a_5891_43370# a_6547_43396# 6.62e-20
C33638 a_15004_44636# a_15095_43370# 9.09e-22
C33639 a_n2293_42834# a_2905_42968# 0.010834f
C33640 a_n2293_43922# a_n1557_42282# 2.21e-19
C33641 a_10193_42453# a_5742_30871# 0.303452f
C33642 a_16922_45042# a_20749_43396# 0.106779f
C33643 a_19279_43940# a_19808_44306# 0.002998f
C33644 a_10057_43914# a_12293_43646# 3.63e-20
C33645 a_18184_42460# a_13678_32519# 0.019189f
C33646 a_n1059_45260# a_8495_42852# 0.00552f
C33647 a_n4209_38216# VREF 0.055795f
C33648 a_n3565_38216# VIN_P 0.029343f
C33649 a_2711_45572# a_6229_45572# 4.93e-19
C33650 a_13483_43940# a_12741_44636# 9.28e-21
C33651 a_18533_43940# a_3090_45724# 5.95e-19
C33652 a_18429_43548# a_13661_43548# 0.010678f
C33653 a_8147_43396# a_4646_46812# 5.39e-20
C33654 a_14537_43646# a_n2293_46634# 0.00342f
C33655 a_15940_43402# a_12549_44172# 1.28e-20
C33656 a_5534_30871# a_4915_47217# 5.12e-19
C33657 a_743_42282# a_n1613_43370# 2.11e-19
C33658 a_9313_44734# a_13259_45724# 0.048952f
C33659 a_2437_43646# EN_OFFSET_CAL 7.51e-19
C33660 a_3357_43084# DATA[3] 0.066637f
C33661 a_7832_46660# VDD 0.077608f
C33662 a_6123_31319# VDAC_Pi 1.96e-19
C33663 a_n784_42308# VDAC_N 0.010218f
C33664 a_1606_42308# a_n4064_37440# 0.002946f
C33665 COMP_P a_22521_40599# 0.204681f
C33666 a_13059_46348# a_13759_46122# 0.249771f
C33667 a_19692_46634# a_6945_45028# 0.669658f
C33668 a_19333_46634# a_10809_44734# 0.011589f
C33669 a_14180_46812# a_2324_44458# 4.9e-20
C33670 a_15227_44166# a_22959_46124# 1.38e-19
C33671 a_10249_46116# a_9823_46482# 1.82e-19
C33672 a_1799_45572# a_n863_45724# 7.63e-20
C33673 a_2107_46812# a_1848_45724# 2.4e-19
C33674 a_2959_46660# a_n2661_45546# 6.8e-21
C33675 a_10428_46928# a_10586_45546# 4.33e-19
C33676 a_171_46873# a_n23_45546# 1.53e-20
C33677 a_n2661_46098# a_n1079_45724# 3.76e-21
C33678 a_n2293_46634# a_2277_45546# 0.001814f
C33679 a_n1853_46287# a_n1991_46122# 0.737461f
C33680 a_n2157_46122# a_n1423_46090# 0.053479f
C33681 a_n2293_46098# a_n1641_46494# 0.006575f
C33682 a_19328_44172# a_15743_43084# 2.2e-21
C33683 a_1209_43370# a_1049_43396# 0.194938f
C33684 a_n97_42460# a_n1557_42282# 0.149645f
C33685 a_n699_43396# a_196_42282# 0.001148f
C33686 a_11341_43940# a_16547_43609# 2.97e-19
C33687 a_n1644_44306# a_n2157_42858# 2.8e-20
C33688 a_453_43940# a_791_42968# 1.04e-20
C33689 a_1414_42308# a_1847_42826# 7.16e-21
C33690 a_15493_43940# a_16137_43396# 0.043956f
C33691 a_11967_42832# a_18599_43230# 0.003648f
C33692 a_15493_43396# a_18783_43370# 0.029898f
C33693 a_458_43396# a_1568_43370# 2.29e-20
C33694 a_n2956_37592# a_n2216_39072# 1.2e-19
C33695 a_4699_43561# VDD 0.262218f
C33696 a_2711_45572# a_18587_45118# 7.13e-22
C33697 a_21513_45002# a_22223_45572# 5.7e-19
C33698 a_20719_45572# a_3357_43084# 2.25e-19
C33699 a_n2104_42282# a_n2312_38680# 2.73e-20
C33700 a_2903_42308# a_768_44030# 2.31e-19
C33701 a_n4318_37592# a_n2442_46660# 0.023729f
C33702 a_20974_43370# a_13259_45724# 2.3e-20
C33703 a_15051_42282# a_10227_46804# 0.361922f
C33704 a_n2302_39866# SMPL_ON_P 5.6e-20
C33705 a_10586_45546# VDD 0.582083f
C33706 a_8696_44636# a_n237_47217# 4e-22
C33707 a_13904_45546# a_13717_47436# 8.89e-22
C33708 a_13527_45546# a_12861_44030# 0.274077f
C33709 a_11823_42460# a_14955_47212# 8.49e-21
C33710 a_12427_45724# a_11599_46634# 1.84e-20
C33711 a_9049_44484# a_10227_46804# 1.51e-20
C33712 a_8049_45260# a_9241_46436# 0.009374f
C33713 a_8034_45724# a_8379_46155# 0.001152f
C33714 a_22223_46124# a_20205_31679# 0.160234f
C33715 a_20708_46348# a_21167_46155# 6.64e-19
C33716 a_6945_45028# a_20692_30879# 6.72e-20
C33717 a_21259_43561# a_4190_30871# 0.198353f
C33718 a_18579_44172# a_13258_32519# 3.63e-20
C33719 a_9145_43396# a_9127_43156# 0.001269f
C33720 a_8685_43396# a_10991_42826# 1.51e-19
C33721 a_n2661_42282# a_5932_42308# 0.070536f
C33722 a_3422_30871# a_19332_42282# 6.32e-20
C33723 a_3877_44458# DATA[3] 1.85e-20
C33724 a_18114_32519# C6_N_btm 2.2e-19
C33725 a_19721_31679# C5_N_btm 1.11e-20
C33726 a_10951_45334# a_n2661_44458# 2.65e-20
C33727 a_16751_45260# a_11691_44458# 1.98e-19
C33728 a_4880_45572# a_3905_42865# 1.35e-19
C33729 a_16019_45002# a_16237_45028# 0.053167f
C33730 a_15861_45028# a_17517_44484# 0.003385f
C33731 a_7418_45067# a_n2661_43370# 4e-19
C33732 a_8696_44636# a_18204_44850# 7.09e-21
C33733 a_5111_44636# a_4743_44484# 0.02485f
C33734 a_5147_45002# a_5343_44458# 0.063193f
C33735 a_3537_45260# a_8103_44636# 0.140404f
C33736 a_n2661_45010# a_n1809_44850# 0.006483f
C33737 a_3232_43370# a_2779_44458# 0.003663f
C33738 a_421_43172# a_n443_42852# 4.81e-19
C33739 a_18599_43230# a_13259_45724# 1.09e-19
C33740 a_8605_42826# a_n357_42282# 0.011429f
C33741 a_8037_42858# a_n755_45592# 0.033004f
C33742 a_2711_45572# a_11415_45002# 0.337384f
C33743 a_13904_45546# a_14035_46660# 8.04e-20
C33744 a_13777_45326# a_12549_44172# 1.49e-20
C33745 a_13556_45296# a_768_44030# 0.267809f
C33746 a_14180_45002# a_12891_46348# 2.92e-20
C33747 a_8696_44636# a_8270_45546# 0.023406f
C33748 a_7499_43078# a_765_45546# 2.08e-20
C33749 a_n37_45144# a_171_46873# 2.73e-19
C33750 a_327_44734# a_n2438_43548# 0.013318f
C33751 a_1667_45002# a_n743_46660# 2.23e-20
C33752 a_2382_45260# a_n1925_46634# 8.42e-21
C33753 a_3429_45260# a_n2293_46634# 0.001376f
C33754 a_413_45260# a_n133_46660# 3.34e-21
C33755 a_626_44172# a_n1613_43370# 0.001807f
C33756 a_16922_45042# a_12861_44030# 0.120012f
C33757 a_11691_44458# a_4915_47217# 0.020788f
C33758 a_n1386_35608# VDD 0.360375f
C33759 a_n1352_44484# a_n746_45260# 0.001882f
C33760 a_n452_44636# a_n971_45724# 1.31e-21
C33761 a_n1641_43230# a_n1630_35242# 6.83e-20
C33762 a_n13_43084# a_n327_42558# 2.86e-20
C33763 a_n1076_43230# a_n3674_37592# 4.57e-20
C33764 a_4361_42308# a_3823_42558# 0.114877f
C33765 a_5534_30871# a_13291_42460# 0.045073f
C33766 a_14543_43071# a_14635_42282# 0.075815f
C33767 a_10341_43396# a_15890_42674# 7.05e-21
C33768 a_743_42282# a_3905_42558# 0.003412f
C33769 a_n2293_42282# a_4149_42891# 1.94e-19
C33770 a_10809_44734# CLK 0.002918f
C33771 a_n3420_39072# VDD 1.01442f
C33772 a_4915_47217# a_4842_47243# 1.81e-19
C33773 a_6151_47436# a_n1613_43370# 0.548675f
C33774 a_n2833_47464# a_n2442_46660# 0.055535f
C33775 a_n2497_47436# a_n2472_46634# 0.009668f
C33776 a_n2288_47178# a_n2661_46634# 1.83e-19
C33777 a_n2109_47186# a_n2956_39768# 4.34e-19
C33778 a_n1151_42308# a_12549_44172# 0.466584f
C33779 a_18479_47436# a_19787_47423# 0.029306f
C33780 a_18780_47178# a_19386_47436# 3.06e-19
C33781 a_16023_47582# a_4883_46098# 5.48e-21
C33782 a_16588_47582# a_13507_46334# 3.49e-21
C33783 a_10227_46804# a_20990_47178# 0.004463f
C33784 a_16241_47178# a_12465_44636# 2.08e-19
C33785 a_11599_46634# a_11453_44696# 0.075707f
C33786 a_21359_45002# a_21398_44850# 0.001485f
C33787 a_12883_44458# a_n2293_43922# 0.06281f
C33788 a_13556_45296# a_13483_43940# 0.001149f
C33789 a_9482_43914# a_14955_43940# 6.17e-19
C33790 a_18989_43940# a_9313_44734# 1.23e-19
C33791 a_18114_32519# a_11967_42832# 0.002218f
C33792 a_n2293_42834# a_5495_43940# 1.87e-21
C33793 a_1307_43914# a_9028_43914# 0.010468f
C33794 a_11823_42460# a_14579_43548# 0.106967f
C33795 a_20193_45348# a_18579_44172# 2.14e-20
C33796 a_n356_44636# a_5891_43370# 4.5e-19
C33797 a_12607_44458# a_13213_44734# 1.94e-19
C33798 a_11691_44458# a_18681_44484# 0.002372f
C33799 a_7499_43078# a_8945_43396# 2.24e-19
C33800 a_n2661_43370# a_2479_44172# 4.26e-20
C33801 a_11827_44484# a_20980_44850# 0.002088f
C33802 a_6171_45002# a_11341_43940# 5.17e-20
C33803 a_n3565_38216# a_n2956_38680# 0.003389f
C33804 a_18175_45572# VDD 0.38478f
C33805 a_17333_42852# RST_Z 1.2e-21
C33806 a_8953_45002# a_3483_46348# 0.121322f
C33807 a_17517_44484# a_19321_45002# 0.264473f
C33808 a_11827_44484# a_19692_46634# 0.04136f
C33809 a_20640_44752# a_12549_44172# 0.004896f
C33810 a_4574_45260# a_5937_45572# 7.5e-21
C33811 a_3537_45260# a_8953_45546# 0.009809f
C33812 a_5111_44636# a_8016_46348# 0.001121f
C33813 a_n913_45002# a_2324_44458# 1.92e-20
C33814 a_5205_44484# a_5164_46348# 7.43e-20
C33815 a_3232_43370# a_6165_46155# 9.41e-20
C33816 a_3357_43084# a_6945_45028# 0.033591f
C33817 a_19479_31679# a_22223_46124# 4.31e-19
C33818 a_16842_45938# a_8049_45260# 1.72e-19
C33819 a_15037_45618# a_13259_45724# 0.098143f
C33820 a_n784_42308# a_5742_30871# 0.550812f
C33821 a_2903_42308# a_6123_31319# 2.22e-20
C33822 a_1606_42308# a_8685_42308# 1.35e-20
C33823 a_16245_42852# a_4958_30871# 6.84e-19
C33824 a_13887_32519# C6_N_btm 1.01e-19
C33825 a_17364_32525# C2_N_btm 1.14e-20
C33826 CAL_P a_22717_37285# 1.35e-20
C33827 a_22609_38406# a_22705_37990# 3.51e-20
C33828 a_12465_44636# a_16721_46634# 9.65e-22
C33829 a_3080_42308# VDAC_N 0.007207f
C33830 a_18597_46090# a_19123_46287# 0.188676f
C33831 a_10227_46804# a_20273_46660# 0.037464f
C33832 a_18479_47436# a_20107_46660# 0.019527f
C33833 a_15811_47375# a_16434_46660# 2.88e-19
C33834 a_6151_47436# a_n2293_46098# 9.86e-20
C33835 a_2063_45854# a_167_45260# 0.359284f
C33836 a_584_46384# a_2521_46116# 4.33e-19
C33837 a_n971_45724# a_5164_46348# 1.88e-20
C33838 a_n237_47217# a_4704_46090# 0.042359f
C33839 a_n2293_46634# a_6755_46942# 1.78e-19
C33840 a_n2661_46634# a_6999_46987# 2.56e-19
C33841 a_5807_45002# a_8846_46660# 6.99e-19
C33842 a_768_44030# a_13607_46688# 2.12e-20
C33843 a_3699_46634# a_4817_46660# 1.58e-19
C33844 a_3524_46660# a_4955_46873# 7.68e-19
C33845 a_2107_46812# a_7411_46660# 7.26e-20
C33846 a_n743_46660# a_10428_46928# 4.37e-20
C33847 a_12549_44172# a_14084_46812# 0.007343f
C33848 a_n699_43396# a_4699_43561# 6.51e-20
C33849 a_742_44458# a_n1557_42282# 6.13e-20
C33850 a_n1761_44111# a_n1644_44306# 0.170098f
C33851 a_2479_44172# a_2998_44172# 0.004129f
C33852 a_14673_44172# a_11341_43940# 0.001734f
C33853 a_11967_42832# a_17737_43940# 0.054562f
C33854 a_4223_44672# a_3080_42308# 2.46e-19
C33855 a_n2065_43946# a_n1453_44318# 0.001881f
C33856 a_5891_43370# a_9165_43940# 8.35e-19
C33857 a_n2661_42834# a_726_44056# 6.09e-19
C33858 a_n1899_43946# a_n3674_39768# 4.83e-19
C33859 a_413_45260# a_2905_42968# 1.46e-20
C33860 a_n1059_45260# a_9127_43156# 0.006366f
C33861 a_n913_45002# a_8387_43230# 0.024148f
C33862 a_n2017_45002# a_8952_43230# 4.34e-20
C33863 a_10440_44484# VDD 0.159539f
C33864 a_n4064_40160# C9_P_btm 0.003109f
C33865 a_22485_44484# a_11415_45002# 3.2e-20
C33866 a_10807_43548# a_3090_45724# 0.031941f
C33867 a_6293_42852# a_768_44030# 5.95e-20
C33868 a_2982_43646# a_13661_43548# 2.6e-20
C33869 a_n2661_43370# a_n443_42852# 0.082119f
C33870 a_22223_45036# a_20205_31679# 2.02e-20
C33871 a_13213_44734# a_10903_43370# 4.28e-19
C33872 a_16547_43609# a_16327_47482# 0.00506f
C33873 a_13749_43396# a_10227_46804# 3.64e-19
C33874 a_15743_43084# a_12861_44030# 0.01437f
C33875 a_743_42282# a_4791_45118# 0.053017f
C33876 a_n3674_39304# SMPL_ON_P 0.040131f
C33877 a_n4064_39616# a_n4064_39072# 0.062881f
C33878 a_n4064_40160# a_n4209_38502# 0.05515f
C33879 a_n4315_30879# a_n3565_38502# 0.085594f
C33880 a_n3420_39616# a_n4251_39392# 8.88e-19
C33881 a_n743_46660# VDD 1.75634f
C33882 a_6123_31319# C9_N_btm 9.33e-20
C33883 a_5934_30871# C7_N_btm 0.007575f
C33884 a_10768_47026# a_3483_46348# 4.61e-20
C33885 a_n2293_46634# a_8049_45260# 1.91e-20
C33886 a_13747_46662# a_14180_46482# 0.008333f
C33887 a_n2661_46098# a_1337_46436# 4.38e-19
C33888 a_2107_46812# a_4365_46436# 1.79e-19
C33889 a_10428_46928# a_11189_46129# 6.48e-21
C33890 a_6755_46942# a_9625_46129# 3.29e-19
C33891 a_10467_46802# a_9290_44172# 2.22e-19
C33892 a_3877_44458# a_6945_45028# 0.001558f
C33893 a_20679_44626# a_4361_42308# 2.91e-20
C33894 a_18989_43940# a_18599_43230# 5.3e-19
C33895 a_9028_43914# a_9396_43370# 3.1e-19
C33896 a_18579_44172# a_20301_43646# 3.55e-20
C33897 a_19862_44208# a_2982_43646# 0.005666f
C33898 a_9313_44734# a_10518_42984# 0.008938f
C33899 a_n2293_43922# a_3935_42891# 1.63e-22
C33900 a_n2661_42834# a_5111_42852# 5.01e-22
C33901 a_n356_44636# a_17595_43084# 2.73e-20
C33902 a_n2293_42834# a_n784_42308# 8.13e-19
C33903 a_1307_43914# a_5421_42558# 4.2e-20
C33904 a_15493_43396# a_3626_43646# 2.49e-20
C33905 a_n1059_45260# a_17124_42282# 0.008817f
C33906 a_2711_45572# a_13159_45002# 9.08e-19
C33907 a_7227_45028# a_7229_43940# 0.019397f
C33908 a_6598_45938# a_6709_45028# 3.05e-21
C33909 a_4880_45572# a_5147_45002# 3.65e-19
C33910 a_13249_42308# a_n2017_45002# 0.030327f
C33911 a_5755_42308# a_4791_45118# 0.003736f
C33912 a_22521_40599# a_22705_37990# 1.29e-19
C33913 a_22469_40625# a_22609_37990# 0.130478f
C33914 CAL_N a_22717_37285# 7.87e-21
C33915 a_n3565_37414# C5_P_btm 1.11e-20
C33916 a_n3420_37440# C7_P_btm 1.33e-20
C33917 a_6886_37412# a_n923_35174# 0.003125f
C33918 a_2982_43646# a_4185_45028# 0.243496f
C33919 a_22400_42852# SMPL_ON_N 3.97e-19
C33920 a_7754_38470# RST_Z 0.034995f
C33921 a_5025_43940# a_526_44458# 1.8e-20
C33922 a_2998_44172# a_n443_42852# 1.29e-19
C33923 a_3499_42826# a_n2661_45546# 5.13e-21
C33924 a_17737_43940# a_13259_45724# 0.016944f
C33925 a_11189_46129# VDD 0.944289f
C33926 a_3638_45822# a_n971_45724# 2.91e-19
C33927 a_7227_45028# a_n237_47217# 1.15e-19
C33928 a_3175_45822# a_2063_45854# 0.002195f
C33929 a_n3565_38502# a_n3420_37440# 0.034147f
C33930 a_n4209_38502# a_n4064_37440# 0.028279f
C33931 a_n4064_38528# a_n4209_37414# 0.027936f
C33932 a_n3420_38528# a_n3565_37414# 0.029229f
C33933 a_9625_46129# a_8049_45260# 0.04571f
C33934 a_8016_46348# a_8379_46155# 0.005265f
C33935 a_8953_45546# a_9241_46436# 2.17e-19
C33936 a_n809_44244# a_n1630_35242# 5.42e-21
C33937 a_10341_43396# a_16547_43609# 0.026476f
C33938 a_6031_43396# a_5649_42852# 4.06e-21
C33939 a_8791_43396# a_743_42282# 2.77e-21
C33940 a_n1557_42282# a_n901_43156# 2.27e-19
C33941 a_n97_42460# a_3935_42891# 5.1e-20
C33942 a_13565_43940# a_13460_43230# 6.29e-20
C33943 a_n1761_44111# a_961_42354# 1.47e-22
C33944 a_8685_43396# a_15231_43396# 0.002861f
C33945 a_12281_43396# a_13837_43396# 7.31e-21
C33946 a_1414_42308# a_n473_42460# 2.2e-21
C33947 a_768_44030# RST_Z 0.05505f
C33948 a_12549_44172# START 8.3e-19
C33949 a_n881_46662# CLK 0.023376f
C33950 a_8128_46384# DATA[3] 1.73e-19
C33951 a_1847_42826# VDD 0.527555f
C33952 a_n2956_37592# a_n2302_37984# 0.005102f
C33953 a_11525_45546# a_n2661_42834# 5.55e-21
C33954 a_11322_45546# a_n2661_43922# 0.001721f
C33955 a_16855_45546# a_14539_43914# 8.46e-20
C33956 a_8696_44636# a_15004_44636# 0.003323f
C33957 a_2711_45572# a_11967_42832# 0.068241f
C33958 a_11652_45724# a_11649_44734# 1.66e-19
C33959 a_2680_45002# a_n2661_43370# 0.006576f
C33960 a_19479_31679# a_22223_45036# 0.01502f
C33961 a_n913_45002# a_16922_45042# 6.18e-19
C33962 a_3357_43084# a_11827_44484# 8.78e-20
C33963 a_6171_45002# a_7418_45394# 1.2e-19
C33964 a_n3565_39304# a_n2956_39768# 0.003389f
C33965 a_15681_43442# a_n443_42852# 0.035093f
C33966 a_18783_43370# a_n357_42282# 5.79e-20
C33967 a_8952_43230# a_526_44458# 0.039329f
C33968 a_13887_32519# a_13259_45724# 0.002751f
C33969 a_n2293_42834# SMPL_ON_P 1.07e-19
C33970 a_501_45348# a_n443_46116# 1.62e-19
C33971 a_7227_45028# a_8270_45546# 1.35e-20
C33972 a_6171_45002# a_16327_47482# 0.001024f
C33973 a_413_45260# a_21496_47436# 8.97e-20
C33974 a_n2810_45028# a_n2312_40392# 0.055228f
C33975 a_2437_43646# a_7989_47542# 9.04e-19
C33976 a_21188_45572# a_12549_44172# 4.02e-21
C33977 a_18799_45938# a_13747_46662# 0.028671f
C33978 a_19256_45572# a_19321_45002# 0.004884f
C33979 a_6812_45938# a_6969_46634# 4.71e-20
C33980 a_10180_45724# a_10150_46912# 7.45e-19
C33981 a_10053_45546# a_10428_46928# 2.44e-21
C33982 a_10193_42453# a_9863_46634# 1.87e-19
C33983 a_19431_45546# a_19594_46812# 2.2e-19
C33984 a_6197_43396# a_7227_42308# 1.57e-20
C33985 a_18783_43370# a_18707_42852# 1.34e-19
C33986 a_13460_43230# a_5534_30871# 0.052631f
C33987 a_n97_42460# a_15890_42674# 0.022679f
C33988 a_3626_43646# a_8791_42308# 0.003196f
C33989 a_2982_43646# a_9803_42558# 1.36e-19
C33990 a_3080_42308# a_5742_30871# 0.097222f
C33991 a_791_42968# a_945_42968# 0.008535f
C33992 a_15743_43084# a_19518_43218# 0.00221f
C33993 a_16823_43084# a_17141_43172# 1.56e-19
C33994 a_17730_32519# C4_N_btm 6.79e-20
C33995 a_4915_47217# a_5129_47502# 0.070911f
C33996 a_n1151_42308# a_6575_47204# 1.72e-19
C33997 a_2124_47436# a_n1435_47204# 2.1e-19
C33998 a_4791_45118# a_6151_47436# 0.019937f
C33999 a_2063_45854# a_11459_47204# 8.65e-20
C34000 a_n443_46116# a_5815_47464# 5.77e-19
C34001 a_15486_42560# VDD 0.275297f
C34002 a_8103_44636# a_8701_44490# 5.82e-19
C34003 a_6298_44484# a_5883_43914# 0.003333f
C34004 a_18479_45785# a_15493_43940# 0.016583f
C34005 a_3065_45002# a_2889_44172# 1.06e-19
C34006 a_2382_45260# a_3600_43914# 0.158274f
C34007 a_n2661_45010# a_1525_44260# 5.65e-20
C34008 en_comp a_n3674_39768# 0.036087f
C34009 a_n2293_45010# a_n822_43940# 4.54e-19
C34010 a_n913_45002# a_n875_44318# 5.75e-19
C34011 a_2680_45002# a_2998_44172# 1.29e-20
C34012 a_10053_45546# VDD 0.150582f
C34013 a_13678_32519# RST_Z 0.048965f
C34014 a_14539_43914# a_13661_43548# 0.193767f
C34015 a_16751_45260# a_15227_44166# 1.7e-20
C34016 a_8103_44636# a_n2293_46634# 7.43e-21
C34017 a_20447_31679# a_21076_30879# 0.055814f
C34018 a_2711_45572# a_13259_45724# 1.26722f
C34019 a_9049_44484# a_8034_45724# 2.06e-20
C34020 a_7230_45938# a_8049_45260# 1.18e-19
C34021 a_413_45260# a_21363_46634# 3.6e-20
C34022 a_15599_45572# a_15682_46116# 0.009928f
C34023 a_15903_45785# a_2324_44458# 0.017867f
C34024 a_8696_44636# a_13759_46122# 1.49e-20
C34025 a_10617_44484# a_11453_44696# 3.76e-20
C34026 a_n2661_43922# a_12465_44636# 0.17969f
C34027 a_n809_44244# a_n971_45724# 0.002895f
C34028 a_2479_44172# a_n2497_47436# 4.48e-20
C34029 a_17333_42852# a_17303_42282# 5.44e-19
C34030 a_17701_42308# a_18057_42282# 4e-19
C34031 a_n4318_38680# a_n3420_39072# 0.310238f
C34032 a_n3674_38216# a_n4318_37592# 2.7294f
C34033 a_n4318_38216# a_n1329_42308# 2.61e-20
C34034 a_n2104_42282# COMP_P 3.78e-19
C34035 a_n3674_39304# a_n2946_39072# 4.03e-21
C34036 a_768_44030# a_2609_46660# 1.29e-19
C34037 a_n2661_46634# a_n2312_38680# 0.106815f
C34038 a_n2442_46660# a_n2293_46634# 0.004958f
C34039 a_n2472_46634# a_n2104_46634# 7.52e-19
C34040 a_n2956_39768# a_n1925_46634# 1.65e-19
C34041 a_n1613_43370# a_3221_46660# 0.003155f
C34042 a_4883_46098# a_8492_46660# 4.2e-20
C34043 a_4915_47217# a_15227_44166# 1.46e-20
C34044 a_n1435_47204# a_11813_46116# 2.37e-20
C34045 a_9482_43914# a_8685_43396# 3.32e-20
C34046 a_19778_44110# a_19741_43940# 0.054731f
C34047 a_12607_44458# a_11341_43940# 8.67e-21
C34048 a_17767_44458# a_15493_43396# 2.64e-21
C34049 a_18287_44626# a_18326_43940# 0.001026f
C34050 a_18248_44752# a_18451_43940# 5.78e-19
C34051 a_11967_42832# a_22485_44484# 3.29e-19
C34052 a_19279_43940# a_21398_44850# 0.183186f
C34053 a_n2661_43922# a_7281_43914# 1.21e-20
C34054 a_n2661_42834# a_7542_44172# 0.019328f
C34055 a_n2293_42834# a_3080_42308# 0.021566f
C34056 a_20640_44752# a_20637_44484# 2.36e-20
C34057 a_6109_44484# a_n2661_42282# 0.003425f
C34058 a_20766_44850# a_3422_30871# 6.2e-20
C34059 a_5883_43914# a_10555_44260# 2.18e-20
C34060 a_1307_43914# a_2437_43396# 2.02e-19
C34061 a_11827_44484# a_18533_44260# 3.57e-19
C34062 a_n2017_45002# a_19700_43370# 4.64e-20
C34063 a_n913_45002# a_15743_43084# 2.14e-19
C34064 a_6171_45002# a_10341_43396# 2.27e-20
C34065 a_6123_31319# RST_Z 0.004252f
C34066 a_5742_30871# a_n1532_35090# 1.92e-19
C34067 a_5934_30871# C3_P_btm 0.011274f
C34068 a_2437_43396# a_n443_46116# 7.55e-19
C34069 a_9313_44734# a_20202_43084# 0.044152f
C34070 a_17767_44458# a_3483_46348# 8.35e-19
C34071 a_10334_44484# a_8016_46348# 0.007545f
C34072 a_n2661_44458# a_2324_44458# 0.134417f
C34073 a_11691_44458# a_10809_44734# 0.354084f
C34074 a_9838_44484# a_8199_44636# 0.024921f
C34075 a_8701_44490# a_8953_45546# 0.005445f
C34076 a_5883_43914# a_5937_45572# 0.454323f
C34077 a_3537_45260# a_1609_45822# 1.84e-20
C34078 a_4574_45260# a_n443_42852# 1.14e-21
C34079 a_7499_43940# a_768_44030# 1.16e-19
C34080 a_14021_43940# a_21588_30879# 1.53e-20
C34081 a_n2661_42282# a_4646_46812# 0.025072f
C34082 a_19332_42282# a_7174_31319# 7.74e-19
C34083 a_5934_30871# a_n4064_38528# 0.004208f
C34084 a_21177_47436# VDD 0.179587f
C34085 a_8128_46384# a_6945_45028# 0.010979f
C34086 a_18597_46090# a_8049_45260# 0.047215f
C34087 a_11599_46634# a_14180_46482# 0.016275f
C34088 a_12861_44030# a_12839_46116# 0.003823f
C34089 a_n971_45724# a_3316_45546# 0.086835f
C34090 a_2063_45854# a_n863_45724# 4.66e-19
C34091 a_n237_47217# a_2957_45546# 5.41e-20
C34092 a_n2497_47436# a_n443_42852# 0.005218f
C34093 a_n1151_42308# a_n2661_45546# 0.044338f
C34094 a_13747_46662# a_13925_46122# 0.020304f
C34095 a_n743_46660# a_7920_46348# 0.006742f
C34096 a_5807_45002# a_14275_46494# 0.013842f
C34097 a_n2661_46634# a_9823_46155# 1.75e-20
C34098 a_n1925_46634# a_8349_46414# 0.006458f
C34099 a_12549_44172# a_19553_46090# 7.25e-21
C34100 a_n2293_46634# a_8953_45546# 0.04453f
C34101 a_6999_46987# a_765_45546# 2.41e-19
C34102 a_12469_46902# a_12925_46660# 4.2e-19
C34103 a_12251_46660# a_12513_46660# 0.001705f
C34104 a_12816_46660# a_12978_47026# 0.006453f
C34105 a_18834_46812# a_15227_44166# 0.231715f
C34106 a_11735_46660# a_14035_46660# 4.06e-21
C34107 a_1799_45572# a_2202_46116# 6.85e-20
C34108 a_n2661_46098# a_1823_45246# 9.15e-19
C34109 a_2107_46812# a_4185_45028# 0.008044f
C34110 a_n984_44318# a_n1557_42282# 2.08e-21
C34111 a_14673_44172# a_10341_43396# 1.61e-19
C34112 a_15493_43940# a_14021_43940# 0.08284f
C34113 a_2479_44172# a_1568_43370# 0.001043f
C34114 a_n699_43396# a_1847_42826# 5.48e-20
C34115 a_2779_44458# a_2905_42968# 2.56e-20
C34116 a_16922_45042# a_20922_43172# 1.86e-19
C34117 a_742_44458# a_3935_42891# 1.81e-19
C34118 a_11827_44484# a_5342_30871# 2.98e-20
C34119 a_18184_42460# a_18083_42858# 0.003624f
C34120 a_10405_44172# a_10555_43940# 0.018661f
C34121 a_10729_43914# a_9801_43940# 7.39e-20
C34122 a_1414_42308# a_4235_43370# 1.4e-19
C34123 a_18494_42460# a_17701_42308# 4.02e-20
C34124 a_n2293_42834# a_7309_43172# 5.7e-19
C34125 a_n1059_45260# a_1755_42282# 0.004197f
C34126 a_n913_45002# a_1606_42308# 0.025848f
C34127 a_n2017_45002# a_2123_42473# 0.0078f
C34128 a_5244_44056# VDD 0.146618f
C34129 a_15143_45578# a_15037_45618# 0.13675f
C34130 a_11823_42460# a_16115_45572# 9.08e-20
C34131 a_11652_45724# a_8696_44636# 3.56e-19
C34132 a_10907_45822# a_10216_45572# 1.14e-19
C34133 a_5829_43940# a_1823_45246# 1.54e-19
C34134 a_20974_43370# a_20202_43084# 0.026132f
C34135 a_n3674_39304# a_n2438_43548# 0.001617f
C34136 a_10991_42826# a_768_44030# 1.43e-20
C34137 a_11341_43940# a_10903_43370# 0.061205f
C34138 a_9248_44260# a_9290_44172# 5.95e-19
C34139 a_17973_43940# a_17715_44484# 0.00355f
C34140 a_1307_43914# CLK 8.72e-21
C34141 a_20841_46902# VDD 0.20446f
C34142 a_n2157_46122# a_n2956_39304# 7.88e-20
C34143 a_n2293_46098# a_n2956_38680# 0.022177f
C34144 a_19123_46287# a_8049_45260# 3.32e-19
C34145 a_13059_46348# a_12379_46436# 9.42e-19
C34146 a_15227_44166# a_20850_46482# 9.67e-19
C34147 a_2804_46116# a_2324_44458# 1.12e-21
C34148 a_8199_44636# a_9823_46155# 0.001773f
C34149 a_8953_45546# a_9625_46129# 0.009628f
C34150 a_8016_46348# a_9290_44172# 0.020766f
C34151 a_4958_30871# a_8530_39574# 1.39e-19
C34152 a_n4064_40160# a_n3607_38304# 5.58e-20
C34153 a_6031_43396# a_8685_43396# 9.68e-21
C34154 a_2982_43646# a_14579_43548# 5.95e-20
C34155 a_n97_42460# a_16547_43609# 0.066612f
C34156 a_n2661_42834# a_n1630_35242# 1.36e-19
C34157 a_11967_42832# a_16877_42852# 0.005423f
C34158 a_6765_43638# a_7274_43762# 2.6e-19
C34159 a_6197_43396# a_6643_43396# 2.28e-19
C34160 a_n2293_43922# a_n3674_37592# 0.062473f
C34161 a_10057_43914# a_5742_30871# 3.08e-19
C34162 a_6151_47436# DATA[3] 0.041263f
C34163 a_15903_45785# a_16922_45042# 5.01e-20
C34164 a_2711_45572# a_18989_43940# 0.006251f
C34165 a_7499_43078# a_5343_44458# 0.050528f
C34166 a_15861_45028# a_15685_45394# 8.17e-20
C34167 a_3065_45002# a_3537_45260# 0.162384f
C34168 a_7871_42858# a_4185_45028# 1.73e-20
C34169 a_18599_43230# a_20202_43084# 5.72e-21
C34170 a_n2302_40160# a_n2312_40392# 0.151095f
C34171 a_n4064_40160# a_n2312_39304# 5.41e-19
C34172 a_6197_43396# a_n2661_45546# 1.24e-21
C34173 a_548_43396# a_n863_45724# 0.001035f
C34174 a_3626_43646# a_n357_42282# 0.020238f
C34175 a_1568_43370# a_n443_42852# 0.038016f
C34176 a_17531_42308# a_12549_44172# 1.47e-21
C34177 a_14456_42282# a_n2293_46634# 3e-20
C34178 a_509_45572# VDD 1.36e-19
C34179 a_11823_42460# a_5807_45002# 0.022934f
C34180 a_6667_45809# a_2107_46812# 4.38e-20
C34181 a_2711_45572# a_1799_45572# 7.16e-20
C34182 a_16855_45546# a_11453_44696# 3.46e-20
C34183 a_18799_45938# a_11599_46634# 0.001679f
C34184 a_18909_45814# a_16327_47482# 0.16767f
C34185 a_2437_43646# a_4915_47217# 0.114772f
C34186 a_2680_45002# a_n2497_47436# 1.29e-19
C34187 a_n955_45028# a_n971_45724# 5.28e-19
C34188 a_3357_43084# a_4700_47436# 6.56e-19
C34189 a_n97_42460# a_n3674_37592# 0.012074f
C34190 a_15743_43084# a_20922_43172# 0.004395f
C34191 a_5649_42852# a_10796_42968# 3.16e-20
C34192 a_4361_42308# a_10341_42308# 0.006315f
C34193 a_743_42282# a_12895_43230# 6.86e-20
C34194 a_11341_43940# a_15959_42545# 1.71e-21
C34195 a_15493_43940# a_15764_42576# 1.53e-21
C34196 a_n4318_39768# a_n4209_39590# 0.105246f
C34197 a_3754_39134# a_3754_38802# 0.296258f
C34198 a_7754_39964# a_7754_38470# 0.241119f
C34199 a_3754_39466# VDAC_Ni 0.001054f
C34200 a_n3420_37984# a_n3607_37440# 2.09e-19
C34201 a_n473_42460# VDD 0.27195f
C34202 a_n2661_43370# a_5518_44484# 0.001247f
C34203 a_22223_45036# a_20193_45348# 2.8e-19
C34204 a_5205_44484# a_n2661_42834# 0.030553f
C34205 a_3232_43370# a_13213_44734# 6.1e-21
C34206 a_22397_42558# a_20202_43084# 1.54e-19
C34207 a_8649_43218# a_n357_42282# 3.99e-19
C34208 a_2123_42473# a_526_44458# 0.012631f
C34209 a_16877_42852# a_13259_45724# 3.34e-20
C34210 a_1755_42282# a_n1925_42282# 0.019802f
C34211 a_10723_42308# a_10903_43370# 1.71e-19
C34212 a_11633_42558# a_9290_44172# 0.014294f
C34213 a_n2661_42834# a_n971_45724# 0.165951f
C34214 a_9313_44734# a_2063_45854# 3.29e-20
C34215 a_5289_44734# a_4791_45118# 7.66e-19
C34216 a_10157_44484# a_10227_46804# 0.008568f
C34217 a_17970_44736# a_12861_44030# 0.001384f
C34218 a_2711_45572# a_18189_46348# 3.03e-20
C34219 a_8568_45546# a_8199_44636# 0.141772f
C34220 a_5907_45546# a_2324_44458# 0.002504f
C34221 a_9049_44484# a_8016_46348# 4.89e-19
C34222 a_11691_44458# a_n881_46662# 4.5e-20
C34223 a_6171_45002# a_8667_46634# 7.94e-23
C34224 a_3357_43084# a_15559_46634# 2.61e-21
C34225 a_7229_43940# a_7715_46873# 2.31e-19
C34226 a_14309_45028# a_13661_43548# 1.43e-19
C34227 a_n2661_43370# a_n2661_46634# 7.12e-19
C34228 a_n2293_42834# a_n2438_43548# 0.138621f
C34229 a_18184_42460# a_12549_44172# 0.03123f
C34230 a_8037_42858# a_8791_42308# 0.002879f
C34231 a_8387_43230# a_8325_42308# 0.003469f
C34232 a_n2293_42282# a_n1630_35242# 0.18361f
C34233 a_133_42852# a_196_42282# 4.15e-19
C34234 a_13291_42460# a_14635_42282# 0.111986f
C34235 a_5649_42852# a_4958_30871# 0.293366f
C34236 a_4361_42308# a_18057_42282# 0.008747f
C34237 a_13678_32519# a_17303_42282# 0.008395f
C34238 a_4190_30871# a_18548_42308# 0.001263f
C34239 a_14401_32519# C6_N_btm 0.054459f
C34240 a_17538_32519# C4_N_btm 3.39e-20
C34241 a_12465_44636# a_19594_46812# 9.01e-20
C34242 a_11453_44696# a_13661_43548# 0.099457f
C34243 a_21496_47436# a_20916_46384# 0.113102f
C34244 a_13507_46334# a_21588_30879# 6.05e-19
C34245 a_16588_47582# a_n743_46660# 1.72e-19
C34246 a_n971_45724# a_8145_46902# 0.051701f
C34247 a_n1741_47186# a_10150_46912# 2.54e-20
C34248 a_n237_47217# a_7715_46873# 0.051915f
C34249 a_n1151_42308# a_5385_46902# 0.0125f
C34250 a_4700_47436# a_3877_44458# 4.34e-21
C34251 a_n443_46116# a_3055_46660# 0.002062f
C34252 a_17719_45144# a_17973_43940# 6.82e-19
C34253 a_1423_45028# a_9801_43940# 5.54e-20
C34254 a_4743_44484# a_3905_42865# 3.75e-22
C34255 a_4223_44672# a_5013_44260# 0.07599f
C34256 a_1307_43914# a_13565_43940# 0.004697f
C34257 a_8696_44636# a_16759_43396# 1.51e-21
C34258 a_n1917_44484# a_n4318_39768# 6.9e-19
C34259 a_n913_45002# a_3539_42460# 0.359316f
C34260 a_n2017_45002# a_n998_43396# 5.23e-20
C34261 a_n2302_38778# a_n2956_38216# 4.36e-19
C34262 a_5111_44636# VDD 1.28013f
C34263 a_14097_32519# EN_VIN_BSTR_N 0.031973f
C34264 COMP_P CAL_P 0.037476f
C34265 a_18114_32519# a_20202_43084# 1.27e-19
C34266 a_18450_45144# a_12741_44636# 4.86e-19
C34267 a_13720_44458# a_13059_46348# 0.008849f
C34268 a_8375_44464# a_3090_45724# 9.88e-21
C34269 a_1115_44172# a_n2438_43548# 5.77e-19
C34270 a_9159_44484# a_8270_45546# 4.45e-19
C34271 a_5205_44484# a_5066_45546# 1.52e-20
C34272 a_n2661_43370# a_8199_44636# 0.126664f
C34273 a_6125_45348# a_2324_44458# 0.001467f
C34274 a_9028_43914# a_n1613_43370# 2.5e-20
C34275 a_15493_43940# a_13507_46334# 0.021188f
C34276 a_n1352_43396# a_n971_45724# 0.005968f
C34277 a_n229_43646# a_n2497_47436# 0.022782f
C34278 a_5379_42460# a_7174_31319# 3.55e-20
C34279 COMP_P a_1736_39587# 0.007099f
C34280 a_n1630_35242# a_n3565_39590# 0.036902f
C34281 a_13575_42558# a_13333_42558# 3.68e-20
C34282 a_n4318_38216# a_n4334_39392# 1.1e-19
C34283 a_n3674_37592# a_n3420_39616# 0.019754f
C34284 a_n1920_47178# VDD 0.229556f
C34285 DATA[4] CLK 1.11e-19
C34286 a_12549_44172# a_12741_44636# 0.090958f
C34287 a_13661_43548# a_17639_46660# 2.94e-20
C34288 a_20916_46384# a_21363_46634# 0.017401f
C34289 a_8145_46902# a_8023_46660# 3.16e-19
C34290 a_7715_46873# a_8270_45546# 2.04e-19
C34291 a_4955_46873# a_3090_45724# 9.92e-20
C34292 a_19321_45002# a_20731_47026# 3.86e-21
C34293 a_5807_45002# a_18280_46660# 3.71e-20
C34294 a_n881_46662# a_n1991_46122# 0.001102f
C34295 a_n1613_43370# a_n1423_46090# 0.15966f
C34296 a_2487_47570# a_167_45260# 9.29e-23
C34297 a_4883_46098# a_5497_46414# 0.007657f
C34298 a_11599_46634# a_13925_46122# 0.549622f
C34299 a_10227_46804# a_10355_46116# 0.022564f
C34300 a_14311_47204# a_14275_46494# 4.74e-21
C34301 a_13717_47436# a_2324_44458# 1.33e-21
C34302 a_12861_44030# a_14840_46494# 7.53e-20
C34303 a_6151_47436# a_6945_45028# 0.335681f
C34304 a_n1151_42308# a_n1533_46116# 0.002268f
C34305 a_584_46384# a_2981_46116# 6.74e-20
C34306 a_n971_45724# a_5066_45546# 0.045749f
C34307 a_7640_43914# a_7287_43370# 0.001047f
C34308 a_14539_43914# a_14579_43548# 0.002303f
C34309 a_14673_44172# a_n97_42460# 1.2e-19
C34310 a_18184_42460# a_21855_43396# 1.51e-19
C34311 a_1307_43914# a_5534_30871# 3.06e-20
C34312 a_18494_42460# a_4361_42308# 0.061307f
C34313 a_10193_42453# a_11323_42473# 0.034215f
C34314 a_10057_43914# a_10849_43646# 0.003423f
C34315 a_n2293_42834# a_2075_43172# 0.005552f
C34316 a_5891_43370# a_6765_43638# 7.33e-21
C34317 a_2711_45572# a_15143_45578# 0.009403f
C34318 a_n2293_42282# a_n971_45724# 6.84e-19
C34319 a_12429_44172# a_12741_44636# 3.86e-19
C34320 a_15682_43940# a_11415_45002# 6.37e-20
C34321 a_1525_44260# a_1138_42852# 2.28e-20
C34322 a_14543_43071# a_4915_47217# 1.12e-21
C34323 a_5883_43914# a_n443_42852# 8.2e-19
C34324 a_10149_43396# a_n2293_46634# 4e-19
C34325 a_17324_43396# a_13661_43548# 9.28e-20
C34326 a_2982_43646# a_5257_43370# 2.26e-20
C34327 a_7112_43396# a_4646_46812# 0.07278f
C34328 a_19319_43548# a_3090_45724# 1.22e-19
C34329 a_2437_43646# DATA[5] 0.059749f
C34330 a_6123_31319# a_7754_39964# 5.24e-20
C34331 a_5934_30871# a_7754_40130# 0.007046f
C34332 a_n1630_35242# a_3726_37500# 0.001279f
C34333 COMP_P CAL_N 0.008927f
C34334 a_491_47026# a_310_45028# 9.66e-21
C34335 a_6755_46942# a_8049_45260# 0.035035f
C34336 a_171_46873# a_n356_45724# 5.68e-21
C34337 a_n2293_46634# a_1609_45822# 0.036096f
C34338 a_n743_46660# a_7_45899# 0.001065f
C34339 a_n2661_46098# a_n2293_45546# 4.48e-20
C34340 a_14035_46660# a_2324_44458# 2.63e-20
C34341 a_19692_46634# a_21137_46414# 0.242332f
C34342 a_13059_46348# a_13351_46090# 0.074689f
C34343 a_765_45546# a_9823_46155# 1.78e-20
C34344 a_19466_46812# a_6945_45028# 2.92e-19
C34345 a_15227_44166# a_10809_44734# 0.034868f
C34346 a_n2157_46122# a_n1991_46122# 0.614266f
C34347 a_n2293_46098# a_n1423_46090# 0.00572f
C34348 a_18451_43940# a_15743_43084# 0.005843f
C34349 a_458_43396# a_1049_43396# 0.052073f
C34350 a_11341_43940# a_16243_43396# 1.07e-19
C34351 a_15493_43396# a_18525_43370# 0.031354f
C34352 a_453_43940# a_685_42968# 1.15e-21
C34353 a_19006_44850# a_18599_43230# 2.2e-20
C34354 a_n97_42460# a_766_43646# 5.09e-19
C34355 a_11967_42832# a_18817_42826# 6.37e-20
C34356 a_9313_44734# a_10793_43218# 1.08e-19
C34357 en_comp comp_n 0.026896f
C34358 a_n2956_37592# a_n2860_39072# 3.22e-20
C34359 a_4235_43370# VDD 0.229422f
C34360 a_7499_43078# a_8560_45348# 0.006911f
C34361 a_21513_45002# a_2437_43646# 0.009475f
C34362 a_21188_45572# a_21297_45572# 0.007416f
C34363 a_21363_45546# a_21542_45572# 0.007399f
C34364 a_21350_45938# a_3357_43084# 3.05e-19
C34365 a_17324_43396# a_4185_45028# 1.18e-21
C34366 a_13678_32519# a_20820_30879# 0.053259f
C34367 a_13467_32519# a_21076_30879# 0.055522f
C34368 a_22223_43396# a_11415_45002# 2.17e-20
C34369 a_n1736_42282# a_n2442_46660# 4.03e-20
C34370 a_n1329_42308# a_n2956_39768# 3.21e-20
C34371 a_n4318_38216# a_n2312_38680# 0.023247f
C34372 a_2713_42308# a_768_44030# 5.49e-20
C34373 a_5837_42852# a_5257_43370# 4.04e-20
C34374 a_14401_32519# a_13259_45724# 4.2e-20
C34375 a_9145_43396# a_2324_44458# 9.23e-23
C34376 a_10341_43396# a_10903_43370# 0.042836f
C34377 a_12281_43396# a_9290_44172# 0.36475f
C34378 a_14113_42308# a_10227_46804# 0.627404f
C34379 a_n4064_39616# SMPL_ON_P 1.56e-20
C34380 a_8379_46155# VDD 2.18e-20
C34381 a_11136_45572# a_n1151_42308# 3.27e-20
C34382 a_11962_45724# a_11599_46634# 1.79e-20
C34383 a_11823_42460# a_14311_47204# 2.5e-21
C34384 a_7499_43078# a_10227_46804# 0.033512f
C34385 a_13163_45724# a_12861_44030# 0.098707f
C34386 a_13527_45546# a_13717_47436# 3.58e-22
C34387 a_2711_45572# a_2747_46873# 3.81e-20
C34388 a_8034_45724# a_8062_46155# 0.002525f
C34389 a_6945_45028# a_20205_31679# 0.00545f
C34390 a_20708_46348# a_20850_46155# 0.005572f
C34391 a_18579_44172# a_19647_42308# 7.92e-19
C34392 a_8685_43396# a_10796_42968# 9.94e-21
C34393 a_n2661_42282# a_6171_42473# 0.013039f
C34394 a_3422_30871# a_18907_42674# 2.69e-20
C34395 a_1568_43370# a_1793_42852# 0.011559f
C34396 a_3877_44458# DATA[2] 0.001477f
C34397 a_18114_32519# C5_N_btm 1.78e-19
C34398 a_19721_31679# C4_N_btm 9.91e-21
C34399 a_8696_44636# a_17517_44484# 0.001184f
C34400 a_10775_45002# a_n2661_44458# 8.26e-21
C34401 a_1307_43914# a_11691_44458# 0.024289f
C34402 a_15861_45028# a_17061_44734# 2.19e-19
C34403 a_4927_45028# a_4223_44672# 2.44e-19
C34404 a_3537_45260# a_6298_44484# 0.001842f
C34405 a_n1059_45260# a_18248_44752# 2.77e-20
C34406 a_n2661_45010# a_n2012_44484# 1.82e-19
C34407 a_3232_43370# a_949_44458# 1.95e-20
C34408 a_5111_44636# a_n699_43396# 0.016349f
C34409 a_18817_42826# a_13259_45724# 2.9e-20
C34410 a_8037_42858# a_n357_42282# 0.048934f
C34411 a_7765_42852# a_n755_45592# 0.00466f
C34412 a_2711_45572# a_20202_43084# 1.42e-19
C34413 a_13904_45546# a_13885_46660# 8.51e-20
C34414 a_13556_45296# a_12549_44172# 0.030045f
C34415 a_13777_45326# a_12891_46348# 0.03955f
C34416 a_9482_43914# a_768_44030# 0.77718f
C34417 a_327_44734# a_n743_46660# 4e-19
C34418 a_n37_45144# a_n133_46660# 4.9e-21
C34419 a_4574_45260# a_n2661_46634# 1.32e-20
C34420 a_7705_45326# a_5807_45002# 8.49e-21
C34421 a_3065_45002# a_n2293_46634# 0.102991f
C34422 a_413_45260# a_n2438_43548# 0.032468f
C34423 a_2437_43646# a_2162_46660# 0.002257f
C34424 a_n2661_45010# a_n2661_46098# 1.31e-20
C34425 a_375_42282# a_n881_46662# 5.71e-20
C34426 a_n1838_35608# VDD 0.523851f
C34427 a_n1352_44484# a_n971_45724# 0.005662f
C34428 a_n1177_44458# a_n746_45260# 0.064145f
C34429 a_743_42282# a_3581_42558# 7.35e-19
C34430 a_n901_43156# a_n3674_37592# 2e-19
C34431 a_n1423_42826# a_n1630_35242# 2.25e-19
C34432 a_n13_43084# a_n784_42308# 1.77e-19
C34433 a_13460_43230# a_14635_42282# 6.39e-20
C34434 a_14543_43071# a_13291_42460# 0.107887f
C34435 a_10341_43396# a_15959_42545# 3.32e-20
C34436 a_5534_30871# a_13003_42852# 0.001789f
C34437 a_n2293_42282# a_3863_42891# 1.73e-19
C34438 a_4361_42308# a_3318_42354# 8.57e-20
C34439 a_n1379_43218# COMP_P 1.55e-21
C34440 a_10809_44734# EN_OFFSET_CAL 0.035912f
C34441 a_n3690_39392# VDD 0.363068f
C34442 a_4915_47217# a_7989_47542# 9.72e-19
C34443 a_5815_47464# a_n1613_43370# 0.360237f
C34444 a_18479_47436# a_19386_47436# 0.219411f
C34445 a_18780_47178# a_18597_46090# 0.175179f
C34446 a_16763_47508# a_13507_46334# 8.88e-21
C34447 a_16327_47482# a_4883_46098# 0.096832f
C34448 a_10227_46804# a_20894_47436# 0.010908f
C34449 a_n443_46116# a_4842_47243# 0.001129f
C34450 a_4791_45118# a_5159_47243# 0.00545f
C34451 a_n1435_47204# a_n89_47570# 2.3e-21
C34452 a_15673_47210# a_12465_44636# 6.52e-19
C34453 a_n2288_47178# a_n2956_39768# 0.001146f
C34454 a_n2497_47436# a_n2661_46634# 0.079801f
C34455 a_n2833_47464# a_n2472_46634# 0.001084f
C34456 a_n1151_42308# a_12891_46348# 0.038292f
C34457 a_2905_45572# a_768_44030# 0.02789f
C34458 a_9482_43914# a_13483_43940# 0.006325f
C34459 a_18374_44850# a_9313_44734# 3.42e-21
C34460 a_12607_44458# a_n2293_43922# 0.078602f
C34461 a_11691_44458# a_18579_44172# 2.18e-19
C34462 a_n2293_42834# a_5013_44260# 3.56e-20
C34463 a_1307_43914# a_8333_44056# 0.006875f
C34464 a_11823_42460# a_13667_43396# 0.107673f
C34465 a_7499_43078# a_8873_43396# 0.001075f
C34466 a_8746_45002# a_10341_43396# 0.002313f
C34467 a_18494_42460# a_20397_44484# 3.54e-19
C34468 a_11827_44484# a_19789_44512# 4.59e-19
C34469 a_3232_43370# a_11341_43940# 0.112367f
C34470 a_16147_45260# VDD 0.197706f
C34471 a_18083_42858# RST_Z 1.06e-20
C34472 a_2437_43646# a_10809_44734# 0.13907f
C34473 a_n1059_45260# a_2324_44458# 4.3e-20
C34474 a_3537_45260# a_5937_45572# 9.77e-19
C34475 a_413_45260# a_11133_46155# 1.62e-21
C34476 a_3357_43084# a_21137_46414# 1.6e-20
C34477 a_22223_45572# a_22223_46124# 0.025171f
C34478 a_12649_45572# a_10586_45546# 6.62e-20
C34479 a_14033_45822# a_13259_45724# 0.004141f
C34480 a_17801_45144# a_3090_45724# 7.84e-20
C34481 a_20362_44736# a_12549_44172# 0.015111f
C34482 a_21359_45002# a_19692_46634# 7.78e-21
C34483 a_8191_45002# a_3483_46348# 0.081038f
C34484 a_11827_44484# a_19466_46812# 1.45e-20
C34485 a_n2661_43370# a_765_45546# 6.55e-22
C34486 a_196_42282# a_5742_30871# 7.34e-20
C34487 a_2713_42308# a_6123_31319# 1.31e-20
C34488 a_5379_42460# a_5932_42308# 0.761308f
C34489 a_1606_42308# a_8325_42308# 1.94e-20
C34490 a_n784_42308# a_11323_42473# 1.56e-20
C34491 a_13887_32519# C5_N_btm 1.01e-19
C34492 a_17364_32525# C1_N_btm 9.59e-21
C34493 a_3080_42308# a_6886_37412# 6.84e-19
C34494 CAL_P a_22705_37990# 1.58e-20
C34495 a_22609_38406# a_22609_37990# 0.32625f
C34496 a_12465_44636# a_16388_46812# 7.04e-20
C34497 a_18597_46090# a_18285_46348# 0.012666f
C34498 a_18479_47436# a_19551_46910# 0.001789f
C34499 a_10227_46804# a_20411_46873# 0.013631f
C34500 a_2063_45854# a_2202_46116# 0.026352f
C34501 a_584_46384# a_167_45260# 0.0321f
C34502 a_n971_45724# a_5068_46348# 3.37e-21
C34503 a_n237_47217# a_4419_46090# 0.049065f
C34504 a_n881_46662# a_15227_44166# 1.74e-19
C34505 a_n2661_46634# a_6682_46987# 4.03e-19
C34506 a_5807_45002# a_8601_46660# 1.44e-19
C34507 a_3524_46660# a_4651_46660# 1.59e-19
C34508 a_3699_46634# a_4955_46873# 2.52e-20
C34509 a_n743_46660# a_10150_46912# 4e-20
C34510 a_12549_44172# a_13607_46688# 0.013421f
C34511 a_2107_46812# a_5257_43370# 0.039927f
C34512 a_895_43940# a_2675_43914# 0.099822f
C34513 a_n2065_43946# a_n1644_44306# 0.090164f
C34514 a_n1761_44111# a_n3674_39768# 7.14e-19
C34515 a_2127_44172# a_2998_44172# 0.001419f
C34516 a_2479_44172# a_2889_44172# 0.002826f
C34517 a_17517_44484# a_20365_43914# 4.82e-21
C34518 a_11967_42832# a_15682_43940# 1.63211f
C34519 a_4223_44672# a_4699_43561# 2.12e-19
C34520 a_10193_42453# a_20753_42852# 0.082713f
C34521 a_n1059_45260# a_8387_43230# 0.005946f
C34522 a_n2017_45002# a_9127_43156# 3.46e-19
C34523 a_n913_45002# a_8605_42826# 0.019641f
C34524 a_10334_44484# VDD 0.19332f
C34525 a_n4064_40160# C10_P_btm 0.460005f
C34526 a_n4064_39616# a_n1532_35090# 1.21e-19
C34527 a_n3420_39616# EN_VIN_BSTR_P 0.06758f
C34528 a_22775_42308# RST_Z 0.001998f
C34529 a_20512_43084# a_11415_45002# 0.001234f
C34530 a_n2012_43396# a_n2438_43548# 0.003029f
C34531 a_10949_43914# a_3090_45724# 0.001234f
C34532 a_6031_43396# a_768_44030# 3.88e-20
C34533 a_8103_44636# a_8049_45260# 0.012205f
C34534 a_6655_43762# a_n881_46662# 2.11e-20
C34535 a_n2293_43922# a_10903_43370# 0.029114f
C34536 a_9313_44734# a_17715_44484# 6.46e-20
C34537 a_n2661_43922# a_12005_46116# 2.87e-22
C34538 a_14579_43548# a_11453_44696# 1.66e-22
C34539 a_10341_43396# a_4883_46098# 4.87e-19
C34540 a_15781_43660# a_10227_46804# 0.002214f
C34541 a_16243_43396# a_16327_47482# 0.295263f
C34542 a_18783_43370# a_12861_44030# 2.29e-20
C34543 a_n1423_42826# a_n971_45724# 1.4e-20
C34544 a_n1021_46688# VDD 0.226043f
C34545 a_6123_31319# C8_N_btm 6.73e-20
C34546 a_5934_30871# C6_N_btm 0.004563f
C34547 a_18285_46348# a_19123_46287# 0.007333f
C34548 a_n1925_46634# a_8034_45724# 0.206805f
C34549 a_12549_44172# a_16375_45002# 0.001412f
C34550 a_5807_45002# a_14371_46494# 0.002046f
C34551 a_10249_46116# a_9625_46129# 0.009289f
C34552 a_6755_46942# a_8953_45546# 0.001323f
C34553 a_10428_46928# a_9290_44172# 1.43e-19
C34554 a_10467_46802# a_10355_46116# 0.008762f
C34555 a_6969_46634# a_5937_45572# 0.001066f
C34556 a_18374_44850# a_18599_43230# 1.49e-21
C34557 a_18989_43940# a_18817_42826# 2.61e-19
C34558 a_20679_44626# a_13467_32519# 4.42e-21
C34559 a_9028_43914# a_8791_43396# 0.001013f
C34560 a_5891_43370# a_10341_42308# 2.08e-19
C34561 a_18579_44172# a_4190_30871# 0.052036f
C34562 a_n2661_43922# a_3935_42891# 1.92e-21
C34563 a_9313_44734# a_10083_42826# 0.013808f
C34564 a_n2293_43922# a_3681_42891# 7.77e-21
C34565 a_n356_44636# a_16795_42852# 8.61e-19
C34566 a_n2293_42834# a_196_42282# 5.62e-20
C34567 a_19328_44172# a_3626_43646# 2.27e-20
C34568 a_n2661_43370# a_n4318_38216# 0.002734f
C34569 a_n2017_45002# a_17124_42282# 0.002905f
C34570 a_16680_45572# a_18596_45572# 3.21e-21
C34571 a_2711_45572# a_13017_45260# 0.050114f
C34572 a_7227_45028# a_7276_45260# 0.098279f
C34573 a_6667_45809# a_6709_45028# 0.001946f
C34574 a_4880_45572# a_4558_45348# 3.7e-19
C34575 a_6511_45714# a_7705_45326# 8.07e-19
C34576 a_5421_42558# a_4791_45118# 0.00311f
C34577 a_22521_40599# a_22609_37990# 0.021352f
C34578 a_22469_40625# a_22705_38406# 1.29e-19
C34579 a_n4209_37414# C4_P_btm 9.91e-21
C34580 a_n3565_37414# C6_P_btm 1.26e-20
C34581 a_3726_37500# a_11530_34132# 3.03e-19
C34582 a_5700_37509# a_n923_35174# 3.61e-19
C34583 a_22765_42852# a_13507_46334# 0.003797f
C34584 a_n97_42460# a_10903_43370# 0.021999f
C34585 a_261_44278# a_n863_45724# 9.97e-19
C34586 a_15682_43940# a_13259_45724# 9.31e-21
C34587 a_2889_44172# a_n443_42852# 1.05e-20
C34588 a_9290_44172# VDD 2.74561f
C34589 a_3775_45552# a_n971_45724# 0.091275f
C34590 a_6598_45938# a_n237_47217# 2.15e-19
C34591 a_2711_45572# a_2063_45854# 0.185507f
C34592 a_8953_45546# a_8049_45260# 0.156816f
C34593 a_10809_44734# a_22959_46124# 0.172346f
C34594 a_8016_46348# a_8062_46155# 0.006879f
C34595 a_7920_46348# a_8379_46155# 6.64e-19
C34596 a_2324_44458# a_n1925_42282# 0.018757f
C34597 a_8199_44636# a_9823_46482# 1.73e-22
C34598 a_n3565_38502# a_n3690_37440# 4.13e-19
C34599 a_n4209_38502# a_n2946_37690# 3.29e-19
C34600 a_n3420_38528# a_n4334_37440# 1.39e-19
C34601 a_2684_37794# VDAC_Ni 0.004723f
C34602 a_n3565_39304# VDAC_P 9.25e-19
C34603 a_n1549_44318# a_n1630_35242# 5.92e-22
C34604 a_6197_43396# a_4361_42308# 4.64e-20
C34605 a_8147_43396# a_743_42282# 2.1e-21
C34606 a_10341_43396# a_16243_43396# 0.058241f
C34607 a_n1557_42282# a_n1641_43230# 7.08e-19
C34608 a_13565_43940# a_13635_43156# 7.88e-21
C34609 a_12281_43396# a_13749_43396# 1.13e-20
C34610 a_8685_43396# a_15125_43396# 8.47e-19
C34611 a_n1761_44111# a_1184_42692# 5.67e-20
C34612 a_12549_44172# RST_Z 9.94e-19
C34613 a_791_42968# VDD 0.128737f
C34614 a_n2810_45028# a_n2302_37984# 0.003394f
C34615 a_n2956_37592# a_n4064_37984# 0.012393f
C34616 a_11322_45546# a_n2661_42834# 4.07e-19
C34617 a_16115_45572# a_14539_43914# 4.47e-19
C34618 a_8696_44636# a_13720_44458# 0.004063f
C34619 a_1307_43914# a_375_42282# 1.11e-20
C34620 a_22223_45572# a_22223_45036# 0.026152f
C34621 a_2382_45260# a_n2661_43370# 0.03415f
C34622 a_3357_43084# a_21359_45002# 6.53e-21
C34623 a_19479_31679# a_11827_44484# 0.01397f
C34624 a_6171_45002# a_6945_45348# 1.2e-19
C34625 a_5193_42852# a_4185_45028# 2.2e-19
C34626 a_18525_43370# a_n357_42282# 3.71e-20
C34627 a_9127_43156# a_526_44458# 0.054699f
C34628 a_14621_43646# a_n443_42852# 0.001398f
C34629 a_375_42282# a_n443_46116# 0.001544f
C34630 a_3495_45348# a_2905_45572# 3.62e-20
C34631 a_413_45260# a_13507_46334# 3.41e-19
C34632 en_comp SMPL_ON_N 8.94e-19
C34633 a_2437_43646# a_n881_46662# 0.084076f
C34634 a_16789_45572# a_5807_45002# 1.08e-19
C34635 a_18596_45572# a_13747_46662# 0.01625f
C34636 a_8746_45002# a_8667_46634# 4.9e-22
C34637 a_19431_45546# a_19321_45002# 0.029441f
C34638 a_6812_45938# a_6755_46942# 2.21e-20
C34639 a_18799_45938# a_13661_43548# 0.004963f
C34640 a_10053_45546# a_10150_46912# 1.88e-20
C34641 a_10180_45724# a_9863_46634# 1.87e-19
C34642 a_1609_45822# a_2277_45546# 2.47e-20
C34643 a_6197_43396# a_6761_42308# 1.61e-19
C34644 a_6031_43396# a_6123_31319# 6.63e-20
C34645 a_13635_43156# a_5534_30871# 0.078849f
C34646 a_13460_43230# a_14543_43071# 0.001783f
C34647 a_n97_42460# a_15959_42545# 0.005005f
C34648 a_2982_43646# a_9223_42460# 1.29e-19
C34649 a_3626_43646# a_8685_42308# 0.002659f
C34650 a_791_42968# a_873_42968# 0.004937f
C34651 a_16823_43084# a_16877_43172# 0.001729f
C34652 a_15743_43084# a_19273_43230# 0.001058f
C34653 a_4520_42826# a_n2293_42282# 3.87e-20
C34654 a_21076_30879# VCM 0.097317f
C34655 a_17730_32519# C3_N_btm 5.52e-20
C34656 a_19237_31679# C1_N_btm 0.001047f
C34657 a_15051_42282# VDD 0.461307f
C34658 a_1431_47204# a_n1435_47204# 0.001005f
C34659 a_n443_46116# a_5129_47502# 0.10632f
C34660 a_4791_45118# a_5815_47464# 0.003581f
C34661 a_n1151_42308# a_7903_47542# 8.5e-20
C34662 a_2063_45854# a_9313_45822# 0.042979f
C34663 a_18175_45572# a_15493_43940# 6.32e-22
C34664 a_5518_44484# a_5883_43914# 5.07e-20
C34665 a_6298_44484# a_8701_44490# 2.01e-20
C34666 a_3065_45002# a_2675_43914# 8.4e-22
C34667 a_2382_45260# a_2998_44172# 0.045272f
C34668 a_3357_43084# a_n2661_42282# 0.028477f
C34669 a_n2956_37592# a_n3674_39768# 0.024317f
C34670 a_n2293_45010# a_261_44278# 1.74e-19
C34671 en_comp a_n4318_39768# 2e-19
C34672 a_961_42354# a_n755_45592# 0.01273f
C34673 a_2351_42308# a_n863_45724# 0.038802f
C34674 a_9049_44484# VDD 0.680993f
C34675 a_20447_31679# a_22959_46660# 3.72e-20
C34676 a_n2661_43370# a_10623_46897# 6.28e-21
C34677 a_1307_43914# a_15227_44166# 0.059667f
C34678 a_14539_43914# a_5807_45002# 0.066683f
C34679 a_6298_44484# a_n2293_46634# 1.21e-19
C34680 a_16112_44458# a_13661_43548# 0.053099f
C34681 a_7499_43078# a_8034_45724# 0.001227f
C34682 a_6812_45938# a_8049_45260# 2.61e-19
C34683 a_413_45260# a_20623_46660# 2.82e-20
C34684 a_15599_45572# a_2324_44458# 0.042604f
C34685 a_8696_44636# a_13351_46090# 5.82e-22
C34686 a_n2661_42834# a_12465_44636# 7.41e-19
C34687 a_13468_44734# a_13507_46334# 1.04e-19
C34688 a_n1549_44318# a_n971_45724# 0.00442f
C34689 a_18083_42858# a_17303_42282# 7.17e-20
C34690 a_n2104_42282# a_n4318_37592# 0.033328f
C34691 a_17701_42308# a_17531_42308# 0.109201f
C34692 a_n3674_39304# a_n3420_39072# 0.065079f
C34693 a_n4318_38216# COMP_P 5.3e-20
C34694 a_n3674_38216# a_n1736_42282# 7.03e-19
C34695 a_9114_42852# a_5934_30871# 5.71e-20
C34696 a_5807_45002# a_2107_46812# 1.5594f
C34697 a_768_44030# a_2443_46660# 2.94e-19
C34698 a_n2661_46634# a_n2104_46634# 0.030211f
C34699 a_n2472_46634# a_n2293_46634# 0.163804f
C34700 a_n2956_39768# a_n2312_38680# 0.076511f
C34701 a_n2840_46634# a_n1925_46634# 5.18e-19
C34702 a_n1613_43370# a_3055_46660# 9.54e-19
C34703 a_4883_46098# a_8667_46634# 2.2e-19
C34704 a_n1435_47204# a_11735_46660# 7.87e-20
C34705 a_n1151_42308# a_12359_47026# 0.002059f
C34706 a_n2497_47436# a_765_45546# 1.79e-20
C34707 a_8975_43940# a_11341_43940# 1.83e-19
C34708 a_18287_44626# a_18079_43940# 0.007509f
C34709 a_18248_44752# a_18326_43940# 7.79e-19
C34710 a_11967_42832# a_20512_43084# 0.106819f
C34711 a_20679_44626# a_22315_44484# 7.27e-21
C34712 a_20835_44721# a_3422_30871# 2.09e-19
C34713 a_n2661_42834# a_7281_43914# 0.010117f
C34714 a_n2293_42834# a_4699_43561# 3.68e-20
C34715 a_20362_44736# a_20637_44484# 0.007416f
C34716 a_5883_43914# a_9895_44260# 2.92e-19
C34717 a_6109_44484# a_6101_44260# 1.75e-20
C34718 a_8953_45002# a_9803_43646# 2.76e-20
C34719 a_3232_43370# a_10341_43396# 2.1e-19
C34720 a_n2017_45002# a_19268_43646# 4.82e-21
C34721 a_n913_45002# a_18783_43370# 2.32e-21
C34722 a_n1059_45260# a_15743_43084# 0.101833f
C34723 a_6123_31319# C2_P_btm 0.01106f
C34724 a_5934_30871# C4_P_btm 0.030578f
C34725 a_3626_43646# a_12861_44030# 3.03e-20
C34726 a_n97_42460# a_4883_46098# 1.42e-20
C34727 a_n4318_39304# a_n2312_39304# 0.023404f
C34728 a_10157_44484# a_8016_46348# 0.016596f
C34729 a_8701_44490# a_5937_45572# 0.022661f
C34730 a_5883_43914# a_8199_44636# 7.86e-19
C34731 a_3537_45260# a_n443_42852# 0.567413f
C34732 a_18579_44172# a_15227_44166# 9.13e-21
C34733 a_6671_43940# a_768_44030# 1.23e-19
C34734 a_19279_43940# a_19692_46634# 8.61e-20
C34735 a_5205_44734# a_n2293_46098# 5.05e-20
C34736 a_16979_44734# a_3483_46348# 0.173123f
C34737 a_n356_44636# a_376_46348# 3.01e-22
C34738 a_20990_47178# VDD 0.210484f
C34739 a_18907_42674# a_7174_31319# 2.21e-20
C34740 a_5742_30871# a_n3420_39072# 0.005978f
C34741 a_17303_42282# a_22775_42308# 0.005701f
C34742 a_18548_42308# a_19511_42282# 3.36e-20
C34743 a_n743_46660# a_6419_46155# 0.00636f
C34744 a_5807_45002# a_14493_46090# 0.006666f
C34745 a_n2661_46634# a_9569_46155# 8.52e-20
C34746 a_n1925_46634# a_8016_46348# 0.014574f
C34747 a_13747_46662# a_13759_46122# 0.02887f
C34748 a_n2293_46634# a_5937_45572# 2.05e-19
C34749 a_13661_43548# a_13925_46122# 2.91e-21
C34750 a_12549_44172# a_18985_46122# 1.04e-20
C34751 a_n1613_43370# a_n2956_39304# 4.39e-21
C34752 a_4883_46098# a_6640_46482# 2.25e-19
C34753 a_18780_47178# a_8049_45260# 2.82e-21
C34754 a_11599_46634# a_12638_46436# 0.006285f
C34755 a_n971_45724# a_3218_45724# 2.69e-19
C34756 a_n785_47204# a_n755_45592# 1.12e-20
C34757 a_n237_47217# a_1848_45724# 0.232571f
C34758 a_327_47204# a_n357_42282# 1.62e-22
C34759 a_584_46384# a_n863_45724# 0.051089f
C34760 a_17609_46634# a_15227_44166# 0.04317f
C34761 a_11735_46660# a_13885_46660# 5.87e-21
C34762 a_12251_46660# a_12347_46660# 0.013793f
C34763 a_12469_46902# a_12513_46660# 3.69e-19
C34764 a_11901_46660# a_12925_46660# 2.36e-20
C34765 a_6682_46987# a_765_45546# 3.8e-19
C34766 a_1799_45572# a_1823_45246# 0.003001f
C34767 a_n2661_46098# a_1138_42852# 0.020229f
C34768 a_2107_46812# a_3699_46348# 0.00528f
C34769 a_2779_44458# a_2075_43172# 1.85e-20
C34770 a_n809_44244# a_n1557_42282# 1.48e-21
C34771 a_2127_44172# a_1568_43370# 3.06e-19
C34772 a_5663_43940# a_n97_42460# 9.61e-20
C34773 a_22223_43948# a_14021_43940# 2.65e-20
C34774 a_895_43940# a_1209_43370# 9.02e-21
C34775 a_n699_43396# a_791_42968# 6.37e-19
C34776 a_11691_44458# a_13635_43156# 2.7e-21
C34777 a_742_44458# a_3681_42891# 4.15e-19
C34778 a_1414_42308# a_4093_43548# 6.35e-21
C34779 a_18184_42460# a_17701_42308# 0.001244f
C34780 a_1307_43914# a_14635_42282# 3.78e-20
C34781 a_16922_45042# a_19987_42826# 0.00105f
C34782 a_n2293_42834# a_6101_43172# 2.77e-19
C34783 a_n1059_45260# a_1606_42308# 0.008752f
C34784 a_n2017_45002# a_1755_42282# 0.012188f
C34785 a_n913_45002# a_1221_42558# 1.43e-20
C34786 a_3905_42865# VDD 0.788273f
C34787 a_14495_45572# a_15037_45618# 0.00244f
C34788 a_11823_42460# a_16333_45814# 1.07e-20
C34789 a_11525_45546# a_8696_44636# 2.88e-21
C34790 a_10193_42453# a_16223_45938# 1.24e-19
C34791 a_8120_45572# a_8192_45572# 0.003395f
C34792 a_5745_43940# a_1823_45246# 9.33e-20
C34793 a_14401_32519# a_20202_43084# 9.39e-20
C34794 a_10796_42968# a_768_44030# 2.7e-22
C34795 a_20512_43084# a_13259_45724# 1.37e-20
C34796 a_17737_43940# a_17715_44484# 0.289085f
C34797 a_20273_46660# VDD 0.247553f
C34798 a_4958_30871# a_7754_38470# 9.47e-20
C34799 a_n4209_39590# a_n3420_37984# 0.032713f
C34800 a_n4064_40160# a_n4251_38304# 0.001069f
C34801 a_n2472_46090# a_n2956_38680# 0.157373f
C34802 a_n2293_46098# a_n2956_39304# 0.001354f
C34803 a_18285_46348# a_8049_45260# 3.95e-19
C34804 a_14035_46660# a_12839_46116# 3.7e-20
C34805 a_15227_44166# a_19443_46116# 7.48e-19
C34806 a_13059_46348# a_12005_46436# 1.79e-21
C34807 a_2698_46116# a_2324_44458# 5.34e-22
C34808 a_5937_45572# a_9625_46129# 1.78e-19
C34809 a_8199_44636# a_9569_46155# 1.7e-19
C34810 a_10807_43548# a_10341_42308# 0.099222f
C34811 a_n97_42460# a_16243_43396# 0.004882f
C34812 a_11967_42832# a_16245_42852# 0.002841f
C34813 a_10949_43914# a_12379_42858# 3.5e-20
C34814 a_n2661_42834# a_564_42282# 1.13e-20
C34815 a_6197_43396# a_7274_43762# 1.46e-19
C34816 a_4915_47217# DATA[5] 0.121371f
C34817 a_5815_47464# DATA[3] 0.00149f
C34818 a_20447_31679# C10_N_btm 2.25e-20
C34819 a_11682_45822# a_11691_44458# 2.81e-20
C34820 a_7230_45938# a_6298_44484# 3.58e-20
C34821 a_2711_45572# a_18374_44850# 5.8e-21
C34822 a_15903_45785# a_16501_45348# 2.45e-20
C34823 a_2437_43646# a_1307_43914# 0.160142f
C34824 a_3065_45002# a_3429_45260# 0.037292f
C34825 a_2680_45002# a_3537_45260# 8.13e-20
C34826 a_n4064_40160# a_n2312_40392# 0.103899f
C34827 a_n4334_40480# a_n2312_39304# 2.31e-19
C34828 a_n144_43396# a_n863_45724# 1.49e-19
C34829 a_2982_43646# a_n755_45592# 0.221452f
C34830 a_1049_43396# a_n443_42852# 0.047375f
C34831 a_17303_42282# a_12549_44172# 4.74e-21
C34832 a_5379_42460# a_4646_46812# 1.84e-21
C34833 a_18817_42826# a_20202_43084# 1.4e-20
C34834 a_n89_45572# VDD 0.001196f
C34835 a_6511_45714# a_2107_46812# 3.47e-20
C34836 a_16115_45572# a_11453_44696# 1.16e-20
C34837 a_18341_45572# a_16327_47482# 0.04767f
C34838 a_18596_45572# a_11599_46634# 0.01377f
C34839 a_16377_45572# a_10227_46804# 1.61e-19
C34840 a_2437_43646# a_n443_46116# 0.410719f
C34841 a_n967_45348# a_n746_45260# 0.028689f
C34842 a_2382_45260# a_n2497_47436# 0.042349f
C34843 a_n2293_45010# a_584_46384# 0.02901f
C34844 a_413_45260# a_n1741_47186# 0.026099f
C34845 a_n659_45366# a_n971_45724# 3.11e-21
C34846 a_3357_43084# a_4007_47204# 1.6e-20
C34847 a_n1177_43370# a_n1630_35242# 5.63e-22
C34848 a_n97_42460# a_n327_42558# 0.020924f
C34849 a_19268_43646# a_19164_43230# 3.42e-20
C34850 a_19700_43370# a_19339_43156# 0.012115f
C34851 a_15743_43084# a_19987_42826# 0.008026f
C34852 a_5649_42852# a_10835_43094# 1.19e-20
C34853 a_4361_42308# a_10922_42852# 4.19e-20
C34854 a_743_42282# a_13113_42826# 3.77e-20
C34855 a_16823_43084# a_5342_30871# 3.63e-37
C34856 a_15493_43940# a_15486_42560# 4.05e-19
C34857 a_11341_43940# a_15803_42450# 1.77e-21
C34858 a_n447_43370# a_n3674_37592# 2.26e-21
C34859 a_n2302_37984# a_n2302_37690# 0.050477f
C34860 VDAC_Pi a_3754_38470# 0.389564f
C34861 a_7754_40130# a_8530_39574# 0.013981f
C34862 a_n961_42308# VDD 0.24416f
C34863 a_11827_44484# a_20193_45348# 0.051742f
C34864 a_n2661_43370# a_5343_44458# 7.17e-19
C34865 a_10193_42453# a_11341_43940# 0.082222f
C34866 a_11823_42460# a_15493_43396# 2.38e-20
C34867 a_6171_45002# a_n2661_43922# 0.020767f
C34868 a_3357_43084# a_19279_43940# 1.53e-20
C34869 a_3232_43370# a_n2293_43922# 9.68e-21
C34870 a_22775_42308# a_20820_30879# 5.97e-21
C34871 a_1755_42282# a_526_44458# 0.006616f
C34872 a_7309_42852# a_n357_42282# 0.016177f
C34873 a_16245_42852# a_13259_45724# 2.29e-20
C34874 a_1606_42308# a_n1925_42282# 0.065478f
C34875 a_11551_42558# a_9290_44172# 0.123803f
C34876 a_5891_43370# a_n1151_42308# 9.29e-22
C34877 a_5205_44734# a_4791_45118# 0.001884f
C34878 a_17767_44458# a_12861_44030# 2.43e-19
C34879 a_n2661_44458# a_n2312_39304# 1.84e-20
C34880 a_7230_45938# a_5937_45572# 7.84e-20
C34881 a_2711_45572# a_17715_44484# 0.009119f
C34882 a_8568_45546# a_8349_46414# 0.001282f
C34883 a_7499_43078# a_8016_46348# 7.22e-19
C34884 a_8162_45546# a_8199_44636# 0.119979f
C34885 a_7276_45260# a_7715_46873# 4.09e-20
C34886 a_7229_43940# a_7411_46660# 3.82e-19
C34887 a_3357_43084# a_15368_46634# 5.03e-20
C34888 a_13807_45067# a_13661_43548# 4.93e-20
C34889 a_n2293_42834# a_n743_46660# 6.42e-20
C34890 a_n2661_43370# a_n2956_39768# 1.14e-19
C34891 a_14309_45028# a_5807_45002# 0.003656f
C34892 a_19778_44110# a_12549_44172# 0.294084f
C34893 a_11823_42460# a_3483_46348# 0.377948f
C34894 a_21855_43396# a_17303_42282# 1.3e-20
C34895 a_8037_42858# a_8685_42308# 3.44e-20
C34896 a_8605_42826# a_8325_42308# 2.47e-19
C34897 a_n2293_42282# a_564_42282# 4.89e-19
C34898 a_4361_42308# a_17531_42308# 0.007428f
C34899 a_13678_32519# a_4958_30871# 0.031033f
C34900 a_743_42282# a_18214_42558# 0.005672f
C34901 a_4190_30871# a_18310_42308# 0.001467f
C34902 a_17538_32519# C3_N_btm 2.76e-20
C34903 a_14401_32519# C5_N_btm 0.001006f
C34904 a_n881_46662# a_7989_47542# 2.79e-20
C34905 a_12465_44636# a_19321_45002# 4.94e-19
C34906 a_11453_44696# a_5807_45002# 0.050036f
C34907 a_13507_46334# a_20916_46384# 0.123008f
C34908 a_21177_47436# a_21588_30879# 3.24e-19
C34909 a_n971_45724# a_7577_46660# 0.523694f
C34910 a_n1741_47186# a_9863_46634# 4.44e-20
C34911 a_n1151_42308# a_4817_46660# 0.029921f
C34912 a_4007_47204# a_3877_44458# 0.002042f
C34913 a_n237_47217# a_7411_46660# 0.033907f
C34914 a_n443_46116# a_3686_47026# 4.1e-19
C34915 a_2063_45854# a_6540_46812# 1.36e-19
C34916 a_17719_45144# a_17737_43940# 2.8e-20
C34917 a_4223_44672# a_5244_44056# 0.019617f
C34918 a_15861_45028# a_16409_43396# 2.62e-21
C34919 a_8696_44636# a_16977_43638# 6.12e-20
C34920 a_1307_43914# a_11257_43940# 7.05e-19
C34921 a_n1699_44726# a_n4318_39768# 3.3e-19
C34922 a_3232_43370# a_n97_42460# 0.113391f
C34923 a_n913_45002# a_3626_43646# 0.104422f
C34924 a_n1059_45260# a_3539_42460# 0.021504f
C34925 a_2382_45260# a_1568_43370# 2.74e-21
C34926 a_n2017_45002# a_n1243_43396# 6.69e-20
C34927 a_3357_43084# a_7112_43396# 2.88e-19
C34928 a_n4064_38528# a_n2956_38216# 3.3e-20
C34929 a_5147_45002# VDD 0.574918f
C34930 a_14097_32519# a_11530_34132# 0.002965f
C34931 a_17969_45144# a_12741_44636# 3.55e-19
C34932 a_13076_44458# a_13059_46348# 7.55e-19
C34933 a_644_44056# a_n2438_43548# 4.81e-19
C34934 a_7640_43914# a_3090_45724# 0.020595f
C34935 a_2479_44172# a_n2293_46634# 0.00465f
C34936 a_8704_45028# a_5937_45572# 0.010036f
C34937 a_5837_45348# a_2324_44458# 3.04e-19
C34938 a_8333_44056# a_n1613_43370# 1.05e-20
C34939 a_22223_43948# a_13507_46334# 0.00424f
C34940 a_n1177_43370# a_n971_45724# 0.014733f
C34941 a_5267_42460# a_7174_31319# 4.88e-21
C34942 COMP_P a_1239_39587# 0.388733f
C34943 a_13070_42354# a_13333_42558# 0.011552f
C34944 a_13575_42558# a_13249_42558# 2.37e-20
C34945 a_6123_31319# a_4958_30871# 0.021709f
C34946 a_n2109_47186# VDD 2.71791f
C34947 a_12891_46348# a_12741_44636# 0.038901f
C34948 a_20916_46384# a_20623_46660# 9.66e-19
C34949 a_10249_46116# a_6755_46942# 0.068878f
C34950 a_7411_46660# a_8270_45546# 1.1e-19
C34951 a_19321_45002# a_20528_46660# 3.62e-19
C34952 a_8145_46902# a_8654_47026# 2.6e-19
C34953 a_7577_46660# a_8023_46660# 2.28e-19
C34954 a_5807_45002# a_17639_46660# 4.64e-19
C34955 a_4651_46660# a_3090_45724# 9.87e-21
C34956 a_n881_46662# a_n1853_46287# 0.229188f
C34957 a_n1613_43370# a_n1991_46122# 0.031697f
C34958 SMPL_ON_N a_4185_45028# 3.43e-19
C34959 a_5649_42852# a_7754_40130# 6.15e-19
C34960 a_4883_46098# a_5204_45822# 0.041898f
C34961 a_14955_47212# a_13925_46122# 4.01e-20
C34962 a_11599_46634# a_13759_46122# 0.262969f
C34963 a_10227_46804# a_9823_46155# 0.004734f
C34964 a_12861_44030# a_15015_46420# 7.95e-20
C34965 a_13717_47436# a_14840_46494# 2.21e-21
C34966 a_4915_47217# a_10809_44734# 0.037616f
C34967 a_5815_47464# a_6945_45028# 9.9e-19
C34968 a_584_46384# a_1431_46436# 3.89e-19
C34969 a_18494_42460# a_13467_32519# 1.67e-19
C34970 a_8975_43940# a_10341_43396# 5.7e-20
C34971 a_7499_43078# a_11633_42558# 2.79e-19
C34972 a_5891_43370# a_6197_43396# 0.003102f
C34973 a_18184_42460# a_4361_42308# 0.058569f
C34974 a_1307_43914# a_14543_43071# 7.06e-21
C34975 a_n2293_42834# a_1847_42826# 0.078127f
C34976 a_n2293_43922# a_4905_42826# 2.78e-20
C34977 a_10193_42453# a_10723_42308# 0.046812f
C34978 a_10057_43914# a_10765_43646# 0.005404f
C34979 a_n1059_45260# a_9061_43230# 1.7e-20
C34980 a_n4209_38216# VIN_P 0.029185f
C34981 a_2711_45572# a_14495_45572# 0.008699f
C34982 a_16979_44734# a_n357_42282# 5e-21
C34983 a_8701_44490# a_n443_42852# 2.96e-20
C34984 a_9885_43396# a_n2293_46634# 1.99e-19
C34985 a_15301_44260# a_13059_46348# 1e-19
C34986 a_17499_43370# a_13661_43548# 8.74e-19
C34987 a_7287_43370# a_4646_46812# 0.07176f
C34988 a_1241_44260# a_1138_42852# 6.56e-19
C34989 a_2437_43646# DATA[4] 0.060047f
C34990 a_1606_42308# a_n3420_37440# 0.001369f
C34991 COMP_P a_11206_38545# 0.002821f
C34992 a_13059_46348# a_12594_46348# 0.03479f
C34993 a_19692_46634# a_20708_46348# 0.318388f
C34994 a_765_45546# a_9569_46155# 2.88e-20
C34995 a_14513_46634# a_14275_46494# 0.001809f
C34996 a_19333_46634# a_6945_45028# 9.77e-20
C34997 a_18834_46812# a_10809_44734# 0.006086f
C34998 a_15227_44166# a_22223_46124# 0.002009f
C34999 a_14035_46660# a_14840_46494# 5.47e-21
C35000 a_2107_46812# a_n755_45592# 4.66e-20
C35001 a_n2293_46634# a_n443_42852# 2.09483f
C35002 a_10249_46116# a_8049_45260# 0.001129f
C35003 a_2609_46660# a_n2661_45546# 1.76e-20
C35004 a_1799_45572# a_n2293_45546# 4.04e-20
C35005 a_948_46660# a_997_45618# 7.48e-19
C35006 a_n133_46660# a_n356_45724# 1.93e-19
C35007 a_n743_46660# a_n310_45899# 1.97e-19
C35008 a_n2661_46098# a_n2956_38216# 0.001609f
C35009 a_288_46660# a_310_45028# 2.47e-19
C35010 a_n2157_46122# a_n1853_46287# 0.617317f
C35011 a_n2293_46098# a_n1991_46122# 0.01544f
C35012 a_15682_43940# a_16867_43762# 0.001981f
C35013 a_18451_43940# a_18783_43370# 0.001344f
C35014 a_458_43396# a_1209_43370# 0.0172f
C35015 a_n97_42460# a_4905_42826# 0.147727f
C35016 a_15493_43396# a_18429_43548# 0.045352f
C35017 a_n3674_39768# a_n2472_42826# 1.25e-19
C35018 a_11341_43940# a_16137_43396# 3.22e-19
C35019 a_11967_42832# a_18249_42858# 0.018824f
C35020 a_n2661_42282# a_743_42282# 0.043675f
C35021 a_9313_44734# a_10553_43218# 7.54e-19
C35022 en_comp a_1736_39043# 2.01e-19
C35023 a_4093_43548# VDD 0.216874f
C35024 a_8568_45546# a_8560_45348# 0.001331f
C35025 a_21188_45572# a_20447_31679# 3.01e-20
C35026 a_17499_43370# a_4185_45028# 9.45e-21
C35027 a_5649_42852# a_11415_45002# 2.71e-20
C35028 a_5193_42852# a_5257_43370# 1.09e-19
C35029 a_n2472_42282# a_n2312_38680# 2.73e-20
C35030 COMP_P a_n2956_39768# 0.003427f
C35031 a_n3674_38216# a_n2442_46660# 0.023932f
C35032 a_21381_43940# a_13259_45724# 9.63e-21
C35033 a_3539_42460# a_n1925_42282# 0.024736f
C35034 a_12293_43646# a_9290_44172# 9.78e-19
C35035 a_13657_42558# a_10227_46804# 8.38e-19
C35036 a_n2946_39866# SMPL_ON_P 1.96e-20
C35037 a_8062_46155# VDD 2.63e-20
C35038 a_8696_44636# a_n971_45724# 0.003003f
C35039 a_11652_45724# a_11599_46634# 5.18e-19
C35040 a_10193_42453# a_16327_47482# 0.163668f
C35041 a_12791_45546# a_12861_44030# 0.248928f
C35042 a_11823_42460# a_13487_47204# 3.88e-21
C35043 a_5066_45546# a_10037_46155# 9.67e-23
C35044 a_21137_46414# a_20205_31679# 2.27e-19
C35045 a_18579_44172# a_19511_42282# 2.1e-20
C35046 a_2982_43646# a_21195_42852# 0.034024f
C35047 a_8685_43396# a_10835_43094# 1.12e-19
C35048 a_16823_43084# a_743_42282# 2.26e-19
C35049 a_n1557_42282# a_n2293_42282# 4.61e-19
C35050 a_n2661_42282# a_5755_42308# 0.002898f
C35051 a_3422_30871# a_18727_42674# 5.4e-20
C35052 a_1568_43370# a_1709_42852# 0.015873f
C35053 a_17678_43396# a_4190_30871# 5.27e-21
C35054 a_3080_42308# a_4156_43218# 0.00153f
C35055 a_18114_32519# C4_N_btm 1.47e-19
C35056 a_19721_31679# C3_N_btm 0.001023f
C35057 a_16019_45002# a_11691_44458# 6.26e-20
C35058 a_8560_45348# a_n2661_43370# 1.75e-19
C35059 a_8696_44636# a_17061_44734# 0.003665f
C35060 a_5111_44636# a_4223_44672# 0.418299f
C35061 a_8953_45002# a_n2661_44458# 6.7e-19
C35062 a_4558_45348# a_4743_44484# 5.35e-20
C35063 a_n1059_45260# a_17970_44736# 3.79e-19
C35064 a_n2017_45002# a_18248_44752# 3.8e-22
C35065 a_9306_43218# a_526_44458# 0.001865f
C35066 a_18249_42858# a_13259_45724# 2.6e-19
C35067 a_7765_42852# a_n357_42282# 0.042157f
C35068 a_7871_42858# a_n755_45592# 0.033537f
C35069 a_9482_43914# a_12549_44172# 0.06308f
C35070 a_13556_45296# a_12891_46348# 0.29495f
C35071 a_13348_45260# a_768_44030# 1.76e-19
C35072 a_11322_45546# a_13059_46348# 2.64e-21
C35073 a_413_45260# a_n743_46660# 0.031499f
C35074 a_n37_45144# a_n2438_43548# 2.58e-21
C35075 a_1667_45002# a_n1925_46634# 4.73e-21
C35076 a_3537_45260# a_n2661_46634# 9.12e-22
C35077 a_n143_45144# a_n133_46660# 1.25e-21
C35078 a_2680_45002# a_n2293_46634# 0.017731f
C35079 a_6709_45028# a_5807_45002# 8.09e-19
C35080 a_n2661_45010# a_1799_45572# 1.31e-20
C35081 a_375_42282# a_n1613_43370# 3.94e-20
C35082 a_n2661_43370# a_10227_46804# 0.033611f
C35083 a_22717_36887# VDD 1.72e-20
C35084 a_n1177_44458# a_n971_45724# 0.007865f
C35085 a_5343_44458# a_n2497_47436# 7.63e-21
C35086 a_743_42282# a_3497_42558# 0.001105f
C35087 a_n1991_42858# a_n1630_35242# 1.18e-19
C35088 a_n1641_43230# a_n3674_37592# 2.78e-20
C35089 a_n901_43156# a_n327_42558# 0.001558f
C35090 a_n1076_43230# a_n784_42308# 9.15e-21
C35091 a_13460_43230# a_13291_42460# 3.16e-19
C35092 a_n13_43084# a_196_42282# 2.75e-19
C35093 a_12281_43396# a_14113_42308# 1.99e-20
C35094 a_10341_43396# a_15803_42450# 3.14e-20
C35095 a_22223_46124# EN_OFFSET_CAL 0.011048f
C35096 a_6945_45028# CLK 0.027466f
C35097 a_n3565_39304# VDD 0.888861f
C35098 a_4915_47217# a_n881_46662# 1.23372f
C35099 a_5129_47502# a_n1613_43370# 0.002387f
C35100 a_18479_47436# a_18597_46090# 0.473843f
C35101 a_10227_46804# a_19787_47423# 0.03269f
C35102 a_16023_47582# a_13507_46334# 1.53e-21
C35103 a_16241_47178# a_4883_46098# 3.3e-21
C35104 a_16327_47482# a_21496_47436# 4.85e-21
C35105 a_4700_47436# a_5159_47243# 6.64e-19
C35106 a_4791_45118# a_4842_47243# 0.006879f
C35107 a_n1435_47204# a_n310_47570# 3.53e-21
C35108 a_15811_47375# a_12465_44636# 5.18e-19
C35109 a_n1151_42308# a_11309_47204# 0.546434f
C35110 a_n2497_47436# a_n2956_39768# 7.4e-19
C35111 a_n2833_47464# a_n2661_46634# 0.011033f
C35112 a_21101_45002# a_20980_44850# 0.001202f
C35113 a_12607_44458# a_n2661_43922# 0.060913f
C35114 a_9482_43914# a_12429_44172# 0.0636f
C35115 a_n2293_42834# a_5244_44056# 6.01e-21
C35116 a_10193_42453# a_10341_43396# 0.064616f
C35117 a_626_44172# a_n2661_42282# 6.14e-21
C35118 a_7499_43078# a_12281_43396# 9.62e-20
C35119 a_11691_44458# a_18245_44484# 8.73e-19
C35120 a_2711_45572# a_16664_43396# 0.001086f
C35121 a_11827_44484# a_20596_44850# 1.17e-19
C35122 a_n4209_38216# a_n2956_38680# 0.001636f
C35123 a_17786_45822# VDD 0.007376f
C35124 a_17701_42308# RST_Z 1.77e-20
C35125 a_8333_44056# a_4791_45118# 4.81e-20
C35126 a_6171_45002# a_5164_46348# 1.28e-19
C35127 a_n2017_45002# a_2324_44458# 5.73e-20
C35128 a_5691_45260# a_5497_46414# 1.88e-19
C35129 a_2437_43646# a_22223_46124# 3.38e-19
C35130 a_3357_43084# a_20708_46348# 0.017189f
C35131 a_22223_45572# a_6945_45028# 3.06e-19
C35132 a_3537_45260# a_8199_44636# 0.199536f
C35133 a_12561_45572# a_10586_45546# 8.99e-20
C35134 a_11823_42460# a_n357_42282# 0.063073f
C35135 a_21101_45002# a_19692_46634# 2.38e-19
C35136 a_15060_45348# a_13059_46348# 0.001051f
C35137 a_20159_44458# a_12549_44172# 0.005504f
C35138 a_17517_44484# a_13747_46662# 0.022087f
C35139 a_7705_45326# a_3483_46348# 8.97e-19
C35140 a_375_42282# a_n2293_46098# 2.05e-20
C35141 a_5379_42460# a_6171_42473# 0.110293f
C35142 a_5267_42460# a_5932_42308# 0.026805f
C35143 a_n784_42308# a_10723_42308# 3.86e-20
C35144 a_4933_42558# a_4921_42308# 0.012385f
C35145 a_13887_32519# C4_N_btm 0.001746f
C35146 a_17364_32525# C0_N_btm 8.17e-21
C35147 a_13678_32519# C7_N_btm 2.68e-20
C35148 a_22469_39537# a_22717_36887# 0.003149f
C35149 CAL_P a_22609_37990# 0.205305f
C35150 a_22609_38406# a_22705_38406# 0.090011f
C35151 a_12465_44636# a_13059_46348# 0.163448f
C35152 a_4883_46098# a_16721_46634# 2.68e-20
C35153 a_18479_47436# a_19123_46287# 8.06e-20
C35154 a_10227_46804# a_20107_46660# 0.312495f
C35155 a_18780_47178# a_18285_46348# 9.29e-19
C35156 a_16327_47482# a_21363_46634# 5.35e-21
C35157 a_n237_47217# a_4185_45028# 0.074951f
C35158 a_2063_45854# a_1823_45246# 0.038948f
C35159 a_n1151_42308# a_472_46348# 1.23e-20
C35160 a_2124_47436# a_167_45260# 1.26e-19
C35161 a_584_46384# a_2202_46116# 0.003336f
C35162 a_n443_46116# a_n1853_46287# 0.013261f
C35163 a_n1741_47186# a_6165_46155# 4.48e-20
C35164 a_12549_44172# a_12816_46660# 0.0037f
C35165 a_n743_46660# a_9863_46634# 0.00299f
C35166 a_n2661_46634# a_6969_46634# 0.006553f
C35167 a_3699_46634# a_4651_46660# 3.85e-19
C35168 a_3524_46660# a_4646_46812# 0.001606f
C35169 a_12891_46348# a_13607_46688# 1.34e-20
C35170 a_2864_46660# a_3877_44458# 1.05e-19
C35171 a_2107_46812# a_5429_46660# 4.28e-19
C35172 a_10193_42453# a_20356_42852# 4.95e-19
C35173 a_n2065_43946# a_n3674_39768# 0.001814f
C35174 a_n1761_44111# a_n4318_39768# 2.23e-20
C35175 a_2127_44172# a_2889_44172# 7.46e-20
C35176 a_1414_42308# a_3600_43914# 0.012293f
C35177 a_2479_44172# a_2675_43914# 0.061502f
C35178 a_17517_44484# a_20269_44172# 5.36e-20
C35179 a_11967_42832# a_14955_43940# 1.47e-21
C35180 a_n699_43396# a_4093_43548# 2.73e-20
C35181 a_4223_44672# a_4235_43370# 5.04e-19
C35182 a_453_43940# a_2998_44172# 1.49e-21
C35183 a_413_45260# a_1847_42826# 2.14e-20
C35184 a_n913_45002# a_8037_42858# 0.316376f
C35185 a_n1059_45260# a_8605_42826# 0.007493f
C35186 a_n2017_45002# a_8387_43230# 4.99e-20
C35187 a_10157_44484# VDD 0.174233f
C35188 a_n4315_30879# C9_P_btm 0.003123f
C35189 a_n3420_39616# a_n923_35174# 0.002953f
C35190 a_21613_42308# RST_Z 2.94e-19
C35191 a_20512_43084# a_20202_43084# 0.130366f
C35192 a_20397_44484# a_12741_44636# 1.18e-19
C35193 a_21145_44484# a_11415_45002# 9.18e-20
C35194 a_10729_43914# a_3090_45724# 0.135702f
C35195 a_19929_45028# a_13259_45724# 2.15e-20
C35196 a_17969_45144# a_16375_45002# 5.89e-19
C35197 a_n2661_43922# a_10903_43370# 0.039051f
C35198 a_13857_44734# a_9290_44172# 1.78e-19
C35199 a_6655_43762# a_n1613_43370# 0.013792f
C35200 a_9885_43646# a_4883_46098# 1.07e-20
C35201 a_15681_43442# a_10227_46804# 0.001396f
C35202 a_16137_43396# a_16327_47482# 2.72e-19
C35203 a_18525_43370# a_12861_44030# 1.13e-19
C35204 a_n1991_42858# a_n971_45724# 8.17e-20
C35205 a_n1545_43230# a_n2497_47436# 1.72e-19
C35206 a_n2946_39866# a_n2946_39072# 0.052227f
C35207 a_1736_39587# a_1343_38525# 0.289453f
C35208 a_n4064_39616# a_n3420_39072# 0.05019f
C35209 a_n3420_39616# a_n4064_39072# 6.32746f
C35210 a_n4315_30879# a_n4209_38502# 0.082287f
C35211 a_n1925_46634# VDD 0.783093f
C35212 a_6123_31319# C7_N_btm 0.005631f
C35213 a_5934_30871# C5_N_btm 0.139996f
C35214 a_19692_46634# a_21542_46660# 4.63e-19
C35215 a_948_46660# a_1337_46116# 1.31e-19
C35216 a_n2661_46098# a_739_46482# 4.97e-19
C35217 a_n1925_46634# a_8283_46482# 5.81e-19
C35218 a_n743_46660# a_5527_46155# 1.92e-19
C35219 a_6755_46942# a_5937_45572# 3.17e-19
C35220 a_10428_46928# a_10355_46116# 0.009109f
C35221 a_10249_46116# a_8953_45546# 3.6e-20
C35222 a_18989_43940# a_18249_42858# 4.24e-19
C35223 a_18287_44626# a_19339_43156# 3.19e-19
C35224 a_11967_42832# a_5649_42852# 1.63e-19
C35225 a_18579_44172# a_21259_43561# 8.21e-19
C35226 a_n2661_42834# a_3935_42891# 3.28e-21
C35227 a_9313_44734# a_8952_43230# 1.48e-19
C35228 a_n2293_43922# a_2905_42968# 1.12e-20
C35229 a_n2661_43922# a_3681_42891# 5.11e-21
C35230 a_20640_44752# a_13467_32519# 1.11e-19
C35231 a_n2293_42834# a_n473_42460# 0.001023f
C35232 a_5111_44636# a_5742_30871# 1.17e-20
C35233 a_n2017_45002# a_16522_42674# 0.002301f
C35234 a_n913_45002# a_13921_42308# 2.11e-20
C35235 a_n1059_45260# a_16104_42674# 4.45e-19
C35236 a_15599_45572# a_17668_45572# 1.29e-20
C35237 a_2711_45572# a_11963_45334# 1.25e-20
C35238 a_16333_45814# a_16789_45572# 4.2e-19
C35239 a_6511_45714# a_6709_45028# 0.001019f
C35240 a_3733_45822# a_3232_43370# 5.07e-20
C35241 a_5337_42558# a_4791_45118# 0.003599f
C35242 a_20753_42852# a_13507_46334# 7.33e-21
C35243 a_14955_43940# a_13259_45724# 8.97e-22
C35244 a_n1441_43940# a_n863_45724# 4.78e-21
C35245 a_2675_43914# a_n443_42852# 6.34e-20
C35246 a_17678_43396# a_15227_44166# 3.54e-19
C35247 a_22521_40599# a_22705_38406# 0.008755f
C35248 a_22469_40625# a_22609_38406# 0.066321f
C35249 CAL_N a_22609_37990# 4.7e-20
C35250 a_n4209_37414# C5_P_btm 1.11e-20
C35251 a_n3565_37414# C7_P_btm 1.43e-20
C35252 a_5088_37509# a_n923_35174# 7.48e-20
C35253 a_3754_38470# RST_Z 0.203816f
C35254 a_10355_46116# VDD 0.222751f
C35255 a_7227_45028# a_n971_45724# 1.87e-20
C35256 a_6667_45809# a_n237_47217# 2.43e-19
C35257 a_2711_45572# a_584_46384# 1.02e-20
C35258 a_n3565_38502# a_n3565_37414# 0.030671f
C35259 a_n4209_38502# a_n3420_37440# 0.033073f
C35260 a_n3420_38528# a_n4209_37414# 0.027951f
C35261 a_2324_44458# a_526_44458# 0.279023f
C35262 a_5937_45572# a_8049_45260# 0.103218f
C35263 a_7920_46348# a_8062_46155# 0.005572f
C35264 a_8016_46348# a_10044_46482# 6.14e-19
C35265 a_21542_46660# a_20692_30879# 3.76e-20
C35266 a_n809_44244# a_n3674_37592# 3.34e-21
C35267 a_6293_42852# a_4361_42308# 1.16e-19
C35268 a_n1557_42282# a_n1423_42826# 9.17e-20
C35269 a_10341_43396# a_16137_43396# 0.021507f
C35270 a_14955_43396# a_16547_43609# 5.64e-21
C35271 a_n356_44636# a_7174_31319# 2.55e-20
C35272 a_8685_43396# a_15037_43396# 1.41e-19
C35273 a_12891_46348# RST_Z 9.63e-21
C35274 a_7989_47542# DATA[4] 1.37e-19
C35275 a_n881_46662# DATA[5] 0.082222f
C35276 a_685_42968# VDD 0.088446f
C35277 a_n2956_37592# a_n2946_37984# 0.004313f
C35278 a_n2810_45028# a_n4064_37984# 0.002525f
C35279 a_16115_45572# a_16112_44458# 7.96e-20
C35280 a_8746_45002# a_n2661_43922# 0.003872f
C35281 a_8696_44636# a_13076_44458# 0.003013f
C35282 a_13249_42308# a_9313_44734# 0.031106f
C35283 a_10193_42453# a_n2293_43922# 0.024214f
C35284 a_1307_43914# a_16751_45260# 1.36e-19
C35285 a_10490_45724# a_n2661_42834# 4.83e-22
C35286 a_2437_43646# a_22223_45036# 3.35e-19
C35287 a_2274_45254# a_n2661_43370# 0.019962f
C35288 a_3357_43084# a_21101_45002# 2.54e-21
C35289 a_21513_45002# a_22959_45036# 7.2e-21
C35290 a_22223_45572# a_11827_44484# 0.00211f
C35291 a_5111_44636# a_n2293_42834# 0.110286f
C35292 a_6171_45002# a_5837_45028# 0.001502f
C35293 a_19479_31679# a_21359_45002# 3.83e-19
C35294 a_4649_42852# a_4185_45028# 0.00531f
C35295 a_9803_42558# a_8270_45546# 2.56e-20
C35296 a_5932_42308# a_3090_45724# 2.53e-20
C35297 a_n4209_39304# a_n2956_39768# 0.001636f
C35298 a_5649_42852# a_13259_45724# 1.92021f
C35299 a_8387_43230# a_526_44458# 0.032585f
C35300 a_14537_43646# a_n443_42852# 0.001647f
C35301 a_413_45260# a_21177_47436# 8.97e-20
C35302 a_1307_43914# a_4915_47217# 5.85e-20
C35303 a_n913_45002# a_n2312_40392# 7.85e-21
C35304 a_3357_43084# a_5063_47570# 1.58e-19
C35305 a_2437_43646# a_n1613_43370# 0.027497f
C35306 a_20623_45572# a_12549_44172# 1.26e-21
C35307 a_18596_45572# a_13661_43548# 7.95e-20
C35308 a_19256_45572# a_13747_46662# 0.040187f
C35309 a_10053_45546# a_9863_46634# 1.27e-19
C35310 a_2711_45572# a_11901_46660# 4.34e-20
C35311 a_n443_42852# a_2277_45546# 1.61e-20
C35312 a_6031_43396# a_7227_42308# 2.05e-20
C35313 a_13635_43156# a_14543_43071# 0.013803f
C35314 a_12895_43230# a_5534_30871# 0.004896f
C35315 a_n97_42460# a_15803_42450# 0.004106f
C35316 a_3626_43646# a_8325_42308# 0.001817f
C35317 a_2982_43646# a_8791_42308# 2.53e-19
C35318 a_685_42968# a_873_42968# 7.47e-21
C35319 a_3935_42891# a_n2293_42282# 8.93e-19
C35320 a_15743_43084# a_18861_43218# 3.78e-19
C35321 a_21076_30879# VREF_GND 0.041931f
C35322 a_n901_46420# DATA[0] 2.21e-19
C35323 a_17730_32519# C2_N_btm 4.56e-20
C35324 a_19237_31679# C0_N_btm 0.040442f
C35325 a_22521_40599# a_22469_40625# 1.99151f
C35326 a_14113_42308# VDD 0.365578f
C35327 a_1239_47204# a_n1435_47204# 2.24e-19
C35328 a_n443_46116# a_4915_47217# 0.395101f
C35329 a_4791_45118# a_5129_47502# 0.240381f
C35330 a_2063_45854# a_11031_47542# 9.91e-19
C35331 a_n1151_42308# a_7227_47204# 1.79e-19
C35332 a_6298_44484# a_8103_44636# 0.016067f
C35333 a_5343_44458# a_5883_43914# 0.042199f
C35334 a_10193_42453# a_n97_42460# 0.304653f
C35335 a_16147_45260# a_15493_43940# 2.22e-19
C35336 a_18479_45785# a_11341_43940# 0.019493f
C35337 a_2680_45002# a_2675_43914# 0.001197f
C35338 a_n2810_45028# a_n3674_39768# 0.023163f
C35339 a_n2293_45010# a_n1441_43940# 0.009441f
C35340 a_n2956_37592# a_n4318_39768# 0.029002f
C35341 a_3357_43084# a_6101_44260# 4.26e-19
C35342 a_2123_42473# a_n863_45724# 0.036254f
C35343 a_961_42354# a_n357_42282# 3.8e-19
C35344 a_1184_42692# a_n755_45592# 0.016193f
C35345 a_7499_43078# VDD 1.87959f
C35346 a_4361_42308# RST_Z 4.9e-19
C35347 a_1423_45028# a_3090_45724# 0.450367f
C35348 a_15004_44636# a_13661_43548# 0.012894f
C35349 a_16019_45002# a_15227_44166# 4.44e-19
C35350 a_949_44458# a_n2438_43548# 1.62911f
C35351 a_2779_44458# a_n743_46660# 1.72e-20
C35352 a_19963_31679# a_21076_30879# 0.055082f
C35353 a_2437_43646# a_n2293_46098# 0.027185f
C35354 a_413_45260# a_20841_46902# 1.91e-20
C35355 a_8696_44636# a_12594_46348# 1.12e-20
C35356 a_n2661_43922# a_4883_46098# 0.022558f
C35357 a_17517_44484# a_11599_46634# 1.5e-21
C35358 a_n1331_43914# a_n971_45724# 0.015263f
C35359 a_453_43940# a_n2497_47436# 0.09742f
C35360 a_n1899_43946# a_n746_45260# 2.35e-20
C35361 a_17595_43084# a_17531_42308# 0.001512f
C35362 a_17701_42308# a_17303_42282# 0.049097f
C35363 a_n2104_42282# a_n1736_42282# 7.52e-19
C35364 a_n3674_39304# a_n3690_39392# 0.071784f
C35365 a_n4318_38216# a_n4318_37592# 0.139499f
C35366 a_n2472_42282# COMP_P 1.38e-19
C35367 a_n2840_46634# a_n2312_38680# 0.040373f
C35368 a_n2472_46634# a_n2442_46660# 0.155358f
C35369 a_n2661_46634# a_n2293_46634# 0.060962f
C35370 a_n1613_43370# a_3686_47026# 2.49e-19
C35371 a_4883_46098# a_7927_46660# 5.28e-21
C35372 a_11459_47204# a_11813_46116# 1.67e-20
C35373 a_n1151_42308# a_12156_46660# 0.003059f
C35374 a_18494_42460# a_19319_43548# 0.016978f
C35375 a_18248_44752# a_18079_43940# 6.24e-19
C35376 a_20766_44850# a_20980_44850# 0.097745f
C35377 a_20679_44626# a_3422_30871# 0.078371f
C35378 a_n2661_42834# a_6453_43914# 0.007635f
C35379 a_n2293_42834# a_4235_43370# 0.009569f
C35380 a_20835_44721# a_21398_44850# 0.049827f
C35381 a_20640_44752# a_22315_44484# 2.12e-19
C35382 a_5883_43914# a_9801_44260# 3.67e-19
C35383 a_10057_43914# a_11341_43940# 1e-19
C35384 a_14539_43914# a_15493_43396# 0.024653f
C35385 a_8953_45002# a_9145_43396# 3.05e-20
C35386 a_n2017_45002# a_15743_43084# 0.049212f
C35387 a_n1059_45260# a_18783_43370# 7.13e-19
C35388 a_5934_30871# C5_P_btm 0.139996f
C35389 a_6123_31319# C3_P_btm 0.011333f
C35390 a_n4318_39304# a_n2312_40392# 0.025248f
C35391 a_4223_44672# a_9290_44172# 7.92e-21
C35392 a_9838_44484# a_8016_46348# 0.004677f
C35393 a_8103_44636# a_5937_45572# 5.28e-21
C35394 a_8701_44490# a_8199_44636# 0.25266f
C35395 a_413_45260# a_509_45572# 3.88e-19
C35396 a_3065_45002# a_1609_45822# 3.61e-21
C35397 a_3232_43370# a_3503_45724# 1.73e-19
C35398 a_n2661_43370# a_8034_45724# 1.49e-20
C35399 a_5829_43940# a_768_44030# 2.06e-19
C35400 a_19279_43940# a_19466_46812# 4.38e-20
C35401 a_20766_44850# a_19692_46634# 1.17e-21
C35402 a_14539_43914# a_3483_46348# 1.24006f
C35403 a_20894_47436# VDD 0.188358f
C35404 a_18727_42674# a_7174_31319# 4.47e-20
C35405 a_17303_42282# a_21613_42308# 0.061584f
C35406 a_5934_30871# a_n3420_38528# 2.14e-19
C35407 a_n743_46660# a_6165_46155# 0.004708f
C35408 a_5807_45002# a_13925_46122# 0.027158f
C35409 a_n2661_46634# a_9625_46129# 3.03e-19
C35410 a_n1925_46634# a_7920_46348# 0.007001f
C35411 a_13661_43548# a_13759_46122# 8.09e-22
C35412 a_n2293_46634# a_8199_44636# 0.029753f
C35413 a_n881_46662# a_10809_44734# 0.026121f
C35414 a_n2312_39304# a_n1925_42282# 6.33e-20
C35415 a_4883_46098# a_6419_46482# 7.98e-20
C35416 a_18479_47436# a_8049_45260# 0.047429f
C35417 a_11599_46634# a_12379_46436# 0.005949f
C35418 a_n971_45724# a_2957_45546# 8.45e-20
C35419 a_2063_45854# a_n2293_45546# 0.002045f
C35420 a_327_47204# a_310_45028# 1.58e-19
C35421 a_2905_45572# a_n2661_45546# 0.003174f
C35422 a_n237_47217# a_997_45618# 1.85e-19
C35423 a_2107_46812# a_3483_46348# 0.100707f
C35424 a_n2661_46098# a_1176_45822# 0.144277f
C35425 a_17609_46634# a_18834_46812# 0.001296f
C35426 a_6969_46634# a_765_45546# 0.001746f
C35427 a_12469_46902# a_12347_46660# 3.16e-19
C35428 a_949_44458# a_2075_43172# 1.09e-20
C35429 a_2779_44458# a_1847_42826# 1.85e-21
C35430 a_n1549_44318# a_n1557_42282# 4.58e-21
C35431 a_453_43940# a_1568_43370# 1.29e-19
C35432 a_5495_43940# a_n97_42460# 3.76e-20
C35433 a_11341_43940# a_14021_43940# 3.06514f
C35434 a_895_43940# a_458_43396# 6.21e-19
C35435 a_1414_42308# a_1756_43548# 6.51e-20
C35436 a_11967_42832# a_8685_43396# 0.005728f
C35437 a_14673_44172# a_14955_43396# 2.24e-22
C35438 a_9313_44734# a_19700_43370# 0.001757f
C35439 a_n699_43396# a_685_42968# 3.03e-20
C35440 a_742_44458# a_2905_42968# 0.15065f
C35441 a_11827_44484# a_5534_30871# 2.07e-22
C35442 a_9672_43914# a_9801_43940# 0.062574f
C35443 a_n2293_42834# a_5837_43172# 1.46e-19
C35444 a_n967_45348# a_n1630_35242# 0.03295f
C35445 a_n2017_45002# a_1606_42308# 0.04498f
C35446 a_n913_45002# a_1149_42558# 4.87e-21
C35447 a_n1059_45260# a_1221_42558# 1.28e-19
C35448 a_3600_43914# VDD 0.22716f
C35449 a_13249_42308# a_15037_45618# 1.93e-21
C35450 a_11823_42460# a_15765_45572# 1.14e-19
C35451 a_11322_45546# a_8696_44636# 6e-19
C35452 a_14495_45572# a_14033_45822# 3.98e-20
C35453 C10_N_btm VCM 10.5945f
C35454 a_5326_44056# a_1823_45246# 7.22e-20
C35455 a_21381_43940# a_20202_43084# 0.108097f
C35456 a_n1076_43230# a_n2438_43548# 2.79e-21
C35457 a_4181_43396# a_3090_45724# 2.49e-22
C35458 a_n2661_42282# a_n2956_38680# 3.65e-20
C35459 a_15682_43940# a_17715_44484# 0.007815f
C35460 a_20411_46873# VDD 0.348821f
C35461 a_n2840_46090# a_n2956_38680# 0.050916f
C35462 a_n2472_46090# a_n2956_39304# 9.6e-19
C35463 a_6755_46942# a_n443_42852# 1.03e-19
C35464 a_2521_46116# a_2324_44458# 1.5e-20
C35465 a_8016_46348# a_9823_46155# 0.048283f
C35466 a_8199_44636# a_9625_46129# 0.011574f
C35467 a_5937_45572# a_8953_45546# 0.3871f
C35468 a_10949_43914# a_10341_42308# 1.01e-22
C35469 a_10807_43548# a_10922_42852# 0.010566f
C35470 a_n97_42460# a_16137_43396# 0.134668f
C35471 a_n2293_43922# a_n784_42308# 1.67292f
C35472 a_n356_44636# a_5932_42308# 0.040714f
C35473 a_18184_42460# a_21887_42336# 1.63e-19
C35474 a_6031_43396# a_6643_43396# 3.82e-19
C35475 a_2479_44172# a_3059_42968# 7.19e-19
C35476 a_11967_42832# a_15953_42852# 2.76e-20
C35477 a_10057_43914# a_10723_42308# 2.38e-19
C35478 a_3626_43646# a_9145_43396# 9.28e-20
C35479 a_4915_47217# DATA[4] 0.069022f
C35480 a_5129_47502# DATA[3] 4.21e-20
C35481 a_5815_47464# DATA[2] 9.97e-21
C35482 a_20447_31679# C9_N_btm 3.26e-20
C35483 a_15781_43660# VDD 0.196099f
C35484 a_8162_45546# a_5343_44458# 7.23e-21
C35485 a_6812_45938# a_6298_44484# 1.87e-20
C35486 a_2711_45572# a_18443_44721# 2.09e-20
C35487 a_15903_45785# a_16405_45348# 4.53e-20
C35488 a_2680_45002# a_3429_45260# 4.16e-19
C35489 a_2382_45260# a_3537_45260# 0.250657f
C35490 a_n1059_45260# a_8953_45002# 8.21e-22
C35491 a_n4315_30879# a_n2312_39304# 0.033437f
C35492 a_n4334_40480# a_n2312_40392# 3.26e-19
C35493 a_2982_43646# a_n357_42282# 0.04908f
C35494 a_1209_43370# a_n443_42852# 0.010053f
C35495 a_8685_43396# a_13259_45724# 0.031693f
C35496 a_18249_42858# a_20202_43084# 2.75e-20
C35497 a_5755_42852# a_4185_45028# 4.48e-21
C35498 a_7871_42858# a_3483_46348# 5.12e-21
C35499 a_n310_45572# VDD 7.01e-20
C35500 a_11962_45724# a_5807_45002# 6.78e-21
C35501 a_6472_45840# a_2107_46812# 4.62e-20
C35502 a_16333_45814# a_11453_44696# 2.89e-21
C35503 a_8696_44636# a_12465_44636# 0.038471f
C35504 a_17478_45572# a_4883_46098# 3.85e-20
C35505 a_19256_45572# a_11599_46634# 0.051691f
C35506 a_18479_45785# a_16327_47482# 0.841261f
C35507 a_16211_45572# a_10227_46804# 3.48e-19
C35508 a_n967_45348# a_n971_45724# 0.581053f
C35509 a_2437_43646# a_4791_45118# 0.00511f
C35510 en_comp a_n746_45260# 2.06e-20
C35511 a_2274_45254# a_n2497_47436# 3.04e-20
C35512 a_n1917_43396# a_n1630_35242# 3.12e-20
C35513 a_104_43370# a_196_42282# 4.54e-20
C35514 a_19268_43646# a_19339_43156# 0.001878f
C35515 a_n97_42460# a_n784_42308# 0.006645f
C35516 a_5649_42852# a_10518_42984# 7.51e-21
C35517 a_4361_42308# a_10991_42826# 2.13e-19
C35518 a_743_42282# a_12545_42858# 8.12e-20
C35519 a_15743_43084# a_19164_43230# 0.0353f
C35520 a_15493_43940# a_15051_42282# 1.93e-19
C35521 a_15559_46634# CLK 2.96e-21
C35522 a_n4064_37984# a_n2302_37690# 2.59e-20
C35523 a_7754_39300# a_7754_38968# 0.296258f
C35524 a_n2302_37984# a_n4064_37440# 2.59e-20
C35525 a_7754_40130# a_7754_38470# 0.111791f
C35526 a_7754_39964# a_3754_38470# 0.081868f
C35527 a_n1329_42308# VDD 0.237697f
C35528 a_21359_45002# a_20193_45348# 3.23e-20
C35529 a_n2661_43370# a_4743_44484# 0.001974f
C35530 a_1423_45028# a_n356_44636# 2.19e-21
C35531 a_11827_44484# a_11691_44458# 0.881979f
C35532 a_18587_45118# a_18545_45144# 7.47e-21
C35533 a_3232_43370# a_n2661_43922# 0.197944f
C35534 a_6171_45002# a_n2661_42834# 0.001465f
C35535 a_21125_42558# a_20202_43084# 0.002691f
C35536 a_1606_42308# a_526_44458# 0.011179f
C35537 a_5837_42852# a_n357_42282# 0.01329f
C35538 a_5742_30871# a_9290_44172# 0.118117f
C35539 CAL_N a_18597_46090# 0.001283f
C35540 a_n2293_43922# SMPL_ON_P 2.28e-19
C35541 a_5883_43914# a_10227_46804# 2.83e-21
C35542 a_16979_44734# a_12861_44030# 5.79e-19
C35543 a_n4318_40392# a_n2312_39304# 0.023465f
C35544 a_n2661_44458# a_n2312_40392# 2.36e-20
C35545 a_7230_45938# a_8199_44636# 8.25e-21
C35546 a_6812_45938# a_5937_45572# 3.01e-19
C35547 a_8162_45546# a_8349_46414# 3.15e-21
C35548 a_4099_45572# a_2324_44458# 1.48e-20
C35549 a_8568_45546# a_8016_46348# 3.81e-20
C35550 a_7229_43940# a_5257_43370# 4.91e-22
C35551 a_3357_43084# a_14976_45028# 3.74e-20
C35552 a_2437_43646# a_16292_46812# 3.48e-20
C35553 a_18911_45144# a_12549_44172# 6.77e-20
C35554 a_12427_45724# a_3483_46348# 1.97e-20
C35555 a_8037_42858# a_8325_42308# 5.53e-19
C35556 a_7871_42858# a_8791_42308# 0.004922f
C35557 a_n2293_42282# a_n3674_37592# 0.08084f
C35558 a_4361_42308# a_17303_42282# 0.050893f
C35559 a_743_42282# a_19332_42282# 0.006778f
C35560 a_13003_42852# a_13291_42460# 2.39e-20
C35561 a_4190_30871# a_18220_42308# 0.00137f
C35562 a_17538_32519# C2_N_btm 2.28e-20
C35563 a_4883_46098# a_19594_46812# 3.17e-19
C35564 a_21177_47436# a_20916_46384# 4.75e-19
C35565 a_20990_47178# a_21588_30879# 2.92e-19
C35566 a_16023_47582# a_n743_46660# 0.004115f
C35567 a_n237_47217# a_5257_43370# 0.022234f
C35568 a_n971_45724# a_7715_46873# 0.029319f
C35569 a_2063_45854# a_5732_46660# 2.69e-20
C35570 a_3785_47178# a_4646_46812# 8.96e-19
C35571 a_n1151_42308# a_4955_46873# 0.261025f
C35572 a_3815_47204# a_3877_44458# 1.11e-19
C35573 a_17613_45144# a_17737_43940# 7.01e-20
C35574 a_n699_43396# a_3600_43914# 1.42e-19
C35575 a_4223_44672# a_3905_42865# 0.019153f
C35576 a_8696_44636# a_16409_43396# 4.05e-20
C35577 a_18479_45785# a_10341_43396# 0.038969f
C35578 a_15861_45028# a_16547_43609# 4.56e-21
C35579 a_1307_43914# a_11173_43940# 3.43e-19
C35580 a_n2267_44484# a_n4318_39768# 4.62e-19
C35581 a_2274_45254# a_1568_43370# 1.33e-21
C35582 a_n1059_45260# a_3626_43646# 0.025708f
C35583 a_n2017_45002# a_3539_42460# 0.042001f
C35584 a_3357_43084# a_7287_43370# 7.22e-20
C35585 a_n2946_38778# a_n2956_38216# 0.004751f
C35586 a_4558_45348# VDD 0.25277f
C35587 a_17896_45144# a_12741_44636# 1.01e-19
C35588 a_18545_45144# a_11415_45002# 1.83e-20
C35589 a_6109_44484# a_3090_45724# 0.001946f
C35590 a_6171_45002# a_5066_45546# 0.002485f
C35591 a_n2661_43370# a_8016_46348# 0.028709f
C35592 a_1307_43914# a_10809_44734# 2.22e-19
C35593 a_7735_45067# a_5937_45572# 6.35e-19
C35594 a_8704_45028# a_8199_44636# 3.64e-19
C35595 a_15493_43396# a_11453_44696# 1.19e-21
C35596 a_11341_43940# a_13507_46334# 0.162723f
C35597 a_14021_43940# a_16327_47482# 0.061511f
C35598 a_n1917_43396# a_n971_45724# 0.001021f
C35599 a_13575_42558# a_14456_42282# 0.008255f
C35600 a_3823_42558# a_7174_31319# 4.88e-21
C35601 a_n3674_38680# a_n4334_39392# 1.52e-19
C35602 a_n3674_37592# a_n3565_39590# 4.6e-20
C35603 a_n1630_35242# a_n4209_39590# 0.12484f
C35604 a_9803_42558# a_10149_42308# 0.013377f
C35605 a_13070_42354# a_13249_42558# 0.010303f
C35606 a_n2288_47178# VDD 0.29372f
C35607 a_768_44030# a_11415_45002# 0.021062f
C35608 a_n2293_46634# a_765_45546# 8.06e-22
C35609 a_20916_46384# a_20841_46902# 2.67e-19
C35610 a_10554_47026# a_6755_46942# 0.005096f
C35611 a_4646_46812# a_3090_45724# 0.199722f
C35612 a_5807_45002# a_16655_46660# 0.006956f
C35613 a_7577_46660# a_8654_47026# 1.46e-19
C35614 a_n881_46662# a_n2157_46122# 0.005335f
C35615 a_n1613_43370# a_n1853_46287# 0.354256f
C35616 a_11453_44696# a_3483_46348# 0.027804f
C35617 a_4883_46098# a_5164_46348# 0.01685f
C35618 a_14955_47212# a_13759_46122# 2.05e-20
C35619 a_11599_46634# a_13351_46090# 0.105205f
C35620 a_14311_47204# a_13925_46122# 1.89e-21
C35621 a_10227_46804# a_9569_46155# 1.63e-20
C35622 a_n1151_42308# a_n967_46494# 4.11e-19
C35623 a_n237_47217# a_1337_46116# 8.45e-19
C35624 a_12861_44030# a_14275_46494# 1.23e-19
C35625 a_13717_47436# a_15015_46420# 4.43e-21
C35626 a_21005_45260# a_20556_43646# 2.16e-21
C35627 a_10057_43914# a_10341_43396# 0.055207f
C35628 a_6109_44484# a_6547_43396# 0.001963f
C35629 a_7499_43078# a_11551_42558# 3.18e-19
C35630 a_n2661_43922# a_4905_42826# 9.3e-21
C35631 a_5891_43370# a_6293_42852# 0.107308f
C35632 a_11827_44484# a_4190_30871# 3.39e-20
C35633 a_1307_43914# a_13460_43230# 1.02e-20
C35634 a_14537_43396# a_15567_42826# 4.38e-22
C35635 a_n2293_42834# a_791_42968# 0.007944f
C35636 a_10193_42453# a_10533_42308# 0.101629f
C35637 a_n1899_43946# a_726_44056# 1.56e-20
C35638 a_18184_42460# a_13467_32519# 0.022572f
C35639 a_n2293_43922# a_3080_42308# 0.084673f
C35640 a_18494_42460# a_19095_43396# 3.48e-20
C35641 a_3232_43370# a_3445_43172# 1.88e-19
C35642 a_2711_45572# a_13249_42308# 0.043493f
C35643 a_13635_43156# a_4915_47217# 1.83e-20
C35644 a_14539_43914# a_n357_42282# 0.028064f
C35645 a_8103_44636# a_n443_42852# 2.86e-19
C35646 a_18797_44260# a_3090_45724# 9.33e-20
C35647 a_15037_44260# a_13059_46348# 7.67e-20
C35648 a_16759_43396# a_13661_43548# 9.73e-21
C35649 a_6547_43396# a_4646_46812# 0.03374f
C35650 a_13483_43940# a_11415_45002# 2.17e-21
C35651 a_20447_31679# RST_Z 0.050985f
C35652 a_2437_43646# DATA[3] 0.075788f
C35653 a_6999_46987# VDD 2.18e-20
C35654 a_19692_46634# a_19900_46494# 0.004501f
C35655 a_765_45546# a_9625_46129# 1.15e-19
C35656 a_14513_46634# a_14493_46090# 0.00967f
C35657 a_14180_46812# a_14275_46494# 0.002474f
C35658 a_15227_44166# a_6945_45028# 0.548194f
C35659 a_17609_46634# a_10809_44734# 0.018125f
C35660 a_13059_46348# a_12005_46116# 3.28e-19
C35661 a_14035_46660# a_15015_46420# 1.29e-20
C35662 a_6123_31319# a_7754_40130# 6.87e-20
C35663 a_n2661_46634# a_2277_45546# 8.59e-21
C35664 a_948_46660# a_n755_45592# 8.59e-22
C35665 a_n743_46660# a_n23_45546# 0.070296f
C35666 a_2443_46660# a_n2661_45546# 1.59e-20
C35667 a_1123_46634# a_997_45618# 1.11e-20
C35668 a_n2438_43548# a_n356_45724# 5.71e-20
C35669 a_n2472_46090# a_n1991_46122# 7.66e-19
C35670 a_n2293_46098# a_n1853_46287# 0.02738f
C35671 COMP_P VDAC_P 0.003408f
C35672 a_1115_44172# a_791_42968# 7.5e-19
C35673 a_15682_43940# a_16664_43396# 0.001235f
C35674 a_18079_43940# a_15743_43084# 6.36e-20
C35675 a_n1177_43370# a_n1557_42282# 4.78e-22
C35676 a_742_44458# a_n784_42308# 4.46e-20
C35677 a_n97_42460# a_3080_42308# 0.353977f
C35678 a_18451_43940# a_18525_43370# 3.66e-19
C35679 a_15493_43396# a_17324_43396# 0.047612f
C35680 a_14021_43940# a_10341_43396# 1.5617f
C35681 a_11967_42832# a_17333_42852# 0.14149f
C35682 a_n3674_39768# a_n2840_42826# 0.001686f
C35683 en_comp a_1239_39043# 0.007802f
C35684 w_11334_34010# CAL_P 0.063131f
C35685 a_1756_43548# VDD 0.138878f
C35686 a_2711_45572# a_17613_45144# 1.8e-20
C35687 a_4808_45572# a_n2661_43370# 2.36e-19
C35688 a_15861_45028# a_6171_45002# 0.09425f
C35689 a_21188_45572# a_22959_45572# 8.11e-21
C35690 a_21363_45546# a_20447_31679# 5.34e-20
C35691 a_17324_43396# a_3483_46348# 1.78e-19
C35692 a_5649_42852# a_20202_43084# 0.011671f
C35693 a_n2104_42282# a_n2442_46660# 4.03e-20
C35694 a_n3674_38680# a_n2312_38680# 0.023204f
C35695 a_n4318_37592# a_n2956_39768# 0.02357f
C35696 a_3539_42460# a_526_44458# 0.213772f
C35697 a_3626_43646# a_n1925_42282# 0.031012f
C35698 a_9885_43396# a_8953_45546# 0.002213f
C35699 a_n3420_39616# SMPL_ON_P 1.92e-20
C35700 a_11823_42460# a_12861_44030# 1.2465f
C35701 a_11525_45546# a_11599_46634# 1.45e-19
C35702 a_5066_45546# a_9751_46155# 6.54e-21
C35703 a_8953_45546# a_n443_42852# 0.134632f
C35704 a_20708_46348# a_20205_31679# 2.2e-19
C35705 a_6945_45028# a_21071_46482# 7.43e-19
C35706 a_2982_43646# a_21356_42826# 0.005304f
C35707 a_8685_43396# a_10518_42984# 4.24e-19
C35708 a_3422_30871# a_18057_42282# 3.03e-20
C35709 a_n97_42460# a_7309_43172# 0.002468f
C35710 a_17433_43396# a_4190_30871# 4.55e-21
C35711 a_1568_43370# a_945_42968# 1.47e-20
C35712 a_3080_42308# a_3935_43218# 4.27e-20
C35713 a_19279_43940# a_13258_32519# 4.56e-21
C35714 a_15743_43084# a_14209_32519# 4.59e-21
C35715 a_18114_32519# C3_N_btm 1.27e-19
C35716 a_19721_31679# C2_N_btm 0.040789f
C35717 a_15595_45028# a_11691_44458# 2.85e-20
C35718 a_8696_44636# a_16241_44734# 0.004986f
C35719 a_3537_45260# a_5343_44458# 0.378482f
C35720 a_8191_45002# a_n2661_44458# 0.001306f
C35721 a_5147_45002# a_4223_44672# 0.047867f
C35722 a_4558_45348# a_n699_43396# 4.82e-22
C35723 a_n1059_45260# a_17767_44458# 2.41e-19
C35724 a_9061_43230# a_526_44458# 8.29e-19
C35725 a_17333_42852# a_13259_45724# 0.077331f
C35726 a_7871_42858# a_n357_42282# 0.035744f
C35727 CAL_N w_11334_34010# 1.49e-19
C35728 a_13348_45260# a_12549_44172# 0.001434f
C35729 a_11823_42460# a_14180_46812# 8.14e-22
C35730 a_9482_43914# a_12891_46348# 0.314487f
C35731 a_n143_45144# a_n2438_43548# 1.67e-20
C35732 a_n37_45144# a_n743_46660# 5.42e-20
C35733 a_327_44734# a_n1925_46634# 2.4e-20
C35734 a_7229_43940# a_5807_45002# 3.1e-20
C35735 a_2382_45260# a_n2293_46634# 0.046113f
C35736 a_1307_43914# a_n881_46662# 1.96e-19
C35737 a_22717_37285# VDD 3.6e-19
C35738 a_4743_44484# a_n2497_47436# 0.003104f
C35739 a_n1533_42852# a_n4318_38216# 4.39e-19
C35740 a_n1853_43023# a_n1630_35242# 1.28e-19
C35741 a_n1423_42826# a_n3674_37592# 4.62e-20
C35742 a_n901_43156# a_n784_42308# 4.44e-19
C35743 a_n13_43084# a_n473_42460# 2.62e-19
C35744 a_13635_43156# a_13291_42460# 0.004222f
C35745 a_4361_42308# a_2713_42308# 2.85e-20
C35746 a_743_42282# a_5379_42460# 0.013947f
C35747 a_12281_43396# a_13657_42558# 1.55e-21
C35748 a_10341_43396# a_15764_42576# 7.76e-21
C35749 a_14209_32519# a_1606_42308# 1.87e-20
C35750 a_n4334_39392# VDD 0.385989f
C35751 a_18143_47464# a_18597_46090# 0.002913f
C35752 a_18479_47436# a_18780_47178# 0.056304f
C35753 a_10227_46804# a_19386_47436# 0.041193f
C35754 a_16327_47482# a_13507_46334# 0.043159f
C35755 a_4700_47436# a_4842_47243# 0.005572f
C35756 a_n443_46116# a_n881_46662# 0.114922f
C35757 a_n1435_47204# a_n2312_39304# 6.02e-19
C35758 a_15507_47210# a_12465_44636# 9.53e-19
C35759 a_2553_47502# a_768_44030# 2.24e-19
C35760 a_n2833_47464# a_n2956_39768# 0.008074f
C35761 a_n237_47217# a_5807_45002# 0.082779f
C35762 a_4915_47217# a_n1613_43370# 0.195064f
C35763 a_21005_45260# a_20980_44850# 5.39e-19
C35764 a_8975_43940# a_n2661_43922# 0.11532f
C35765 a_18287_44626# a_9313_44734# 6.97e-21
C35766 a_20193_45348# a_19279_43940# 0.021458f
C35767 a_18184_42460# a_22315_44484# 1.48e-22
C35768 a_n2661_43370# a_1414_42308# 9.45e-21
C35769 a_n2293_42834# a_3905_42865# 0.039227f
C35770 a_9482_43914# a_11750_44172# 0.020902f
C35771 a_2711_45572# a_19700_43370# 0.016505f
C35772 a_18494_42460# a_3422_30871# 7.81e-19
C35773 a_18479_45785# a_n97_42460# 0.072469f
C35774 a_11691_44458# a_18005_44484# 0.001888f
C35775 a_12607_44458# a_n2661_42834# 5.21e-19
C35776 a_11827_44484# a_18753_44484# 0.001286f
C35777 a_14456_42282# a_n443_42852# 7.8e-21
C35778 a_17595_43084# RST_Z 2.39e-21
C35779 a_3232_43370# a_5164_46348# 5.59e-20
C35780 a_413_45260# a_9290_44172# 3.87e-22
C35781 a_3357_43084# a_19900_46494# 7.4e-21
C35782 a_2437_43646# a_6945_45028# 2.26888f
C35783 a_14976_45348# a_13059_46348# 0.001245f
C35784 a_n356_44636# a_4646_46812# 1.8e-20
C35785 a_n2293_43922# a_n2438_43548# 0.575621f
C35786 a_19615_44636# a_12549_44172# 0.157395f
C35787 a_11967_42832# a_768_44030# 1.22e-21
C35788 a_21101_45002# a_19466_46812# 2.51e-20
C35789 a_17517_44484# a_13661_43548# 0.01824f
C35790 a_11827_44484# a_15227_44166# 0.084637f
C35791 a_21005_45260# a_19692_46634# 4.64e-19
C35792 a_6709_45028# a_3483_46348# 0.002873f
C35793 a_2351_42308# a_5934_30871# 1.01e-20
C35794 a_3905_42558# a_4921_42308# 4.04e-22
C35795 a_5379_42460# a_5755_42308# 0.004559f
C35796 a_n784_42308# a_10533_42308# 2.26e-20
C35797 a_3823_42558# a_5932_42308# 4.34e-21
C35798 a_13678_32519# C6_N_btm 1.22e-19
C35799 a_13887_32519# C3_N_btm 0.030933f
C35800 a_14209_32519# C1_N_btm 4.13e-20
C35801 a_22469_39537# a_22717_37285# 0.002793f
C35802 a_4883_46098# a_16388_46812# 0.041939f
C35803 a_18597_46090# a_765_45546# 1.63e-19
C35804 a_18479_47436# a_18285_46348# 7.49e-21
C35805 a_12861_44030# a_18280_46660# 0.140921f
C35806 a_n237_47217# a_3699_46348# 0.044064f
C35807 a_n443_46116# a_n2157_46122# 3.46e-20
C35808 a_584_46384# a_1823_45246# 0.094654f
C35809 a_1431_47204# a_167_45260# 5.7e-22
C35810 a_2124_47436# a_2202_46116# 4.23e-20
C35811 a_2063_45854# a_1138_42852# 2.69e-19
C35812 a_5807_45002# a_8270_45546# 0.029164f
C35813 a_12891_46348# a_12816_46660# 0.024711f
C35814 a_n743_46660# a_8492_46660# 1.3e-20
C35815 a_n2661_46634# a_6755_46942# 1.40968f
C35816 a_3699_46634# a_4646_46812# 2.69e-19
C35817 a_3524_46660# a_3877_44458# 0.008528f
C35818 a_12549_44172# a_12991_46634# 0.010497f
C35819 a_2609_46660# a_4817_46660# 0.00171f
C35820 a_2107_46812# a_5263_46660# 8.47e-19
C35821 a_n971_45724# a_4419_46090# 2.52e-19
C35822 a_10193_42453# a_20256_42852# 4.84e-19
C35823 a_2479_44172# a_895_43940# 0.318312f
C35824 a_1414_42308# a_2998_44172# 0.447595f
C35825 a_n2472_43914# a_n3674_39768# 0.162742f
C35826 a_n2065_43946# a_n4318_39768# 3.52e-21
C35827 a_2127_44172# a_2675_43914# 0.090298f
C35828 a_11967_42832# a_13483_43940# 1.65e-20
C35829 a_5891_43370# a_7499_43940# 7.45e-20
C35830 a_17517_44484# a_19862_44208# 2.23e-19
C35831 a_n699_43396# a_1756_43548# 0.004876f
C35832 a_742_44458# a_3080_42308# 5.11e-20
C35833 a_4223_44672# a_4093_43548# 1.33e-19
C35834 a_10057_43914# a_n97_42460# 4.56e-21
C35835 a_n1059_45260# a_8037_42858# 0.048776f
C35836 a_327_44734# a_685_42968# 4.03e-22
C35837 a_n913_45002# a_7765_42852# 4.6e-19
C35838 a_9838_44484# VDD 0.242131f
C35839 a_n4315_30879# C10_P_btm 1.5848f
C35840 a_n3420_39616# a_n1532_35090# 1.07e-19
C35841 a_21887_42336# RST_Z 1.97e-20
C35842 a_17517_44484# a_4185_45028# 0.006178f
C35843 a_21073_44484# a_11415_45002# 4.79e-20
C35844 a_648_43396# a_768_44030# 5.84e-19
C35845 a_10405_44172# a_3090_45724# 0.126512f
C35846 a_18545_45144# a_13259_45724# 2.48e-21
C35847 a_17896_45144# a_16375_45002# 3.43e-20
C35848 a_n2661_42834# a_10903_43370# 0.269313f
C35849 a_6452_43396# a_n1613_43370# 3.31e-19
C35850 a_14205_43396# a_12465_44636# 8.42e-21
C35851 a_10341_43396# a_13507_46334# 0.030637f
C35852 a_14621_43646# a_10227_46804# 3.58e-19
C35853 a_18429_43548# a_12861_44030# 3.85e-19
C35854 a_n1853_43023# a_n971_45724# 0.02483f
C35855 a_n901_43156# SMPL_ON_P 4.04e-21
C35856 a_10907_45822# CLK 0.035046f
C35857 a_1239_39587# a_1343_38525# 0.011696f
C35858 a_n3565_39590# a_n2302_39072# 8.95e-20
C35859 a_7174_31319# a_1177_38525# 1.57e-19
C35860 a_n2312_38680# VDD 0.540248f
C35861 a_6123_31319# C6_N_btm 6.31e-19
C35862 a_5934_30871# C4_N_btm 0.030578f
C35863 a_19692_46634# a_21297_46660# 5.35e-19
C35864 a_768_44030# a_13259_45724# 0.315247f
C35865 a_1123_46634# a_1337_46116# 1.76e-19
C35866 a_n2661_46634# a_8049_45260# 0.027919f
C35867 a_n2661_46098# a_518_46482# 0.001429f
C35868 a_5807_45002# a_12638_46436# 0.006618f
C35869 a_n743_46660# a_5210_46155# 1.05e-19
C35870 a_10150_46912# a_10355_46116# 7.72e-19
C35871 a_6755_46942# a_8199_44636# 3.74e-19
C35872 a_18287_44626# a_18599_43230# 2.95e-19
C35873 a_20835_44721# a_20556_43646# 9.48e-20
C35874 a_11967_42832# a_13678_32519# 1.08e-19
C35875 a_20679_44626# a_21487_43396# 5.88e-19
C35876 a_8333_44056# a_8147_43396# 0.011009f
C35877 a_n2661_43922# a_2905_42968# 2.14e-21
C35878 a_9313_44734# a_9127_43156# 0.001322f
C35879 a_14021_43940# a_n97_42460# 0.002657f
C35880 a_18374_44850# a_18249_42858# 3.5e-21
C35881 a_n2661_42834# a_3681_42891# 1.08e-21
C35882 a_n356_44636# a_15567_42826# 1.19e-20
C35883 a_n2293_42834# a_n961_42308# 0.001885f
C35884 a_18494_42460# a_18504_43218# 8.04e-19
C35885 a_n2017_45002# a_16104_42674# 0.004413f
C35886 a_2711_45572# a_11787_45002# 2.49e-20
C35887 a_15765_45572# a_16789_45572# 2.36e-20
C35888 a_17478_45572# a_18341_45572# 5.87e-19
C35889 a_6472_45840# a_6709_45028# 8.56e-19
C35890 a_6598_45938# a_5205_44484# 5.22e-19
C35891 a_6511_45714# a_7229_43940# 6.9e-21
C35892 a_11823_42460# a_n913_45002# 0.281323f
C35893 a_3638_45822# a_3232_43370# 1.51e-20
C35894 a_4921_42308# a_4791_45118# 0.172224f
C35895 a_22469_40625# CAL_P 0.001716f
C35896 a_22521_40599# a_22609_38406# 0.032572f
C35897 CAL_N a_22705_38406# 4.85e-21
C35898 a_n4209_37414# C6_P_btm 1.26e-20
C35899 a_n3565_37414# C8_P_btm 1.71e-20
C35900 a_4338_37500# a_n923_35174# 1.22e-19
C35901 a_3353_43940# a_526_44458# 0.002743f
C35902 a_13483_43940# a_13259_45724# 0.002807f
C35903 a_895_43940# a_n443_42852# 6.44e-19
C35904 a_17433_43396# a_15227_44166# 1.76e-19
C35905 a_5755_42852# a_5257_43370# 7.53e-19
C35906 a_9823_46155# VDD 0.102474f
C35907 a_6511_45714# a_n237_47217# 3.49e-19
C35908 a_6598_45938# a_n971_45724# 2.89e-20
C35909 a_n3565_38502# a_n4334_37440# 4.13e-19
C35910 a_n4209_38502# a_n3690_37440# 3.34e-19
C35911 a_n4209_39304# VDAC_P 0.001867f
C35912 a_6945_45028# a_22959_46124# 4.91e-20
C35913 a_8199_44636# a_8049_45260# 0.069189f
C35914 a_22223_46124# a_10809_44734# 0.005525f
C35915 a_765_45546# a_2277_45546# 3.26e-20
C35916 a_n1899_43946# a_n1630_35242# 1.8e-21
C35917 a_n809_44244# a_n327_42558# 7.98e-21
C35918 a_6031_43396# a_4361_42308# 3.96e-20
C35919 a_7287_43370# a_743_42282# 2.89e-20
C35920 a_2982_43646# a_20749_43396# 0.00204f
C35921 a_n1557_42282# a_n1991_42858# 1.42e-19
C35922 a_175_44278# a_196_42282# 4.29e-21
C35923 a_9313_44734# a_17124_42282# 4.54e-20
C35924 a_15095_43370# a_16547_43609# 2.35e-21
C35925 a_10807_43548# a_11554_42852# 0.002521f
C35926 a_10341_43396# a_13943_43396# 7.41e-20
C35927 a_7989_47542# DATA[3] 2.61e-19
C35928 a_n881_46662# DATA[4] 0.087677f
C35929 a_421_43172# VDD 1.56e-19
C35930 a_n2956_37592# a_n3420_37984# 0.001223f
C35931 a_10193_42453# a_n2661_43922# 0.025533f
C35932 a_15765_45572# a_14539_43914# 1.95e-20
C35933 a_16333_45814# a_16112_44458# 4.95e-21
C35934 a_8746_45002# a_n2661_42834# 1.37e-19
C35935 a_8696_44636# a_12883_44458# 0.002403f
C35936 a_2437_43646# a_11827_44484# 0.013953f
C35937 a_1667_45002# a_n2661_43370# 0.01f
C35938 a_3232_43370# a_5837_45028# 0.01175f
C35939 a_3357_43084# a_21005_45260# 1.78e-20
C35940 a_21513_45002# a_22223_45036# 7.29e-20
C35941 a_5147_45002# a_n2293_42834# 1.41e-21
C35942 a_19479_31679# a_21101_45002# 5.63e-19
C35943 a_9223_42460# a_8270_45546# 2.21e-19
C35944 a_17324_43396# a_n357_42282# 1.48e-20
C35945 a_8605_42826# a_526_44458# 0.021896f
C35946 a_13678_32519# a_13259_45724# 0.013938f
C35947 a_10149_43396# a_n443_42852# 8.96e-19
C35948 a_3537_45260# a_10227_46804# 2.05e-20
C35949 a_1307_43914# a_n443_46116# 0.442637f
C35950 a_2809_45028# a_n971_45724# 0.037351f
C35951 a_n2017_45002# a_n2312_39304# 9.89e-22
C35952 a_413_45260# a_20990_47178# 1.26e-19
C35953 a_3357_43084# a_4842_47570# 1.16e-19
C35954 a_19256_45572# a_13661_43548# 0.00171f
C35955 a_16223_45938# a_n743_46660# 1.43e-19
C35956 a_19431_45546# a_13747_46662# 0.02276f
C35957 a_2711_45572# a_11813_46116# 1.5e-19
C35958 a_n443_42852# a_1609_45822# 1.4e-19
C35959 a_n356_45724# a_603_45572# 6.01e-19
C35960 a_21076_30879# VREF 0.417978f
C35961 a_16137_43396# a_20256_42852# 1.75e-20
C35962 a_6031_43396# a_6761_42308# 3.22e-19
C35963 a_13635_43156# a_13460_43230# 0.234322f
C35964 a_13113_42826# a_5534_30871# 0.024339f
C35965 a_n97_42460# a_15764_42576# 0.174403f
C35966 a_2982_43646# a_8685_42308# 1.03e-19
C35967 a_3681_42891# a_n2293_42282# 0.012859f
C35968 CAL_N a_22469_40625# 0.007453f
C35969 a_3422_30871# C10_N_btm 0.002966f
C35970 a_17730_32519# C1_N_btm 3.84e-20
C35971 a_13657_42558# VDD 0.195727f
C35972 a_1209_47178# a_n1435_47204# 5.76e-19
C35973 a_4791_45118# a_4915_47217# 0.226891f
C35974 a_2063_45854# a_9863_47436# 0.12173f
C35975 a_18175_45572# a_11341_43940# 1.54e-21
C35976 a_5343_44458# a_8701_44490# 8.47e-20
C35977 a_2382_45260# a_2675_43914# 1.8e-20
C35978 a_n2810_45028# a_n4318_39768# 0.027945f
C35979 a_3065_45002# a_2479_44172# 5.13e-21
C35980 a_3357_43084# a_5841_44260# 2.14e-21
C35981 a_1576_42282# a_n755_45592# 0.025747f
C35982 a_1755_42282# a_n863_45724# 0.050501f
C35983 a_1184_42692# a_n357_42282# 2.11e-19
C35984 a_8568_45546# VDD 0.182812f
C35985 a_13467_32519# RST_Z 0.048761f
C35986 a_n2661_43370# a_10428_46928# 2.58e-21
C35987 a_15595_45028# a_15227_44166# 0.007902f
C35988 a_949_44458# a_n743_46660# 3.73e-20
C35989 a_742_44458# a_n2438_43548# 0.171623f
C35990 a_5343_44458# a_n2293_46634# 0.026475f
C35991 a_13720_44458# a_13661_43548# 0.122691f
C35992 a_20447_31679# a_20820_30879# 0.053904f
C35993 a_21542_45572# a_11415_45002# 5.19e-19
C35994 a_8162_45546# a_8034_45724# 0.14162f
C35995 a_8746_45002# a_5066_45546# 1.34e-19
C35996 a_6171_45002# a_13059_46348# 0.070496f
C35997 a_413_45260# a_20273_46660# 2.73e-21
C35998 a_8696_44636# a_12005_46116# 7.73e-21
C35999 a_n2661_42834# a_4883_46098# 0.019268f
C36000 a_n1761_44111# a_n746_45260# 2.69e-20
C36001 a_n1899_43946# a_n971_45724# 0.021838f
C36002 a_1414_42308# a_n2497_47436# 0.005579f
C36003 a_17595_43084# a_17303_42282# 1.12e-19
C36004 a_n2104_42282# a_n3674_38216# 0.155459f
C36005 a_n2472_42282# a_n4318_37592# 0.030006f
C36006 a_8495_42852# a_8515_42308# 2.45e-19
C36007 a_n3674_39304# a_n3565_39304# 0.128699f
C36008 a_17701_42308# a_4958_30871# 0.007602f
C36009 a_n4318_38680# a_n4334_39392# 1.76e-19
C36010 a_n4318_38216# a_n1736_42282# 1.83e-19
C36011 a_n3674_38680# COMP_P 2.55e-20
C36012 a_n2661_46634# a_n2442_46660# 0.063483f
C36013 a_n2956_39768# a_n2293_46634# 3.22e-21
C36014 a_768_44030# a_1799_45572# 9.95e-20
C36015 a_n881_46662# a_1302_46660# 1.67e-19
C36016 a_11459_47204# a_11735_46660# 0.010464f
C36017 a_18184_42460# a_19319_43548# 0.032261f
C36018 a_20679_44626# a_21398_44850# 0.086708f
C36019 a_n2661_43922# a_5495_43940# 2.85e-20
C36020 a_17970_44736# a_18079_43940# 4.64e-19
C36021 a_n2661_42834# a_5663_43940# 0.01057f
C36022 a_1307_43914# a_9396_43370# 4.91e-20
C36023 a_n2293_42834# a_4093_43548# 0.00711f
C36024 a_20835_44721# a_20980_44850# 0.057222f
C36025 a_20159_44458# a_20397_44484# 0.007399f
C36026 a_20640_44752# a_3422_30871# 0.006762f
C36027 a_5883_43914# a_9248_44260# 0.003192f
C36028 a_n1059_45260# a_18525_43370# 0.001977f
C36029 a_n2017_45002# a_18783_43370# 1.92e-20
C36030 a_n2661_43370# VDD 1.53673f
C36031 a_5934_30871# C6_P_btm 0.004563f
C36032 a_6123_31319# C4_P_btm 0.132906f
C36033 a_2982_43646# a_12861_44030# 2.08e-20
C36034 a_8685_43396# a_2063_45854# 9.17e-20
C36035 a_n97_42460# a_13507_46334# 1.31e-19
C36036 a_5883_43914# a_8016_46348# 2.29e-20
C36037 a_8103_44636# a_8199_44636# 0.256009f
C36038 a_6298_44484# a_5937_45572# 0.036004f
C36039 a_2680_45002# a_1609_45822# 1.31e-20
C36040 a_3232_43370# a_3316_45546# 2.28e-19
C36041 a_3065_45002# a_n443_42852# 0.022494f
C36042 a_2382_45260# a_2277_45546# 0.00187f
C36043 a_5745_43940# a_768_44030# 9.71e-20
C36044 a_20835_44721# a_19692_46634# 1.53e-19
C36045 a_14673_44172# a_13059_46348# 0.108306f
C36046 a_n356_44636# a_n901_46420# 9.91e-21
C36047 a_19787_47423# VDD 0.256911f
C36048 a_18057_42282# a_7174_31319# 2.5e-20
C36049 a_17303_42282# a_21887_42336# 0.001033f
C36050 a_5932_42308# a_1177_38525# 1.83e-19
C36051 a_19332_42282# a_13258_32519# 7.57e-19
C36052 a_5742_30871# a_n3565_39304# 5.51e-21
C36053 a_n743_46660# a_5497_46414# 0.005602f
C36054 a_5807_45002# a_13759_46122# 0.022269f
C36055 a_n2661_46634# a_8953_45546# 8.33e-19
C36056 a_n1925_46634# a_6419_46155# 4.08e-20
C36057 a_12549_44172# a_17957_46116# 8.35e-19
C36058 a_13747_46662# a_12594_46348# 1.1e-19
C36059 a_n2312_40392# a_n1925_42282# 0.002171f
C36060 a_4883_46098# a_5066_45546# 0.00636f
C36061 a_11599_46634# a_12005_46436# 2.27e-19
C36062 a_13487_47204# a_14180_46482# 1.57e-20
C36063 a_n237_47217# a_n755_45592# 0.286948f
C36064 a_n971_45724# a_1848_45724# 6.57e-22
C36065 a_327_47204# a_n1099_45572# 1.03e-21
C36066 a_584_46384# a_n2293_45546# 0.029113f
C36067 a_n785_47204# a_310_45028# 9.87e-21
C36068 a_2107_46812# a_3147_46376# 0.010901f
C36069 a_n2661_46098# a_1208_46090# 0.023477f
C36070 a_6755_46942# a_765_45546# 0.002909f
C36071 a_12469_46902# a_12978_47026# 2.6e-19
C36072 a_11901_46660# a_12347_46660# 2.28e-19
C36073 a_11735_46660# a_12925_46660# 2.56e-19
C36074 a_949_44458# a_1847_42826# 3.24e-19
C36075 a_1414_42308# a_1568_43370# 0.01352f
C36076 a_5013_44260# a_n97_42460# 1.01e-19
C36077 a_21115_43940# a_14021_43940# 1.8e-20
C36078 a_1467_44172# a_1756_43548# 0.100052f
C36079 a_9313_44734# a_19268_43646# 1.06e-20
C36080 a_n2661_44458# a_7765_42852# 5.2e-21
C36081 a_742_44458# a_2075_43172# 0.002798f
C36082 a_n3674_39768# a_n2433_43396# 0.002677f
C36083 a_n1644_44306# a_n4318_39304# 1.35e-19
C36084 a_n2293_42834# a_5457_43172# 1.98e-19
C36085 a_n913_45002# a_961_42354# 4.8e-20
C36086 en_comp a_n1630_35242# 2.31448f
C36087 a_n1059_45260# a_1149_42558# 1.69e-19
C36088 a_n2017_45002# a_1221_42558# 4.86e-19
C36089 a_2998_44172# VDD 0.362233f
C36090 C9_N_btm VCM 6.06251f
C36091 C10_N_btm VREF_GND 10.3207f
C36092 a_11823_42460# a_15903_45785# 2.67e-19
C36093 a_9241_45822# a_9159_45572# 5.37e-19
C36094 a_13249_42308# a_14033_45822# 0.006215f
C36095 a_5025_43940# a_1823_45246# 8.65e-20
C36096 a_19319_43548# a_12741_44636# 3.83e-20
C36097 a_n4318_38680# a_n2312_38680# 0.023332f
C36098 a_n901_43156# a_n2438_43548# 3.58e-21
C36099 a_n2661_42282# a_n2956_39304# 5.57e-20
C36100 a_20107_46660# VDD 0.442554f
C36101 a_n2840_46090# a_n2956_39304# 0.158668f
C36102 a_765_45546# a_8049_45260# 6.27e-19
C36103 a_3483_46348# a_13925_46122# 2.92e-19
C36104 a_167_45260# a_2324_44458# 0.001084f
C36105 a_8349_46414# a_9625_46129# 7.25e-20
C36106 a_8199_44636# a_8953_45546# 0.71291f
C36107 a_8016_46348# a_9569_46155# 0.044705f
C36108 a_n4064_40160# a_n4064_37984# 0.067467f
C36109 a_10807_43548# a_10991_42826# 0.01427f
C36110 a_11750_44172# a_10796_42968# 1.07e-21
C36111 a_n2293_43922# a_196_42282# 1.63e-19
C36112 a_n356_44636# a_6171_42473# 1.17e-19
C36113 a_10057_43914# a_10533_42308# 7.44e-20
C36114 a_18494_42460# a_7174_31319# 0.023968f
C36115 a_18184_42460# a_21335_42336# 8.18e-20
C36116 a_11967_42832# a_15597_42852# 0.004349f
C36117 a_6293_42852# a_5837_43396# 3.72e-20
C36118 a_4915_47217# DATA[3] 0.07179f
C36119 a_5129_47502# DATA[2] 8.34e-20
C36120 a_19963_31679# C10_N_btm 2.25e-20
C36121 a_20447_31679# C8_N_btm 5.41e-20
C36122 a_15681_43442# VDD 0.159054f
C36123 a_2711_45572# a_18287_44626# 1.79e-20
C36124 a_7499_43078# a_4223_44672# 0.02232f
C36125 a_15903_45785# a_16321_45348# 1.49e-19
C36126 a_2680_45002# a_3065_45002# 0.13328f
C36127 a_2382_45260# a_3429_45260# 0.011518f
C36128 a_2274_45254# a_3537_45260# 3.29e-20
C36129 a_n4315_30879# a_n2312_40392# 0.389397f
C36130 a_458_43396# a_n443_42852# 0.023429f
C36131 a_5111_42852# a_4185_45028# 0.001197f
C36132 a_22315_44484# RST_Z 5.65e-20
C36133 a_2307_45899# VDD 7.28e-19
C36134 a_11652_45724# a_5807_45002# 7.11e-20
C36135 a_6194_45824# a_2107_46812# 1.15e-20
C36136 a_15765_45572# a_11453_44696# 5.36e-20
C36137 a_15861_45028# a_4883_46098# 3.69e-21
C36138 a_18175_45572# a_16327_47482# 0.346603f
C36139 a_19431_45546# a_11599_46634# 0.056971f
C36140 a_2437_43646# a_4700_47436# 0.007905f
C36141 a_1667_45002# a_n2497_47436# 9.11e-20
C36142 a_n2661_45010# a_584_46384# 0.017317f
C36143 a_3357_43084# a_3785_47178# 9.76e-20
C36144 a_413_45260# a_n2109_47186# 0.027314f
C36145 en_comp a_n971_45724# 5.07e-20
C36146 a_n1177_43370# a_n3674_37592# 4.34e-22
C36147 a_n97_42460# a_196_42282# 0.002328f
C36148 a_15743_43084# a_19339_43156# 0.128224f
C36149 a_5649_42852# a_10083_42826# 3.09e-20
C36150 a_4361_42308# a_10796_42968# 1.44e-19
C36151 a_743_42282# a_12089_42308# 0.016016f
C36152 a_11341_43940# a_15486_42560# 2.91e-21
C36153 a_n3674_39768# a_n4064_40160# 0.139482f
C36154 a_15493_43940# a_14113_42308# 1.63e-20
C36155 a_15368_46634# CLK 5.78e-20
C36156 a_n4064_37984# a_n4064_37440# 0.061238f
C36157 VDAC_Pi VDAC_Ni 3.18068f
C36158 COMP_P VDD 3.48893f
C36159 a_21101_45002# a_20193_45348# 1.15e-19
C36160 a_n2661_43370# a_n699_43396# 8.19e-19
C36161 a_9482_43914# a_5891_43370# 0.005232f
C36162 a_18315_45260# a_18545_45144# 0.004937f
C36163 a_5691_45260# a_n2661_43922# 5.88e-20
C36164 a_3232_43370# a_n2661_42834# 0.127534f
C36165 a_3357_43084# a_20835_44721# 5.14e-21
C36166 a_6171_45002# a_11649_44734# 8.52e-20
C36167 a_5193_42852# a_n357_42282# 0.00356f
C36168 a_11323_42473# a_9290_44172# 0.006277f
C36169 a_14539_43914# a_12861_44030# 0.02276f
C36170 a_n2661_43922# SMPL_ON_P 0.002089f
C36171 a_n4318_40392# a_n2312_40392# 0.025284f
C36172 a_13076_44458# a_11599_46634# 8.18e-23
C36173 a_5437_45600# a_5937_45572# 3.8e-19
C36174 a_8162_45546# a_8016_46348# 0.001995f
C36175 a_2711_45572# a_15682_46116# 0.001308f
C36176 a_6171_45002# a_7577_46660# 3.93e-21
C36177 a_3357_43084# a_3090_45724# 0.546562f
C36178 a_20731_45938# a_19692_46634# 3.6e-19
C36179 a_n2293_42834# a_n1925_46634# 0.004172f
C36180 a_15685_45394# a_13661_43548# 4.18e-20
C36181 a_18587_45118# a_12549_44172# 5.24e-21
C36182 a_7871_42858# a_8685_42308# 1.33e-20
C36183 a_8952_43230# a_5934_30871# 0.001535f
C36184 a_4361_42308# a_4958_30871# 0.087697f
C36185 a_743_42282# a_18907_42674# 0.00626f
C36186 a_4190_30871# a_18214_42558# 0.078091f
C36187 a_13467_32519# a_17303_42282# 0.040387f
C36188 a_17538_32519# C1_N_btm 1.92e-20
C36189 a_2747_46873# a_768_44030# 0.00308f
C36190 a_n1613_43370# a_n881_46662# 1.06426f
C36191 a_12465_44636# a_13747_46662# 0.039773f
C36192 a_20990_47178# a_20916_46384# 4.4e-19
C36193 a_4883_46098# a_19321_45002# 0.026904f
C36194 a_20894_47436# a_21588_30879# 1.66e-19
C36195 a_13507_46334# a_20843_47204# 4.38e-21
C36196 a_16327_47482# a_n743_46660# 0.53683f
C36197 a_10227_46804# a_n2293_46634# 0.032913f
C36198 a_n971_45724# a_7411_46660# 0.567031f
C36199 a_n1741_47186# a_8667_46634# 4.44e-20
C36200 a_n1151_42308# a_4651_46660# 0.028941f
C36201 a_3785_47178# a_3877_44458# 5.26e-20
C36202 a_2063_45854# a_5907_46634# 1.01e-19
C36203 a_14797_45144# a_15037_43940# 1.29e-20
C36204 a_n699_43396# a_2998_44172# 0.127437f
C36205 a_15861_45028# a_16243_43396# 5.52e-22
C36206 a_4223_44672# a_3600_43914# 0.00242f
C36207 a_n2293_43922# a_13296_44484# 3.07e-19
C36208 a_n2433_44484# a_n3674_39768# 0.003677f
C36209 a_8696_44636# a_16547_43609# 2.74e-20
C36210 a_1307_43914# a_10867_43940# 0.001506f
C36211 a_n2129_44697# a_n4318_39768# 1.04e-19
C36212 a_n913_45002# a_2982_43646# 0.498826f
C36213 a_n967_45348# a_n1557_42282# 0.092498f
C36214 a_n2017_45002# a_3626_43646# 0.023645f
C36215 a_3357_43084# a_6547_43396# 8.19e-19
C36216 a_n3420_38528# a_n2956_38216# 8.07e-19
C36217 a_n2302_38778# a_n2810_45572# 0.001992f
C36218 a_4574_45260# VDD 0.122256f
C36219 COMP_P a_22469_39537# 0.0359f
C36220 a_13807_45067# a_3483_46348# 2.62e-19
C36221 a_17801_45144# a_12741_44636# 3.91e-19
C36222 a_15433_44458# a_6755_46942# 0.006016f
C36223 a_12607_44458# a_13059_46348# 0.033056f
C36224 a_n984_44318# a_n2438_43548# 2.41e-21
C36225 a_3232_43370# a_5066_45546# 0.00301f
C36226 a_8953_45002# a_526_44458# 1.35e-19
C36227 a_3537_45260# a_8034_45724# 1.54e-20
C36228 a_n2661_43370# a_7920_46348# 1.68e-20
C36229 a_7418_45067# a_5937_45572# 9.73e-20
C36230 a_n1190_43762# a_n2497_47436# 4.44e-19
C36231 a_n1699_43638# a_n971_45724# 0.001253f
C36232 a_3318_42354# a_7174_31319# 4.88e-21
C36233 a_n3674_38680# a_n4209_39304# 8.12e-21
C36234 a_9803_42558# a_9885_42308# 0.003935f
C36235 a_n3674_37592# a_n4334_39616# 6.44e-20
C36236 a_n2497_47436# VDD 1.33346f
C36237 a_12549_44172# a_11415_45002# 0.028008f
C36238 a_3877_44458# a_3090_45724# 0.23348f
C36239 a_20916_46384# a_20273_46660# 2.16e-19
C36240 a_10554_47026# a_10249_46116# 0.023301f
C36241 a_10623_46897# a_6755_46942# 0.008749f
C36242 a_7927_46660# a_8035_47026# 0.057222f
C36243 a_7411_46660# a_8023_46660# 3.82e-19
C36244 a_5807_45002# a_16434_46660# 9.16e-19
C36245 a_n881_46662# a_n2293_46098# 0.291354f
C36246 a_n1613_43370# a_n2157_46122# 0.296124f
C36247 a_4883_46098# a_5068_46348# 0.031466f
C36248 a_n1151_42308# a_n1379_46482# 3.56e-19
C36249 a_n237_47217# a_835_46155# 3.57e-20
C36250 a_12861_44030# a_14493_46090# 7.43e-20
C36251 a_13487_47204# a_13925_46122# 1.5e-19
C36252 a_4915_47217# a_6945_45028# 0.207881f
C36253 a_14311_47204# a_13759_46122# 2.53e-21
C36254 a_10227_46804# a_9625_46129# 4.82e-19
C36255 a_11599_46634# a_12594_46348# 0.085826f
C36256 a_20567_45036# a_20556_43646# 6.02e-22
C36257 a_21359_45002# a_4190_30871# 3.76e-20
C36258 a_10440_44484# a_10341_43396# 2.81e-20
C36259 a_10057_43914# a_9885_43646# 8.16e-19
C36260 a_n2661_43370# a_n4318_38680# 0.001014f
C36261 a_n2661_43922# a_3080_42308# 3.25e-20
C36262 a_n2661_42834# a_4905_42826# 3.66e-20
C36263 a_5891_43370# a_6031_43396# 0.01824f
C36264 a_11827_44484# a_21259_43561# 4.17e-22
C36265 a_n2293_42834# a_685_42968# 0.006422f
C36266 a_1307_43914# a_13635_43156# 2.74e-20
C36267 a_14537_43396# a_5342_30871# 1.75e-19
C36268 a_7499_43078# a_5742_30871# 0.019993f
C36269 a_2711_45572# a_17124_42282# 1.5e-21
C36270 a_11691_44458# a_16823_43084# 5.66e-20
C36271 a_3232_43370# a_n2293_42282# 0.00771f
C36272 a_n1059_45260# a_7309_42852# 0.006756f
C36273 a_2382_45260# a_3059_42968# 6.58e-20
C36274 a_2711_45572# a_13904_45546# 0.021385f
C36275 a_5495_43940# a_5164_46348# 9.57e-20
C36276 a_15433_44458# a_8049_45260# 4.08e-21
C36277 a_6298_44484# a_n443_42852# 2.15e-20
C36278 a_15037_43940# a_14976_45028# 3.42e-20
C36279 a_14761_44260# a_13059_46348# 8.03e-20
C36280 a_16977_43638# a_13661_43548# 1.71e-20
C36281 a_6765_43638# a_4646_46812# 0.043651f
C36282 a_12429_44172# a_11415_45002# 1.15e-21
C36283 a_10949_43914# a_12741_44636# 7.98e-20
C36284 a_2437_43646# DATA[2] 0.046972f
C36285 a_22959_45572# RST_Z 0.001363f
C36286 a_6682_46987# VDD 6.34e-20
C36287 a_7174_31319# C10_N_btm 1.34e-19
C36288 a_n4064_40160# C0_P_btm 3.38e-19
C36289 a_n743_46660# a_n356_45724# 0.223429f
C36290 a_n2661_46098# a_n2661_45546# 0.011799f
C36291 a_10623_46897# a_8049_45260# 9.22e-20
C36292 a_1123_46634# a_n755_45592# 1.46e-19
C36293 a_948_46660# a_n357_42282# 1.33e-19
C36294 a_n2293_46634# a_n906_45572# 5.29e-19
C36295 a_19466_46812# a_19900_46494# 2.79e-19
C36296 a_13059_46348# a_10903_43370# 0.11738f
C36297 a_15227_44166# a_21137_46414# 0.081665f
C36298 a_19692_46634# a_20075_46420# 5.36e-19
C36299 a_765_45546# a_8953_45546# 3.61e-19
C36300 a_14513_46634# a_13925_46122# 2.11e-19
C36301 a_14180_46812# a_14493_46090# 1.41e-20
C36302 a_18834_46812# a_6945_45028# 1.91e-20
C36303 a_16292_46812# a_10809_44734# 0.005743f
C36304 a_14035_46660# a_14275_46494# 3.12e-19
C36305 a_n2472_46090# a_n1853_46287# 8.45e-19
C36306 a_n2293_46098# a_n2157_46122# 0.015455f
C36307 a_644_44056# a_791_42968# 3.17e-20
C36308 a_18326_43940# a_18525_43370# 0.003065f
C36309 a_n1917_43396# a_n1557_42282# 7.04e-19
C36310 a_n97_42460# a_4699_43561# 0.025323f
C36311 a_15493_43940# a_15781_43660# 0.049304f
C36312 a_18451_43940# a_18429_43548# 0.001082f
C36313 a_15493_43396# a_17499_43370# 0.038093f
C36314 a_11967_42832# a_18083_42858# 0.472348f
C36315 a_18588_44850# a_18249_42858# 1.79e-21
C36316 a_n4318_39768# a_n2840_42826# 5.83e-21
C36317 a_1568_43370# VDD 0.433732f
C36318 a_7499_43078# a_n2293_42834# 0.352878f
C36319 a_8696_44636# a_6171_45002# 0.070776f
C36320 a_21188_45572# a_19963_31679# 4.63e-19
C36321 a_20731_45938# a_3357_43084# 0.005715f
C36322 a_20841_45814# a_21297_45572# 4.2e-19
C36323 a_13678_32519# a_20202_43084# 0.027425f
C36324 a_13467_32519# a_20820_30879# 0.053319f
C36325 a_5342_30871# a_3090_45724# 0.001809f
C36326 a_n2840_42282# a_n2312_38680# 2.73e-20
C36327 a_n1736_42282# a_n2956_39768# 3.63e-20
C36328 a_n4318_38216# a_n2442_46660# 0.023718f
C36329 COMP_P a_22612_30879# 3.57e-19
C36330 a_3626_43646# a_526_44458# 0.022127f
C36331 a_1241_43940# a_n755_45592# 3.29e-21
C36332 a_11322_45546# a_11599_46634# 1.09e-19
C36333 a_12427_45724# a_12861_44030# 0.002445f
C36334 a_13163_45724# a_13381_47204# 4.49e-21
C36335 a_11823_42460# a_13717_47436# 1.19e-20
C36336 a_2324_44458# a_n863_45724# 0.01106f
C36337 a_5937_45572# a_n443_42852# 5.42e-20
C36338 a_15743_43084# a_22591_43396# 0.016556f
C36339 a_8685_43396# a_10083_42826# 0.007757f
C36340 a_2982_43646# a_20922_43172# 0.004571f
C36341 a_16823_43084# a_4190_30871# 0.004047f
C36342 a_3626_43646# a_19164_43230# 2.65e-20
C36343 a_3422_30871# a_17531_42308# 2.58e-20
C36344 a_4235_43370# a_4156_43218# 9.61e-19
C36345 a_1568_43370# a_873_42968# 1.46e-20
C36346 a_3080_42308# a_3445_43172# 2.6e-22
C36347 a_18114_32519# C2_N_btm 1.17e-19
C36348 a_16855_45546# a_17061_44734# 2.71e-21
C36349 a_15415_45028# a_11691_44458# 0.002488f
C36350 a_16751_45260# a_11827_44484# 7.2e-21
C36351 a_8696_44636# a_14673_44172# 0.017655f
C36352 a_8560_45348# a_8704_45028# 6.84e-19
C36353 a_4574_45260# a_n699_43396# 1.24e-19
C36354 a_3537_45260# a_4743_44484# 0.01411f
C36355 a_4558_45348# a_4223_44672# 7.57e-20
C36356 a_7705_45326# a_n2661_44458# 1.38e-20
C36357 a_n1059_45260# a_16979_44734# 4.85e-22
C36358 a_n913_45002# a_14539_43914# 0.003048f
C36359 a_3357_43084# a_n356_44636# 3.56e-20
C36360 a_8649_43218# a_526_44458# 0.002066f
C36361 a_18083_42858# a_13259_45724# 0.002348f
C36362 a_5755_42852# a_n755_45592# 6.41e-21
C36363 a_7227_42852# a_n357_42282# 0.185359f
C36364 a_11823_42460# a_14035_46660# 0.003215f
C36365 a_13159_45002# a_12549_44172# 4.23e-20
C36366 a_13348_45260# a_12891_46348# 0.097519f
C36367 a_13017_45260# a_768_44030# 0.031385f
C36368 a_n143_45144# a_n743_46660# 0.00133f
C36369 a_3065_45002# a_n2661_46634# 3.58e-21
C36370 a_2274_45254# a_n2293_46634# 0.018017f
C36371 a_7276_45260# a_5807_45002# 1.33e-20
C36372 a_413_45260# a_n1925_46634# 0.02974f
C36373 a_16019_45002# a_n881_46662# 5.4e-20
C36374 a_1307_43914# a_n1613_43370# 0.056988f
C36375 a_11827_44484# a_4915_47217# 0.002572f
C36376 a_22705_37990# VDD 0.085164f
C36377 a_n699_43396# a_n2497_47436# 0.355158f
C36378 a_n2267_44484# a_n746_45260# 0.003717f
C36379 a_n2157_42858# a_n1630_35242# 2.26e-19
C36380 a_n1991_42858# a_n3674_37592# 6.3e-20
C36381 a_12895_43230# a_13291_42460# 0.002402f
C36382 a_743_42282# a_5267_42460# 0.010719f
C36383 a_10341_43396# a_15486_42560# 4.67e-21
C36384 a_9145_43396# a_13657_42308# 1.47e-19
C36385 a_6945_45028# DATA[5] 0.047689f
C36386 a_n4209_39304# VDD 0.984278f
C36387 a_18143_47464# a_18780_47178# 0.001596f
C36388 a_10227_46804# a_18597_46090# 0.07604f
C36389 a_n443_46116# a_n1613_43370# 0.410263f
C36390 a_13717_47436# a_22959_47212# 8.82e-19
C36391 a_16241_47178# a_13507_46334# 6.13e-21
C36392 a_15811_47375# a_4883_46098# 1.03e-21
C36393 a_12861_44030# a_11453_44696# 0.173308f
C36394 a_4791_45118# a_n881_46662# 0.429542f
C36395 a_n1435_47204# a_n2312_40392# 0.002491f
C36396 a_11599_46634# a_12465_44636# 0.018625f
C36397 a_n2833_47464# a_n2840_46634# 0.019713f
C36398 a_2063_45854# a_768_44030# 0.027746f
C36399 a_4915_47217# a_3411_47243# 2.39e-21
C36400 a_11823_42460# a_9145_43396# 0.146085f
C36401 a_10057_43914# a_n2661_43922# 0.034016f
C36402 a_8975_43940# a_n2661_42834# 0.083892f
C36403 a_18248_44752# a_9313_44734# 1.88e-21
C36404 a_20193_45348# a_20766_44850# 4.03e-19
C36405 a_5837_45028# a_5495_43940# 4.33e-21
C36406 a_9482_43914# a_10807_43548# 0.002194f
C36407 a_13017_45260# a_13483_43940# 3.52e-21
C36408 a_10193_42453# a_14955_43396# 4.69e-21
C36409 a_2711_45572# a_19268_43646# 3.71e-19
C36410 a_375_42282# a_n2661_42282# 2.72e-19
C36411 a_18184_42460# a_3422_30871# 0.649102f
C36412 a_7499_43078# a_10849_43646# 0.003558f
C36413 a_18450_45144# a_11967_42832# 1.01e-19
C36414 a_11827_44484# a_18681_44484# 7.17e-19
C36415 a_22775_42308# a_13259_45724# 0.007982f
C36416 a_13575_42558# a_n443_42852# 2.2e-21
C36417 a_21513_45002# a_6945_45028# 1.8e-20
C36418 a_3357_43084# a_20075_46420# 4.81e-21
C36419 a_5111_44636# a_5497_46414# 3.91e-19
C36420 a_4927_45028# a_5204_45822# 4.9e-19
C36421 a_5691_45260# a_5164_46348# 0.00167f
C36422 a_3537_45260# a_8016_46348# 5.67e-20
C36423 a_2437_43646# a_21137_46414# 3.15e-23
C36424 a_14815_43914# a_n2293_46634# 0.057388f
C36425 a_11967_42832# a_12549_44172# 0.193926f
C36426 a_11691_44458# a_15368_46634# 0.002402f
C36427 a_17517_44484# a_5807_45002# 1.9e-19
C36428 a_7229_43940# a_3483_46348# 0.03702f
C36429 a_n2661_43922# a_n2438_43548# 0.06887f
C36430 a_20567_45036# a_19692_46634# 5.15e-19
C36431 a_1307_43914# a_n2293_46098# 0.107603f
C36432 a_2123_42473# a_5934_30871# 1.01e-20
C36433 a_16877_42852# a_17124_42282# 4.18e-19
C36434 a_3318_42354# a_5932_42308# 4.34e-21
C36435 a_5379_42460# a_5421_42558# 0.002327f
C36436 a_5267_42460# a_5755_42308# 0.055455f
C36437 a_13678_32519# C5_N_btm 1.22e-19
C36438 CAL_P a_22609_38406# 2.83e-19
C36439 a_22469_39537# a_22705_37990# 3.12e-20
C36440 a_4883_46098# a_13059_46348# 0.097406f
C36441 a_13507_46334# a_16721_46634# 0.00543f
C36442 a_18597_46090# a_17339_46660# 0.018491f
C36443 a_10227_46804# a_19123_46287# 9.33e-20
C36444 a_11599_46634# a_20528_46660# 2.63e-20
C36445 a_18143_47464# a_18285_46348# 2.02e-19
C36446 a_16327_47482# a_20841_46902# 8.93e-20
C36447 a_18780_47178# a_765_45546# 2.8e-19
C36448 a_12861_44030# a_17639_46660# 0.033515f
C36449 a_n443_46116# a_n2293_46098# 0.251135f
C36450 a_584_46384# a_1138_42852# 0.491749f
C36451 a_n971_45724# a_4185_45028# 4.59e-19
C36452 a_n237_47217# a_3483_46348# 0.090759f
C36453 a_n1151_42308# a_n1076_46494# 0.023834f
C36454 a_1239_47204# a_167_45260# 2.52e-21
C36455 a_2124_47436# a_1823_45246# 9.81e-21
C36456 a_2063_45854# a_1176_45822# 2.25e-19
C36457 a_n1741_47186# a_5204_45822# 4.65e-20
C36458 a_12549_44172# a_12251_46660# 0.001402f
C36459 a_n2661_46634# a_10249_46116# 0.055133f
C36460 a_12891_46348# a_12991_46634# 0.018656f
C36461 a_n743_46660# a_8667_46634# 9.34e-20
C36462 a_3699_46634# a_3877_44458# 0.087244f
C36463 a_2443_46660# a_4817_46660# 2.35e-21
C36464 a_2864_46660# a_3055_46660# 4.61e-19
C36465 a_2959_46660# a_4646_46812# 8.56e-21
C36466 a_5807_45002# a_8189_46660# 7.17e-19
C36467 a_10193_42453# a_19326_42852# 1.39e-19
C36468 a_n2840_43914# a_n3674_39768# 0.022122f
C36469 a_2127_44172# a_895_43940# 0.132679f
C36470 a_1414_42308# a_2889_44172# 0.128883f
C36471 a_1467_44172# a_2998_44172# 1.71e-20
C36472 a_11967_42832# a_12429_44172# 6.2e-19
C36473 a_5891_43370# a_6671_43940# 1.15e-20
C36474 a_n699_43396# a_1568_43370# 0.004191f
C36475 a_n2472_43914# a_n4318_39768# 3.22e-19
C36476 a_n913_45002# a_7871_42858# 0.005608f
C36477 a_n2017_45002# a_8037_42858# 6.62e-20
C36478 a_n1059_45260# a_7765_42852# 0.004965f
C36479 a_5883_43914# VDD 0.859221f
C36480 a_21335_42336# RST_Z 1.97e-20
C36481 a_20637_44484# a_11415_45002# 2.19e-20
C36482 a_9672_43914# a_3090_45724# 0.004104f
C36483 a_5343_44458# a_8049_45260# 3.51e-20
C36484 a_18450_45144# a_13259_45724# 3.75e-19
C36485 a_9313_44734# a_2324_44458# 0.001086f
C36486 a_14358_43442# a_12465_44636# 3.52e-20
C36487 a_14537_43646# a_10227_46804# 2.7e-19
C36488 a_n2157_42858# a_n971_45724# 2.88e-19
C36489 a_10210_45822# CLK 5.07e-19
C36490 a_n3420_39616# a_n3420_39072# 0.115485f
C36491 a_n3565_39590# a_n4064_39072# 0.033734f
C36492 a_n4064_39616# a_n3565_39304# 0.028003f
C36493 a_n2104_46634# VDD 0.286113f
C36494 a_5932_42308# C10_N_btm 1.34e-19
C36495 a_6123_31319# C5_N_btm 0.022099f
C36496 a_5934_30871# C3_N_btm 0.011274f
C36497 a_8270_45546# a_3483_46348# 0.058754f
C36498 a_765_45546# a_18285_46348# 5.85e-19
C36499 a_12549_44172# a_13259_45724# 0.110646f
C36500 a_2107_46812# a_3873_46454# 4.52e-19
C36501 a_5807_45002# a_12379_46436# 0.006522f
C36502 a_6755_46942# a_8349_46414# 0.001141f
C36503 a_9863_46634# a_10355_46116# 0.00109f
C36504 a_10150_46912# a_9823_46155# 5.05e-19
C36505 a_10249_46116# a_8199_44636# 0.002313f
C36506 a_20679_44626# a_20556_43646# 1.59e-20
C36507 a_11967_42832# a_21855_43396# 0.002687f
C36508 a_18248_44752# a_18599_43230# 2.16e-21
C36509 a_18989_43940# a_18083_42858# 9.56e-20
C36510 a_20640_44752# a_21487_43396# 1.18e-19
C36511 a_19279_43940# a_4190_30871# 4.5e-20
C36512 a_n2661_42834# a_2905_42968# 6.38e-21
C36513 a_18443_44721# a_18249_42858# 3.84e-21
C36514 a_n2293_43922# a_1847_42826# 1.69e-20
C36515 a_1307_43914# a_3905_42558# 4.45e-19
C36516 a_n356_44636# a_5342_30871# 0.133551f
C36517 a_n2293_42834# a_n1329_42308# 0.002332f
C36518 a_5891_43370# a_10796_42968# 8.14e-20
C36519 a_18184_42460# a_18504_43218# 3.21e-21
C36520 a_n2661_42282# a_6655_43762# 4.97e-19
C36521 a_22591_44484# a_15743_43084# 1.16e-20
C36522 a_20512_43084# a_19700_43370# 7.17e-19
C36523 a_17478_45572# a_18479_45785# 3.4e-19
C36524 a_2711_45572# a_10951_45334# 5.77e-20
C36525 a_15861_45028# a_18341_45572# 9.93e-20
C36526 a_6511_45714# a_7276_45260# 1.03e-19
C36527 a_7227_45028# a_6171_45002# 0.029883f
C36528 a_6667_45809# a_5205_44484# 1.28e-19
C36529 a_3775_45552# a_3232_43370# 1.51e-20
C36530 a_6598_45938# a_6431_45366# 0.001277f
C36531 a_11823_42460# a_n1059_45260# 0.100641f
C36532 a_4933_42558# a_4791_45118# 0.001758f
C36533 a_22521_40599# CAL_P 6.35e-19
C36534 CAL_N a_22609_38406# 0.204621f
C36535 a_n4209_37414# C7_P_btm 1.43e-20
C36536 a_n3565_37414# C9_P_btm 3.18e-20
C36537 a_3726_37500# a_n923_35174# 0.029905f
C36538 VDAC_Ni RST_Z 1.24e-19
C36539 a_n1441_43940# a_n2293_45546# 1.11e-19
C36540 a_2479_44172# a_n443_42852# 0.035023f
C36541 a_16823_43084# a_15227_44166# 0.022136f
C36542 a_5111_42852# a_5257_43370# 0.013892f
C36543 a_743_42282# a_3090_45724# 1.62e-19
C36544 a_9569_46155# VDD 0.19288f
C36545 a_6472_45840# a_n237_47217# 4e-19
C36546 a_6667_45809# a_n971_45724# 9.13e-19
C36547 a_765_45546# a_1609_45822# 0.021736f
C36548 a_9625_46129# a_8034_45724# 1.73e-19
C36549 a_8349_46414# a_8049_45260# 2.39e-20
C36550 a_8199_44636# a_8781_46436# 2.2e-19
C36551 a_6945_45028# a_10809_44734# 0.953135f
C36552 a_n3565_38502# a_n4209_37414# 0.029366f
C36553 a_n4209_38502# a_n3565_37414# 0.030019f
C36554 a_21076_30879# a_20692_30879# 0.117886f
C36555 a_n1761_44111# a_n1630_35242# 0.060838f
C36556 a_n809_44244# a_n784_42308# 1.32e-20
C36557 a_6547_43396# a_743_42282# 3.34e-20
C36558 a_15095_43370# a_16243_43396# 2.69e-21
C36559 a_n97_42460# a_1847_42826# 2.77e-20
C36560 a_13565_43940# a_12545_42858# 1.31e-20
C36561 a_n1557_42282# a_n1853_43023# 1.74e-20
C36562 a_14205_43396# a_16547_43609# 8.78e-22
C36563 a_14955_43396# a_16137_43396# 7.94e-20
C36564 a_10807_43548# a_11301_43218# 0.001467f
C36565 a_10341_43396# a_13837_43396# 7.41e-20
C36566 a_8685_43396# a_16664_43396# 1.93e-19
C36567 a_n881_46662# DATA[3] 0.001196f
C36568 a_133_43172# VDD 8.22e-19
C36569 a_n2956_37592# a_n3690_38304# 1.91e-20
C36570 a_n2810_45028# a_n3420_37984# 5.66e-21
C36571 a_10193_42453# a_n2661_42834# 0.034215f
C36572 a_16019_45002# a_1307_43914# 0.01609f
C36573 a_8696_44636# a_12607_44458# 0.005383f
C36574 a_10180_45724# a_n2661_43922# 1.65e-19
C36575 a_327_44734# a_n2661_43370# 0.035472f
C36576 a_3357_43084# a_20567_45036# 4.77e-19
C36577 a_21513_45002# a_11827_44484# 0.010541f
C36578 a_5691_45260# a_5837_45028# 0.171361f
C36579 a_6709_45028# a_6517_45366# 5.76e-19
C36580 a_19479_31679# a_21005_45260# 3.22e-19
C36581 a_5755_42308# a_3090_45724# 1.13e-20
C36582 a_n2302_39866# a_n2312_38680# 1.63e-19
C36583 a_17499_43370# a_n357_42282# 1.53e-19
C36584 a_8037_42858# a_526_44458# 0.01672f
C36585 a_9885_43396# a_n443_42852# 0.001051f
C36586 a_413_45260# a_20894_47436# 8.97e-20
C36587 a_1423_45028# a_n1151_42308# 1.11e-19
C36588 a_1307_43914# a_4791_45118# 0.027544f
C36589 a_n2017_45002# a_n2312_40392# 1.3e-21
C36590 a_n913_45002# a_11453_44696# 1.71e-20
C36591 a_19431_45546# a_13661_43548# 4.64e-19
C36592 a_6472_45840# a_8270_45546# 1.23e-19
C36593 a_19256_45572# a_5807_45002# 0.015716f
C36594 a_18341_45572# a_19321_45002# 0.001456f
C36595 a_18691_45572# a_13747_46662# 0.030666f
C36596 a_2711_45572# a_11735_46660# 1.14e-19
C36597 a_20273_45572# a_12549_44172# 1.54e-20
C36598 a_n356_45724# a_509_45572# 9.76e-19
C36599 a_16137_43396# a_19326_42852# 1.63e-20
C36600 a_2905_42968# a_n2293_42282# 0.001495f
C36601 a_12545_42858# a_5534_30871# 0.17182f
C36602 a_2982_43646# a_8325_42308# 1.03e-19
C36603 a_n97_42460# a_15486_42560# 0.055334f
C36604 a_12895_43230# a_13460_43230# 7.99e-20
C36605 a_3626_43646# a_4169_42308# 6.63e-19
C36606 a_20820_30879# VCM 0.05604f
C36607 a_21076_30879# VIN_N 0.068195f
C36608 a_3422_30871# C9_N_btm 0.003737f
C36609 a_17730_32519# C0_N_btm 3.27e-20
C36610 CAL_N a_22521_40599# 0.006786f
C36611 a_13333_42558# VDD 0.008231f
C36612 a_327_47204# a_n1435_47204# 0.001005f
C36613 a_4700_47436# a_4915_47217# 0.07122f
C36614 a_2063_45854# a_9067_47204# 1.79e-19
C36615 a_n1151_42308# a_6491_46660# 1.03e-19
C36616 a_3785_47178# a_6151_47436# 4.24e-20
C36617 a_4791_45118# a_n443_46116# 0.115639f
C36618 a_5343_44458# a_8103_44636# 0.001348f
C36619 a_10907_45822# a_11257_43940# 8.34e-20
C36620 a_16147_45260# a_11341_43940# 2.74e-20
C36621 a_16922_45042# a_9313_44734# 5.83e-19
C36622 a_3537_45260# a_1414_42308# 1.29e-19
C36623 a_2274_45254# a_2675_43914# 1.86e-20
C36624 a_413_45260# a_3600_43914# 2.35e-19
C36625 a_2680_45002# a_2479_44172# 1.33e-19
C36626 a_n913_45002# a_n3674_39768# 2.02e-20
C36627 a_1067_42314# a_n755_45592# 0.047422f
C36628 a_1576_42282# a_n357_42282# 1.92e-19
C36629 a_1606_42308# a_n863_45724# 0.20593f
C36630 a_8162_45546# VDD 0.266272f
C36631 a_15415_45028# a_15227_44166# 0.222342f
C36632 a_4743_44484# a_n2293_46634# 2.4e-20
C36633 a_18989_43940# a_12549_44172# 0.016062f
C36634 a_13720_44458# a_5807_45002# 0.001051f
C36635 a_742_44458# a_n743_46660# 3.66e-22
C36636 a_n2661_44458# a_2107_46812# 0.02628f
C36637 a_21542_45572# a_20202_43084# 7.05e-19
C36638 a_19963_31679# a_12741_44636# 2.28e-21
C36639 a_21297_45572# a_11415_45002# 2.47e-19
C36640 a_413_45260# a_20411_46873# 1.63e-20
C36641 a_15037_45618# a_2324_44458# 1.52e-19
C36642 a_8696_44636# a_10903_43370# 0.031601f
C36643 a_n998_44484# a_n1613_43370# 0.002879f
C36644 a_1467_44172# a_n2497_47436# 0.046456f
C36645 a_n2065_43946# a_n746_45260# 2.94e-21
C36646 a_n1761_44111# a_n971_45724# 0.084835f
C36647 a_16795_42852# a_17303_42282# 0.010298f
C36648 a_17595_43084# a_4958_30871# 9.74e-19
C36649 a_8495_42852# a_5934_30871# 8.72e-19
C36650 a_n3674_39304# a_n4334_39392# 0.060327f
C36651 a_n4318_38216# a_n3674_38216# 2.91597f
C36652 a_n3674_38680# a_n4318_37592# 0.084223f
C36653 a_n2840_42282# COMP_P 7.51e-20
C36654 a_n2840_46634# a_n2293_46634# 2.97e-19
C36655 a_n2661_46634# a_n2472_46634# 0.0842f
C36656 a_n2956_39768# a_n2442_46660# 6.5214f
C36657 a_n881_46662# a_1057_46660# 1.39e-19
C36658 a_n1613_43370# a_1302_46660# 0.001965f
C36659 a_4883_46098# a_7577_46660# 7.2e-20
C36660 a_10227_46804# a_6755_46942# 0.778648f
C36661 a_19778_44110# a_19319_43548# 0.003354f
C36662 a_17970_44736# a_17973_43940# 0.002178f
C36663 a_20679_44626# a_20980_44850# 9.73e-19
C36664 a_20640_44752# a_21398_44850# 0.056391f
C36665 a_17767_44458# a_18079_43940# 3.68e-19
C36666 a_n2661_43922# a_5013_44260# 7.36e-20
C36667 a_n2661_42834# a_5495_43940# 0.009774f
C36668 a_n2293_42834# a_1756_43548# 1.53e-20
C36669 a_1307_43914# a_8791_43396# 4.19e-20
C36670 a_1423_45028# a_6197_43396# 4.8e-22
C36671 a_16922_45042# a_20974_43370# 0.077191f
C36672 a_20766_44850# a_20596_44850# 2.6e-19
C36673 a_20362_44736# a_3422_30871# 3.94e-20
C36674 a_n913_45002# a_17324_43396# 7.64e-21
C36675 a_n1059_45260# a_18429_43548# 0.002978f
C36676 a_5111_44636# a_10341_43396# 0.009186f
C36677 a_5934_30871# C7_P_btm 0.007575f
C36678 a_6123_31319# C5_P_btm 0.022099f
C36679 a_5343_44458# a_8953_45546# 0.002817f
C36680 a_11827_44484# a_10809_44734# 0.029958f
C36681 a_6298_44484# a_8199_44636# 0.002319f
C36682 a_5518_44484# a_5937_45572# 4.36e-19
C36683 a_20193_45348# a_19900_46494# 8.77e-21
C36684 a_2382_45260# a_1609_45822# 0.001939f
C36685 a_7229_43940# a_n357_42282# 1.8e-20
C36686 a_2274_45254# a_2277_45546# 0.011988f
C36687 a_8560_45348# a_8049_45260# 8.56e-19
C36688 a_14581_44484# a_13059_46348# 7.41e-20
C36689 a_3820_44260# a_3877_44458# 4.75e-19
C36690 a_15301_44260# a_13661_43548# 4.13e-19
C36691 a_19279_43940# a_15227_44166# 1.77e-21
C36692 a_20679_44626# a_19692_46634# 0.010957f
C36693 a_15004_44636# a_3483_46348# 1.48e-20
C36694 a_19386_47436# VDD 0.121241f
C36695 a_19332_42282# a_19647_42308# 0.084365f
C36696 a_17531_42308# a_7174_31319# 2.13e-20
C36697 a_18214_42558# a_19511_42282# 9.74e-21
C36698 a_17303_42282# a_21335_42336# 2.99e-19
C36699 a_6123_31319# a_n3420_38528# 0.003315f
C36700 a_5934_30871# a_n3565_38502# 4.1e-21
C36701 a_15368_46634# a_15227_44166# 0.002374f
C36702 a_10249_46116# a_765_45546# 0.005411f
C36703 a_11901_46660# a_12978_47026# 1.46e-19
C36704 a_3090_45724# a_19466_46812# 1.49e-19
C36705 a_n2661_46634# a_5937_45572# 2.16e-19
C36706 a_n743_46660# a_5204_45822# 0.034798f
C36707 a_5807_45002# a_13351_46090# 0.002035f
C36708 a_n1925_46634# a_6165_46155# 6.31e-20
C36709 a_n2293_46634# a_8016_46348# 4.84e-19
C36710 a_13661_43548# a_12594_46348# 1.57e-21
C36711 a_12549_44172# a_18189_46348# 2.08e-19
C36712 a_n881_46662# a_6945_45028# 0.239384f
C36713 a_4883_46098# a_5431_46482# 2.13e-19
C36714 a_10227_46804# a_8049_45260# 0.058336f
C36715 a_n971_45724# a_997_45618# 4.51e-22
C36716 a_n746_45260# a_n755_45592# 0.172774f
C36717 a_327_47204# a_380_45546# 1.52e-21
C36718 a_n237_47217# a_n357_42282# 4.85e-21
C36719 a_n785_47204# a_n1099_45572# 1.19e-20
C36720 a_n23_47502# a_310_45028# 6.86e-20
C36721 a_n2661_46098# a_805_46414# 0.044109f
C36722 a_2107_46812# a_2804_46116# 0.008475f
C36723 a_1799_45572# a_1208_46090# 0.008066f
C36724 a_949_44458# a_791_42968# 3.01e-19
C36725 a_n1899_43946# a_n1557_42282# 1.37e-19
C36726 a_5244_44056# a_n97_42460# 2.33e-20
C36727 a_14673_44172# a_14205_43396# 7.49e-20
C36728 a_20935_43940# a_14021_43940# 7.94e-20
C36729 a_742_44458# a_1847_42826# 0.372436f
C36730 a_1467_44172# a_1568_43370# 0.055004f
C36731 a_9313_44734# a_15743_43084# 1.48048f
C36732 a_n2661_44458# a_7871_42858# 6.62e-21
C36733 a_n356_44636# a_743_42282# 0.063042f
C36734 a_9028_43914# a_9420_43940# 0.016359f
C36735 a_n3674_39768# a_n4318_39304# 2.75695f
C36736 a_1414_42308# a_1049_43396# 0.003017f
C36737 a_n2293_42834# a_5193_43172# 2.71e-19
C36738 a_n1059_45260# a_961_42354# 0.07089f
C36739 a_n967_45348# a_n3674_37592# 0.002659f
C36740 a_n913_45002# a_1184_42692# 0.031137f
C36741 a_3357_43084# a_3823_42558# 3.77e-19
C36742 a_n2956_37592# a_n1630_35242# 5.5e-19
C36743 a_n2017_45002# a_1149_42558# 4.17e-19
C36744 a_2889_44172# VDD 0.1447f
C36745 a_13527_45546# a_15037_45618# 2.92e-22
C36746 a_11823_42460# a_15599_45572# 3.42e-19
C36747 a_8746_45002# a_8696_44636# 0.058163f
C36748 a_10193_42453# a_15861_45028# 0.432483f
C36749 a_13904_45546# a_14033_45822# 0.062574f
C36750 C8_N_btm VCM 2.61094f
C36751 C9_N_btm VREF_GND 5.18245f
C36752 C10_N_btm VREF 14.773f
C36753 a_3992_43940# a_1823_45246# 1.48e-19
C36754 a_10083_42826# a_768_44030# 3.74e-20
C36755 a_n3674_39304# a_n2312_38680# 0.023501f
C36756 a_n1641_43230# a_n2438_43548# 4.44e-20
C36757 a_11341_43940# a_9290_44172# 0.040892f
C36758 a_19551_46910# VDD 0.226848f
C36759 a_17339_46660# a_8049_45260# 0.023006f
C36760 a_14180_46812# a_14180_46482# 6.29e-19
C36761 a_8270_45546# a_n357_42282# 5.72e-20
C36762 a_15227_44166# a_19597_46482# 6.67e-19
C36763 a_3483_46348# a_13759_46122# 6.81e-19
C36764 a_8016_46348# a_9625_46129# 0.128435f
C36765 a_8199_44636# a_5937_45572# 0.573373f
C36766 a_n4315_30879# a_n2302_37984# 6.48e-20
C36767 a_7174_31319# VDAC_Pi 2.22e-19
C36768 a_n4064_40160# a_n2946_37984# 2.04e-20
C36769 a_10405_44172# a_10341_42308# 5.11e-21
C36770 a_10949_43914# a_10991_42826# 3.02e-20
C36771 a_10807_43548# a_10796_42968# 0.030352f
C36772 a_11750_44172# a_10835_43094# 2e-20
C36773 a_8791_43396# a_9396_43370# 0.011032f
C36774 a_20974_43370# a_15743_43084# 6.72e-19
C36775 a_18184_42460# a_7174_31319# 0.007789f
C36776 a_n2293_43922# a_n473_42460# 8.65e-20
C36777 a_n356_44636# a_5755_42308# 2.77e-19
C36778 a_3905_42865# a_4156_43218# 7.76e-19
C36779 a_2982_43646# a_9145_43396# 1.33e-20
C36780 a_4915_47217# DATA[2] 9.44e-19
C36781 a_n443_46116# DATA[3] 1.57e-20
C36782 a_19963_31679# C9_N_btm 1.91e-20
C36783 a_20447_31679# C7_N_btm 7.54e-20
C36784 a_14621_43646# VDD 0.008139f
C36785 a_2711_45572# a_18248_44752# 8.88e-20
C36786 a_2382_45260# a_3065_45002# 0.632538f
C36787 a_413_45260# a_4558_45348# 4.69e-20
C36788 a_n229_43646# a_n443_42852# 0.001316f
C36789 a_3539_42460# a_n863_45724# 8.25e-22
C36790 a_5742_30871# a_n2312_38680# 4.94e-21
C36791 a_4520_42826# a_4185_45028# 0.012305f
C36792 a_3422_30871# RST_Z 0.0872f
C36793 a_1990_45899# VDD 0.001563f
C36794 a_15143_45578# a_12549_44172# 2.08e-21
C36795 a_5907_45546# a_2107_46812# 1.16e-20
C36796 a_15903_45785# a_11453_44696# 0.003342f
C36797 a_17478_45572# a_13507_46334# 1.05e-20
C36798 a_8696_44636# a_4883_46098# 0.023202f
C36799 a_18691_45572# a_11599_46634# 0.034093f
C36800 a_16147_45260# a_16327_47482# 0.017922f
C36801 a_14127_45572# a_10227_46804# 2.84e-19
C36802 a_18799_45938# a_12861_44030# 6.19e-20
C36803 a_2437_43646# a_4007_47204# 0.007098f
C36804 a_327_44734# a_n2497_47436# 1.11e-19
C36805 a_15682_43940# a_17124_42282# 8.07e-20
C36806 a_n2267_43396# a_n1630_35242# 2.12e-20
C36807 a_n1917_43396# a_n3674_37592# 1.93e-20
C36808 a_n97_42460# a_n473_42460# 0.096579f
C36809 a_15743_43084# a_18599_43230# 0.001457f
C36810 a_n1076_43230# a_791_42968# 4.35e-20
C36811 a_n13_43084# a_685_42968# 0.002159f
C36812 a_5649_42852# a_8952_43230# 3.14e-21
C36813 a_4361_42308# a_10835_43094# 2.74e-20
C36814 a_743_42282# a_12379_42858# 2.73e-19
C36815 a_11341_43940# a_15051_42282# 3.24e-20
C36816 a_n3674_39768# a_n4334_40480# 0.004086f
C36817 a_n4318_39768# a_n4064_40160# 0.293052f
C36818 a_8685_43396# a_10553_43218# 1.84e-19
C36819 a_19692_46634# SINGLE_ENDED 4.63e-20
C36820 a_14976_45028# CLK 4.29e-20
C36821 a_n2946_37984# a_n4064_37440# 3.78e-20
C36822 a_n4064_37984# a_n2946_37690# 3.78e-20
C36823 a_7754_39964# VDAC_Ni 0.207118f
C36824 VDAC_Pi a_7754_38636# 1.59e-19
C36825 a_7754_40130# a_3754_38470# 0.191861f
C36826 a_n4318_37592# VDD 0.919667f
C36827 a_21101_45002# a_11691_44458# 1.41e-20
C36828 a_11827_44484# a_22959_45036# 4.91e-20
C36829 a_21005_45260# a_20193_45348# 3.32e-20
C36830 a_n2661_43370# a_4223_44672# 0.001914f
C36831 a_626_44172# a_n356_44636# 0.249281f
C36832 a_10193_42453# a_20623_43914# 0.001477f
C36833 a_18315_45260# a_18450_45144# 0.008535f
C36834 a_13249_42308# a_14955_43940# 6.27e-21
C36835 a_5691_45260# a_n2661_42834# 1.59e-21
C36836 a_3357_43084# a_20679_44626# 5.72e-21
C36837 a_5111_44636# a_n2293_43922# 4.86e-20
C36838 a_3232_43370# a_11649_44734# 0.011508f
C36839 a_21363_45546# a_3422_30871# 9.12e-20
C36840 a_22775_42308# a_20202_43084# 1.98e-19
C36841 a_961_42354# a_n1925_42282# 8.52e-20
C36842 a_4649_42852# a_n357_42282# 0.00298f
C36843 a_10723_42308# a_9290_44172# 8.75e-19
C36844 a_n2661_42834# SMPL_ON_P 0.002304f
C36845 a_n2661_43922# a_n1741_47186# 1.28e-19
C36846 a_n2661_44458# a_11453_44696# 0.174607f
C36847 a_2711_45572# a_2324_44458# 0.804101f
C36848 a_8162_45546# a_7920_46348# 2.96e-19
C36849 a_11827_44484# a_n881_46662# 2.46e-20
C36850 a_20731_45938# a_19466_46812# 1.24e-20
C36851 a_6171_45002# a_7715_46873# 3.86e-20
C36852 a_3357_43084# a_15009_46634# 1.23e-20
C36853 a_2437_43646# a_15368_46634# 1.64e-19
C36854 a_3232_43370# a_7577_46660# 6.76e-22
C36855 a_5205_44484# a_5257_43370# 0.021038f
C36856 a_15060_45348# a_13661_43548# 6.77e-19
C36857 a_18479_45785# a_16388_46812# 3.13e-19
C36858 a_11652_45724# a_3483_46348# 0.035818f
C36859 a_4361_42308# a_16269_42308# 2.5e-19
C36860 a_7871_42858# a_8325_42308# 7.98e-19
C36861 a_9127_43156# a_5934_30871# 0.003851f
C36862 a_n2293_42282# a_n784_42308# 0.055588f
C36863 a_8387_43230# a_8515_42308# 7.06e-20
C36864 a_4190_30871# a_19332_42282# 0.154377f
C36865 a_743_42282# a_18727_42674# 0.006169f
C36866 a_13467_32519# a_4958_30871# 0.031235f
C36867 a_17538_32519# C0_N_btm 1.63e-20
C36868 a_12465_44636# a_13661_43548# 0.106973f
C36869 a_13507_46334# a_19594_46812# 0.007313f
C36870 a_20894_47436# a_20916_46384# 4.94e-19
C36871 a_16241_47178# a_n743_46660# 0.001102f
C36872 a_n1435_47204# a_1983_46706# 5.62e-21
C36873 a_n971_45724# a_5257_43370# 0.001362f
C36874 a_2063_45854# a_5167_46660# 6.73e-19
C36875 a_n1151_42308# a_4646_46812# 0.330834f
C36876 a_17023_45118# a_15682_43940# 8.14e-19
C36877 a_16922_45042# a_17737_43940# 6.1e-19
C36878 a_n2661_44458# a_n3674_39768# 0.037999f
C36879 a_n2433_44484# a_n4318_39768# 0.00138f
C36880 a_n699_43396# a_2889_44172# 0.006735f
C36881 a_14537_43396# a_15037_43940# 0.018234f
C36882 a_n2293_43922# a_12829_44484# 0.009626f
C36883 a_4223_44672# a_2998_44172# 0.035464f
C36884 a_13249_42308# a_5649_42852# 3.17e-20
C36885 a_1307_43914# a_10651_43940# 0.001528f
C36886 a_5111_44636# a_n97_42460# 0.211832f
C36887 a_n1059_45260# a_2982_43646# 0.020128f
C36888 en_comp a_n1557_42282# 4.48e-20
C36889 a_3357_43084# a_6765_43638# 3.46e-19
C36890 a_n4064_38528# a_n2810_45572# 2.53e-19
C36891 a_3537_45260# VDD 3.9063f
C36892 COMP_P a_22821_38993# 2.95e-19
C36893 a_16981_45144# a_12741_44636# 5.15e-19
C36894 a_1414_42308# a_n2293_46634# 0.260739f
C36895 a_n809_44244# a_n2438_43548# 3.12e-21
C36896 a_14815_43914# a_6755_46942# 1.72e-19
C36897 a_5691_45260# a_5066_45546# 1.08e-20
C36898 a_n2661_43370# a_6419_46155# 1.94e-20
C36899 a_1307_43914# a_6945_45028# 3.38e-20
C36900 a_11173_44260# a_10227_46804# 3.86e-20
C36901 a_n2129_43609# a_n746_45260# 1.13e-21
C36902 a_n1809_43762# a_n2497_47436# 0.005726f
C36903 a_n2267_43396# a_n971_45724# 3.28e-19
C36904 a_13070_42354# a_13575_42558# 1e-19
C36905 a_2903_42308# a_7174_31319# 9.76e-21
C36906 COMP_P a_n2302_39866# 1.42e-19
C36907 a_n3674_37592# a_n4209_39590# 3.94e-20
C36908 a_9223_42460# a_9885_42308# 9.07e-20
C36909 a_n2833_47464# VDD 0.461379f
C36910 C2_P_btm VCM 0.716172f
C36911 DATA[3] DATA[4] 0.001426f
C36912 a_12891_46348# a_11415_45002# 0.059955f
C36913 a_12549_44172# a_20202_43084# 0.028142f
C36914 a_20843_47204# a_20841_46902# 0.002074f
C36915 a_13661_43548# a_20528_46660# 1.2e-20
C36916 a_n743_46660# a_16721_46634# 0.038286f
C36917 a_10467_46802# a_6755_46942# 0.256039f
C36918 a_10623_46897# a_10249_46116# 0.032312f
C36919 a_8145_46902# a_8035_47026# 0.097745f
C36920 a_7927_46660# a_7832_46660# 0.049827f
C36921 a_20916_46384# a_20411_46873# 0.004811f
C36922 a_n881_46662# a_n2472_46090# 1.56e-19
C36923 a_n1613_43370# a_n2293_46098# 0.037934f
C36924 a_n1151_42308# a_n1545_46494# 4.22e-19
C36925 a_n237_47217# a_518_46155# 5.8e-20
C36926 a_584_46384# a_739_46482# 0.004982f
C36927 a_9313_45822# a_2324_44458# 0.004416f
C36928 a_13487_47204# a_13759_46122# 1.3e-19
C36929 a_12861_44030# a_13925_46122# 0.012485f
C36930 a_11599_46634# a_12005_46116# 0.27095f
C36931 a_4883_46098# a_4704_46090# 0.1774f
C36932 a_10334_44484# a_10341_43396# 4.4e-19
C36933 a_13720_44458# a_13667_43396# 2.79e-20
C36934 a_20159_44458# a_19319_43548# 6.17e-19
C36935 a_6109_44484# a_6197_43396# 0.001019f
C36936 a_14539_43914# a_9145_43396# 0.008138f
C36937 a_n2661_43370# a_n3674_39304# 0.002283f
C36938 a_n2661_43922# a_4699_43561# 3.07e-20
C36939 a_n2661_42834# a_3080_42308# 2.61e-19
C36940 a_18184_42460# a_21487_43396# 5.5e-20
C36941 a_10193_42453# a_9885_42558# 0.006254f
C36942 a_7499_43078# a_11323_42473# 5.37e-19
C36943 a_11691_44458# a_17021_43396# 1.04e-20
C36944 a_2711_45572# a_16522_42674# 8.16e-20
C36945 a_18114_32519# a_15743_43084# 1.84e-21
C36946 a_n2293_42834# a_421_43172# 2.71e-19
C36947 a_n1059_45260# a_5837_42852# 0.005989f
C36948 a_2382_45260# a_2987_42968# 6.35e-20
C36949 a_11541_44484# VDD 0.004886f
C36950 a_2711_45572# a_13527_45546# 0.006151f
C36951 a_n2293_42282# SMPL_ON_P 1.31e-19
C36952 a_n2661_43922# a_10586_45546# 6.49e-20
C36953 a_15004_44636# a_n357_42282# 2.78e-22
C36954 a_9145_43396# a_2107_46812# 1.58e-19
C36955 a_14485_44260# a_13059_46348# 1.96e-19
C36956 a_12281_43396# a_n2293_46634# 0.007661f
C36957 a_15037_43940# a_3090_45724# 0.007895f
C36958 a_16409_43396# a_13661_43548# 0.001637f
C36959 a_16867_43762# a_12549_44172# 7.49e-20
C36960 a_6197_43396# a_4646_46812# 0.601282f
C36961 a_11750_44172# a_11415_45002# 6.76e-21
C36962 a_2437_43646# DATA[1] 0.014934f
C36963 a_3357_43084# SINGLE_ENDED 0.131897f
C36964 a_19963_31679# RST_Z 0.050135f
C36965 a_n4334_38304# a_n3565_38216# 0.001004f
C36966 a_6969_46634# VDD 0.154507f
C36967 a_7174_31319# C9_N_btm 9.33e-20
C36968 a_n4064_40160# C1_P_btm 1.21e-19
C36969 a_5932_42308# VDAC_Pi 2.52e-19
C36970 COMP_P VDAC_N 0.003716f
C36971 a_6755_46942# a_8034_45724# 4.79e-20
C36972 a_n743_46660# a_3503_45724# 1.13e-21
C36973 a_10467_46802# a_8049_45260# 1.3e-20
C36974 a_1799_45572# a_n2661_45546# 0.003948f
C36975 a_n2661_46634# a_n443_42852# 3.69e-19
C36976 a_n2293_46634# a_n1013_45572# 0.001008f
C36977 a_765_45546# a_5937_45572# 9.62e-20
C36978 a_15227_44166# a_20708_46348# 0.106656f
C36979 a_19466_46812# a_20075_46420# 0.007984f
C36980 a_19692_46634# a_19335_46494# 0.002287f
C36981 a_14513_46634# a_13759_46122# 3.91e-20
C36982 a_14180_46812# a_13925_46122# 4.05e-19
C36983 a_13885_46660# a_14275_46494# 5.27e-19
C36984 a_17609_46634# a_6945_45028# 4.21e-20
C36985 a_15559_46634# a_10809_44734# 0.004011f
C36986 a_14035_46660# a_14493_46090# 2.33e-20
C36987 a_n2840_46090# a_n1853_46287# 2.2e-19
C36988 a_n2472_46090# a_n2157_46122# 0.080495f
C36989 a_18326_43940# a_18429_43548# 9.67e-19
C36990 a_644_44056# a_685_42968# 2.21e-19
C36991 a_17737_43940# a_15743_43084# 1.41e-19
C36992 a_n97_42460# a_4235_43370# 0.003683f
C36993 a_14021_43940# a_14955_43396# 0.01294f
C36994 a_15493_43940# a_15681_43442# 0.03571f
C36995 a_15493_43396# a_16759_43396# 0.029803f
C36996 a_11967_42832# a_17701_42308# 0.030406f
C36997 a_n1699_43638# a_n1557_42282# 3.96e-21
C36998 a_1049_43396# VDD 0.196328f
C36999 a_20273_45572# a_21297_45572# 2.36e-20
C37000 a_2711_45572# a_16922_45042# 1.19e-19
C37001 a_8696_44636# a_3232_43370# 0.169534f
C37002 a_16680_45572# a_6171_45002# 7.1e-19
C37003 a_21188_45572# a_22591_45572# 1.52e-20
C37004 a_21363_45546# a_19963_31679# 2.99e-19
C37005 a_20528_45572# a_3357_43084# 5.18e-19
C37006 a_21855_43396# a_20202_43084# 3.14e-20
C37007 a_15279_43071# a_3090_45724# 4.84e-21
C37008 a_n2472_42282# a_n2442_46660# 4.03e-20
C37009 a_n3674_38216# a_n2956_39768# 0.023755f
C37010 COMP_P a_21588_30879# 0.001821f
C37011 a_2982_43646# a_n1925_42282# 0.036209f
C37012 a_10341_43396# a_9290_44172# 0.157042f
C37013 a_9885_43396# a_8199_44636# 0.002068f
C37014 a_14456_42282# a_10227_46804# 6.75e-20
C37015 a_n3565_39590# SMPL_ON_P 0.001613f
C37016 a_7227_45028# a_4883_46098# 1.07e-19
C37017 a_10490_45724# a_11599_46634# 1.42e-20
C37018 a_11962_45724# a_12861_44030# 0.184706f
C37019 a_8697_45822# a_6151_47436# 1.19e-20
C37020 a_10907_45822# a_4915_47217# 2e-21
C37021 a_8034_45724# a_8049_45260# 0.141057f
C37022 a_8199_44636# a_n443_42852# 0.021145f
C37023 a_19900_46494# a_20062_46116# 0.006453f
C37024 a_18985_46122# a_21167_46155# 1.63e-20
C37025 a_n4064_37440# C1_P_btm 0.031032f
C37026 a_19700_43370# a_5649_42852# 1.35e-22
C37027 a_8685_43396# a_8952_43230# 0.003917f
C37028 a_2982_43646# a_19987_42826# 7.49e-20
C37029 a_15743_43084# a_13887_32519# 0.075021f
C37030 a_n2661_42282# a_4921_42308# 0.001195f
C37031 a_3422_30871# a_17303_42282# 0.063198f
C37032 a_3626_43646# a_19339_43156# 0.001776f
C37033 a_n97_42460# a_5837_43172# 0.006105f
C37034 a_4235_43370# a_3935_43218# 3.44e-20
C37035 a_1568_43370# a_133_42852# 1.19e-20
C37036 a_3080_42308# a_n2293_42282# 0.122474f
C37037 a_18114_32519# C1_N_btm 1.21e-19
C37038 a_14797_45144# a_11691_44458# 1.53e-19
C37039 a_1307_43914# a_11827_44484# 0.025083f
C37040 a_n2293_42834# a_n2661_43370# 0.038946f
C37041 a_3537_45260# a_n699_43396# 0.025655f
C37042 a_4574_45260# a_4223_44672# 9.56e-20
C37043 a_6709_45028# a_n2661_44458# 2.58e-21
C37044 a_n1059_45260# a_14539_43914# 0.029964f
C37045 a_3065_45002# a_5343_44458# 3.26e-21
C37046 a_7309_42852# a_526_44458# 8.78e-19
C37047 a_17701_42308# a_13259_45724# 0.137488f
C37048 a_5111_42852# a_n755_45592# 2.12e-20
C37049 a_5755_42852# a_n357_42282# 0.179701f
C37050 a_1755_42282# a_1823_45246# 9.08e-19
C37051 a_13017_45260# a_12549_44172# 8.3e-19
C37052 a_13159_45002# a_12891_46348# 0.031652f
C37053 a_11963_45334# a_768_44030# 2.59e-20
C37054 a_10193_42453# a_13059_46348# 6.88e-21
C37055 a_12016_45572# a_11813_46116# 7.88e-20
C37056 a_6171_45002# a_13747_46662# 1.31e-19
C37057 a_n467_45028# a_n743_46660# 0.001437f
C37058 a_n37_45144# a_n1925_46634# 1.2e-20
C37059 a_5205_44484# a_5807_45002# 3.77e-19
C37060 a_1667_45002# a_n2293_46634# 0.009008f
C37061 a_15595_45028# a_n881_46662# 7.5e-20
C37062 a_13807_45067# a_12861_44030# 7.89e-20
C37063 a_22609_37990# VDD 0.079488f
C37064 a_n2129_44697# a_n746_45260# 0.17701f
C37065 a_4223_44672# a_n2497_47436# 0.047068f
C37066 a_n2267_44484# a_n971_45724# 4.09e-19
C37067 a_n2472_42826# a_n1630_35242# 2.09e-20
C37068 a_n1853_43023# a_n3674_37592# 8.55e-20
C37069 a_n901_43156# a_n473_42460# 0.006054f
C37070 a_n1736_43218# a_n1736_42282# 8.52e-19
C37071 a_n1076_43230# a_n961_42308# 2.85e-19
C37072 a_743_42282# a_3823_42558# 0.015894f
C37073 a_13113_42826# a_13291_42460# 1.73e-19
C37074 a_10341_43396# a_15051_42282# 4.87e-20
C37075 a_n4318_38680# a_n4318_37592# 0.027855f
C37076 a_13460_43230# a_13569_43230# 0.007416f
C37077 a_13635_43156# a_13814_43218# 0.007399f
C37078 a_12895_43230# a_13003_42852# 0.057222f
C37079 a_3080_42308# a_n3565_39590# 4.45e-21
C37080 a_6945_45028# DATA[4] 0.0111f
C37081 a_1343_38525# VDD 3.25389f
C37082 a_10227_46804# a_18780_47178# 0.050298f
C37083 a_18143_47464# a_18479_47436# 0.238309f
C37084 a_17591_47464# a_18597_46090# 8.92e-19
C37085 a_4791_45118# a_n1613_43370# 0.223884f
C37086 a_15507_47210# a_4883_46098# 4.76e-22
C37087 a_13717_47436# a_11453_44696# 0.041574f
C37088 a_15673_47210# a_13507_46334# 0.001528f
C37089 a_14955_47212# a_12465_44636# 0.002323f
C37090 a_n1151_42308# a_9804_47204# 0.108722f
C37091 a_584_46384# a_768_44030# 0.105366f
C37092 a_n971_45724# a_5807_45002# 0.0339f
C37093 a_10440_44484# a_n2661_43922# 0.006052f
C37094 a_10057_43914# a_n2661_42834# 0.053564f
C37095 a_13249_42308# a_8685_43396# 0.03355f
C37096 a_20193_45348# a_20835_44721# 1.49e-19
C37097 a_11827_44484# a_18579_44172# 0.045146f
C37098 a_9482_43914# a_10949_43914# 0.025292f
C37099 a_2711_45572# a_15743_43084# 0.075024f
C37100 a_8975_43940# a_11649_44734# 3.69e-19
C37101 a_n2293_42834# a_2998_44172# 6.49e-20
C37102 a_7499_43078# a_10765_43646# 0.002149f
C37103 a_21613_42308# a_13259_45724# 0.077442f
C37104 a_13070_42354# a_n443_42852# 7.16e-20
C37105 a_16842_45938# VDD 4.6e-19
C37106 a_3537_45260# a_7920_46348# 5.32e-20
C37107 a_413_45260# a_9823_46155# 2.74e-21
C37108 a_3357_43084# a_19335_46494# 2.49e-21
C37109 a_5147_45002# a_5497_46414# 4.57e-19
C37110 a_4927_45028# a_5164_46348# 0.09665f
C37111 a_5111_44636# a_5204_45822# 8.78e-19
C37112 a_20193_45348# a_3090_45724# 1.53e-20
C37113 a_11967_42832# a_12891_46348# 3.62e-21
C37114 a_14673_44172# a_13747_46662# 4.77e-21
C37115 a_n2661_42834# a_n2438_43548# 0.057776f
C37116 a_19006_44850# a_12549_44172# 5.76e-20
C37117 a_16241_44734# a_13661_43548# 0.047309f
C37118 a_11691_44458# a_14976_45028# 6.38e-19
C37119 a_18494_42460# a_19692_46634# 6.49e-19
C37120 a_7276_45260# a_3483_46348# 0.003843f
C37121 a_n2661_43922# a_n743_46660# 1.41e-20
C37122 a_1755_42282# a_5934_30871# 3.43e-20
C37123 a_2351_42308# a_6123_31319# 8.95e-21
C37124 a_1606_42308# a_8515_42308# 1.34e-20
C37125 a_2903_42308# a_5932_42308# 8.68e-21
C37126 a_5267_42460# a_5421_42558# 0.010303f
C37127 a_5379_42460# a_5337_42558# 8.44e-19
C37128 COMP_P a_5742_30871# 0.1094f
C37129 a_13678_32519# C4_N_btm 1.42e-19
C37130 a_13467_32519# C7_N_btm 1.83e-20
C37131 a_13887_32519# C1_N_btm 8.65e-20
C37132 a_22469_39537# a_22609_37990# 0.490939f
C37133 a_12549_44172# a_12469_46902# 0.00102f
C37134 a_n2661_46634# a_10554_47026# 0.009556f
C37135 a_3177_46902# a_4646_46812# 2.63e-20
C37136 a_2443_46660# a_4955_46873# 4.31e-21
C37137 a_n1925_46634# a_8492_46660# 9.51e-19
C37138 a_2609_46660# a_4651_46660# 1.13e-19
C37139 a_2959_46660# a_3877_44458# 2.53e-19
C37140 a_12891_46348# a_12251_46660# 0.003575f
C37141 a_5807_45002# a_8023_46660# 0.001248f
C37142 a_2107_46812# a_3878_46660# 3.62e-19
C37143 a_n881_46662# a_15559_46634# 3.94e-20
C37144 a_11453_44696# a_14035_46660# 1.53e-20
C37145 a_3080_42308# a_3726_37500# 0.004001f
C37146 a_13507_46334# a_16388_46812# 0.083261f
C37147 a_18143_47464# a_17829_46910# 2.74e-19
C37148 a_18479_47436# a_765_45546# 1.7e-19
C37149 a_10227_46804# a_18285_46348# 5.46e-20
C37150 a_12861_44030# a_16655_46660# 6.9e-19
C37151 a_n237_47217# a_3147_46376# 0.052931f
C37152 a_584_46384# a_1176_45822# 0.039976f
C37153 a_n971_45724# a_3699_46348# 0.013334f
C37154 a_n1151_42308# a_n901_46420# 0.002158f
C37155 a_1209_47178# a_167_45260# 2.76e-21
C37156 a_4791_45118# a_n2293_46098# 0.411939f
C37157 a_2063_45854# a_1208_46090# 4.06e-19
C37158 a_n2109_47186# a_5497_46414# 0.017063f
C37159 a_n1741_47186# a_5164_46348# 3.78e-20
C37160 a_n2840_43914# a_n4318_39768# 0.170372f
C37161 a_2127_44172# a_2479_44172# 0.168988f
C37162 a_453_43940# a_895_43940# 0.420851f
C37163 a_1414_42308# a_2675_43914# 0.305556f
C37164 a_1115_44172# a_2998_44172# 6.12e-20
C37165 a_17517_44484# a_15493_43396# 7.93e-20
C37166 a_7640_43914# a_7499_43940# 0.049504f
C37167 a_n699_43396# a_1049_43396# 0.006702f
C37168 a_5891_43370# a_5829_43940# 1.98e-19
C37169 a_742_44458# a_4235_43370# 3.35e-20
C37170 a_n1059_45260# a_7871_42858# 0.032582f
C37171 a_n2017_45002# a_7765_42852# 7.13e-20
C37172 a_8701_44490# VDD 0.164475f
C37173 a_7174_31319# RST_Z 0.216004f
C37174 a_4958_30871# VCM 0.642743f
C37175 a_n2216_37984# a_n2956_38216# 8.63e-19
C37176 a_17517_44484# a_3483_46348# 0.004031f
C37177 a_20397_44484# a_11415_45002# 2.5e-20
C37178 a_9028_43914# a_3090_45724# 0.00399f
C37179 a_17969_45144# a_13259_45724# 8.9e-19
C37180 a_n2293_43922# a_9290_44172# 0.369185f
C37181 a_8791_43396# a_n1613_43370# 4.34e-20
C37182 a_9145_43396# a_11453_44696# 2.08e-20
C37183 a_14579_43548# a_12465_44636# 1.92e-21
C37184 a_n1423_42826# SMPL_ON_P 8.78e-21
C37185 a_n3674_39304# a_n2497_47436# 4.4e-20
C37186 a_n4334_39616# a_n4064_39072# 7.91e-19
C37187 a_n3690_39616# a_n3420_39072# 8.87e-19
C37188 a_n2946_39866# a_n3565_39304# 0.001251f
C37189 a_n2302_39866# a_n4209_39304# 0.001254f
C37190 a_n4209_39590# a_n2302_39072# 0.00133f
C37191 a_n4064_39616# a_n4334_39392# 0.001768f
C37192 a_n3420_39616# a_n3690_39392# 0.018295f
C37193 a_n3565_39590# a_n2946_39072# 0.001251f
C37194 a_n2293_46634# VDD 1.52629f
C37195 a_5932_42308# C9_N_btm 9.33e-20
C37196 a_6123_31319# C4_N_btm 0.132906f
C37197 a_5934_30871# C2_N_btm 0.011047f
C37198 a_17339_46660# a_18285_46348# 0.184197f
C37199 a_765_45546# a_17829_46910# 0.069261f
C37200 a_12891_46348# a_13259_45724# 1.04614f
C37201 a_2107_46812# a_n1925_42282# 0.006094f
C37202 a_n2661_46098# a_n722_46482# 0.001878f
C37203 a_5807_45002# a_12005_46436# 8.93e-20
C37204 a_6755_46942# a_8016_46348# 0.002347f
C37205 a_9863_46634# a_9823_46155# 9.52e-19
C37206 a_2747_46873# a_n2661_45546# 1.72e-21
C37207 a_20679_44626# a_743_42282# 7.32e-21
C37208 a_20640_44752# a_20556_43646# 1.74e-20
C37209 a_11967_42832# a_4361_42308# 0.012085f
C37210 a_18287_44626# a_18249_42858# 2.07e-21
C37211 a_18248_44752# a_18817_42826# 8.42e-22
C37212 a_22485_44484# a_15743_43084# 0.003457f
C37213 a_19279_43940# a_21259_43561# 5.61e-22
C37214 a_n2661_43922# a_1847_42826# 3.92e-22
C37215 a_3499_42826# a_3457_43396# 0.005429f
C37216 a_5891_43370# a_10835_43094# 1.38e-20
C37217 a_n2293_42834# COMP_P 8.54e-19
C37218 a_n2661_42282# a_6452_43396# 0.011968f
C37219 a_1307_43914# a_3581_42558# 4.31e-20
C37220 a_20512_43084# a_19268_43646# 2.18e-19
C37221 en_comp a_15890_42674# 1.81e-20
C37222 a_17478_45572# a_18175_45572# 0.001484f
C37223 a_2711_45572# a_10775_45002# 1.05e-19
C37224 a_15599_45572# a_16789_45572# 2.56e-19
C37225 a_8696_44636# a_18341_45572# 1.27e-19
C37226 a_15861_45028# a_18479_45785# 3.3e-20
C37227 a_6598_45938# a_6171_45002# 0.002784f
C37228 a_6511_45714# a_5205_44484# 5.08e-20
C37229 a_6667_45809# a_6431_45366# 0.002877f
C37230 a_6472_45840# a_7276_45260# 6.14e-21
C37231 a_11823_42460# a_n2017_45002# 0.098619f
C37232 a_7227_45028# a_3232_43370# 9.21e-19
C37233 a_3905_42558# a_4791_45118# 8.4e-21
C37234 CAL_N CAL_P 5.91728f
C37235 a_n3565_37414# C10_P_btm 1.19e-19
C37236 a_n4209_37414# C8_P_btm 1.65e-20
C37237 a_n97_42460# a_9290_44172# 0.351467f
C37238 a_9248_44260# a_8049_45260# 1.1e-21
C37239 a_2127_44172# a_n443_42852# 5.26e-20
C37240 a_n2293_42282# a_n2438_43548# 1.27e-19
C37241 a_9625_46129# VDD 0.996485f
C37242 a_6194_45824# a_n237_47217# 2.56e-20
C37243 a_6511_45714# a_n971_45724# 0.001043f
C37244 a_22959_46660# a_20692_30879# 0.004672f
C37245 a_21076_30879# a_20205_31679# 0.055235f
C37246 a_765_45546# a_n443_42852# 0.232932f
C37247 a_8016_46348# a_8049_45260# 0.09608f
C37248 a_8953_45546# a_8034_45724# 2.24e-19
C37249 a_21137_46414# a_10809_44734# 1.12e-20
C37250 a_6945_45028# a_22223_46124# 0.17119f
C37251 a_n4209_38502# a_n4334_37440# 3.34e-19
C37252 a_2684_37794# a_3754_38802# 9.44e-20
C37253 a_n1613_43370# DATA[3] 3.98e-19
C37254 a_15095_43370# a_16137_43396# 1.7e-19
C37255 a_n2065_43946# a_n1630_35242# 4.6e-22
C37256 a_n1557_42282# a_n2157_42858# 0.007773f
C37257 a_n97_42460# a_791_42968# 0.039538f
C37258 a_n1761_44111# a_564_42282# 1.16e-19
C37259 a_10807_43548# a_11229_43218# 6.49e-19
C37260 a_10341_43396# a_13749_43396# 9.69e-20
C37261 a_n881_46662# DATA[2] 2.22e-20
C37262 a_22612_30879# a_22609_37990# 1.7e-20
C37263 a_n1533_42852# VDD 0.142813f
C37264 a_15599_45572# a_14539_43914# 2.3e-21
C37265 a_8696_44636# a_8975_43940# 0.003372f
C37266 a_15595_45028# a_1307_43914# 4.87e-19
C37267 a_10180_45724# a_n2661_42834# 5.55e-20
C37268 a_2711_45572# a_16789_44484# 2.48e-19
C37269 a_413_45260# a_n2661_43370# 1.31746f
C37270 a_21513_45002# a_21359_45002# 0.289039f
C37271 a_19479_31679# a_20567_45036# 3.97e-20
C37272 a_8685_42308# a_8270_45546# 2.23e-21
C37273 a_n2216_39866# a_n2442_46660# 0.003462f
C37274 a_4361_42308# a_13259_45724# 0.054653f
C37275 a_16759_43396# a_n357_42282# 0.007988f
C37276 a_7765_42852# a_526_44458# 0.023934f
C37277 a_8945_43396# a_n443_42852# 3.77e-20
C37278 a_n1059_45260# a_11453_44696# 1.65e-20
C37279 a_6171_45002# a_11599_46634# 3.62e-19
C37280 a_413_45260# a_19787_47423# 8.86e-20
C37281 a_n2293_42834# a_n2497_47436# 0.010004f
C37282 a_2437_43646# a_5063_47570# 8.52e-19
C37283 a_17478_45572# a_n743_46660# 9.46e-19
C37284 a_18479_45785# a_19321_45002# 0.114441f
C37285 a_20107_45572# a_12549_44172# 2.47e-19
C37286 a_18909_45814# a_13747_46662# 0.025022f
C37287 a_19431_45546# a_5807_45002# 0.01527f
C37288 a_18691_45572# a_13661_43548# 0.020905f
C37289 a_7499_43078# a_8492_46660# 1.8e-19
C37290 a_509_45822# a_n443_42852# 0.035689f
C37291 a_6293_42852# a_5932_42308# 8.47e-19
C37292 a_12089_42308# a_5534_30871# 0.012295f
C37293 a_3457_43396# a_3318_42354# 8.91e-20
C37294 a_6197_43396# a_6171_42473# 5.91e-20
C37295 a_n97_42460# a_15051_42282# 0.049661f
C37296 a_13113_42826# a_13460_43230# 0.051162f
C37297 a_1847_42826# a_3445_43172# 4.44e-21
C37298 a_15743_43084# a_16877_42852# 1.77e-20
C37299 a_3626_43646# a_3905_42308# 0.002949f
C37300 a_20820_30879# VREF_GND 0.02097f
C37301 a_3422_30871# C8_N_btm 4.06e-19
C37302 a_13249_42558# VDD 0.009141f
C37303 a_n785_47204# a_n1435_47204# 9.32e-19
C37304 a_n1151_42308# a_6545_47178# 0.01616f
C37305 a_2063_45854# a_6575_47204# 0.002711f
C37306 a_3785_47178# a_5815_47464# 2.66e-19
C37307 a_4007_47204# a_4915_47217# 0.001046f
C37308 a_4700_47436# a_n443_46116# 0.255594f
C37309 a_19431_45546# a_19478_44306# 9.3e-21
C37310 a_5343_44458# a_6298_44484# 0.128602f
C37311 a_17668_45572# a_17737_43940# 2.42e-20
C37312 a_19256_45572# a_15493_43396# 2.21e-21
C37313 a_4223_44672# a_5883_43914# 0.967973f
C37314 a_15861_45028# a_14021_43940# 3.03e-20
C37315 a_2680_45002# a_2127_44172# 2.9e-20
C37316 a_413_45260# a_2998_44172# 0.161528f
C37317 a_3429_45260# a_1414_42308# 1.27e-22
C37318 a_3357_43084# a_3499_42826# 0.134316f
C37319 a_2382_45260# a_2479_44172# 0.00555f
C37320 a_n2017_45002# a_n1644_44306# 0.00478f
C37321 a_n2293_45010# a_n1287_44306# 8.54e-19
C37322 a_1221_42558# a_n863_45724# 0.003967f
C37323 a_1067_42314# a_n357_42282# 5.85e-20
C37324 a_n1630_35242# a_n755_45592# 0.044103f
C37325 a_7230_45938# VDD 0.077608f
C37326 a_n452_44636# a_n743_46660# 3.36e-20
C37327 a_14797_45144# a_15227_44166# 0.011685f
C37328 a_n699_43396# a_n2293_46634# 0.016884f
C37329 a_18374_44850# a_12549_44172# 2.67e-20
C37330 a_19963_31679# a_20820_30879# 0.057032f
C37331 a_19479_31679# a_21076_30879# 0.054875f
C37332 a_20447_31679# a_11415_45002# 2.6e-19
C37333 a_21297_45572# a_20202_43084# 2.32e-19
C37334 a_413_45260# a_20107_46660# 1.46e-20
C37335 a_15037_45618# a_14840_46494# 1.08e-19
C37336 a_10907_45822# a_10809_44734# 0.003912f
C37337 a_n1243_44484# a_n1613_43370# 6.03e-19
C37338 a_15463_44811# a_10227_46804# 1.33e-19
C37339 a_14673_44172# a_11599_46634# 3.2e-21
C37340 a_n2065_43946# a_n971_45724# 0.016306f
C37341 a_1115_44172# a_n2497_47436# 0.069778f
C37342 a_16795_42852# a_4958_30871# 0.001047f
C37343 a_n2840_42282# a_n4318_37592# 0.037154f
C37344 a_n2472_42282# a_n3674_38216# 0.040147f
C37345 a_n3674_39304# a_n4209_39304# 0.059449f
C37346 a_n4318_38216# a_n2104_42282# 7.75e-19
C37347 a_14097_32519# a_n784_42308# 0.005039f
C37348 a_9306_43218# a_5934_30871# 4.18e-20
C37349 a_n2840_46634# a_n2442_46660# 0.007415f
C37350 a_n2956_39768# a_n2472_46634# 5e-19
C37351 a_n1613_43370# a_1057_46660# 2.95e-19
C37352 a_4883_46098# a_7715_46873# 0.01159f
C37353 a_10227_46804# a_10249_46116# 0.137273f
C37354 a_6151_47436# a_15009_46634# 0.00896f
C37355 a_4915_47217# a_15368_46634# 4.4e-21
C37356 a_18587_45118# a_18533_43940# 6.8e-22
C37357 a_17970_44736# a_17737_43940# 1.63e-19
C37358 a_17767_44458# a_17973_43940# 0.012863f
C37359 a_n2661_43922# a_5244_44056# 2.61e-20
C37360 a_n2661_42834# a_5013_44260# 0.021017f
C37361 a_n2661_43370# a_n2012_43396# 1.88e-20
C37362 a_n2293_42834# a_1568_43370# 0.037512f
C37363 a_1307_43914# a_8147_43396# 2.66e-20
C37364 a_n2293_43922# a_3905_42865# 2.09e-20
C37365 a_20640_44752# a_20980_44850# 0.027606f
C37366 a_19778_44110# a_19808_44306# 0.004261f
C37367 a_20159_44458# a_3422_30871# 2.52e-20
C37368 a_16922_45042# a_14401_32519# 1.06e-19
C37369 a_5111_44636# a_9885_43646# 0.010527f
C37370 a_n1059_45260# a_17324_43396# 0.003177f
C37371 a_n913_45002# a_17499_43370# 2.4e-20
C37372 a_8704_45028# VDD 0.004293f
C37373 a_5934_30871# C8_P_btm 1.41e-19
C37374 a_6123_31319# C6_P_btm 6.31e-19
C37375 a_5932_42308# RST_Z 0.005263f
C37376 a_20692_30879# C10_N_btm 2.44e-19
C37377 a_8791_43396# a_4791_45118# 1.84e-20
C37378 a_11827_44484# a_22223_46124# 4.45e-19
C37379 a_5343_44458# a_5937_45572# 0.024374f
C37380 a_8103_44636# a_8016_46348# 8.07e-22
C37381 a_20193_45348# a_20075_46420# 4.06e-21
C37382 a_2382_45260# a_n443_42852# 0.020006f
C37383 a_2274_45254# a_1609_45822# 0.11737f
C37384 a_8488_45348# a_8049_45260# 7.56e-19
C37385 a_15037_44260# a_13661_43548# 0.003411f
C37386 a_14021_43940# a_19321_45002# 1.97e-19
C37387 a_20766_44850# a_15227_44166# 3.54e-21
C37388 a_20640_44752# a_19692_46634# 0.001236f
C37389 a_13720_44458# a_3483_46348# 0.010665f
C37390 a_18597_46090# VDD 0.930122f
C37391 a_19332_42282# a_19511_42282# 0.174683f
C37392 a_17303_42282# a_7174_31319# 0.027048f
C37393 a_18214_42558# a_18548_42308# 2.43e-19
C37394 a_5742_30871# a_n4209_39304# 6.2e-21
C37395 a_n2661_46098# a_472_46348# 0.065456f
C37396 a_2107_46812# a_2698_46116# 0.00811f
C37397 a_14976_45028# a_15227_44166# 0.035507f
C37398 a_12251_46660# a_12359_47026# 0.057222f
C37399 a_11735_46660# a_12347_46660# 3.82e-19
C37400 a_6755_46942# a_15312_46660# 2.66e-21
C37401 a_13747_46662# a_10903_43370# 0.027209f
C37402 a_n743_46660# a_5164_46348# 0.031878f
C37403 a_12549_44172# a_17715_44484# 0.03426f
C37404 a_5807_45002# a_12594_46348# 0.001952f
C37405 a_n2661_46634# a_8199_44636# 2.29e-19
C37406 a_n1925_46634# a_5497_46414# 6.78e-20
C37407 a_n1613_43370# a_6945_45028# 0.049203f
C37408 a_4883_46098# a_5210_46482# 2.25e-19
C37409 a_17591_47464# a_8049_45260# 1.43e-20
C37410 a_12861_44030# a_12638_46436# 6.45e-19
C37411 a_n746_45260# a_n357_42282# 0.002027f
C37412 a_2063_45854# a_n2661_45546# 0.038547f
C37413 a_n971_45724# a_n755_45592# 0.347347f
C37414 a_3905_42865# a_n97_42460# 0.071125f
C37415 a_14673_44172# a_14358_43442# 0.00447f
C37416 a_20623_43914# a_14021_43940# 1.48e-19
C37417 a_453_43940# a_458_43396# 9.25e-20
C37418 a_1467_44172# a_1049_43396# 0.002443f
C37419 a_1115_44172# a_1568_43370# 1.06e-19
C37420 a_9313_44734# a_18783_43370# 8.63e-20
C37421 a_11827_44484# a_13635_43156# 3.57e-21
C37422 a_n1761_44111# a_n1557_42282# 0.018977f
C37423 a_n4318_39768# a_n4318_39304# 0.042825f
C37424 a_9028_43914# a_9165_43940# 0.126609f
C37425 a_1414_42308# a_1209_43370# 0.003338f
C37426 a_742_44458# a_791_42968# 3.18e-19
C37427 a_n2293_42834# a_4743_43172# 2.14e-19
C37428 a_n3674_39768# a_n2840_43370# 0.006059f
C37429 a_3357_43084# a_3318_42354# 2.7e-19
C37430 a_n1059_45260# a_1184_42692# 0.019924f
C37431 a_n967_45348# a_n327_42558# 5.76e-21
C37432 a_n913_45002# a_1576_42282# 0.001393f
C37433 a_n2017_45002# a_961_42354# 0.00519f
C37434 a_n2810_45028# a_n1630_35242# 4.11e-19
C37435 en_comp a_n3674_37592# 0.050998f
C37436 a_2675_43914# VDD 0.200923f
C37437 a_13163_45724# a_15037_45618# 7.32e-23
C37438 a_10193_42453# a_8696_44636# 0.225102f
C37439 a_8697_45822# a_8791_45572# 1.26e-19
C37440 C7_N_btm VCM 1.58335f
C37441 C8_N_btm VREF_GND 2.58605f
C37442 C9_N_btm VREF 7.369471f
C37443 C10_N_btm VIN_N 3.66034f
C37444 a_3737_43940# a_1823_45246# 8.92e-19
C37445 a_8952_43230# a_768_44030# 2.43e-19
C37446 a_9803_43646# a_8270_45546# 0.066865f
C37447 a_n1423_42826# a_n2438_43548# 9.01e-21
C37448 a_15433_44458# a_n443_42852# 1.08e-21
C37449 a_15682_43940# a_2324_44458# 0.321744f
C37450 a_9895_44260# a_8199_44636# 0.002714f
C37451 a_9248_44260# a_8953_45546# 4.19e-20
C37452 a_19123_46287# VDD 0.336379f
C37453 a_n4315_30879# a_n4064_37984# 0.034375f
C37454 a_n4064_40160# a_n3420_37984# 0.053114f
C37455 a_19692_46634# a_19240_46482# 4.58e-21
C37456 a_14035_46660# a_14180_46482# 0.157972f
C37457 a_19466_46812# a_19431_46494# 0.001367f
C37458 a_1823_45246# a_2324_44458# 0.069409f
C37459 a_3483_46348# a_13351_46090# 1.87e-20
C37460 a_8016_46348# a_8953_45546# 0.060003f
C37461 a_8349_46414# a_5937_45572# 6.5e-20
C37462 a_10949_43914# a_10796_42968# 9.1e-19
C37463 a_10057_43914# a_9885_42558# 4.04e-21
C37464 a_10807_43548# a_10835_43094# 0.02952f
C37465 a_19741_43940# a_19700_43370# 5.56e-19
C37466 a_10729_43914# a_10991_42826# 1.29e-20
C37467 a_14401_32519# a_15743_43084# 0.017308f
C37468 a_n2661_42834# a_196_42282# 1.99e-22
C37469 a_n2293_43922# a_n961_42308# 1.63e-19
C37470 a_18494_42460# a_20107_42308# 0.035023f
C37471 a_18184_42460# a_20712_42282# 3.18e-19
C37472 a_3905_42865# a_3935_43218# 0.004982f
C37473 a_n443_46116# DATA[2] 0.006001f
C37474 a_4791_45118# DATA[3] 5.9e-20
C37475 a_20447_31679# C6_N_btm 0.001141f
C37476 a_19963_31679# C8_N_btm 1.65e-20
C37477 a_14537_43646# VDD 0.008942f
C37478 a_8162_45546# a_4223_44672# 4.14e-21
C37479 a_2711_45572# a_17970_44736# 6.8e-21
C37480 a_2382_45260# a_2680_45002# 0.023953f
C37481 a_413_45260# a_4574_45260# 7.73e-20
C37482 a_3626_43646# a_n863_45724# 1.16e-20
C37483 a_15567_42826# a_12741_44636# 1.49e-21
C37484 a_3422_30871# C2_P_btm 9.13e-20
C37485 a_2277_45546# VDD 0.209584f
C37486 a_14495_45572# a_12549_44172# 4.78e-19
C37487 a_5263_45724# a_2107_46812# 7.2e-22
C37488 a_13249_42308# a_768_44030# 0.012496f
C37489 a_15599_45572# a_11453_44696# 4.53e-20
C37490 a_18909_45814# a_11599_46634# 0.042943f
C37491 a_17786_45822# a_16327_47482# 1.4e-20
C37492 a_14033_45572# a_10227_46804# 2.4e-19
C37493 a_18596_45572# a_12861_44030# 0.007922f
C37494 a_3357_43084# a_n1151_42308# 0.028306f
C37495 a_2437_43646# a_3815_47204# 0.012198f
C37496 a_n745_45366# a_n746_45260# 0.119822f
C37497 a_413_45260# a_n2497_47436# 0.028795f
C37498 a_n1177_43370# a_n784_42308# 2.67e-21
C37499 a_15743_43084# a_18817_42826# 0.003018f
C37500 a_18783_43370# a_18599_43230# 6.07e-19
C37501 a_n1076_43230# a_685_42968# 4.61e-19
C37502 a_5649_42852# a_9127_43156# 8.16e-20
C37503 a_743_42282# a_10341_42308# 0.020229f
C37504 a_19268_43646# a_18249_42858# 7.34e-20
C37505 a_n3674_39768# a_n4315_30879# 7.29e-19
C37506 a_n13_43084# a_421_43172# 0.003935f
C37507 a_n4318_39768# a_n4334_40480# 0.002408f
C37508 a_14401_32519# a_1606_42308# 0.001872f
C37509 a_3080_42308# a_14097_32519# 1.75e-20
C37510 a_8685_43396# a_8495_42852# 2.66e-19
C37511 a_19692_46634# START 1.28e-19
C37512 a_3090_45724# CLK 0.001129f
C37513 a_n3420_37984# a_n4064_37440# 7.43287f
C37514 a_n2946_37984# a_n2946_37690# 0.050477f
C37515 a_n4064_37984# a_n3420_37440# 0.053897f
C37516 a_7754_39964# a_7754_38636# 0.005394f
C37517 a_n1736_42282# VDD 0.227152f
C37518 a_11827_44484# a_22223_45036# 0.179208f
C37519 a_20567_45036# a_20193_45348# 0.037561f
C37520 a_n2661_43370# a_2779_44458# 1.59e-19
C37521 a_7499_43078# a_11341_43940# 0.00321f
C37522 a_13249_42308# a_13483_43940# 0.193724f
C37523 a_10193_42453# a_20365_43914# 1.25e-20
C37524 a_16922_45042# a_20205_45028# 0.0038f
C37525 a_n2293_42834# a_5883_43914# 0.015714f
C37526 a_21363_45546# a_21398_44850# 1.78e-21
C37527 a_5111_44636# a_n2661_43922# 0.061031f
C37528 a_8953_45002# a_9313_44734# 0.001727f
C37529 a_21513_45002# a_19279_43940# 0.003201f
C37530 a_3357_43084# a_20640_44752# 4.03e-21
C37531 a_3232_43370# a_9159_44484# 0.005178f
C37532 a_15890_42674# a_4185_45028# 6.54e-20
C37533 a_21613_42308# a_20202_43084# 0.07574f
C37534 a_13258_32519# a_21076_30879# 0.059077f
C37535 a_4149_42891# a_n357_42282# 2.65e-19
C37536 a_1184_42692# a_n1925_42282# 5.67e-20
C37537 a_961_42354# a_526_44458# 2.74e-21
C37538 a_1709_42852# a_n443_42852# 5.75e-21
C37539 a_13622_42852# a_13259_45724# 1.68e-19
C37540 a_10533_42308# a_9290_44172# 0.001105f
C37541 a_12607_44458# a_11599_46634# 1.01e-22
C37542 a_4880_45572# a_5937_45572# 1.79e-19
C37543 a_n913_45002# a_8270_45546# 1.44e-20
C37544 a_20528_45572# a_19466_46812# 0.157758f
C37545 a_6171_45002# a_7411_46660# 4.46e-21
C37546 a_2437_43646# a_14976_45028# 1.11e-19
C37547 a_3232_43370# a_7715_46873# 1.19e-20
C37548 a_21188_45572# a_19692_46634# 7.15e-19
C37549 a_14976_45348# a_13661_43548# 9.13e-21
C37550 a_18175_45572# a_16388_46812# 1.3e-20
C37551 a_17719_45144# a_12549_44172# 2.85e-20
C37552 a_11525_45546# a_3483_46348# 2.41e-19
C37553 a_4361_42308# a_16197_42308# 1.2e-19
C37554 a_21487_43396# a_17303_42282# 4.02e-21
C37555 a_8605_42826# a_8515_42308# 0.001559f
C37556 a_8387_43230# a_5934_30871# 0.001004f
C37557 a_n2293_42282# a_196_42282# 4.89e-19
C37558 a_5649_42852# a_17124_42282# 1.31e-19
C37559 a_743_42282# a_18057_42282# 0.008889f
C37560 a_4190_30871# a_18907_42674# 0.040515f
C37561 a_14401_32519# C1_N_btm 6.64e-20
C37562 a_12465_44636# a_5807_45002# 0.59474f
C37563 a_4883_46098# a_13747_46662# 0.050962f
C37564 a_20990_47178# a_20843_47204# 0.003683f
C37565 a_13507_46334# a_19321_45002# 0.034054f
C37566 a_21177_47436# a_19594_46812# 4.79e-20
C37567 a_15673_47210# a_n743_46660# 0.002403f
C37568 a_n1435_47204# a_2107_46812# 5.14e-20
C37569 a_n1151_42308# a_3877_44458# 0.019733f
C37570 a_3160_47472# a_4646_46812# 2.88e-21
C37571 a_n443_46116# a_3067_47026# 0.030121f
C37572 a_16922_45042# a_15682_43940# 0.001439f
C37573 a_2779_44458# a_2998_44172# 0.007931f
C37574 a_n699_43396# a_2675_43914# 0.015641f
C37575 a_n4318_40392# a_n3674_39768# 0.026429f
C37576 a_n2293_43922# a_12553_44484# 1.41e-19
C37577 a_742_44458# a_3905_42865# 0.002336f
C37578 a_n2661_44458# a_n4318_39768# 8.38e-19
C37579 a_8696_44636# a_16137_43396# 2.49e-20
C37580 a_1307_43914# a_10555_43940# 0.001112f
C37581 a_5147_45002# a_n97_42460# 0.085495f
C37582 a_3357_43084# a_6197_43396# 0.001107f
C37583 a_n2017_45002# a_2982_43646# 0.023101f
C37584 a_n3565_38502# a_n2956_38216# 0.072968f
C37585 a_3429_45260# VDD 0.142923f
C37586 COMP_P a_22545_38993# 4.2e-21
C37587 a_16886_45144# a_12741_44636# 4.07e-19
C37588 a_n1549_44318# a_n2438_43548# 3.51e-20
C37589 a_1467_44172# a_n2293_46634# 3.1e-20
C37590 a_4927_45028# a_5066_45546# 0.001602f
C37591 a_8560_45348# a_5937_45572# 0.045711f
C37592 a_n2661_43370# a_6165_46155# 9.24e-21
C37593 a_6756_44260# a_n1613_43370# 0.00105f
C37594 a_18326_43940# a_11453_44696# 3.74e-20
C37595 a_10555_44260# a_10227_46804# 1.96e-19
C37596 a_n2129_43609# a_n971_45724# 0.173854f
C37597 a_n2012_43396# a_n2497_47436# 1.4e-19
C37598 a_2713_42308# a_7174_31319# 4.88e-21
C37599 a_n1630_35242# a_n2302_40160# 1.59e-19
C37600 w_11334_34010# VDD 1.90683f
C37601 a_5342_30871# C10_N_btm 2.16e-19
C37602 C2_P_btm VREF_GND 0.671742f
C37603 C3_P_btm VCM 0.716273f
C37604 a_4883_46098# a_4419_46090# 0.006295f
C37605 a_n2661_46634# a_765_45546# 1.82448f
C37606 a_11309_47204# a_11415_45002# 0.001299f
C37607 a_20916_46384# a_20107_46660# 8.05e-20
C37608 a_n743_46660# a_16388_46812# 0.035819f
C37609 a_10623_46897# a_10554_47026# 0.209641f
C37610 a_10428_46928# a_6755_46942# 0.155315f
C37611 a_10467_46802# a_10249_46116# 0.12624f
C37612 a_7577_46660# a_8035_47026# 0.027606f
C37613 a_3055_46660# a_3090_45724# 9.03e-20
C37614 a_19321_45002# a_20623_46660# 3.43e-19
C37615 a_13747_46662# a_21188_46660# 2.57e-20
C37616 a_n1613_43370# a_n2472_46090# 3.22e-20
C37617 a_4791_45118# a_6945_45028# 0.493927f
C37618 a_12861_44030# a_13759_46122# 0.032694f
C37619 a_13717_47436# a_13925_46122# 5.15e-19
C37620 a_10227_46804# a_5937_45572# 2.11e-20
C37621 a_11599_46634# a_10903_43370# 0.439916f
C37622 a_19615_44636# a_19319_43548# 0.001036f
C37623 a_n2661_42834# a_4699_43561# 6.89e-20
C37624 a_6109_44484# a_6293_42852# 3.01e-21
C37625 a_14537_43396# a_5534_30871# 2.84e-19
C37626 a_13556_45296# a_15567_42826# 4.05e-21
C37627 a_18494_42460# a_743_42282# 0.476713f
C37628 a_7499_43078# a_10723_42308# 0.029878f
C37629 a_9313_44734# a_3626_43646# 2.37e-19
C37630 a_11691_44458# a_16855_43396# 4.36e-20
C37631 a_11967_42832# a_18533_43940# 4.96e-19
C37632 a_n2293_42834# a_133_43172# 4.3e-19
C37633 a_n1059_45260# a_5193_42852# 0.004497f
C37634 a_n4064_38528# VCM 0.007464f
C37635 a_2711_45572# a_13163_45724# 0.006905f
C37636 a_17364_32525# SMPL_ON_N 0.029237f
C37637 a_n2661_42834# a_10586_45546# 3.13e-20
C37638 a_5343_44458# a_n443_42852# 0.057128f
C37639 a_12293_43646# a_n2293_46634# 0.001258f
C37640 a_16547_43609# a_13661_43548# 1.23e-19
C37641 a_16664_43396# a_12549_44172# 9.47e-20
C37642 a_6293_42852# a_4646_46812# 0.030189f
C37643 a_14021_43940# a_13059_46348# 0.082427f
C37644 a_2437_43646# DATA[0] 9.16e-20
C37645 a_3357_43084# START 0.045418f
C37646 a_22591_45572# RST_Z 5.34e-19
C37647 a_n4209_38216# a_n3565_38216# 6.80743f
C37648 a_6755_46942# VDD 1.05713f
C37649 a_7174_31319# C8_N_btm 7.53e-20
C37650 a_n1630_35242# a_n2302_37690# 1.59e-19
C37651 a_5934_30871# a_2113_38308# 6.72e-20
C37652 COMP_P a_6886_37412# 0.00104f
C37653 a_n743_46660# a_3316_45546# 2.86e-19
C37654 a_n2661_46098# a_n2840_45546# 3.06e-19
C37655 a_10428_46928# a_8049_45260# 2.57e-20
C37656 a_33_46660# a_997_45618# 7.11e-21
C37657 a_15227_44166# a_19900_46494# 0.053335f
C37658 a_14035_46660# a_13925_46122# 0.207108f
C37659 a_19692_46634# a_19553_46090# 1.1e-19
C37660 a_19466_46812# a_19335_46494# 0.017838f
C37661 a_14180_46812# a_13759_46122# 0.001754f
C37662 a_13885_46660# a_14493_46090# 0.001138f
C37663 a_16292_46812# a_6945_45028# 3.43e-20
C37664 a_15368_46634# a_10809_44734# 0.002169f
C37665 a_765_45546# a_8199_44636# 8.72e-20
C37666 a_n2840_46090# a_n2157_46122# 7.58e-21
C37667 a_n2472_46090# a_n2293_46098# 0.176709f
C37668 a_15682_43940# a_15743_43084# 6.12e-19
C37669 a_n2267_43396# a_n1557_42282# 1.4e-20
C37670 a_n97_42460# a_4093_43548# 0.028602f
C37671 a_14021_43940# a_15095_43370# 0.001284f
C37672 a_11341_43940# a_15781_43660# 4.59e-21
C37673 a_15493_43396# a_16977_43638# 0.018523f
C37674 a_11967_42832# a_17595_43084# 0.0964f
C37675 a_3499_42826# a_743_42282# 1.89e-19
C37676 a_14539_43914# a_18861_43218# 4.42e-20
C37677 a_5891_43370# a_9114_42852# 1.43e-19
C37678 en_comp a_n2302_39072# 4.43e-20
C37679 a_1209_43370# VDD 0.191694f
C37680 a_8162_45546# a_n2293_42834# 0.001469f
C37681 a_10907_45822# a_1307_43914# 5.29e-20
C37682 a_2711_45572# a_16501_45348# 4.66e-19
C37683 a_20107_45572# a_21297_45572# 2.56e-19
C37684 a_21188_45572# a_3357_43084# 0.057919f
C37685 a_20623_45572# a_19963_31679# 8.99e-21
C37686 a_4361_42308# a_20202_43084# 0.472299f
C37687 a_16977_43638# a_3483_46348# 4.05e-19
C37688 a_5534_30871# a_3090_45724# 0.001578f
C37689 a_n2104_42282# a_n2956_39768# 3.63e-20
C37690 a_n3674_38680# a_n2442_46660# 0.023617f
C37691 a_2982_43646# a_526_44458# 0.048644f
C37692 a_726_44056# a_n357_42282# 4.98e-19
C37693 a_9885_43646# a_9290_44172# 0.008596f
C37694 a_10149_43396# a_8016_46348# 1.24e-19
C37695 a_13575_42558# a_10227_46804# 0.001718f
C37696 a_8049_45260# VDD 1.89366f
C37697 a_6598_45938# a_4883_46098# 6.94e-20
C37698 a_6977_45572# a_6545_47178# 9.76e-20
C37699 a_11136_45572# a_2063_45854# 0.054713f
C37700 a_8034_45724# a_8781_46436# 0.009374f
C37701 a_5066_45546# a_10586_45546# 9.49e-20
C37702 a_2324_44458# a_n2293_45546# 9.66e-19
C37703 a_20708_46348# a_20850_46482# 0.007833f
C37704 a_18985_46122# a_20850_46155# 4.3e-20
C37705 a_n3420_37440# C0_P_btm 0.033333f
C37706 a_15743_43084# a_22223_43396# 0.004521f
C37707 a_8685_43396# a_9127_43156# 0.01312f
C37708 a_2982_43646# a_19164_43230# 1.37e-20
C37709 a_3422_30871# a_4958_30871# 0.101017f
C37710 a_n97_42460# a_5457_43172# 4.93e-20
C37711 a_18114_32519# C0_N_btm 3.38e-19
C37712 a_3059_42968# VDD 8.13e-19
C37713 a_14537_43396# a_11691_44458# 0.092307f
C37714 a_16019_45002# a_11827_44484# 4.4e-20
C37715 a_3537_45260# a_4223_44672# 0.1907f
C37716 a_7229_43940# a_n2661_44458# 0.028622f
C37717 a_n2017_45002# a_14539_43914# 0.01532f
C37718 a_5837_42852# a_526_44458# 0.057897f
C37719 a_17595_43084# a_13259_45724# 0.118887f
C37720 a_5111_42852# a_n357_42282# 0.011577f
C37721 a_4520_42826# a_n755_45592# 2.49e-20
C37722 a_1606_42308# a_1823_45246# 6.6e-20
C37723 VDAC_P w_1575_34946# 0.037571f
C37724 a_n3607_37440# SMPL_ON_P 7.77e-21
C37725 a_11787_45002# a_768_44030# 3.39e-21
C37726 a_13017_45260# a_12891_46348# 0.210934f
C37727 a_6431_45366# a_5807_45002# 0.018543f
C37728 a_2437_43646# a_3524_46660# 1.78e-20
C37729 a_2382_45260# a_n2661_46634# 2.63e-21
C37730 a_n143_45144# a_n1925_46634# 1.28e-21
C37731 a_327_44734# a_n2293_46634# 0.024588f
C37732 a_6171_45002# a_13661_43548# 0.032575f
C37733 a_15415_45028# a_n881_46662# 3.95e-20
C37734 a_22705_38406# VDD 0.085998f
C37735 a_n2661_44458# a_n237_47217# 1.04e-19
C37736 a_n2129_44697# a_n971_45724# 0.017407f
C37737 a_n2433_44484# a_n746_45260# 2.7e-20
C37738 a_2779_44458# a_n2497_47436# 0.034441f
C37739 a_14955_43396# a_15486_42560# 1.53e-19
C37740 a_n2840_42826# a_n1630_35242# 2.09e-20
C37741 a_n2157_42858# a_n3674_37592# 0.001748f
C37742 a_n901_43156# a_n961_42308# 0.002229f
C37743 a_12545_42858# a_13291_42460# 1.52e-19
C37744 a_13113_42826# a_13003_42852# 0.097745f
C37745 a_743_42282# a_3318_42354# 0.01411f
C37746 a_10341_43396# a_14113_42308# 1.45e-20
C37747 a_n3674_39304# a_n4318_37592# 0.023516f
C37748 a_5649_42852# a_1755_42282# 0.023826f
C37749 a_6945_45028# DATA[3] 0.014238f
C37750 a_n2956_39304# CLK_DATA 0.003272f
C37751 a_n3607_39616# VDD 2.79e-20
C37752 a_10227_46804# a_18479_47436# 1.40697f
C37753 a_n443_46116# a_3094_47243# 4.19e-19
C37754 a_4700_47436# a_n1613_43370# 5.19e-21
C37755 a_13717_47436# SMPL_ON_N 0.132417f
C37756 a_15811_47375# a_13507_46334# 0.002419f
C37757 a_11599_46634# a_4883_46098# 0.261488f
C37758 a_16327_47482# a_20894_47436# 4.5e-21
C37759 a_4007_47204# a_n881_46662# 4.68e-20
C37760 a_n1151_42308# a_8128_46384# 0.328697f
C37761 a_14311_47204# a_12465_44636# 0.004308f
C37762 a_2063_45854# a_12891_46348# 4.37e-20
C37763 a_4915_47217# a_5063_47570# 0.003687f
C37764 a_10334_44484# a_n2661_43922# 0.008746f
C37765 a_10440_44484# a_n2661_42834# 7.54e-20
C37766 a_7499_43078# a_10341_43396# 0.061281f
C37767 a_20193_45348# a_20679_44626# 0.017743f
C37768 a_n2293_42834# a_2889_44172# 3.27e-21
C37769 a_9482_43914# a_10729_43914# 0.047853f
C37770 a_10193_42453# a_14205_43396# 5.63e-21
C37771 a_2711_45572# a_18783_43370# 6.16e-20
C37772 a_16922_45042# a_20512_43084# 0.055985f
C37773 a_1307_43914# a_n2661_42282# 0.042336f
C37774 a_8975_43940# a_9159_44484# 0.00805f
C37775 a_11827_44484# a_18245_44484# 1.94e-19
C37776 a_21887_42336# a_13259_45724# 6.84e-19
C37777 a_19237_31679# SMPL_ON_N 0.029331f
C37778 a_n2661_42282# a_n443_46116# 2.25e-20
C37779 a_3232_43370# a_4419_46090# 4.56e-21
C37780 a_5111_44636# a_5164_46348# 0.024532f
C37781 a_5147_45002# a_5204_45822# 3.69e-19
C37782 a_3357_43084# a_19553_46090# 4.81e-21
C37783 a_413_45260# a_9569_46155# 1.76e-20
C37784 en_comp a_10903_43370# 4.34e-21
C37785 a_n2661_45010# a_2324_44458# 0.001752f
C37786 a_13711_45394# a_13059_46348# 6.86e-19
C37787 a_6171_45002# a_4185_45028# 2.76e-20
C37788 a_n2661_44458# a_8270_45546# 0.019483f
C37789 a_18588_44850# a_12549_44172# 1.05e-20
C37790 a_18494_42460# a_19466_46812# 1.2e-19
C37791 a_18184_42460# a_19692_46634# 1.68e-19
C37792 a_14673_44172# a_13661_43548# 0.36897f
C37793 a_5205_44484# a_3483_46348# 0.065176f
C37794 a_11691_44458# a_3090_45724# 0.245063f
C37795 a_21005_45260# a_15227_44166# 3.8e-19
C37796 a_2123_42473# a_6123_31319# 8.95e-21
C37797 a_1606_42308# a_5934_30871# 0.095492f
C37798 a_5379_42460# a_4921_42308# 0.033756f
C37799 a_2713_42308# a_5932_42308# 4.34e-21
C37800 a_5267_42460# a_5337_42558# 0.011552f
C37801 a_13467_32519# C6_N_btm 1.49e-19
C37802 a_13678_32519# C3_N_btm 0.001771f
C37803 a_22521_39511# a_22717_37285# 2.12e-20
C37804 a_12549_44172# a_11901_46660# 0.001645f
C37805 a_n2661_46634# a_10623_46897# 0.006678f
C37806 a_2443_46660# a_4651_46660# 1.35e-19
C37807 a_3524_46660# a_3686_47026# 0.006453f
C37808 a_2959_46660# a_3221_46660# 0.001705f
C37809 a_12891_46348# a_12469_46902# 0.009064f
C37810 a_2609_46660# a_4646_46812# 4.37e-20
C37811 a_3177_46902# a_3877_44458# 3.33e-19
C37812 a_2107_46812# a_3633_46660# 2.47e-19
C37813 a_11309_47204# a_12251_46660# 1.48e-19
C37814 a_n881_46662# a_15368_46634# 0.023127f
C37815 a_13507_46334# a_13059_46348# 0.192049f
C37816 a_10227_46804# a_17829_46910# 4.34e-19
C37817 a_18479_47436# a_17339_46660# 3.12e-20
C37818 a_11599_46634# a_21188_46660# 3.88e-21
C37819 a_16327_47482# a_20411_46873# 5.72e-19
C37820 a_18143_47464# a_765_45546# 0.001396f
C37821 a_12861_44030# a_16434_46660# 0.001465f
C37822 a_n237_47217# a_2804_46116# 0.039625f
C37823 a_n971_45724# a_3483_46348# 0.211534f
C37824 a_584_46384# a_1208_46090# 0.034313f
C37825 a_1431_47204# a_1138_42852# 1.47e-19
C37826 a_n1151_42308# a_n1641_46494# 0.003575f
C37827 a_2063_45854# a_805_46414# 8.93e-20
C37828 a_n2109_47186# a_5204_45822# 7.25e-19
C37829 a_n1741_47186# a_5068_46348# 1.28e-20
C37830 a_949_44458# a_1756_43548# 0.001231f
C37831 a_1414_42308# a_895_43940# 0.208524f
C37832 a_17517_44484# a_19328_44172# 7.19e-21
C37833 a_n699_43396# a_1209_43370# 0.004475f
C37834 a_5891_43370# a_5745_43940# 2.82e-19
C37835 a_742_44458# a_4093_43548# 2.85e-20
C37836 a_18989_43940# a_18533_43940# 0.001685f
C37837 a_453_43940# a_2479_44172# 0.003275f
C37838 a_11967_42832# a_10807_43548# 1.1e-20
C37839 a_10193_42453# a_22400_42852# 3.3e-21
C37840 a_n2293_43922# a_12710_44260# 9.27e-19
C37841 a_n913_45002# a_5755_42852# 1.7e-20
C37842 a_n1059_45260# a_7227_42852# 0.005565f
C37843 a_n2017_45002# a_7871_42858# 1.28e-19
C37844 a_22469_40625# VDD 0.564837f
C37845 a_8103_44636# VDD 0.124028f
C37846 a_7174_31319# C2_P_btm 1.86e-20
C37847 a_n3565_39590# a_n1386_35608# 1.44e-19
C37848 a_20712_42282# RST_Z 4.07e-20
C37849 a_4958_30871# VREF_GND 0.054206f
C37850 a_n2860_37984# a_n2956_38216# 0.001353f
C37851 a_17061_44734# a_3483_46348# 0.009179f
C37852 a_22315_44484# a_11415_45002# 0.001541f
C37853 a_8333_44056# a_3090_45724# 0.001679f
C37854 a_7499_43940# a_4646_46812# 0.002542f
C37855 a_n2661_43370# a_n23_45546# 3.29e-20
C37856 a_17896_45144# a_13259_45724# 9.29e-19
C37857 a_n2661_43922# a_9290_44172# 0.029391f
C37858 a_8147_43396# a_n1613_43370# 3.58e-19
C37859 a_13667_43396# a_12465_44636# 2.31e-21
C37860 a_15781_43660# a_16327_47482# 7.49e-21
C37861 a_16759_43396# a_12861_44030# 2.75e-20
C37862 a_4361_42308# a_2063_45854# 1.32e-20
C37863 a_n13_43084# a_n2497_47436# 1.74e-20
C37864 a_743_42282# a_n1151_42308# 1.08e-19
C37865 a_1239_39587# a_1736_39587# 0.105143f
C37866 a_n3690_39616# a_n3690_39392# 0.052468f
C37867 a_n3420_39616# a_n3565_39304# 0.035199f
C37868 a_n4064_39616# a_n4209_39304# 0.029393f
C37869 a_n3565_39590# a_n3420_39072# 0.033891f
C37870 a_n4209_39590# a_n4064_39072# 0.03458f
C37871 a_n2442_46660# VDD 0.693209f
C37872 a_5932_42308# C8_N_btm 1.4e-19
C37873 a_6123_31319# C3_N_btm 0.011333f
C37874 a_5934_30871# C1_N_btm 0.011025f
C37875 a_19692_46634# a_12741_44636# 0.022879f
C37876 a_17339_46660# a_17829_46910# 1.33e-19
C37877 a_2107_46812# a_526_44458# 0.008773f
C37878 a_n743_46660# a_5066_45546# 0.124676f
C37879 a_22612_30879# a_8049_45260# 7.79e-20
C37880 a_n2661_46098# a_n967_46494# 8.5e-19
C37881 a_6755_46942# a_7920_46348# 1.43e-19
C37882 a_10623_46897# a_8199_44636# 3.42e-19
C37883 a_10150_46912# a_9625_46129# 2.39e-19
C37884 a_10249_46116# a_8016_46348# 0.001301f
C37885 a_10227_46804# a_n443_42852# 0.043674f
C37886 a_9313_44734# a_8037_42858# 5.36e-20
C37887 a_18248_44752# a_18249_42858# 1.79e-20
C37888 a_18287_44626# a_17333_42852# 2.93e-20
C37889 a_20835_44721# a_4190_30871# 1.12e-20
C37890 a_5891_43370# a_10518_42984# 0.001688f
C37891 a_17737_43940# a_3626_43646# 5.73e-21
C37892 a_18579_44172# a_16823_43084# 1.17e-21
C37893 a_n2293_42834# a_n4318_37592# 0.003537f
C37894 a_n2661_42834# a_1847_42826# 6.72e-21
C37895 a_n2293_43922# a_685_42968# 8.95e-21
C37896 a_20512_43084# a_15743_43084# 0.761578f
C37897 a_14539_43914# a_19164_43230# 7.82e-21
C37898 a_n356_44636# a_5534_30871# 0.054103f
C37899 a_3499_42826# a_2813_43396# 2.45e-19
C37900 a_11967_42832# a_13467_32519# 3.36e-21
C37901 a_3537_45260# a_5742_30871# 3.39e-20
C37902 en_comp a_15959_42545# 3.92e-20
C37903 a_11173_44260# VDD 0.005546f
C37904 a_16680_45572# a_18341_45572# 6.97e-20
C37905 a_17478_45572# a_16147_45260# 0.050291f
C37906 a_8696_44636# a_18479_45785# 1.47e-20
C37907 a_15861_45028# a_18175_45572# 8.48e-20
C37908 a_6472_45840# a_5205_44484# 2.12e-20
C37909 a_6511_45714# a_6431_45366# 6.29e-19
C37910 a_6667_45809# a_6171_45002# 0.004899f
C37911 a_2711_45572# a_8953_45002# 0.003719f
C37912 a_14097_32519# a_13507_46334# 0.001207f
C37913 a_22959_43948# a_8049_45260# 1.04e-19
C37914 a_2253_43940# a_526_44458# 9.54e-20
C37915 a_7542_44172# a_n357_42282# 2.72e-19
C37916 a_453_43940# a_n443_42852# 0.005083f
C37917 a_4190_30871# a_3090_45724# 1.55e-21
C37918 a_3539_42460# a_1823_45246# 0.678673f
C37919 a_11206_38545# CAL_P 0.234643f
C37920 a_22469_40625# a_22469_39537# 0.604831f
C37921 a_n4209_37414# C9_P_btm 1.91e-20
C37922 a_19721_31679# a_21589_35634# 1.38e-20
C37923 a_8953_45546# VDD 1.32809f
C37924 a_5907_45546# a_n237_47217# 1.7e-19
C37925 a_6472_45840# a_n971_45724# 5.6e-19
C37926 a_n4209_38502# a_n4209_37414# 0.028607f
C37927 a_12741_44636# a_20692_30879# 7.57e-19
C37928 a_22959_46660# a_20205_31679# 0.00182f
C37929 a_765_45546# a_509_45822# 0.008717f
C37930 a_5937_45572# a_8034_45724# 0.052916f
C37931 a_7920_46348# a_8049_45260# 0.003857f
C37932 a_20708_46348# a_10809_44734# 1.69e-21
C37933 a_n809_44244# a_n473_42460# 1.26e-20
C37934 a_6197_43396# a_743_42282# 3.82e-20
C37935 a_10341_43396# a_15781_43660# 0.011941f
C37936 a_14021_43940# a_22959_42860# 3.35e-19
C37937 a_n97_42460# a_685_42968# 0.034735f
C37938 a_13565_43940# a_12379_42858# 1.27e-20
C37939 a_n984_44318# a_n961_42308# 1.84e-20
C37940 a_n1761_44111# a_n3674_37592# 0.002395f
C37941 a_1568_43370# a_n13_43084# 1.85e-20
C37942 a_14579_43548# a_16547_43609# 5.47e-21
C37943 a_n1613_43370# DATA[2] 3.98e-20
C37944 a_n881_46662# DATA[1] 8.44e-22
C37945 a_21588_30879# a_22609_37990# 1.43e-20
C37946 a_n722_43218# VDD 1.22e-19
C37947 a_15599_45572# a_16112_44458# 7.05e-19
C37948 a_15595_45028# a_16019_45002# 0.017418f
C37949 a_15415_45028# a_1307_43914# 1.07e-19
C37950 a_8696_44636# a_10057_43914# 0.001707f
C37951 a_9482_43914# a_1423_45028# 0.014596f
C37952 a_7499_43078# a_n2293_43922# 1.48e-19
C37953 a_9049_44484# a_n2661_43922# 0.003185f
C37954 a_8746_45002# a_10617_44484# 0.01623f
C37955 a_2711_45572# a_16335_44484# 0.001233f
C37956 a_n37_45144# a_n2661_43370# 0.007073f
C37957 a_5111_44636# a_5837_45028# 0.019542f
C37958 a_3537_45260# a_n2293_42834# 0.195818f
C37959 a_4927_45028# a_5093_45028# 0.143754f
C37960 a_21513_45002# a_21101_45002# 0.003301f
C37961 a_n2946_39866# a_n2312_38680# 3.47e-20
C37962 a_n2860_39866# a_n2442_46660# 6.14e-19
C37963 a_16977_43638# a_n357_42282# 6.48e-19
C37964 a_7871_42858# a_526_44458# 0.031818f
C37965 a_13467_32519# a_13259_45724# 0.030863f
C37966 a_8873_43396# a_n443_42852# 8.24e-20
C37967 a_17701_42308# a_17715_44484# 0.002546f
C37968 a_413_45260# a_19386_47436# 1.03e-19
C37969 a_8953_45002# a_9313_45822# 0.001732f
C37970 a_626_44172# a_n1151_42308# 3.18e-21
C37971 a_2437_43646# a_4842_47570# 8.98e-19
C37972 a_15861_45028# a_n743_46660# 0.005332f
C37973 a_18341_45572# a_13747_46662# 0.554429f
C37974 a_18691_45572# a_5807_45002# 0.001465f
C37975 a_18175_45572# a_19321_45002# 0.01259f
C37976 a_8568_45546# a_8492_46660# 2.74e-20
C37977 a_18909_45814# a_13661_43548# 0.006912f
C37978 a_7499_43078# a_8667_46634# 1.51e-19
C37979 a_6293_42852# a_6171_42473# 0.00101f
C37980 a_6031_43396# a_5932_42308# 3.68e-19
C37981 a_1847_42826# a_n2293_42282# 4.45e-19
C37982 a_12379_42858# a_5534_30871# 0.128429f
C37983 a_12545_42858# a_13460_43230# 0.118423f
C37984 a_n97_42460# a_14113_42308# 0.356407f
C37985 a_3539_42460# a_5934_30871# 1.41e-20
C37986 a_3626_43646# a_8515_42308# 0.003306f
C37987 a_15743_43084# a_16245_42852# 4.92e-19
C37988 a_20820_30879# VREF 0.195875f
C37989 a_n1853_46287# DATA[0] 2.73e-20
C37990 a_3422_30871# C7_N_btm 2.94e-19
C37991 a_11206_38545# CAL_N 0.050483f
C37992 a_14456_42282# VDD 0.265543f
C37993 a_n23_47502# a_n1435_47204# 4.14e-19
C37994 a_n1151_42308# a_6151_47436# 0.026437f
C37995 a_2063_45854# a_7903_47542# 1.25e-20
C37996 a_3785_47178# a_5129_47502# 4.3e-19
C37997 a_3815_47204# a_4915_47217# 2.1e-19
C37998 a_4700_47436# a_4791_45118# 0.31818f
C37999 a_4007_47204# a_n443_46116# 0.006041f
C38000 a_19431_45546# a_15493_43396# 1.48e-19
C38001 a_8696_44636# a_14021_43940# 2.1e-19
C38002 a_5343_44458# a_5518_44484# 0.054464f
C38003 a_7499_43078# a_n97_42460# 0.212833f
C38004 a_2711_45572# a_3626_43646# 0.072582f
C38005 a_3065_45002# a_1414_42308# 4.93e-19
C38006 a_413_45260# a_2889_44172# 0.127135f
C38007 a_n2293_45010# a_n1453_44318# 0.001505f
C38008 a_n2017_45002# a_n3674_39768# 2.64e-19
C38009 a_1149_42558# a_n863_45724# 0.002168f
C38010 a_564_42282# a_n755_45592# 0.036154f
C38011 a_n1630_35242# a_n357_42282# 0.086672f
C38012 a_6812_45938# VDD 0.132317f
C38013 a_17364_32525# a_18194_35068# 9.45e-20
C38014 a_22469_40625# a_22612_30879# 7.32e-20
C38015 a_n2661_43370# a_8492_46660# 1.86e-21
C38016 a_3357_43084# a_12741_44636# 0.036536f
C38017 a_14537_43396# a_15227_44166# 0.105881f
C38018 a_18443_44721# a_12549_44172# 1.36e-19
C38019 a_4223_44672# a_n2293_46634# 3.24e-21
C38020 a_12607_44458# a_13661_43548# 0.00102f
C38021 a_20447_31679# a_20202_43084# 8.03e-21
C38022 a_16751_45260# a_14976_45028# 1.25e-20
C38023 a_22591_45572# a_20820_30879# 9.76e-21
C38024 a_22959_45572# a_11415_45002# 0.001334f
C38025 a_19963_31679# a_22591_46660# 1.81e-20
C38026 a_15037_45618# a_15015_46420# 0.001025f
C38027 a_12016_45572# a_2324_44458# 2.57e-19
C38028 a_15146_44811# a_10227_46804# 6.31e-20
C38029 a_17517_44484# a_12861_44030# 0.069119f
C38030 a_644_44056# a_n2497_47436# 0.016428f
C38031 a_16414_43172# a_4958_30871# 8.46e-19
C38032 a_n2472_42282# a_n2104_42282# 7.52e-19
C38033 a_n3674_38680# a_n3674_38216# 0.059687f
C38034 a_9061_43230# a_5934_30871# 5.05e-21
C38035 a_n2956_39768# a_n2661_46634# 0.006224f
C38036 a_n2840_46634# a_n2472_46634# 7.52e-19
C38037 a_n1613_43370# a_3067_47026# 0.013046f
C38038 a_4883_46098# a_7411_46660# 4.36e-20
C38039 a_10227_46804# a_10554_47026# 0.166977f
C38040 a_2063_45854# a_12359_47026# 9.65e-22
C38041 a_n1741_47186# a_13059_46348# 0.001771f
C38042 a_4915_47217# a_14976_45028# 3.23e-21
C38043 a_11031_47542# a_11186_47026# 2.5e-19
C38044 a_6151_47436# a_14084_46812# 5.28e-21
C38045 a_17767_44458# a_17737_43940# 0.004352f
C38046 a_11967_42832# a_22315_44484# 6.72e-19
C38047 a_n2661_43922# a_3905_42865# 3.56e-19
C38048 a_n2661_42834# a_5244_44056# 0.00436f
C38049 a_n2293_42834# a_1049_43396# 0.001716f
C38050 a_1307_43914# a_7112_43396# 3.85e-21
C38051 a_19279_43940# a_18579_44172# 0.372064f
C38052 a_16922_45042# a_21381_43940# 0.003996f
C38053 a_n913_45002# a_16759_43396# 3.29e-21
C38054 a_n2017_45002# a_17324_43396# 1.13e-19
C38055 a_n1059_45260# a_17499_43370# 0.385066f
C38056 a_7735_45067# VDD 2.18e-20
C38057 a_5934_30871# C9_P_btm 1.37e-19
C38058 a_6123_31319# C7_P_btm 0.005631f
C38059 a_5932_42308# C2_P_btm 0.011289f
C38060 a_20692_30879# C9_N_btm 1.64e-19
C38061 a_20205_31679# C10_N_btm 2.25e-20
C38062 a_11827_44484# a_6945_45028# 8.14e-20
C38063 a_5343_44458# a_8199_44636# 7.94e-19
C38064 a_5205_44484# a_n357_42282# 3.84e-20
C38065 a_2274_45254# a_n443_42852# 1.98e-21
C38066 a_1667_45002# a_1609_45822# 0.001741f
C38067 a_8137_45348# a_8049_45260# 2.64e-19
C38068 a_15493_43940# a_n2293_46634# 0.003183f
C38069 a_14761_44260# a_13661_43548# 5.06e-19
C38070 a_3992_43940# a_768_44030# 0.006422f
C38071 a_20362_44736# a_19692_46634# 3.19e-21
C38072 a_20835_44721# a_15227_44166# 4.95e-20
C38073 a_13076_44458# a_3483_46348# 4.08e-21
C38074 a_18780_47178# VDD 0.245515f
C38075 a_4958_30871# a_7174_31319# 0.107892f
C38076 a_17303_42282# a_20712_42282# 3.71e-19
C38077 a_5742_30871# a_1343_38525# 1.5e-19
C38078 a_18907_42674# a_19511_42282# 0.001351f
C38079 a_5934_30871# a_n4209_38502# 6.81e-22
C38080 a_6123_31319# a_n3565_38502# 3.8e-21
C38081 a_1983_46706# a_167_45260# 2.62e-20
C38082 a_1799_45572# a_472_46348# 5.48e-20
C38083 a_n2661_46098# a_376_46348# 0.060405f
C38084 a_2107_46812# a_2521_46116# 0.008501f
C38085 a_1110_47026# a_1176_45822# 6.94e-20
C38086 a_3090_45724# a_15227_44166# 0.428743f
C38087 a_12469_46902# a_12359_47026# 0.097745f
C38088 a_12251_46660# a_12156_46660# 0.049827f
C38089 a_6755_46942# a_14447_46660# 0.001822f
C38090 a_n743_46660# a_5068_46348# 0.005784f
C38091 a_12549_44172# a_17583_46090# 3.17e-20
C38092 a_5807_45002# a_12005_46116# 0.004606f
C38093 a_n1925_46634# a_5204_45822# 2.89e-19
C38094 a_13661_43548# a_10903_43370# 9.73e-19
C38095 a_11599_46634# a_11608_46482# 7.81e-19
C38096 a_584_46384# a_n2661_45546# 0.100439f
C38097 a_n746_45260# a_310_45028# 0.378188f
C38098 a_n971_45724# a_n357_42282# 0.271282f
C38099 a_n452_47436# a_n755_45592# 1.25e-21
C38100 a_742_44458# a_685_42968# 9.87e-20
C38101 a_1115_44172# a_1049_43396# 3.25e-19
C38102 a_1467_44172# a_1209_43370# 0.004302f
C38103 a_3600_43914# a_n97_42460# 3.85e-21
C38104 a_20365_43914# a_14021_43940# 0.003393f
C38105 a_14673_44172# a_14579_43548# 2.2e-20
C38106 a_n4318_39768# a_n2840_43370# 7.62e-19
C38107 a_9313_44734# a_18525_43370# 8.26e-20
C38108 a_n356_44636# a_4190_30871# 0.04771f
C38109 a_14537_43396# a_14635_42282# 4.55e-19
C38110 a_n2293_42834# a_4649_43172# 2.27e-19
C38111 a_n967_45348# a_n784_42308# 0.007598f
C38112 a_n913_45002# a_1067_42314# 9.28e-20
C38113 a_n1059_45260# a_1576_42282# 0.003521f
C38114 a_n2017_45002# a_1184_42692# 0.040166f
C38115 a_n2956_37592# a_n3674_37592# 0.025613f
C38116 a_895_43940# VDD 0.318652f
C38117 a_10193_42453# a_16680_45572# 1.46e-20
C38118 a_8697_45822# a_8697_45572# 6.96e-20
C38119 a_10180_45724# a_8696_44636# 0.002551f
C38120 C7_N_btm VREF_GND 1.61142f
C38121 C6_N_btm VCM 0.877241f
C38122 C8_N_btm VREF 3.6701f
C38123 C9_N_btm VIN_N 1.82823f
C38124 a_3353_43940# a_1823_45246# 4.96e-20
C38125 a_15301_44260# a_3483_46348# 6.81e-19
C38126 a_19319_43548# a_11415_45002# 2.49e-20
C38127 a_n1991_42858# a_n2438_43548# 9.37e-19
C38128 a_9145_43396# a_8270_45546# 0.02247f
C38129 a_9127_43156# a_768_44030# 1.24e-19
C38130 a_n4318_38680# a_n2442_46660# 0.023781f
C38131 a_6655_43762# a_3090_45724# 0.002552f
C38132 a_14815_43914# a_n443_42852# 8.61e-20
C38133 a_14955_43940# a_2324_44458# 0.029449f
C38134 a_10555_44260# a_8016_46348# 0.007104f
C38135 a_9801_44260# a_8199_44636# 6.23e-19
C38136 a_22959_42860# a_13507_46334# 0.004407f
C38137 a_18285_46348# VDD 0.259614f
C38138 a_n4064_40160# a_n3690_38304# 3.42e-19
C38139 a_19466_46812# a_19240_46482# 0.003742f
C38140 a_3483_46348# a_12594_46348# 0.011082f
C38141 a_4185_45028# a_10903_43370# 1.24e-19
C38142 a_1138_42852# a_2324_44458# 9.6e-21
C38143 a_21542_46660# a_10809_44734# 4.32e-19
C38144 a_8016_46348# a_5937_45572# 0.021789f
C38145 a_8349_46414# a_8199_44636# 0.032352f
C38146 a_10729_43914# a_10796_42968# 7.16e-21
C38147 a_10949_43914# a_10835_43094# 4.11e-21
C38148 a_8147_43396# a_8791_43396# 0.001846f
C38149 a_10807_43548# a_10518_42984# 7.97e-19
C38150 a_n97_42460# a_15781_43660# 0.001962f
C38151 a_21381_43940# a_15743_43084# 0.02274f
C38152 a_18184_42460# a_20107_42308# 0.013525f
C38153 a_18494_42460# a_13258_32519# 0.298557f
C38154 a_n2293_43922# a_n1329_42308# 4.07e-19
C38155 a_6547_43396# a_6655_43762# 0.057222f
C38156 a_11967_42832# a_18695_43230# 0.001256f
C38157 a_4791_45118# DATA[2] 7.19e-19
C38158 a_4700_47436# DATA[3] 3.7e-20
C38159 a_20447_31679# C5_N_btm 0.040445f
C38160 a_19479_31679# C10_N_btm 2.25e-20
C38161 a_19963_31679# C7_N_btm 1.43e-20
C38162 a_2274_45254# a_2680_45002# 0.076507f
C38163 a_413_45260# a_3537_45260# 3.32e-19
C38164 a_4361_42308# a_17715_44484# 6.15e-21
C38165 a_n1557_42282# a_n755_45592# 0.199254f
C38166 a_5742_30871# a_n2293_46634# 2.68e-19
C38167 a_14635_42282# a_3090_45724# 0.007468f
C38168 a_5342_30871# a_12741_44636# 1.14e-22
C38169 a_3422_30871# C3_P_btm 1.1e-19
C38170 a_19237_31679# a_18194_35068# 7.27e-20
C38171 a_1609_45822# VDD 0.270106f
C38172 a_13249_42308# a_12549_44172# 0.066967f
C38173 a_13904_45546# a_768_44030# 0.005947f
C38174 a_10490_45724# a_5807_45002# 4.75e-23
C38175 a_3775_45552# a_n743_46660# 3.52e-20
C38176 a_4099_45572# a_2107_46812# 4.87e-20
C38177 a_10193_42453# a_13747_46662# 7.93e-21
C38178 a_3260_45572# a_n2293_46634# 3.64e-19
C38179 a_8696_44636# a_13507_46334# 3.72e-19
C38180 a_18341_45572# a_11599_46634# 0.588263f
C38181 a_16377_45572# a_16327_47482# 0.001903f
C38182 a_2437_43646# a_3785_47178# 0.015875f
C38183 a_n745_45366# a_n971_45724# 1.48e-20
C38184 a_n913_45002# a_n746_45260# 0.051081f
C38185 a_n37_45144# a_n2497_47436# 2.82e-20
C38186 a_n967_45348# SMPL_ON_P 5.24e-20
C38187 a_19692_46634# RST_Z 3.49e-20
C38188 a_15682_43940# a_16104_42674# 1.03e-20
C38189 a_n2433_43396# a_n1630_35242# 2.03e-20
C38190 a_n2267_43396# a_n3674_37592# 1.26e-20
C38191 a_18525_43370# a_18599_43230# 4.07e-19
C38192 a_15743_43084# a_18249_42858# 0.002881f
C38193 a_18783_43370# a_18817_42826# 0.012757f
C38194 a_n901_43156# a_685_42968# 1.06e-20
C38195 a_5649_42852# a_8387_43230# 1.14e-20
C38196 a_4361_42308# a_10083_42826# 1.21e-19
C38197 a_743_42282# a_10922_42852# 1.14e-20
C38198 a_n1809_43762# a_n1736_42282# 1.55e-20
C38199 a_3422_30871# a_n4064_38528# 0.031148f
C38200 a_n13_43084# a_133_43172# 0.013377f
C38201 a_n3674_39304# a_n1533_42852# 8.15e-22
C38202 a_n4318_39768# a_n4315_30879# 0.002449f
C38203 a_8685_43396# a_9306_43218# 1.84e-19
C38204 a_19466_46812# START 9.72e-20
C38205 a_15009_46634# CLK 1.39e-20
C38206 a_n3690_38304# a_n4064_37440# 6.81e-20
C38207 a_n3420_37984# a_n2946_37690# 2.59e-20
C38208 a_n4064_37984# a_n3690_37440# 6.81e-20
C38209 a_n2946_37984# a_n3420_37440# 2.59e-20
C38210 a_n3674_38216# VDD 0.309006f
C38211 a_18494_42460# a_20193_45348# 0.116597f
C38212 a_n2661_43370# a_949_44458# 6.02e-19
C38213 a_375_42282# a_n356_44636# 0.015238f
C38214 a_13904_45546# a_13483_43940# 2.98e-21
C38215 a_10193_42453# a_20269_44172# 3.41e-21
C38216 a_17719_45144# a_17969_45144# 0.008267f
C38217 a_16922_45042# a_19929_45028# 0.003656f
C38218 a_13249_42308# a_12429_44172# 5.54e-19
C38219 a_5111_44636# a_n2661_42834# 0.04935f
C38220 a_5147_45002# a_n2661_43922# 0.029995f
C38221 a_3232_43370# a_10617_44484# 0.020516f
C38222 a_15959_42545# a_4185_45028# 1.27e-19
C38223 a_21887_42336# a_20202_43084# 0.082645f
C38224 a_3863_42891# a_n357_42282# 3.29e-19
C38225 a_1184_42692# a_526_44458# 6.23e-19
C38226 a_1576_42282# a_n1925_42282# 1.31e-19
C38227 a_945_42968# a_n443_42852# 9.8e-19
C38228 a_8483_43230# a_n755_45592# 2.93e-19
C38229 a_10545_42558# a_9290_44172# 6.22e-19
C38230 CAL_N a_10227_46804# 7.26e-19
C38231 a_13720_44458# a_12861_44030# 4.84e-19
C38232 a_3363_44484# a_n971_45724# 4.12e-21
C38233 a_556_44484# a_n746_45260# 0.045671f
C38234 a_5891_43370# a_2063_45854# 1.78e-19
C38235 a_2711_45572# a_15015_46420# 1.15e-20
C38236 a_4808_45572# a_5937_45572# 6.9e-20
C38237 a_21188_45572# a_19466_46812# 4.5e-20
C38238 a_n1059_45260# a_8270_45546# 5.56e-20
C38239 a_6171_45002# a_5257_43370# 3.04e-19
C38240 a_21363_45546# a_19692_46634# 8.99e-19
C38241 a_413_45260# a_6969_46634# 2.65e-20
C38242 a_3357_43084# a_13607_46688# 1.82e-20
C38243 a_2437_43646# a_3090_45724# 1.6e-19
C38244 a_3232_43370# a_7411_46660# 8.54e-22
C38245 a_20731_45938# a_15227_44166# 3.88e-19
C38246 a_n2293_42834# a_n2293_46634# 0.027042f
C38247 a_17613_45144# a_12549_44172# 7.44e-21
C38248 a_11322_45546# a_3483_46348# 0.554731f
C38249 a_4361_42308# a_15761_42308# 1.23e-19
C38250 a_8605_42826# a_5934_30871# 6.8e-19
C38251 a_n2293_42282# a_n473_42460# 2.57e-19
C38252 a_8037_42858# a_8515_42308# 6.68e-20
C38253 a_4190_30871# a_18727_42674# 0.035226f
C38254 a_743_42282# a_17531_42308# 0.007539f
C38255 a_20692_30879# RST_Z 0.051046f
C38256 a_4883_46098# a_13661_43548# 0.032161f
C38257 a_20990_47178# a_19594_46812# 9.2e-20
C38258 a_20894_47436# a_20843_47204# 0.134298f
C38259 a_10227_46804# a_n2661_46634# 0.030546f
C38260 a_15811_47375# a_n743_46660# 8.06e-19
C38261 a_n1435_47204# a_948_46660# 7.47e-21
C38262 a_n1741_47186# a_7577_46660# 1.46e-20
C38263 a_2063_45854# a_4817_46660# 8.38e-20
C38264 a_2905_45572# a_4646_46812# 2.42e-21
C38265 a_n443_46116# a_2864_46660# 0.006317f
C38266 a_3160_47472# a_3877_44458# 2.11e-19
C38267 a_n1151_42308# a_3221_46660# 8.15e-21
C38268 a_n2840_44458# a_n3674_39768# 0.005491f
C38269 a_2779_44458# a_2889_44172# 0.005445f
C38270 a_n699_43396# a_895_43940# 0.001028f
C38271 a_n4318_40392# a_n4318_39768# 2.73673f
C38272 a_n2661_43922# a_12553_44484# 0.009634f
C38273 a_1307_43914# a_9801_43940# 0.004166f
C38274 a_n2661_43370# a_11341_43940# 8.02e-20
C38275 a_3357_43084# a_6293_42852# 0.001183f
C38276 a_n2810_45028# a_n1557_42282# 9.47e-21
C38277 a_3065_45002# VDD 0.501045f
C38278 COMP_P a_22521_39511# 1.79e-19
C38279 a_16237_45028# a_12741_44636# 0.00167f
C38280 a_n356_44636# a_15227_44166# 8.76e-20
C38281 a_4181_44734# a_3090_45724# 0.003724f
C38282 a_n1331_43914# a_n2438_43548# 7.33e-21
C38283 a_5111_44636# a_5066_45546# 7.73e-19
C38284 a_8560_45348# a_8199_44636# 0.03862f
C38285 a_n2661_43370# a_5497_46414# 4.83e-21
C38286 a_n2661_42282# a_n1613_43370# 0.017743f
C38287 a_18079_43940# a_11453_44696# 1.52e-19
C38288 a_15493_43940# a_18597_46090# 0.024181f
C38289 a_n2433_43396# a_n971_45724# 8.25e-19
C38290 a_104_43370# a_n2497_47436# 0.001117f
C38291 a_12563_42308# a_13070_42354# 0.001596f
C38292 a_n1630_35242# a_n4064_40160# 1.13e-19
C38293 a_n4318_37592# a_n4064_39616# 0.021014f
C38294 a_5932_42308# a_4958_30871# 0.01835f
C38295 a_n3674_37592# a_n4251_40480# 9.61e-20
C38296 w_1575_34946# VDD 1.58877f
C38297 a_5342_30871# C9_N_btm 5.28e-19
C38298 C3_P_btm VREF_GND 0.67174f
C38299 C4_P_btm VCM 0.716447f
C38300 C2_P_btm VREF 0.987884f
C38301 a_n743_46660# a_13059_46348# 0.060636f
C38302 a_10150_46912# a_6755_46942# 0.006336f
C38303 a_7577_46660# a_7832_46660# 0.056391f
C38304 a_10428_46928# a_10249_46116# 0.704177f
C38305 a_10467_46802# a_10554_47026# 0.07009f
C38306 a_5257_43370# a_6903_46660# 3.74e-20
C38307 a_19594_46812# a_20273_46660# 1.32e-19
C38308 a_13747_46662# a_21363_46634# 8.65e-20
C38309 a_12465_44636# a_3483_46348# 0.210833f
C38310 a_4883_46098# a_4185_45028# 7.37e-19
C38311 a_n237_47217# a_n1925_42282# 0.109762f
C38312 a_13717_47436# a_13759_46122# 3.79e-20
C38313 a_12861_44030# a_13351_46090# 1.04e-19
C38314 a_11599_46634# a_11387_46155# 0.035936f
C38315 a_10227_46804# a_8199_44636# 0.460391f
C38316 a_18494_42460# a_20301_43646# 0.006153f
C38317 a_15004_44636# a_9145_43396# 3.39e-20
C38318 a_9482_43914# a_15567_42826# 1.86e-19
C38319 a_11967_42832# a_19319_43548# 5.45e-20
C38320 a_6109_44484# a_6031_43396# 0.007586f
C38321 a_n2661_43922# a_4093_43548# 4.66e-20
C38322 a_14537_43396# a_14543_43071# 9.84e-19
C38323 a_18184_42460# a_743_42282# 0.126294f
C38324 a_1307_43914# a_12545_42858# 4.9e-21
C38325 a_13556_45296# a_5342_30871# 1.19e-20
C38326 a_7499_43078# a_10533_42308# 0.225871f
C38327 a_16922_45042# a_5649_42852# 8.28e-21
C38328 a_n2293_42834# a_n1533_42852# 0.003489f
C38329 a_n1059_45260# a_4649_42852# 0.003629f
C38330 a_n4064_38528# VREF_GND 0.034351f
C38331 a_15463_44811# VDD 6.37e-19
C38332 a_2711_45572# a_12791_45546# 0.008464f
C38333 a_4743_44484# a_n443_42852# 1.62e-20
C38334 a_10849_43646# a_n2293_46634# 0.001727f
C38335 a_11257_43940# a_3090_45724# 6.36e-20
C38336 a_13829_44260# a_13059_46348# 0.002505f
C38337 a_16243_43396# a_13661_43548# 0.001958f
C38338 a_6031_43396# a_4646_46812# 0.849684f
C38339 a_19700_43370# a_12549_44172# 7.13e-19
C38340 a_n2661_42282# a_n2293_46098# 0.182071f
C38341 a_10949_43914# a_11415_45002# 1.43e-20
C38342 a_3357_43084# RST_Z 0.031959f
C38343 a_n4209_38216# a_n4334_38304# 0.253307f
C38344 a_10249_46116# VDD 1.03004f
C38345 a_7174_31319# C7_N_btm 9.97e-20
C38346 a_n2840_46090# a_n2293_46098# 0.003755f
C38347 a_n743_46660# a_3218_45724# 1.78e-20
C38348 a_383_46660# a_310_45028# 4.66e-21
C38349 a_10150_46912# a_8049_45260# 2.18e-20
C38350 a_601_46902# a_n357_42282# 7.55e-20
C38351 a_15227_44166# a_20075_46420# 0.060002f
C38352 a_13059_46348# a_11189_46129# 6.1e-21
C38353 a_14035_46660# a_13759_46122# 0.162408f
C38354 a_19466_46812# a_19553_46090# 0.001855f
C38355 a_19692_46634# a_18985_46122# 4.31e-19
C38356 a_19333_46634# a_19335_46494# 4.28e-19
C38357 a_15559_46634# a_6945_45028# 1.52e-20
C38358 a_13885_46660# a_13925_46122# 0.004214f
C38359 a_14976_45028# a_10809_44734# 0.001621f
C38360 a_n1630_35242# a_n4064_37440# 2.18e-20
C38361 a_1606_42308# a_8530_39574# 0.006802f
C38362 a_n97_42460# a_1756_43548# 0.052563f
C38363 a_14021_43940# a_14205_43396# 0.008914f
C38364 a_11341_43940# a_15681_43442# 1.37e-20
C38365 a_15493_43396# a_16409_43396# 0.566182f
C38366 a_11967_42832# a_16795_42852# 0.061673f
C38367 a_n2129_43609# a_n1557_42282# 9.91e-21
C38368 a_n356_44636# a_14635_42282# 1.57e-19
C38369 a_14539_43914# a_17749_42852# 0.002266f
C38370 a_n2956_37592# a_n2302_39072# 0.005021f
C38371 a_458_43396# VDD 0.431902f
C38372 a_2711_45572# a_16405_45348# 5.81e-19
C38373 a_16115_45572# a_6171_45002# 3.23e-20
C38374 a_20841_45814# a_19963_31679# 5.16e-20
C38375 a_21188_45572# a_19479_31679# 3.41e-20
C38376 a_21363_45546# a_3357_43084# 0.061421f
C38377 a_16409_43396# a_3483_46348# 3.88e-19
C38378 a_16243_43396# a_4185_45028# 8.86e-21
C38379 a_13467_32519# a_20202_43084# 0.333168f
C38380 a_1755_42282# a_768_44030# 2.83e-20
C38381 a_14543_43071# a_3090_45724# 0.003291f
C38382 a_n2840_42282# a_n2442_46660# 4.03e-20
C38383 a_n4318_38216# a_n2956_39768# 0.023554f
C38384 a_5934_30871# a_n2312_39304# 5.64e-21
C38385 a_13070_42354# a_10227_46804# 7.16e-20
C38386 a_n4209_39590# SMPL_ON_P 0.007959f
C38387 a_6667_45809# a_4883_46098# 6.08e-20
C38388 a_10193_42453# a_11599_46634# 0.100544f
C38389 a_6977_45572# a_6151_47436# 9.54e-19
C38390 a_6905_45572# a_6545_47178# 1.54e-20
C38391 a_11064_45572# a_2063_45854# 0.001139f
C38392 a_5066_45546# a_8379_46155# 0.001042f
C38393 a_8062_46482# a_8049_45260# 2.78e-21
C38394 a_8016_46348# a_n443_42852# 1.96e-19
C38395 a_n3420_37440# C1_P_btm 0.001902f
C38396 a_15743_43084# a_5649_42852# 0.024346f
C38397 a_8685_43396# a_8387_43230# 0.002391f
C38398 a_3626_43646# a_18817_42826# 1.64e-20
C38399 a_2982_43646# a_19339_43156# 6.56e-21
C38400 a_16823_43084# a_17678_43396# 0.001907f
C38401 a_4235_43370# a_n2293_42282# 7.36e-20
C38402 a_16333_45814# a_16241_44734# 1.85e-20
C38403 a_6511_45714# a_6453_43914# 4.5e-21
C38404 a_15595_45028# a_11827_44484# 9.92e-21
C38405 a_3065_45002# a_n699_43396# 0.020711f
C38406 a_7276_45260# a_n2661_44458# 1.14e-20
C38407 a_n913_45002# a_13720_44458# 3.43e-23
C38408 a_2437_43646# a_n356_44636# 1.45e-20
C38409 a_2382_45260# a_5343_44458# 1e-19
C38410 a_n1736_43218# a_n443_42852# 5.95e-22
C38411 a_16795_42852# a_13259_45724# 2.94e-19
C38412 a_5193_42852# a_526_44458# 0.058324f
C38413 a_4520_42826# a_n357_42282# 0.005592f
C38414 a_3935_42891# a_n755_45592# 3.21e-22
C38415 a_17303_42282# a_19692_46634# 6.55e-21
C38416 VDAC_N w_11334_34010# 0.049022f
C38417 a_10951_45334# a_768_44030# 7.27e-21
C38418 a_6171_45002# a_5807_45002# 0.193427f
C38419 a_2437_43646# a_3699_46634# 5.21e-20
C38420 a_413_45260# a_n2293_46634# 0.497204f
C38421 a_n967_45348# a_n2438_43548# 4.25e-21
C38422 a_14797_45144# a_n881_46662# 1.1e-19
C38423 a_15685_45394# a_12861_44030# 5.1e-20
C38424 a_22609_38406# VDD 0.317066f
C38425 a_n2661_44458# a_n746_45260# 0.079054f
C38426 a_n2433_44484# a_n971_45724# 4.54e-20
C38427 a_949_44458# a_n2497_47436# 0.127971f
C38428 a_n2472_42826# a_n3674_37592# 0.00166f
C38429 a_14955_43396# a_15051_42282# 2.17e-19
C38430 a_n1076_43230# COMP_P 1.14e-20
C38431 a_12379_42858# a_14635_42282# 3.89e-21
C38432 a_743_42282# a_2903_42308# 0.010301f
C38433 a_12281_43396# a_13575_42558# 5.62e-20
C38434 a_15095_43370# a_15486_42560# 0.001728f
C38435 a_n4318_38680# a_n3674_38216# 0.023866f
C38436 a_12545_42858# a_13003_42852# 0.027606f
C38437 a_5534_30871# a_12800_43218# 1.43e-19
C38438 a_12089_42308# a_13291_42460# 1.22e-19
C38439 a_n1853_43023# a_n784_42308# 8.46e-21
C38440 a_3080_42308# a_n4209_39590# 7.41e-22
C38441 a_n4251_39616# VDD 3.95e-19
C38442 a_3422_30871# a_7754_40130# 4.49e-20
C38443 a_16327_47482# a_19787_47423# 2.23e-19
C38444 a_10227_46804# a_18143_47464# 0.112443f
C38445 a_17591_47464# a_18479_47436# 6.29e-19
C38446 a_n443_46116# a_5063_47570# 0.006259f
C38447 a_4007_47204# a_n1613_43370# 7.26e-20
C38448 a_13487_47204# a_12465_44636# 0.001864f
C38449 a_15507_47210# a_13507_46334# 1.32e-19
C38450 a_14955_47212# a_4883_46098# 1.4e-20
C38451 a_13717_47436# a_22731_47423# 0.109987f
C38452 a_n1151_42308# a_5159_47243# 2.93e-19
C38453 a_3815_47204# a_n881_46662# 0.001037f
C38454 a_2063_45854# a_11309_47204# 0.141276f
C38455 a_11963_45334# a_11750_44172# 5.86e-21
C38456 a_10157_44484# a_n2661_43922# 0.00841f
C38457 a_10334_44484# a_n2661_42834# 5.65e-20
C38458 a_20193_45348# a_20640_44752# 0.017592f
C38459 a_16979_44734# a_9313_44734# 1.28e-21
C38460 a_n2293_42834# a_2675_43914# 1.48e-20
C38461 a_9482_43914# a_10405_44172# 0.01085f
C38462 a_7499_43078# a_9885_43646# 2.67e-20
C38463 a_10193_42453# a_14358_43442# 2.71e-21
C38464 a_2711_45572# a_18525_43370# 7.09e-20
C38465 a_8975_43940# a_10617_44484# 0.025058f
C38466 a_1307_43914# a_6101_44260# 7.06e-19
C38467 a_626_44172# a_2537_44260# 4.41e-22
C38468 a_11827_44484# a_18005_44484# 3.81e-19
C38469 a_21335_42336# a_13259_45724# 5.02e-20
C38470 a_n2216_38778# a_n2956_38680# 0.001511f
C38471 a_5342_30871# RST_Z 0.048618f
C38472 a_10807_43548# a_2063_45854# 0.094631f
C38473 a_n2661_42282# a_4791_45118# 9.1e-19
C38474 a_5147_45002# a_5164_46348# 0.060833f
C38475 a_2437_43646# a_20075_46420# 1.37e-20
C38476 a_3357_43084# a_18985_46122# 2.92e-20
C38477 a_413_45260# a_9625_46129# 4.85e-21
C38478 a_5111_44636# a_5068_46348# 2.11e-19
C38479 a_8696_44636# a_10586_45546# 1.39e-19
C38480 a_13490_45394# a_13059_46348# 4.86e-19
C38481 a_n2293_43922# a_n2312_38680# 3.87e-20
C38482 a_14673_44172# a_5807_45002# 0.001217f
C38483 a_3232_43370# a_4185_45028# 0.018743f
C38484 a_19113_45348# a_3090_45724# 0.128103f
C38485 a_20567_45036# a_15227_44166# 2.08e-20
C38486 a_18184_42460# a_19466_46812# 0.006722f
C38487 a_6431_45366# a_3483_46348# 0.002186f
C38488 a_19778_44110# a_19692_46634# 1.92e-20
C38489 a_1755_42282# a_6123_31319# 0.033073f
C38490 a_5267_42460# a_4921_42308# 0.04229f
C38491 a_1606_42308# a_7963_42308# 1.34e-20
C38492 a_13467_32519# C5_N_btm 1.49e-19
C38493 a_13678_32519# C2_N_btm 0.03058f
C38494 a_22469_39537# a_22609_38406# 0.198764f
C38495 a_22459_39145# a_22717_36887# 0.011525f
C38496 a_22521_39511# a_22705_37990# 0.004065f
C38497 a_768_44030# a_11735_46660# 2.94e-21
C38498 a_12891_46348# a_11901_46660# 0.028795f
C38499 a_n2661_46634# a_10467_46802# 0.033928f
C38500 a_n1925_46634# a_7927_46660# 0.009262f
C38501 a_n743_46660# a_7577_46660# 6.2e-20
C38502 a_2959_46660# a_3055_46660# 0.013793f
C38503 a_3177_46902# a_3221_46660# 3.69e-19
C38504 a_2609_46660# a_3877_44458# 4.32e-19
C38505 a_2443_46660# a_4646_46812# 2.79e-21
C38506 a_12549_44172# a_11813_46116# 2.08e-20
C38507 a_5807_45002# a_6903_46660# 5.51e-19
C38508 a_n881_46662# a_14976_45028# 0.020069f
C38509 a_12465_44636# a_14513_46634# 0.01549f
C38510 a_16327_47482# a_20107_46660# 0.007614f
C38511 a_17591_47464# a_17829_46910# 8.36e-19
C38512 a_10227_46804# a_765_45546# 0.038035f
C38513 a_11599_46634# a_21363_46634# 5.21e-21
C38514 a_18143_47464# a_17339_46660# 6.71e-19
C38515 a_2063_45854# a_472_46348# 3.39e-19
C38516 a_n237_47217# a_2698_46116# 0.032015f
C38517 a_584_46384# a_805_46414# 0.135394f
C38518 a_n971_45724# a_3147_46376# 0.001884f
C38519 a_1239_47204# a_1138_42852# 9.6e-21
C38520 a_4007_47204# a_n2293_46098# 1.9e-21
C38521 a_n1151_42308# a_n1423_46090# 0.009064f
C38522 a_1209_47178# a_1823_45246# 4.52e-19
C38523 a_n2109_47186# a_5164_46348# 0.603312f
C38524 a_949_44458# a_1568_43370# 6.56e-19
C38525 a_18374_44850# a_18533_43940# 8.18e-21
C38526 a_453_43940# a_2127_44172# 0.007699f
C38527 a_1467_44172# a_895_43940# 0.017277f
C38528 a_1414_42308# a_2479_44172# 0.110442f
C38529 a_n699_43396# a_458_43396# 0.064001f
C38530 a_742_44458# a_1756_43548# 0.152145f
C38531 a_11967_42832# a_10949_43914# 2.29e-20
C38532 a_10193_42453# a_20836_43172# 0.009033f
C38533 a_6109_44484# a_6671_43940# 0.008633f
C38534 a_18989_43940# a_19319_43548# 3.72e-20
C38535 a_n2661_43370# a_10341_43396# 2.26e-20
C38536 a_13490_45067# a_9145_43396# 5.1e-21
C38537 a_n913_45002# a_5111_42852# 2.26e-19
C38538 a_n1059_45260# a_5755_42852# 0.005901f
C38539 a_22521_40599# VDD 0.804442f
C38540 a_6298_44484# VDD 1.21616f
C38541 a_7174_31319# C3_P_btm 3.5e-20
C38542 a_n3565_39590# a_n1838_35608# 2.37e-19
C38543 a_n4209_39590# a_n1532_35090# 1.12e-19
C38544 a_20107_42308# RST_Z 4.07e-20
C38545 a_3422_30871# a_11415_45002# 0.002932f
C38546 a_15493_43940# a_6755_46942# 0.001348f
C38547 a_n1917_43396# a_n2438_43548# 2.8e-19
C38548 a_n2012_43396# a_n2293_46634# 1.17e-21
C38549 a_n2661_43370# a_n356_45724# 7.45e-20
C38550 a_4223_44672# a_8049_45260# 1.63e-20
C38551 a_16237_45028# a_16375_45002# 0.035582f
C38552 a_17801_45144# a_13259_45724# 3.04e-19
C38553 a_n2661_42834# a_9290_44172# 0.046011f
C38554 a_7112_43396# a_n1613_43370# 0.245085f
C38555 a_16977_43638# a_12861_44030# 5.41e-21
C38556 a_4361_42308# a_584_46384# 6.47e-21
C38557 a_n1076_43230# a_n2497_47436# 2.48e-20
C38558 a_n1853_43023# SMPL_ON_P 8.05e-21
C38559 a_n3565_39590# a_n3690_39392# 7.97e-20
C38560 a_n3690_39616# a_n3565_39304# 7.97e-20
C38561 a_n2946_39866# a_n4209_39304# 5.32e-20
C38562 a_n3420_39616# a_n4334_39392# 0.014828f
C38563 a_n4209_39590# a_n2946_39072# 5.32e-20
C38564 a_n4064_40160# a_n3607_39392# 5.58e-20
C38565 a_n2472_46634# VDD 0.287589f
C38566 a_5932_42308# C7_N_btm 0.003981f
C38567 a_6123_31319# C2_N_btm 0.01106f
C38568 a_5934_30871# C0_N_btm 0.015126f
C38569 a_19466_46812# a_12741_44636# 0.043645f
C38570 a_17339_46660# a_765_45546# 0.244447f
C38571 a_n2661_46634# a_8034_45724# 1.89e-20
C38572 a_21588_30879# a_8049_45260# 7.12e-20
C38573 a_2107_46812# a_2981_46116# 0.002293f
C38574 a_n2661_46098# a_n1379_46482# 0.002086f
C38575 a_9863_46634# a_9625_46129# 0.001647f
C38576 a_10467_46802# a_8199_44636# 3.56e-19
C38577 a_6755_46942# a_6419_46155# 7.31e-19
C38578 a_n2312_39304# a_n2293_45546# 6.75e-19
C38579 a_12465_44636# a_n357_42282# 1.28e-20
C38580 a_18287_44626# a_18083_42858# 4.69e-21
C38581 a_18248_44752# a_17333_42852# 4.89e-19
C38582 a_20679_44626# a_4190_30871# 8.87e-19
C38583 a_20159_44458# a_20556_43646# 7.51e-20
C38584 a_5891_43370# a_10083_42826# 0.016347f
C38585 a_15682_43940# a_3626_43646# 5.73e-21
C38586 a_20835_44721# a_21259_43561# 7.23e-22
C38587 a_n2661_43922# a_685_42968# 1.03e-21
C38588 a_n2661_42834# a_791_42968# 1.41e-20
C38589 a_n356_44636# a_14543_43071# 1.16e-21
C38590 a_n2293_42834# a_n1736_42282# 0.002516f
C38591 a_n699_43396# a_2987_42968# 8.45e-20
C38592 a_1307_43914# a_5379_42460# 2.61e-20
C38593 a_20512_43084# a_18783_43370# 8.84e-20
C38594 a_5111_44636# a_9885_42558# 3.55e-21
C38595 en_comp a_15803_42450# 8.24e-20
C38596 a_10555_44260# VDD 0.004772f
C38597 a_16680_45572# a_18479_45785# 5.64e-19
C38598 a_15861_45028# a_16147_45260# 0.146279f
C38599 a_8696_44636# a_18175_45572# 3.95e-21
C38600 a_17478_45572# a_17786_45822# 0.017351f
C38601 a_16855_45546# a_18341_45572# 7.24e-20
C38602 a_6511_45714# a_6171_45002# 0.012882f
C38603 a_6472_45840# a_6431_45366# 4.9e-19
C38604 a_6194_45824# a_5205_44484# 1.42e-21
C38605 a_2711_45572# a_8191_45002# 0.003439f
C38606 a_10193_42453# en_comp 1.87e-19
C38607 a_22400_42852# a_13507_46334# 0.235269f
C38608 a_5742_30871# w_11334_34010# 1.73e-19
C38609 a_22469_40625# a_22821_38993# 0.002743f
C38610 VDAC_P CAL_P 6.16e-21
C38611 a_22521_40599# a_22469_39537# 0.380006f
C38612 a_n4209_37414# C10_P_btm 2.25e-20
C38613 a_15493_43940# a_8049_45260# 4.49e-20
C38614 a_1443_43940# a_526_44458# 0.001014f
C38615 a_1414_42308# a_n443_42852# 0.193113f
C38616 a_17486_43762# a_15227_44166# 1.43e-19
C38617 a_3626_43646# a_1823_45246# 0.033967f
C38618 a_4905_42826# a_4185_45028# 0.039846f
C38619 a_19721_31679# a_19864_35138# 1.22e-21
C38620 a_5937_45572# VDD 2.20055f
C38621 a_5263_45724# a_n237_47217# 1.16e-19
C38622 a_20820_30879# a_20692_30879# 8.973741f
C38623 a_12741_44636# a_20205_31679# 0.003338f
C38624 a_8199_44636# a_8034_45724# 0.127067f
C38625 a_21137_46414# a_6945_45028# 0.042885f
C38626 a_19900_46494# a_10809_44734# 3.7e-20
C38627 a_n809_44244# a_n961_42308# 2.8e-19
C38628 a_6293_42852# a_743_42282# 1.73e-19
C38629 a_10341_43396# a_15681_43442# 0.008134f
C38630 a_8685_43396# a_15743_43084# 1.67e-19
C38631 a_n97_42460# a_421_43172# 0.003376f
C38632 a_n1761_44111# a_n327_42558# 0.004022f
C38633 a_n356_44636# a_19511_42282# 5.6e-21
C38634 a_n881_46662# DATA[0] 0.003238f
C38635 a_n1613_43370# DATA[1] 7.06e-20
C38636 a_22612_30879# a_22609_38406# 8.17e-21
C38637 a_n967_43230# VDD 2.82e-20
C38638 a_14797_45144# a_1307_43914# 6.81e-21
C38639 a_14537_43396# a_16751_45260# 0.011362f
C38640 a_8696_44636# a_10440_44484# 0.00348f
C38641 a_7499_43078# a_n2661_43922# 0.087751f
C38642 a_11823_42460# a_9313_44734# 0.0934f
C38643 a_2711_45572# a_16241_44484# 0.001104f
C38644 a_n143_45144# a_n2661_43370# 0.002979f
C38645 a_5111_44636# a_5093_45028# 0.021262f
C38646 a_4927_45028# a_5009_45028# 0.096132f
C38647 a_5147_45002# a_5837_45028# 0.001063f
C38648 a_21513_45002# a_21005_45260# 3.98e-19
C38649 a_3357_43084# a_19778_44110# 1.15e-19
C38650 a_8483_43230# a_3483_46348# 1.15e-21
C38651 a_n2302_39866# a_n2442_46660# 0.161638f
C38652 a_4921_42308# a_3090_45724# 0.001886f
C38653 a_n3420_39616# a_n2312_38680# 1.39e-19
C38654 a_16409_43396# a_n357_42282# 1.19e-20
C38655 a_7227_42852# a_526_44458# 0.062474f
C38656 a_12281_43396# a_n443_42852# 0.030395f
C38657 a_17595_43084# a_17715_44484# 7.53e-21
C38658 a_n2661_45010# a_n2312_39304# 1.13e-20
C38659 a_413_45260# a_18597_46090# 1.48e-19
C38660 a_14537_43396# a_4915_47217# 5.76e-19
C38661 a_5837_45028# a_n2109_47186# 0.001685f
C38662 a_2304_45348# a_2063_45854# 0.001671f
C38663 a_16147_45260# a_19321_45002# 1.91e-21
C38664 a_8696_44636# a_n743_46660# 0.032893f
C38665 a_18479_45785# a_13747_46662# 0.020713f
C38666 a_18909_45814# a_5807_45002# 0.001758f
C38667 a_18341_45572# a_13661_43548# 0.037017f
C38668 a_21076_30879# EN_OFFSET_CAL 0.2809f
C38669 a_13113_42826# a_12895_43230# 0.209641f
C38670 a_12379_42858# a_14543_43071# 5.72e-21
C38671 a_12545_42858# a_13635_43156# 0.041762f
C38672 a_6031_43396# a_6171_42473# 2.49e-21
C38673 a_2813_43396# a_2903_42308# 6.21e-21
C38674 a_3626_43646# a_5934_30871# 0.192998f
C38675 a_n97_42460# a_13657_42558# 0.011259f
C38676 a_15743_43084# a_15953_42852# 0.006469f
C38677 a_2982_43646# a_3905_42308# 4.18e-19
C38678 a_20820_30879# VIN_N 0.049556f
C38679 VDAC_P CAL_N 2.76e-19
C38680 a_3422_30871# C6_N_btm 2.2e-19
C38681 a_13575_42558# VDD 0.182133f
C38682 a_n237_47217# a_n1435_47204# 0.001134f
C38683 a_3785_47178# a_4915_47217# 0.006427f
C38684 a_n1151_42308# a_5815_47464# 0.001311f
C38685 a_4007_47204# a_4791_45118# 0.002181f
C38686 a_3815_47204# a_n443_46116# 9.13e-19
C38687 a_4743_44484# a_5518_44484# 1.16e-19
C38688 a_4223_44672# a_8103_44636# 1.47e-19
C38689 a_n2661_43370# a_n2293_43922# 0.001105f
C38690 a_2274_45254# a_2127_44172# 5.57e-20
C38691 a_2680_45002# a_1414_42308# 6.45e-20
C38692 a_413_45260# a_2675_43914# 0.048283f
C38693 a_n913_45002# a_7542_44172# 9.32e-22
C38694 a_n2293_45010# a_n1644_44306# 3.56e-19
C38695 a_327_44734# a_895_43940# 3.3e-19
C38696 a_n2017_45002# a_n4318_39768# 9.4e-20
C38697 a_564_42282# a_n357_42282# 0.026735f
C38698 a_961_42354# a_n863_45724# 0.038222f
C38699 a_n3674_37592# a_n755_45592# 0.063692f
C38700 a_17364_32525# EN_VIN_BSTR_N 0.959329f
C38701 a_743_42282# RST_Z 2.55e-19
C38702 a_22521_40599# a_22612_30879# 9.6e-20
C38703 a_22469_40625# a_21588_30879# 6.62e-20
C38704 a_14180_45002# a_15227_44166# 2.28e-19
C38705 a_2779_44458# a_n2293_46634# 0.004655f
C38706 a_18287_44626# a_12549_44172# 0.006594f
C38707 a_19963_31679# a_11415_45002# 0.033926f
C38708 a_1307_43914# a_14976_45028# 4.47e-20
C38709 a_n1917_44484# a_n2438_43548# 2.8e-19
C38710 a_12607_44458# a_5807_45002# 5.72e-21
C38711 a_2437_43646# a_21076_30879# 3e-20
C38712 a_9049_44484# a_5066_45546# 3.93e-19
C38713 a_413_45260# a_19123_46287# 4.85e-21
C38714 a_11778_45572# a_2324_44458# 8.28e-19
C38715 a_15433_44458# a_10227_46804# 0.001023f
C38716 a_17061_44734# a_12861_44030# 1.88e-19
C38717 a_175_44278# a_n2497_47436# 0.05097f
C38718 a_15567_42826# a_4958_30871# 7.19e-21
C38719 a_n2472_42282# a_n4318_38216# 0.157105f
C38720 a_n2840_42282# a_n3674_38216# 0.03703f
C38721 a_n2840_46634# a_n2661_46634# 0.180867f
C38722 a_n881_46662# a_3524_46660# 2.99e-19
C38723 a_n1613_43370# a_2864_46660# 0.014165f
C38724 a_4883_46098# a_5257_43370# 0.026597f
C38725 a_2063_45854# a_12156_46660# 2.28e-19
C38726 a_4915_47217# a_3090_45724# 2.35e-20
C38727 a_6151_47436# a_13607_46688# 2.73e-20
C38728 a_10227_46804# a_10623_46897# 0.180903f
C38729 a_11967_42832# a_3422_30871# 0.139082f
C38730 a_n2661_43922# a_3600_43914# 8.69e-19
C38731 a_n2661_42834# a_3905_42865# 0.018962f
C38732 a_n2661_43370# a_n97_42460# 6.42e-21
C38733 a_n2293_42834# a_1209_43370# 0.001969f
C38734 a_1307_43914# a_7287_43370# 1.2e-19
C38735 a_20640_44752# a_20596_44850# 1.46e-19
C38736 a_17517_44484# a_19237_31679# 0.00388f
C38737 a_10193_42453# a_22165_42308# 2.46e-21
C38738 a_n913_45002# a_16977_43638# 1.48e-21
C38739 a_n1059_45260# a_16759_43396# 1.17e-19
C38740 a_n2017_45002# a_17499_43370# 4.8e-19
C38741 en_comp a_16137_43396# 1.88e-20
C38742 a_7418_45067# VDD 0.001744f
C38743 a_5934_30871# C10_P_btm 1.89e-19
C38744 a_6123_31319# C8_P_btm 6.73e-20
C38745 a_5932_42308# C3_P_btm 0.121156f
C38746 a_20205_31679# C9_N_btm 1.91e-20
C38747 a_20692_30879# C8_N_btm 1.15e-19
C38748 a_9803_43646# a_n971_45724# 5.86e-21
C38749 a_7112_43396# a_4791_45118# 1.4e-19
C38750 a_6298_44484# a_7920_46348# 1.48e-19
C38751 a_21359_45002# a_6945_45028# 1.23e-21
C38752 a_4223_44672# a_8953_45546# 5.72e-21
C38753 a_17896_45144# a_17715_44484# 3.62e-20
C38754 a_1667_45002# a_n443_42852# 3.6e-19
C38755 a_413_45260# a_2277_45546# 1.14e-20
C38756 a_n2293_42834# a_8049_45260# 0.224469f
C38757 a_14485_44260# a_13661_43548# 4.85e-19
C38758 a_3737_43940# a_768_44030# 0.038628f
C38759 a_20159_44458# a_19692_46634# 0.001725f
C38760 a_5663_43940# a_5257_43370# 0.014098f
C38761 a_14021_43940# a_13747_46662# 1.12e-19
C38762 a_20362_44736# a_19466_46812# 3.02e-19
C38763 a_20679_44626# a_15227_44166# 1.44e-21
C38764 a_18479_47436# VDD 1.47669f
C38765 a_17303_42282# a_20107_42308# 3.68e-19
C38766 a_18727_42674# a_19511_42282# 5.06e-19
C38767 a_n2661_46098# a_n1076_46494# 0.037593f
C38768 a_1983_46706# a_2202_46116# 0.001054f
C38769 a_2107_46812# a_167_45260# 0.012514f
C38770 a_10467_46802# a_765_45546# 0.003784f
C38771 a_11901_46660# a_12359_47026# 0.034619f
C38772 a_6755_46942# a_14226_46660# 0.001921f
C38773 a_768_44030# a_2324_44458# 0.047942f
C38774 a_n743_46660# a_4704_46090# 0.011859f
C38775 a_12549_44172# a_15682_46116# 6.67e-19
C38776 a_5807_45002# a_10903_43370# 0.002924f
C38777 a_n2661_46634# a_8016_46348# 1.16e-19
C38778 a_n1925_46634# a_5164_46348# 2.7e-19
C38779 a_n746_45260# a_n1099_45572# 0.015931f
C38780 a_n815_47178# a_n755_45592# 2.36e-20
C38781 a_n237_47217# a_380_45546# 6.95e-20
C38782 a_n971_45724# a_310_45028# 4.56e-21
C38783 a_n2293_42834# a_3059_42968# 1.04e-19
C38784 a_18989_43940# a_19095_43396# 2.42e-19
C38785 a_2998_44172# a_n97_42460# 4.27e-19
C38786 a_20269_44172# a_14021_43940# 5.52e-20
C38787 a_1115_44172# a_1209_43370# 1.17e-19
C38788 a_9313_44734# a_18429_43548# 3.66e-20
C38789 a_8333_44056# a_8487_44056# 0.008678f
C38790 a_14537_43396# a_13291_42460# 2.95e-20
C38791 a_n967_45348# a_196_42282# 3.02e-20
C38792 a_n1059_45260# a_1067_42314# 0.006623f
C38793 a_n2293_45010# a_961_42354# 2.42e-20
C38794 a_n2017_45002# a_1576_42282# 0.008099f
C38795 a_n2810_45028# a_n3674_37592# 0.025732f
C38796 a_n913_45002# a_n1630_35242# 3.81e-19
C38797 en_comp a_n784_42308# 0.025103f
C38798 a_2479_44172# VDD 0.431428f
C38799 a_11823_42460# a_15037_45618# 0.099829f
C38800 a_10193_42453# a_16855_45546# 3.49e-20
C38801 a_10907_45822# a_11280_45822# 0.001255f
C38802 C6_N_btm VREF_GND 0.836236f
C38803 C5_N_btm VCM 0.719982f
C38804 C7_N_btm VREF 1.818f
C38805 C8_N_btm VIN_N 0.907642f
C38806 a_3052_44056# a_1823_45246# 2.45e-20
C38807 a_19319_43548# a_20202_43084# 2.44e-19
C38808 a_15037_44260# a_3483_46348# 6.29e-19
C38809 a_8387_43230# a_768_44030# 1.54e-20
C38810 a_n3674_39304# a_n2442_46660# 0.024039f
C38811 a_n1853_43023# a_n2438_43548# 0.001525f
C38812 a_6452_43396# a_3090_45724# 0.001752f
C38813 a_3905_42865# a_5066_45546# 0.001745f
C38814 a_3422_30871# a_13259_45724# 0.587088f
C38815 a_14112_44734# a_n443_42852# 2.65e-20
C38816 a_13483_43940# a_2324_44458# 3.39e-21
C38817 a_22223_42860# a_13507_46334# 0.049534f
C38818 a_17829_46910# VDD 0.37446f
C38819 a_21076_30879# a_22959_46124# 5.19e-19
C38820 a_765_45546# a_8034_45724# 1.01e-21
C38821 a_19466_46812# a_16375_45002# 5.87e-21
C38822 a_15227_44166# a_19431_46494# 0.001203f
C38823 a_3483_46348# a_12005_46116# 4.4e-21
C38824 a_21297_46660# a_10809_44734# 2.09e-19
C38825 a_7920_46348# a_5937_45572# 4.23e-21
C38826 a_8016_46348# a_8199_44636# 0.33718f
C38827 a_7174_31319# a_7754_40130# 0.005009f
C38828 a_n4315_30879# a_n3420_37984# 0.034791f
C38829 a_10949_43914# a_10518_42984# 2.24e-21
C38830 a_6765_43638# a_6655_43762# 0.097745f
C38831 a_10729_43914# a_10835_43094# 4.2e-21
C38832 a_10405_44172# a_10796_42968# 1.23e-20
C38833 a_18184_42460# a_13258_32519# 0.038977f
C38834 a_n2661_42834# a_n961_42308# 1.03e-20
C38835 a_n2293_43922# COMP_P 0.151768f
C38836 a_n356_44636# a_4921_42308# 8e-19
C38837 a_18494_42460# a_19647_42308# 0.030348f
C38838 a_6547_43396# a_6452_43396# 0.049827f
C38839 a_11967_42832# a_18504_43218# 0.015494f
C38840 a_3905_42865# a_n2293_42282# 4.89e-19
C38841 a_19741_43940# a_15743_43084# 4.79e-20
C38842 a_4700_47436# DATA[2] 0.001637f
C38843 a_n443_46116# DATA[0] 4.31e-19
C38844 a_n1151_42308# CLK 0.022274f
C38845 a_6151_47436# RST_Z 0.010195f
C38846 a_19479_31679# C9_N_btm 1.91e-20
C38847 a_19963_31679# C6_N_btm 1.26e-20
C38848 a_11525_45546# a_n2661_44458# 1.89e-19
C38849 a_2711_45572# a_16979_44734# 6.79e-20
C38850 a_2274_45254# a_2382_45260# 0.130215f
C38851 a_413_45260# a_3429_45260# 4.84e-19
C38852 a_n913_45002# a_5205_44484# 4.56e-21
C38853 a_766_43646# a_n755_45592# 3.04e-19
C38854 a_2982_43646# a_n863_45724# 2.39e-20
C38855 a_n1557_42282# a_n357_42282# 0.384406f
C38856 a_5742_30871# a_n2442_46660# 8.02e-21
C38857 a_15803_42450# a_13661_43548# 3.06e-22
C38858 a_13291_42460# a_3090_45724# 0.002769f
C38859 a_3422_30871# C4_P_btm 1.36e-19
C38860 a_19237_31679# EN_VIN_BSTR_N 0.069167f
C38861 a_n443_42852# VDD 3.69394f
C38862 a_13527_45546# a_768_44030# 1.49e-20
C38863 a_8746_45002# a_5807_45002# 7.32e-20
C38864 a_13904_45546# a_12549_44172# 5.84e-19
C38865 a_13249_42308# a_12891_46348# 0.166217f
C38866 a_10193_42453# a_13661_43548# 0.211481f
C38867 a_7227_45028# a_n743_46660# 0.001306f
C38868 a_2211_45572# a_n2293_46634# 3.32e-19
C38869 a_15765_45572# a_12465_44636# 2.53e-21
C38870 a_18479_45785# a_11599_46634# 0.028968f
C38871 a_16211_45572# a_16327_47482# 1.79e-19
C38872 a_19431_45546# a_12861_44030# 1.85e-20
C38873 a_n913_45002# a_n971_45724# 0.101346f
C38874 a_2437_43646# a_3381_47502# 0.004114f
C38875 a_n1059_45260# a_n746_45260# 0.138039f
C38876 a_n143_45144# a_n2497_47436# 1.83e-21
C38877 en_comp SMPL_ON_P 0.034192f
C38878 a_18783_43370# a_18249_42858# 3.47e-20
C38879 a_15743_43084# a_17333_42852# 2.59e-20
C38880 a_4361_42308# a_8952_43230# 1.43e-20
C38881 a_743_42282# a_10991_42826# 1.68e-19
C38882 a_5649_42852# a_8605_42826# 9.36e-21
C38883 a_19268_43646# a_18083_42858# 1.18e-19
C38884 a_15493_43396# a_15890_42674# 1.56e-21
C38885 a_n4318_39304# a_n1630_35242# 2.74e-20
C38886 a_n97_42460# COMP_P 7.27e-21
C38887 a_5829_43940# a_5932_42308# 1.65e-20
C38888 a_15231_43396# a_5342_30871# 2.63e-19
C38889 a_8685_43396# a_9061_43230# 7.37e-20
C38890 a_19466_46812# RST_Z 2.04e-20
C38891 a_15227_44166# SINGLE_ENDED 3.5e-21
C38892 a_19333_46634# START 3.38e-20
C38893 a_n3420_37984# a_n3420_37440# 0.132162f
C38894 a_n4064_37984# a_n3565_37414# 0.029309f
C38895 VDAC_Pi a_3754_38802# 0.00191f
C38896 a_n2104_42282# VDD 0.280329f
C38897 a_18184_42460# a_20193_45348# 0.074414f
C38898 a_21359_45002# a_11827_44484# 0.005947f
C38899 a_n2661_43370# a_742_44458# 2.53e-19
C38900 a_n2293_42834# a_8103_44636# 0.006106f
C38901 a_10193_42453# a_19862_44208# 0.099944f
C38902 a_17719_45144# a_17896_45144# 0.004187f
C38903 a_16922_45042# a_18545_45144# 0.001431f
C38904 a_18494_42460# a_11691_44458# 1.03e-19
C38905 a_13249_42308# a_11750_44172# 3.55e-20
C38906 a_n1059_45260# a_17517_44484# 1.46e-20
C38907 a_5147_45002# a_n2661_42834# 0.060392f
C38908 a_4558_45348# a_n2661_43922# 6.4e-20
C38909 a_20623_45572# a_20980_44850# 1.83e-20
C38910 a_15803_42450# a_4185_45028# 2.86e-19
C38911 a_21335_42336# a_20202_43084# 0.227943f
C38912 a_8483_43230# a_n357_42282# 7.88e-19
C38913 a_8292_43218# a_n755_45592# 0.010247f
C38914 a_18504_43218# a_13259_45724# 9.31e-20
C38915 a_1067_42314# a_n1925_42282# 5.5e-20
C38916 a_1576_42282# a_526_44458# 2.98e-20
C38917 a_873_42968# a_n443_42852# 5.2e-19
C38918 a_9885_42558# a_9290_44172# 0.021204f
C38919 a_5742_30871# a_8953_45546# 1.11e-19
C38920 a_13076_44458# a_12861_44030# 0.01178f
C38921 a_n2293_43922# a_n2497_47436# 9.38e-20
C38922 a_2711_45572# a_14275_46494# 1.13e-20
C38923 a_6812_45938# a_6419_46155# 7.41e-19
C38924 a_21363_45546# a_19466_46812# 9.08e-21
C38925 a_n2017_45002# a_8270_45546# 4.47e-21
C38926 a_3232_43370# a_5257_43370# 0.022872f
C38927 a_413_45260# a_6755_46942# 6.02e-20
C38928 a_3357_43084# a_12816_46660# 5.53e-21
C38929 a_2437_43646# a_15009_46634# 7.72e-21
C38930 a_20623_45572# a_19692_46634# 5.14e-19
C38931 a_14403_45348# a_5807_45002# 0.002634f
C38932 a_16147_45260# a_13059_46348# 1.3e-19
C38933 a_17023_45118# a_12549_44172# 5.36e-21
C38934 a_10193_42453# a_4185_45028# 3.16135f
C38935 a_10490_45724# a_3483_46348# 0.207668f
C38936 a_4361_42308# a_15521_42308# 1.42e-19
C38937 a_8037_42858# a_5934_30871# 7.18e-19
C38938 a_n2293_42282# a_n961_42308# 4.89e-19
C38939 a_743_42282# a_17303_42282# 0.034786f
C38940 a_4190_30871# a_18057_42282# 0.02374f
C38941 a_20205_31679# RST_Z 0.049474f
C38942 a_4883_46098# a_5807_45002# 1.76125f
C38943 a_13507_46334# a_13747_46662# 0.049663f
C38944 a_20990_47178# a_19321_45002# 1.58e-19
C38945 a_20894_47436# a_19594_46812# 7.48e-20
C38946 a_18597_46090# a_20916_46384# 6.92e-19
C38947 a_15507_47210# a_n743_46660# 0.003069f
C38948 a_n1435_47204# a_1123_46634# 6.22e-20
C38949 a_n1741_47186# a_7715_46873# 2.98e-19
C38950 a_2063_45854# a_4955_46873# 0.002567f
C38951 a_n443_46116# a_3524_46660# 0.049574f
C38952 a_2905_45572# a_3877_44458# 6.4e-20
C38953 a_3160_47472# a_3221_46660# 8.54e-19
C38954 a_13777_45326# a_13565_43940# 1.03e-20
C38955 a_n2840_44458# a_n4318_39768# 0.007737f
C38956 a_2779_44458# a_2675_43914# 1.27e-19
C38957 a_13556_45296# a_15037_43940# 0.001578f
C38958 a_n699_43396# a_2479_44172# 0.063139f
C38959 a_742_44458# a_2998_44172# 1.08e-19
C38960 a_13249_42308# a_4361_42308# 0.009442f
C38961 a_n2661_43922# a_12189_44484# 1.22e-19
C38962 a_n2661_42834# a_12553_44484# 4.92e-20
C38963 a_1307_43914# a_9420_43940# 9.31e-19
C38964 a_327_44734# a_458_43396# 1.92e-21
C38965 a_4574_45260# a_n97_42460# 9.85e-22
C38966 a_3357_43084# a_6031_43396# 0.001792f
C38967 en_comp a_3080_42308# 1.28517f
C38968 a_n4209_38502# a_n2956_38216# 0.023653f
C38969 a_2680_45002# VDD 0.145087f
C38970 a_20193_45348# a_12741_44636# 0.012699f
C38971 a_13720_44458# a_14035_46660# 7.64e-21
C38972 a_5663_43940# a_5807_45002# 2.36e-20
C38973 a_n1899_43946# a_n2438_43548# 8.61e-19
C38974 a_413_45260# a_8049_45260# 0.140877f
C38975 a_5147_45002# a_5066_45546# 5.3e-19
C38976 a_5111_44636# a_5431_46482# 6.74e-20
C38977 a_n2661_43370# a_5204_45822# 4.54e-21
C38978 a_8488_45348# a_8199_44636# 0.001482f
C38979 a_n2293_42834# a_8953_45546# 4.91e-20
C38980 a_17973_43940# a_11453_44696# 1.73e-21
C38981 a_n97_42460# a_n2497_47436# 0.026966f
C38982 a_n3674_37592# a_n2302_40160# 6.29e-20
C38983 a_5534_30871# C10_N_btm 1.08e-19
C38984 a_5342_30871# C8_N_btm 0.093874f
C38985 C4_P_btm VREF_GND 0.671882f
C38986 C5_P_btm VCM 0.719982f
C38987 C3_P_btm VREF 0.984942f
C38988 a_19594_46812# a_20411_46873# 1.02e-20
C38989 a_10428_46928# a_10554_47026# 0.181217f
C38990 a_9863_46634# a_6755_46942# 0.014818f
C38991 a_7411_46660# a_8035_47026# 9.73e-19
C38992 a_7715_46873# a_7832_46660# 0.157972f
C38993 a_10467_46802# a_10623_46897# 0.107482f
C38994 a_10150_46912# a_10249_46116# 0.066949f
C38995 a_5257_43370# a_6682_46660# 1.27e-19
C38996 a_19321_45002# a_20273_46660# 0.001516f
C38997 a_4883_46098# a_3699_46348# 2.14e-19
C38998 a_n971_45724# a_3873_46454# 6.84e-19
C38999 a_n2109_47186# a_5066_45546# 0.02651f
C39000 a_n237_47217# a_526_44458# 0.198088f
C39001 a_12861_44030# a_12594_46348# 0.43362f
C39002 a_18494_42460# a_4190_30871# 0.242908f
C39003 a_9838_44484# a_9885_43646# 4.23e-22
C39004 a_13720_44458# a_9145_43396# 6.13e-21
C39005 a_n2661_43922# a_1756_43548# 5.14e-21
C39006 a_n2661_42834# a_4093_43548# 1.69e-19
C39007 a_9313_44734# a_2982_43646# 0.027994f
C39008 a_9482_43914# a_5342_30871# 5.46e-21
C39009 a_10193_42453# a_9803_42558# 0.20198f
C39010 a_18184_42460# a_20301_43646# 6.85e-19
C39011 a_7499_43078# a_10545_42558# 0.003046f
C39012 a_11827_44484# a_16823_43084# 4.84e-20
C39013 a_n2293_42834# a_n722_43218# 2.66e-19
C39014 a_n1059_45260# a_4149_42891# 4.67e-19
C39015 a_15146_44811# VDD 6.34e-20
C39016 a_n3420_38528# VCM 0.00888f
C39017 a_n4064_38528# VREF 2.95e-20
C39018 a_2711_45572# a_11823_42460# 0.065343f
C39019 a_14209_32519# SMPL_ON_N 0.02932f
C39020 a_19279_43940# a_6945_45028# 1.94e-21
C39021 a_n699_43396# a_n443_42852# 0.333516f
C39022 a_10765_43646# a_n2293_46634# 0.001573f
C39023 a_13565_44260# a_13059_46348# 8.69e-19
C39024 a_11173_43940# a_3090_45724# 1.22e-19
C39025 a_16137_43396# a_13661_43548# 2.21e-19
C39026 a_19268_43646# a_12549_44172# 3.27e-20
C39027 a_4905_42826# a_5257_43370# 0.254437f
C39028 a_6101_44260# a_n2293_46098# 1.56e-19
C39029 a_10729_43914# a_11415_45002# 1.25e-20
C39030 a_19479_31679# RST_Z 0.049574f
C39031 a_2437_43646# SINGLE_ENDED 0.117817f
C39032 a_10554_47026# VDD 0.205847f
C39033 a_7174_31319# C6_N_btm 2.51e-19
C39034 a_n2840_46090# a_n2472_46090# 7.52e-19
C39035 a_383_46660# a_n1099_45572# 9.12e-21
C39036 a_n2293_46634# a_n23_45546# 2.45e-19
C39037 a_n743_46660# a_2957_45546# 2.2e-20
C39038 a_n2438_43548# a_1848_45724# 1.12e-20
C39039 a_171_46873# a_n755_45592# 1.47e-22
C39040 a_9863_46634# a_8049_45260# 1.3e-20
C39041 a_33_46660# a_n357_42282# 9.6e-20
C39042 a_n133_46660# a_997_45618# 3.7e-20
C39043 a_2107_46812# a_n863_45724# 3.26e-20
C39044 a_8270_45546# a_526_44458# 0.007312f
C39045 a_15227_44166# a_19335_46494# 0.024137f
C39046 a_14035_46660# a_13351_46090# 1.44e-19
C39047 a_19333_46634# a_19553_46090# 0.001209f
C39048 a_765_45546# a_8016_46348# 6.75e-20
C39049 a_19692_46634# a_18819_46122# 2.56e-19
C39050 a_19466_46812# a_18985_46122# 0.033782f
C39051 a_13885_46660# a_13759_46122# 0.002423f
C39052 a_15368_46634# a_6945_45028# 3.82e-19
C39053 a_3090_45724# a_10809_44734# 0.002539f
C39054 a_13059_46348# a_9290_44172# 2.64e-19
C39055 a_6123_31319# a_2113_38308# 7.39e-20
C39056 a_n1630_35242# a_n2946_37690# 1.09e-19
C39057 a_1606_42308# a_7754_38470# 1.54e-19
C39058 a_n97_42460# a_1568_43370# 0.074153f
C39059 a_14021_43940# a_14358_43442# 0.007211f
C39060 a_18079_43940# a_17499_43370# 0.001409f
C39061 a_15493_43396# a_16547_43609# 0.022221f
C39062 a_20974_43370# a_2982_43646# 0.051776f
C39063 a_11967_42832# a_16414_43172# 0.058563f
C39064 a_17517_44484# a_19987_42826# 6.08e-21
C39065 a_n2433_43396# a_n1557_42282# 2.44e-21
C39066 a_n356_44636# a_13291_42460# 1.18e-19
C39067 a_14539_43914# a_17665_42852# 0.003264f
C39068 a_n2810_45028# a_n2302_39072# 4.97e-19
C39069 a_n2956_37592# a_n4064_39072# 0.010695f
C39070 a_n229_43646# VDD 0.278436f
C39071 a_20273_45572# a_19963_31679# 0.001592f
C39072 a_2711_45572# a_16321_45348# 7.82e-19
C39073 a_20528_45572# a_2437_43646# 8.27e-22
C39074 a_21188_45572# a_22223_45572# 9.49e-20
C39075 a_20623_45572# a_3357_43084# 0.041244f
C39076 a_8696_44636# a_5111_44636# 3.25e-20
C39077 a_16333_45814# a_6171_45002# 3.41e-19
C39078 a_21487_43396# a_11415_45002# 1.71e-21
C39079 a_16137_43396# a_4185_45028# 1.37e-19
C39080 a_16547_43609# a_3483_46348# 5.46e-20
C39081 a_1606_42308# a_768_44030# 0.00182f
C39082 a_13460_43230# a_3090_45724# 0.004635f
C39083 a_n2472_42282# a_n2956_39768# 3.63e-20
C39084 a_1987_43646# a_526_44458# 3.41e-20
C39085 a_13667_43396# a_10903_43370# 7.81e-20
C39086 a_5934_30871# a_n2312_40392# 8.24e-21
C39087 a_9223_42460# a_4883_46098# 2.45e-19
C39088 a_6633_46155# VDD 6.34e-20
C39089 a_6511_45714# a_4883_46098# 6.24e-20
C39090 a_6905_45572# a_6151_47436# 0.003156f
C39091 a_11322_45546# a_12861_44030# 7.65e-19
C39092 a_5066_45546# a_8062_46155# 9.9e-19
C39093 a_19553_46090# a_20062_46116# 2.6e-19
C39094 a_n3565_37414# C0_P_btm 0.040442f
C39095 a_19700_43370# a_4361_42308# 7.65e-21
C39096 a_18783_43370# a_5649_42852# 1.76e-21
C39097 a_3626_43646# a_18249_42858# 4.73e-20
C39098 a_11967_42832# a_7174_31319# 5.83e-20
C39099 a_2982_43646# a_18599_43230# 2.4e-20
C39100 a_15743_43084# a_13678_32519# 0.020598f
C39101 a_16823_43084# a_17433_43396# 8.76e-19
C39102 a_4093_43548# a_n2293_42282# 5.81e-20
C39103 a_8685_43396# a_8605_42826# 0.001894f
C39104 a_1793_42852# VDD 6.57e-19
C39105 a_13777_45326# a_11691_44458# 5.49e-20
C39106 a_15415_45028# a_11827_44484# 5.8e-21
C39107 a_5205_44484# a_n2661_44458# 0.072981f
C39108 a_3065_45002# a_4223_44672# 0.001102f
C39109 a_2382_45260# a_4743_44484# 5.73e-20
C39110 a_2680_45002# a_n699_43396# 2.59e-19
C39111 a_15597_42852# a_2324_44458# 3.41e-19
C39112 a_16414_43172# a_13259_45724# 3.58e-20
C39113 a_4649_42852# a_526_44458# 0.028795f
C39114 a_3935_42891# a_n357_42282# 0.007216f
C39115 a_3681_42891# a_n755_45592# 1.63e-20
C39116 a_n784_42308# a_4185_45028# 7.16e-20
C39117 a_1221_42558# a_1138_42852# 6.61e-20
C39118 a_10775_45002# a_768_44030# 1.05e-21
C39119 en_comp a_n2438_43548# 0.915368f
C39120 a_n37_45144# a_n2293_46634# 0.006632f
C39121 a_3232_43370# a_5807_45002# 0.091049f
C39122 a_14537_43396# a_n881_46662# 1.17e-21
C39123 CAL_P VDD 22.4716f
C39124 a_n2661_44458# a_n971_45724# 0.051008f
C39125 a_742_44458# a_n2497_47436# 0.153038f
C39126 a_n1736_43218# a_n4318_38216# 3.63e-19
C39127 a_15095_43370# a_15051_42282# 0.003143f
C39128 a_14955_43396# a_14113_42308# 1.29e-21
C39129 a_n901_43156# COMP_P 8.12e-21
C39130 a_n1641_43230# a_n1329_42308# 0.004511f
C39131 a_12379_42858# a_13291_42460# 6.47e-20
C39132 a_743_42282# a_2713_42308# 0.024879f
C39133 a_12281_43396# a_13070_42354# 5.19e-19
C39134 a_17364_32525# a_n1630_35242# 1.85e-20
C39135 a_13113_42826# a_13569_43230# 4.2e-19
C39136 a_n3674_39304# a_n3674_38216# 0.023464f
C39137 a_13678_32519# a_1606_42308# 6.06e-20
C39138 a_n4318_39304# a_n3607_39392# 8.54e-20
C39139 a_1736_39587# VDD 3.14139f
C39140 a_12861_44030# a_12465_44636# 0.242761f
C39141 a_13717_47436# a_22223_47212# 0.00262f
C39142 a_14311_47204# a_4883_46098# 1.02e-20
C39143 a_11599_46634# a_13507_46334# 0.259318f
C39144 a_3815_47204# a_n1613_43370# 0.001154f
C39145 a_n443_46116# a_4842_47570# 0.001342f
C39146 a_16327_47482# a_19386_47436# 3.57e-20
C39147 a_17591_47464# a_18143_47464# 0.003298f
C39148 a_n1151_42308# a_4842_47243# 8.14e-19
C39149 a_3785_47178# a_n881_46662# 6.74e-19
C39150 a_20107_45572# a_19319_43548# 3.02e-20
C39151 a_11787_45002# a_11750_44172# 8e-19
C39152 a_10057_43914# a_10617_44484# 0.033364f
C39153 a_9838_44484# a_n2661_43922# 0.006262f
C39154 a_9482_43914# a_9672_43914# 0.122568f
C39155 a_10157_44484# a_n2661_42834# 6.22e-20
C39156 a_20193_45348# a_20362_44736# 0.013057f
C39157 a_11827_44484# a_19279_43940# 0.078733f
C39158 a_n2661_43370# a_n984_44318# 7.79e-21
C39159 a_n2293_42834# a_895_43940# 7.7e-20
C39160 a_5093_45028# a_3905_42865# 2.69e-19
C39161 a_14539_43914# a_9313_44734# 0.016028f
C39162 a_10193_42453# a_14579_43548# 5.04e-21
C39163 a_2711_45572# a_18429_43548# 2.62e-20
C39164 a_n356_44636# a_700_44734# 4.08e-19
C39165 a_626_44172# a_2253_44260# 6.94e-21
C39166 a_19778_44110# a_19789_44512# 7.63e-19
C39167 a_6171_45002# a_15493_43396# 1.54e-20
C39168 a_7174_31319# a_13259_45724# 0.033027f
C39169 a_15890_42674# a_n357_42282# 1.81e-20
C39170 a_n2860_38778# a_n2956_38680# 0.001355f
C39171 a_5342_30871# C2_P_btm 7.86e-20
C39172 a_17730_32519# SMPL_ON_N 0.029186f
C39173 a_10949_43914# a_2063_45854# 0.129837f
C39174 a_2437_43646# a_19335_46494# 5.23e-21
C39175 a_3357_43084# a_18819_46122# 3.26e-20
C39176 a_5147_45002# a_5068_46348# 5.26e-21
C39177 a_4558_45348# a_5164_46348# 0.002407f
C39178 a_413_45260# a_8953_45546# 4.56e-21
C39179 a_5691_45260# a_4185_45028# 1.6e-19
C39180 a_13940_44484# a_13661_43548# 0.002141f
C39181 a_9313_44734# a_2107_46812# 0.023852f
C39182 a_n2661_43922# a_n2312_38680# 1.97e-21
C39183 a_18494_42460# a_15227_44166# 3.03e-20
C39184 a_19778_44110# a_19466_46812# 0.116901f
C39185 a_3232_43370# a_3699_46348# 6.75e-20
C39186 a_6171_45002# a_3483_46348# 0.153232f
C39187 a_1606_42308# a_6123_31319# 1.43958f
C39188 a_3823_42558# a_4921_42308# 0.001205f
C39189 a_n784_42308# a_9803_42558# 2.06e-20
C39190 a_16877_43172# a_4958_30871# 1.48e-19
C39191 a_13467_32519# C4_N_btm 1.74e-19
C39192 a_4190_30871# C10_N_btm 0.446355f
C39193 a_13678_32519# C1_N_btm 1.26e-19
C39194 a_22821_38993# a_22609_38406# 8.2e-19
C39195 a_22469_39537# CAL_P 0.024901f
C39196 a_22521_39511# a_22609_37990# 0.333805f
C39197 a_22459_39145# a_22717_37285# 0.012249f
C39198 a_12549_44172# a_11735_46660# 1.77e-19
C39199 a_n2661_46634# a_10428_46928# 0.052586f
C39200 a_n1925_46634# a_8145_46902# 0.005351f
C39201 a_n743_46660# a_7715_46873# 0.003347f
C39202 a_2443_46660# a_3877_44458# 2.31e-19
C39203 a_3177_46902# a_3055_46660# 3.16e-19
C39204 a_12891_46348# a_11813_46116# 1.48e-19
C39205 a_5807_45002# a_6682_46660# 6.46e-19
C39206 a_2107_46812# a_5072_46660# 8.97e-19
C39207 a_11309_47204# a_11901_46660# 0.001315f
C39208 a_n881_46662# a_3090_45724# 0.107805f
C39209 a_12465_44636# a_14180_46812# 0.026945f
C39210 a_16327_47482# a_19551_46910# 1.05e-19
C39211 a_17591_47464# a_765_45546# 0.004682f
C39212 a_11599_46634# a_20623_46660# 4.44e-20
C39213 a_10227_46804# a_17339_46660# 2.73e-20
C39214 a_n971_45724# a_2804_46116# 1.43e-19
C39215 a_n237_47217# a_2521_46116# 0.039248f
C39216 a_584_46384# a_472_46348# 0.31609f
C39217 a_n1151_42308# a_n1991_46122# 0.027139f
C39218 a_1209_47178# a_1138_42852# 1.18e-20
C39219 a_1239_47204# a_1176_45822# 4.07e-21
C39220 a_3815_47204# a_n2293_46098# 2.35e-20
C39221 a_2063_45854# a_376_46348# 3.28e-20
C39222 a_n2109_47186# a_5068_46348# 1.71e-20
C39223 a_n1741_47186# a_4419_46090# 4.26e-20
C39224 a_949_44458# a_1049_43396# 0.001408f
C39225 a_18443_44721# a_18533_43940# 6.51e-20
C39226 a_1115_44172# a_895_43940# 0.029554f
C39227 a_1414_42308# a_2127_44172# 0.091064f
C39228 a_5883_43914# a_n97_42460# 5.99e-19
C39229 a_n699_43396# a_n229_43646# 0.043893f
C39230 a_742_44458# a_1568_43370# 0.525694f
C39231 a_1467_44172# a_2479_44172# 2.93e-20
C39232 a_18989_43940# a_19808_44306# 1.9e-20
C39233 a_13249_42308# a_13622_42852# 1.85e-19
C39234 a_n913_45002# a_4520_42826# 0.001583f
C39235 a_n1059_45260# a_5111_42852# 0.005242f
C39236 a_n2017_45002# a_5755_42852# 1.59e-20
C39237 CAL_N VDD 26.069302f
C39238 a_5518_44484# VDD 0.40715f
C39239 a_4958_30871# VIN_N 0.025339f
C39240 a_7174_31319# C4_P_btm 2.64e-20
C39241 a_n4209_39590# a_n1386_35608# 1.02e-19
C39242 a_13258_32519# RST_Z 0.059424f
C39243 a_14673_44172# a_3483_46348# 0.026455f
C39244 a_3422_30871# a_20202_43084# 0.527141f
C39245 a_21398_44850# a_11415_45002# 9.56e-19
C39246 a_5829_43940# a_4646_46812# 2.16e-19
C39247 a_n1699_43638# a_n2438_43548# 4.93e-19
C39248 a_5343_44458# a_8034_45724# 2.52e-21
C39249 a_n2661_43370# a_3503_45724# 3.04e-20
C39250 a_6547_43396# a_n881_46662# 1.22e-20
C39251 a_7287_43370# a_n1613_43370# 0.337957f
C39252 a_16409_43396# a_12861_44030# 9.01e-20
C39253 a_n901_43156# a_n2497_47436# 0.006149f
C39254 a_n2157_42858# SMPL_ON_P 6.32e-21
C39255 a_n3565_39590# a_n3565_39304# 0.046203f
C39256 a_n3420_39616# a_n4209_39304# 0.05141f
C39257 a_n4209_39590# a_n3420_39072# 0.034738f
C39258 a_n4064_39616# a_n3607_39616# 7.1e-19
C39259 a_n4064_40160# a_n4251_39392# 0.001069f
C39260 a_n2661_46634# VDD 2.23057f
C39261 a_5934_30871# C0_dummy_N_btm 1.48e-19
C39262 a_6123_31319# C1_N_btm 0.011005f
C39263 a_5932_42308# C6_N_btm 3.73e-19
C39264 a_20916_46384# a_8049_45260# 0.003776f
C39265 a_n2661_46098# a_n1545_46494# 0.004305f
C39266 a_n1925_46634# a_5066_45546# 0.195997f
C39267 a_5807_45002# a_11608_46482# 5.69e-19
C39268 a_2107_46812# a_1431_46436# 1.17e-19
C39269 a_10428_46928# a_8199_44636# 5.81e-19
C39270 a_n2312_39304# a_n2956_38216# 0.060648f
C39271 a_18248_44752# a_18083_42858# 1.84e-20
C39272 a_20640_44752# a_4190_30871# 5.05e-22
C39273 a_20679_44626# a_21259_43561# 9.33e-20
C39274 a_11967_42832# a_21487_43396# 1.24e-20
C39275 a_n2661_42834# a_685_42968# 1.91e-21
C39276 a_5891_43370# a_8952_43230# 0.016573f
C39277 a_9313_44734# a_7871_42858# 1.01e-19
C39278 a_17970_44736# a_17333_42852# 5.58e-21
C39279 a_14539_43914# a_18599_43230# 1.28e-19
C39280 a_n2293_42834# a_n3674_38216# 0.001875f
C39281 a_1307_43914# a_5267_42460# 9.19e-21
C39282 en_comp a_15764_42576# 5.59e-20
C39283 a_3065_45002# a_5742_30871# 1.24e-20
C39284 a_16680_45572# a_18175_45572# 4.94e-20
C39285 a_8696_44636# a_16147_45260# 0.284694f
C39286 a_16855_45546# a_18479_45785# 1.38e-20
C39287 a_16020_45572# a_16211_45572# 4.61e-19
C39288 a_6511_45714# a_3232_43370# 5.46e-20
C39289 a_6472_45840# a_6171_45002# 0.005155f
C39290 a_5907_45546# a_5205_44484# 2.98e-20
C39291 a_2711_45572# a_7705_45326# 0.001295f
C39292 a_11322_45546# a_n913_45002# 4.81e-21
C39293 a_20753_42852# a_18597_46090# 3.09e-19
C39294 a_8325_42308# a_n971_45724# 4.93e-20
C39295 a_5379_42460# a_4791_45118# 0.197725f
C39296 a_5742_30871# w_1575_34946# 0.032598f
C39297 CAL_N a_22469_39537# 0.024229f
C39298 a_22521_40599# a_22821_38993# 0.002401f
C39299 a_22469_40625# a_22545_38993# 9.26e-21
C39300 a_8912_37509# CAL_P 0.007121f
C39301 a_n1453_44318# a_n2293_45546# 1.08e-19
C39302 a_1467_44172# a_n443_42852# 0.008372f
C39303 a_2998_44172# a_3503_45724# 3.02e-21
C39304 a_15940_43402# a_15227_44166# 6.38e-19
C39305 a_3080_42308# a_4185_45028# 0.030391f
C39306 a_3540_43646# a_1823_45246# 8.6e-19
C39307 a_20193_45348# RST_Z 6.04e-20
C39308 a_8199_44636# VDD 1.43837f
C39309 a_6598_45938# a_n1741_47186# 1.67e-22
C39310 a_4099_45572# a_n237_47217# 1.6e-19
C39311 a_20820_30879# a_20205_31679# 0.087297f
C39312 a_20202_43084# a_21167_46155# 2.55e-19
C39313 a_22591_46660# a_20692_30879# 0.001224f
C39314 a_8349_46414# a_8034_45724# 0.05863f
C39315 a_20708_46348# a_6945_45028# 0.002334f
C39316 a_20075_46420# a_10809_44734# 2.78e-20
C39317 a_6031_43396# a_743_42282# 4.36e-20
C39318 a_14955_43396# a_15781_43660# 1.56e-19
C39319 a_3626_43646# a_5649_42852# 0.032897f
C39320 a_19237_31679# a_n1630_35242# 7.69e-20
C39321 a_n1761_44111# a_n784_42308# 0.034368f
C39322 a_n97_42460# a_133_43172# 0.002798f
C39323 a_14579_43548# a_16137_43396# 6.3e-20
C39324 a_n356_44636# a_18548_42308# 4.18e-20
C39325 a_14021_43940# a_22165_42308# 6.79e-20
C39326 a_10341_43396# a_14621_43646# 4.92e-19
C39327 a_5063_47570# DATA[3] 3.18e-20
C39328 a_n1613_43370# DATA[0] 0.001615f
C39329 a_21588_30879# a_22609_38406# 6.34e-21
C39330 a_n1379_43218# VDD 1.08e-19
C39331 a_15037_45618# a_14539_43914# 4.54e-21
C39332 a_15415_45028# a_15595_45028# 0.185422f
C39333 a_14537_43396# a_1307_43914# 0.0516f
C39334 a_8696_44636# a_10334_44484# 0.001709f
C39335 a_7499_43078# a_n2661_42834# 0.089963f
C39336 a_21513_45002# a_20567_45036# 2e-19
C39337 a_19479_31679# a_19778_44110# 1.24e-19
C39338 a_6431_45366# a_6517_45366# 0.006584f
C39339 a_3065_45002# a_n2293_42834# 0.021132f
C39340 a_n467_45028# a_n2661_43370# 0.016799f
C39341 a_5111_44636# a_5009_45028# 8.57e-19
C39342 a_5147_45002# a_5093_45028# 0.008723f
C39343 a_21363_45546# a_20193_45348# 1.77e-22
C39344 a_n4064_39616# a_n2442_46660# 0.224005f
C39345 a_4933_42558# a_3090_45724# 1.87e-19
C39346 a_n2216_39866# a_n2956_39768# 0.001489f
C39347 a_16547_43609# a_n357_42282# 0.004365f
C39348 a_5755_42852# a_526_44458# 0.054788f
C39349 a_12293_43646# a_n443_42852# 7.27e-19
C39350 a_2437_43646# a_2266_47243# 4.08e-19
C39351 a_n2661_45010# a_n2312_40392# 1.45e-20
C39352 en_comp a_13507_46334# 1.11e-19
C39353 a_413_45260# a_18780_47178# 2.11e-19
C39354 a_14180_45002# a_4915_47217# 0.007501f
C39355 a_375_42282# a_n1151_42308# 1.19e-19
C39356 a_16680_45572# a_n743_46660# 0.011176f
C39357 a_18341_45572# a_5807_45002# 0.0023f
C39358 a_18175_45572# a_13747_46662# 0.03273f
C39359 a_18479_45785# a_13661_43548# 0.087389f
C39360 a_7_45899# a_n443_42852# 5.72e-19
C39361 a_685_42968# a_n2293_42282# 2.16e-20
C39362 a_12545_42858# a_12895_43230# 0.215953f
C39363 a_12379_42858# a_13460_43230# 0.102325f
C39364 a_15743_43084# a_15597_42852# 0.055955f
C39365 a_3539_42460# a_6123_31319# 9e-21
C39366 a_3626_43646# a_7963_42308# 0.003306f
C39367 a_2982_43646# a_8515_42308# 1.02e-19
C39368 a_n97_42460# a_13333_42558# 1.53e-20
C39369 a_22959_46660# EN_OFFSET_CAL 0.050989f
C39370 a_3422_30871# C5_N_btm 1.71e-19
C39371 VDAC_P a_11206_38545# 0.101449f
C39372 a_8912_37509# CAL_N 0.017398f
C39373 a_13070_42354# VDD 0.18656f
C39374 a_n1741_47186# a_11599_46634# 0.164599f
C39375 a_n746_45260# a_n1435_47204# 5.74e-19
C39376 a_n1151_42308# a_5129_47502# 0.002765f
C39377 a_3381_47502# a_4915_47217# 9.99e-20
C39378 a_4007_47204# a_4700_47436# 0.010942f
C39379 a_3785_47178# a_n443_46116# 0.040847f
C39380 a_3815_47204# a_4791_45118# 6.07e-20
C39381 a_4743_44484# a_5343_44458# 4.42e-19
C39382 a_4223_44672# a_6298_44484# 3.26e-19
C39383 a_n2661_43370# a_n2661_43922# 0.13591f
C39384 a_2711_45572# a_2982_43646# 9.28e-19
C39385 a_18479_45785# a_19862_44208# 2.98e-20
C39386 a_2382_45260# a_1414_42308# 0.005789f
C39387 a_n1059_45260# a_7542_44172# 5.06e-21
C39388 a_413_45260# a_895_43940# 0.001706f
C39389 a_n2293_45010# a_n3674_39768# 6.8e-20
C39390 a_2437_43646# a_3499_42826# 1.38e-20
C39391 a_10149_42308# a_526_44458# 1.05e-19
C39392 a_n327_42558# a_n755_45592# 0.003126f
C39393 a_1184_42692# a_n863_45724# 0.563857f
C39394 a_n3674_37592# a_n357_42282# 0.327427f
C39395 a_6428_45938# VDD 4.6e-19
C39396 a_17364_32525# a_11530_34132# 0.007158f
C39397 a_22521_40599# a_21588_30879# 8.64e-20
C39398 a_18479_45785# a_4185_45028# 9.87e-21
C39399 a_22591_45572# a_11415_45002# 0.02488f
C39400 a_15415_45028# a_15559_46634# 3.5e-19
C39401 a_3357_43084# a_22591_46660# 3.95e-20
C39402 a_1307_43914# a_3090_45724# 2.66267f
C39403 a_13777_45326# a_15227_44166# 4.73e-20
C39404 a_949_44458# a_n2293_46634# 4.57e-19
C39405 a_18248_44752# a_12549_44172# 2.68e-19
C39406 a_19479_31679# a_20820_30879# 0.052973f
C39407 a_19963_31679# a_20202_43084# 5.55e-20
C39408 a_16019_45002# a_14976_45028# 2.19e-19
C39409 a_n1699_44726# a_n2438_43548# 3.52e-19
C39410 a_2437_43646# a_22959_46660# 8.36e-21
C39411 a_7499_43078# a_5066_45546# 0.002848f
C39412 a_6171_45002# a_14513_46634# 1.88e-21
C39413 a_413_45260# a_18285_46348# 1.46e-20
C39414 a_8696_44636# a_9290_44172# 0.032264f
C39415 a_11688_45572# a_2324_44458# 7.44e-19
C39416 a_n23_44458# a_n1613_43370# 2.25e-20
C39417 a_14815_43914# a_10227_46804# 0.004604f
C39418 a_n984_44318# a_n2497_47436# 8.35e-19
C39419 a_5342_30871# a_4958_30871# 10.9366f
C39420 a_n3674_38680# a_n4318_38216# 2.82961f
C39421 a_17701_42308# a_17124_42282# 5.83e-19
C39422 a_n3674_39304# a_n4251_39616# 5.77e-20
C39423 a_13747_46662# a_n743_46660# 0.042998f
C39424 a_n2840_46634# a_n2956_39768# 0.156182f
C39425 a_n881_46662# a_3699_46634# 0.001985f
C39426 a_n1613_43370# a_3524_46660# 0.28004f
C39427 a_n443_46116# a_3090_45724# 0.011392f
C39428 a_4915_47217# a_15009_46634# 1.25e-20
C39429 a_6151_47436# a_12816_46660# 6.67e-20
C39430 a_10227_46804# a_10467_46802# 0.678578f
C39431 a_17517_44484# a_22959_44484# 0.00251f
C39432 a_n2661_43922# a_2998_44172# 0.003621f
C39433 a_5708_44484# a_5495_43940# 1.89e-19
C39434 a_n2661_42834# a_3600_43914# 0.012088f
C39435 a_16979_44734# a_15682_43940# 0.001729f
C39436 a_n2293_42834# a_458_43396# 0.003568f
C39437 a_1307_43914# a_6547_43396# 1.88e-19
C39438 a_20362_44736# a_20596_44850# 0.006453f
C39439 a_11967_42832# a_21398_44850# 0.01381f
C39440 a_14539_43914# a_17737_43940# 5.43e-19
C39441 a_n2017_45002# a_16759_43396# 1.39e-21
C39442 a_n913_45002# a_16409_43396# 9.35e-21
C39443 a_n1059_45260# a_16977_43638# 1.07e-19
C39444 a_3537_45260# a_10341_43396# 4.95e-20
C39445 a_8953_45002# a_8685_43396# 6.4e-21
C39446 a_6123_31319# C9_P_btm 9.33e-20
C39447 a_5932_42308# C4_P_btm 0.032349f
C39448 a_20205_31679# C8_N_btm 1.65e-20
C39449 a_20692_30879# C7_N_btm 0.001136f
C39450 a_17538_32519# SMPL_ON_N 0.029166f
C39451 a_9145_43396# a_n971_45724# 2.62e-19
C39452 a_7287_43370# a_4791_45118# 3.82e-21
C39453 a_3232_43370# a_n755_45592# 4.34e-19
C39454 a_327_44734# a_n443_42852# 0.005815f
C39455 a_413_45260# a_1609_45822# 0.001816f
C39456 a_6298_44484# a_6419_46155# 4.03e-19
C39457 a_20567_45036# a_10809_44734# 5.98e-22
C39458 a_21359_45002# a_21137_46414# 8.41e-21
C39459 a_4223_44672# a_5937_45572# 0.016442f
C39460 a_17801_45144# a_17715_44484# 2.78e-19
C39461 a_7639_45394# a_8049_45260# 2.57e-19
C39462 a_3353_43940# a_768_44030# 4.43e-19
C39463 a_14485_44260# a_5807_45002# 1.16e-20
C39464 a_11341_43940# a_n2293_46634# 0.487839f
C39465 a_18579_44172# a_3090_45724# 0.16932f
C39466 a_5495_43940# a_5257_43370# 0.009999f
C39467 a_14021_43940# a_13661_43548# 0.103152f
C39468 a_20159_44458# a_19466_46812# 1.25e-19
C39469 a_20640_44752# a_15227_44166# 3.05e-21
C39470 a_12607_44458# a_3483_46348# 0.001786f
C39471 a_18143_47464# VDD 0.388551f
C39472 a_18057_42282# a_19511_42282# 1.23e-20
C39473 a_17303_42282# a_13258_32519# 0.064259f
C39474 a_6123_31319# a_n4209_38502# 6.28e-22
C39475 a_n2661_46098# a_n901_46420# 0.054328f
C39476 a_1983_46706# a_1823_45246# 0.005043f
C39477 a_2107_46812# a_2202_46116# 0.008835f
C39478 a_948_46660# a_167_45260# 8.29e-21
C39479 a_3090_45724# a_17609_46634# 9.39e-20
C39480 a_11901_46660# a_12156_46660# 0.06121f
C39481 a_15368_46634# a_15559_46634# 0.022471f
C39482 a_10428_46928# a_765_45546# 0.003387f
C39483 a_11186_47026# a_10933_46660# 4.61e-19
C39484 a_14976_45028# a_16292_46812# 1.49e-19
C39485 a_12549_44172# a_2324_44458# 0.506903f
C39486 a_5807_45002# a_11387_46155# 0.005659f
C39487 a_n1925_46634# a_5068_46348# 4.81e-20
C39488 a_11599_46634# a_10586_45546# 1.89e-19
C39489 a_n2497_47436# a_3503_45724# 4.5e-21
C39490 a_n971_45724# a_n1099_45572# 0.508925f
C39491 a_n746_45260# a_380_45546# 0.003276f
C39492 a_n237_47217# a_n452_45724# 6.22e-21
C39493 a_1431_47204# a_n2661_45546# 3.64e-21
C39494 a_n743_46660# a_4419_46090# 0.032595f
C39495 a_2889_44172# a_n97_42460# 2.34e-20
C39496 a_19862_44208# a_14021_43940# 0.021104f
C39497 a_9313_44734# a_17324_43396# 2.24e-20
C39498 a_11827_44484# a_12545_42858# 1.69e-22
C39499 a_8333_44056# a_8415_44056# 0.004999f
C39500 a_n967_45348# a_n473_42460# 9.24e-19
C39501 a_n913_45002# a_564_42282# 1.62e-19
C39502 a_n1059_45260# a_n1630_35242# 0.007613f
C39503 a_n2017_45002# a_1067_42314# 0.01039f
C39504 a_2127_44172# VDD 0.138239f
C39505 C5_N_btm VREF_GND 0.676559f
C39506 C4_N_btm VCM 0.716447f
C39507 C6_N_btm VREF 1.41944f
C39508 C7_N_btm VIN_N 1.52449f
C39509 a_11823_42460# a_14033_45822# 0.093809f
C39510 a_10193_42453# a_16115_45572# 0.001215f
C39511 a_8336_45822# a_8192_45572# 6.84e-19
C39512 a_9049_44484# a_8696_44636# 0.043734f
C39513 a_14021_43940# a_4185_45028# 0.038946f
C39514 a_n2157_42858# a_n2438_43548# 0.266513f
C39515 a_9396_43370# a_3090_45724# 0.003506f
C39516 a_14673_44172# a_n357_42282# 4.84e-20
C39517 a_12429_44172# a_2324_44458# 1.55e-21
C39518 a_22165_42308# a_13507_46334# 0.126777f
C39519 a_765_45546# VDD 2.19953f
C39520 a_22959_46660# a_22959_46124# 0.026152f
C39521 a_15227_44166# a_19240_46482# 2.61e-19
C39522 a_21076_30879# a_10809_44734# 0.002069f
C39523 a_3483_46348# a_10903_43370# 0.404121f
C39524 a_7920_46348# a_8199_44636# 5.3e-19
C39525 a_6419_46155# a_5937_45572# 1.25e-20
C39526 a_8016_46348# a_8349_46414# 0.232167f
C39527 a_4007_47204# DATA[2] 0.337596f
C39528 a_10729_43914# a_10518_42984# 4.92e-21
C39529 a_10057_43914# a_9803_42558# 5.35e-21
C39530 a_3626_43646# a_8685_43396# 8.81e-20
C39531 a_10405_44172# a_10835_43094# 2.45e-20
C39532 a_18494_42460# a_19511_42282# 0.047119f
C39533 a_8975_43940# a_9223_42460# 8.9e-22
C39534 a_18184_42460# a_19647_42308# 0.034507f
C39535 a_20193_45348# a_17303_42282# 0.013391f
C39536 a_6197_43396# a_6655_43762# 0.027317f
C39537 a_11967_42832# a_17141_43172# 0.001676f
C39538 a_n2293_43922# a_n4318_37592# 0.019728f
C39539 a_19479_31679# C8_N_btm 1.65e-20
C39540 a_19963_31679# C5_N_btm 1.11e-20
C39541 a_11322_45546# a_n2661_44458# 0.005353f
C39542 a_4880_45572# a_4743_44484# 7.1e-20
C39543 a_2711_45572# a_14539_43914# 0.199754f
C39544 a_413_45260# a_3065_45002# 0.027891f
C39545 a_1667_45002# a_2382_45260# 3.51e-19
C39546 a_n1059_45260# a_5205_44484# 3.03e-20
C39547 a_22465_38105# SMPL_ON_N 0.001357f
C39548 a_766_43646# a_n357_42282# 0.004396f
C39549 a_2896_43646# a_n863_45724# 1.77e-20
C39550 a_4905_42826# a_n755_45592# 7.37e-20
C39551 a_3422_30871# C5_P_btm 1.71e-19
C39552 a_17730_32519# a_18194_35068# 1.21e-19
C39553 a_509_45822# VDD 0.190119f
C39554 a_13527_45546# a_12549_44172# 0.09647f
C39555 a_10193_42453# a_5807_45002# 5.69e-19
C39556 a_3775_45552# a_n1925_46634# 4.34e-21
C39557 a_6598_45938# a_n743_46660# 0.001817f
C39558 a_2711_45572# a_2107_46812# 0.034922f
C39559 a_13163_45724# a_768_44030# 3.17e-20
C39560 a_1990_45572# a_n2293_46634# 1.08e-19
C39561 a_15037_45618# a_11453_44696# 1.16e-20
C39562 a_16855_45546# a_13507_46334# 2.29e-21
C39563 a_18175_45572# a_11599_46634# 0.844188f
C39564 a_18691_45572# a_12861_44030# 0.007387f
C39565 a_n2956_37592# SMPL_ON_P 0.03953f
C39566 a_n467_45028# a_n2497_47436# 2.36e-19
C39567 a_n2017_45002# a_n746_45260# 2.03e-19
C39568 a_2437_43646# a_n1151_42308# 0.036608f
C39569 a_n1059_45260# a_n971_45724# 0.322275f
C39570 a_n2433_43396# a_n3674_37592# 5.99e-20
C39571 a_n1177_43370# a_n961_42308# 1.24e-19
C39572 a_18525_43370# a_18249_42858# 0.002332f
C39573 a_15743_43084# a_18083_42858# 0.00444f
C39574 a_5649_42852# a_8037_42858# 2.33e-20
C39575 a_4361_42308# a_9127_43156# 2.94e-19
C39576 a_743_42282# a_10796_42968# 1e-19
C39577 a_15493_43396# a_15959_42545# 8.88e-21
C39578 a_3422_30871# a_n3420_38528# 0.031237f
C39579 a_n1736_43218# a_n1545_43230# 4.61e-19
C39580 a_n4318_38680# a_n1379_43218# 1.55e-20
C39581 a_8685_43396# a_8649_43218# 7.48e-20
C39582 a_15125_43396# a_5342_30871# 3.56e-20
C39583 a_19333_46634# RST_Z 1.4e-20
C39584 a_13607_46688# CLK 2.1e-20
C39585 a_15227_44166# START 0.001035f
C39586 a_3754_39964# VDAC_Ni 7.07e-21
C39587 VDAC_Pi a_7754_38968# 8.23e-20
C39588 a_n4064_37984# a_n4334_37440# 9.42e-19
C39589 a_n3420_37984# a_n3690_37440# 0.017537f
C39590 a_3754_39466# a_3754_39134# 0.296258f
C39591 a_n2302_37984# a_n4209_37414# 9.15e-19
C39592 a_n2946_37984# a_n3565_37414# 9.15e-19
C39593 a_n3690_38304# a_n3420_37440# 7.84e-19
C39594 a_n4318_38216# VDD 0.538766f
C39595 a_21513_45002# a_20679_44626# 0.001342f
C39596 a_3537_45260# a_n2293_43922# 1.59e-19
C39597 a_5691_45260# a_5708_44484# 5.85e-20
C39598 a_4558_45348# a_n2661_42834# 8.96e-21
C39599 a_4574_45260# a_n2661_43922# 9.45e-20
C39600 a_18184_42460# a_11691_44458# 2.38e-19
C39601 a_16922_45042# a_18450_45144# 0.002084f
C39602 a_19778_44110# a_20193_45348# 0.020562f
C39603 a_17719_45144# a_17801_45144# 0.00659f
C39604 a_10193_42453# a_19478_44306# 4.96e-20
C39605 a_1307_43914# a_n356_44636# 0.013327f
C39606 a_n2293_42834# a_6298_44484# 0.002718f
C39607 a_n2661_43370# a_n452_44636# 0.002717f
C39608 a_21101_45002# a_11827_44484# 0.006993f
C39609 a_7174_31319# a_20202_43084# 5.3e-20
C39610 a_15764_42576# a_4185_45028# 1.97e-19
C39611 a_13258_32519# a_20820_30879# 0.056725f
C39612 a_133_42852# a_n443_42852# 0.004247f
C39613 a_n1630_35242# a_n1925_42282# 0.049072f
C39614 a_8292_43218# a_n357_42282# 0.002687f
C39615 a_19721_31679# SMPL_ON_N 0.029197f
C39616 a_n2661_44458# a_12465_44636# 3.22e-19
C39617 a_12883_44458# a_12861_44030# 0.041056f
C39618 a_n356_44636# a_n443_46116# 0.004124f
C39619 a_n2661_43922# a_n2497_47436# 0.095407f
C39620 a_7640_43914# a_2063_45854# 1.19e-20
C39621 a_20841_45814# a_19692_46634# 0.003435f
C39622 a_3357_43084# a_12991_46634# 5.11e-20
C39623 a_413_45260# a_10249_46116# 4.88e-20
C39624 a_5691_45260# a_5257_43370# 0.009554f
C39625 a_20623_45572# a_19466_46812# 2.08e-19
C39626 a_2711_45572# a_14493_46090# 7.68e-21
C39627 a_13711_45394# a_13661_43548# 4.59e-20
C39628 a_14309_45348# a_5807_45002# 7.13e-19
C39629 a_1423_45028# a_1799_45572# 2.07e-20
C39630 a_16922_45042# a_12549_44172# 0.803336f
C39631 a_8746_45002# a_3483_46348# 0.605995f
C39632 a_4361_42308# a_17124_42282# 0.008373f
C39633 a_4190_30871# a_17531_42308# 3.05e-20
C39634 a_743_42282# a_4958_30871# 0.063224f
C39635 a_7871_42858# a_8515_42308# 2.54e-20
C39636 a_8037_42858# a_7963_42308# 8.28e-20
C39637 a_n2293_42282# a_n1329_42308# 4.66e-19
C39638 a_13507_46334# a_13661_43548# 0.038602f
C39639 a_20894_47436# a_19321_45002# 1.6e-20
C39640 a_19787_47423# a_19594_46812# 0.108653f
C39641 a_11599_46634# a_n743_46660# 0.248412f
C39642 a_18479_47436# a_21588_30879# 2.9e-20
C39643 a_n1435_47204# a_383_46660# 4.95e-20
C39644 a_9313_45822# a_2107_46812# 0.298046f
C39645 a_n1741_47186# a_7411_46660# 8.61e-20
C39646 a_2063_45854# a_4651_46660# 1.12e-19
C39647 a_n443_46116# a_3699_46634# 0.036317f
C39648 a_n971_45724# a_3878_46660# 0.00101f
C39649 a_13556_45296# a_13565_43940# 4.17e-20
C39650 a_9482_43914# a_15037_43940# 1.66e-20
C39651 a_n699_43396# a_2127_44172# 7.77e-20
C39652 a_742_44458# a_2889_44172# 2.44e-20
C39653 a_n2661_42834# a_12189_44484# 0.010003f
C39654 a_1307_43914# a_9165_43940# 0.003526f
C39655 a_n2661_43922# a_11909_44484# 2.94e-20
C39656 a_3537_45260# a_n97_42460# 0.74108f
C39657 a_413_45260# a_458_43396# 1.25e-20
C39658 a_n913_45002# a_n1557_42282# 0.015193f
C39659 a_n3565_38502# a_n2810_45572# 0.409424f
C39660 a_2382_45260# VDD 1.6285f
C39661 COMP_P a_22459_39145# 0.032214f
C39662 a_11691_44458# a_12741_44636# 0.81445f
C39663 a_14403_45348# a_3483_46348# 2.17e-20
C39664 a_5495_43940# a_5807_45002# 3.78e-19
C39665 a_n1761_44111# a_n2438_43548# 0.001148f
C39666 a_4558_45348# a_5066_45546# 0.009388f
C39667 a_n2661_43370# a_5164_46348# 0.010428f
C39668 a_n2293_42834# a_5937_45572# 0.097247f
C39669 a_8137_45348# a_8199_44636# 1.55e-21
C39670 a_17737_43940# a_11453_44696# 2.12e-20
C39671 a_19862_44208# a_13507_46334# 5.48e-20
C39672 a_15493_43940# a_18479_47436# 0.05409f
C39673 a_11341_43940# a_18597_46090# 0.033543f
C39674 a_n447_43370# a_n2497_47436# 0.192476f
C39675 a_n2267_43396# SMPL_ON_P 0.001234f
C39676 a_n2840_43370# a_n971_45724# 3.49e-20
C39677 a_n3674_37592# a_n4064_40160# 0.022617f
C39678 a_n4318_37592# a_n3420_39616# 0.020563f
C39679 a_n1630_35242# a_n4315_30879# 0.129428f
C39680 a_n3674_38216# a_n4064_39616# 0.020042f
C39681 a_5342_30871# C7_N_btm 5.39e-19
C39682 a_5534_30871# C9_N_btm 7.29e-20
C39683 C2_P_btm VIN_P 0.502408f
C39684 C5_P_btm VREF_GND 0.676559f
C39685 C6_P_btm VCM 0.877162f
C39686 RST_Z CLK 0.064624f
C39687 C4_P_btm VREF 0.98728f
C39688 a_19594_46812# a_20107_46660# 0.001514f
C39689 a_13661_43548# a_20623_46660# 4.62e-21
C39690 a_19321_45002# a_20411_46873# 7.75e-19
C39691 a_10428_46928# a_10623_46897# 0.21686f
C39692 a_9863_46634# a_10249_46116# 0.027588f
C39693 a_8492_46660# a_6755_46942# 0.024647f
C39694 a_7411_46660# a_7832_46660# 0.086708f
C39695 a_10150_46912# a_10554_47026# 0.051162f
C39696 a_n237_47217# a_2981_46116# 0.024703f
C39697 a_n746_45260# a_526_44458# 0.096099f
C39698 a_n971_45724# a_n1925_42282# 5.37e-19
C39699 a_13487_47204# a_10903_43370# 1.95e-20
C39700 a_13717_47436# a_12594_46348# 4.38e-22
C39701 a_n1435_47204# a_13351_46090# 4.5e-21
C39702 a_10227_46804# a_8016_46348# 0.093061f
C39703 a_11599_46634# a_11189_46129# 0.0158f
C39704 a_13507_46334# a_4185_45028# 0.479559f
C39705 a_4883_46098# a_3483_46348# 0.813604f
C39706 a_n1059_45260# a_3863_42891# 4.31e-19
C39707 a_n913_45002# a_8483_43230# 2.14e-19
C39708 a_n2293_42834# a_n967_43230# 7.58e-20
C39709 a_13076_44458# a_9145_43396# 1.6e-19
C39710 a_11967_42832# a_18797_44260# 3.24e-19
C39711 a_7499_43078# a_9885_42558# 0.020607f
C39712 a_10193_42453# a_9223_42460# 6.94e-19
C39713 a_1307_43914# a_12379_42858# 2.23e-20
C39714 a_18184_42460# a_4190_30871# 0.630738f
C39715 a_n356_44636# a_9396_43370# 1.18e-20
C39716 a_n2661_43922# a_1568_43370# 4.28e-22
C39717 a_n2661_42834# a_1756_43548# 9.68e-20
C39718 a_13556_45296# a_5534_30871# 1.32e-21
C39719 a_15433_44458# VDD 0.201121f
C39720 a_n3420_38528# VREF_GND 0.047244f
C39721 a_2711_45572# a_12427_45724# 0.014959f
C39722 a_4808_45572# a_4880_45572# 0.003395f
C39723 a_949_44458# a_2277_45546# 6.13e-20
C39724 a_4223_44672# a_n443_42852# 0.001694f
C39725 a_10617_44484# a_10586_45546# 9.55e-19
C39726 a_12710_44260# a_13059_46348# 1.05e-20
C39727 a_10341_43396# a_n2293_46634# 2.04894f
C39728 a_10867_43940# a_3090_45724# 0.00115f
C39729 a_3080_42308# a_5257_43370# 0.00466f
C39730 a_15743_43084# a_12549_44172# 0.021095f
C39731 a_5841_44260# a_n2293_46098# 8.09e-20
C39732 a_5013_44260# a_4185_45028# 3.66e-19
C39733 a_5663_43940# a_3483_46348# 0.00218f
C39734 a_22223_45572# RST_Z 7.78e-20
C39735 a_2437_43646# START 0.12936f
C39736 a_10623_46897# VDD 0.189083f
C39737 a_7174_31319# C5_N_btm 3.27e-20
C39738 a_n3674_37592# a_n4064_37440# 0.651412f
C39739 a_n1630_35242# a_n3420_37440# 6.45e-19
C39740 a_383_46660# a_380_45546# 1.76e-21
C39741 a_n2293_46634# a_n356_45724# 6.18e-19
C39742 a_n743_46660# a_1848_45724# 0.003213f
C39743 a_n2438_43548# a_997_45618# 0.008987f
C39744 a_8492_46660# a_8049_45260# 4.06e-21
C39745 a_33_46660# a_310_45028# 3.11e-20
C39746 a_n133_46660# a_n755_45592# 2.19e-22
C39747 a_948_46660# a_n863_45724# 1.85e-20
C39748 a_14035_46660# a_12594_46348# 9.29e-22
C39749 a_15227_44166# a_19553_46090# 0.047784f
C39750 a_19466_46812# a_18819_46122# 0.02948f
C39751 a_19333_46634# a_18985_46122# 0.002899f
C39752 a_14976_45028# a_6945_45028# 2.34e-19
C39753 a_15009_46634# a_10809_44734# 0.00292f
C39754 a_5891_43370# a_8495_42852# 3.14e-20
C39755 a_17973_43940# a_17499_43370# 0.018568f
C39756 a_n97_42460# a_1049_43396# 0.195034f
C39757 a_14021_43940# a_14579_43548# 1.31e-19
C39758 a_17737_43940# a_17324_43396# 0.001548f
C39759 a_15493_43396# a_16243_43396# 0.041358f
C39760 a_11967_42832# a_15567_42826# 0.067391f
C39761 a_n4318_40392# a_n1630_35242# 1.96e-19
C39762 a_14401_32519# a_2982_43646# 4.51e-20
C39763 a_n2956_37592# a_n2946_39072# 2.49e-19
C39764 a_n1655_43396# VDD 8.44e-20
C39765 a_20273_45572# a_22591_45572# 4.71e-20
C39766 a_21188_45572# a_2437_43646# 0.00191f
C39767 a_20841_45814# a_3357_43084# 0.047766f
C39768 a_20107_45572# a_19963_31679# 3.1e-20
C39769 a_15765_45572# a_6171_45002# 0.001099f
C39770 a_2711_45572# a_14309_45028# 0.028068f
C39771 a_16243_43396# a_3483_46348# 0.001863f
C39772 a_21487_43396# a_20202_43084# 0.019942f
C39773 a_13635_43156# a_3090_45724# 0.00703f
C39774 a_n3674_38680# a_n2956_39768# 0.023454f
C39775 a_15493_43940# a_n443_42852# 0.301211f
C39776 a_1443_43940# a_n863_45724# 0.005869f
C39777 a_1891_43646# a_526_44458# 4.7e-19
C39778 a_10695_43548# a_10903_43370# 0.041719f
C39779 a_14205_43396# a_9290_44172# 0.010382f
C39780 a_6123_31319# a_n2312_39304# 5.16e-21
C39781 a_n4064_39616# w_1575_34946# 0.027505f
C39782 a_6347_46155# VDD 2.18e-20
C39783 a_2711_45572# a_11453_44696# 0.033654f
C39784 a_6472_45840# a_4883_46098# 4.6e-20
C39785 a_6469_45572# a_6151_47436# 6.03e-19
C39786 a_10490_45724# a_12861_44030# 2.29e-20
C39787 a_8192_45572# a_n1151_42308# 9.32e-20
C39788 a_2324_44458# a_n2661_45546# 0.019247f
C39789 a_10903_43370# a_n357_42282# 0.028411f
C39790 a_18985_46122# a_20062_46116# 1.46e-19
C39791 a_n3565_37414# C1_P_btm 0.001047f
C39792 a_18579_44172# a_18727_42674# 4.15e-22
C39793 a_2982_43646# a_18817_42826# 3.67e-20
C39794 a_3626_43646# a_17333_42852# 2.21e-20
C39795 a_8685_43396# a_8037_42858# 0.001875f
C39796 a_15743_43084# a_21855_43396# 0.001426f
C39797 a_19268_43646# a_4361_42308# 4.9e-21
C39798 a_1709_42852# VDD 0.001589f
C39799 a_3775_45552# a_3600_43914# 9.84e-21
C39800 a_13556_45296# a_11691_44458# 0.399095f
C39801 a_14797_45144# a_11827_44484# 5.28e-21
C39802 a_5837_45028# a_n2661_43370# 0.005758f
C39803 a_8488_45348# a_8560_45348# 0.003395f
C39804 a_8696_44636# a_12553_44484# 8.86e-20
C39805 a_3065_45002# a_2779_44458# 0.001276f
C39806 a_6431_45366# a_n2661_44458# 7.71e-21
C39807 a_2382_45260# a_n699_43396# 0.075387f
C39808 a_2905_42968# a_n755_45592# 4.85e-20
C39809 a_3681_42891# a_n357_42282# 0.005491f
C39810 a_4149_42891# a_526_44458# 2.3e-20
C39811 a_17538_32519# a_18194_35068# 1.07e-19
C39812 a_6886_37412# w_1575_34946# 0.001151f
C39813 a_16223_45938# a_6755_46942# 0.002064f
C39814 a_327_44734# a_n2661_46634# 5.27e-21
C39815 a_5691_45260# a_5807_45002# 0.19412f
C39816 a_n143_45144# a_n2293_46634# 0.00576f
C39817 a_8953_45002# a_768_44030# 3.3e-19
C39818 a_n2956_37592# a_n2438_43548# 0.004958f
C39819 a_n967_45348# a_n1021_46688# 5.18e-21
C39820 a_22876_39857# VDD 3.12e-19
C39821 a_n452_44636# a_n2497_47436# 0.001121f
C39822 a_n2267_44484# SMPL_ON_P 5.37e-21
C39823 a_n1641_43230# COMP_P 8.01e-19
C39824 a_n1991_42858# a_n961_42308# 0.001344f
C39825 a_12379_42858# a_13003_42852# 9.73e-19
C39826 a_n1423_42826# a_n1329_42308# 0.001077f
C39827 a_12281_43396# a_12563_42308# 0.173003f
C39828 a_n4318_38680# a_n4318_38216# 0.055776f
C39829 a_12895_43230# a_13157_43218# 0.001705f
C39830 a_12545_42858# a_13569_43230# 2.36e-20
C39831 a_4361_42308# a_1755_42282# 0.015476f
C39832 a_15095_43370# a_14113_42308# 6.79e-20
C39833 a_2982_43646# a_21421_42336# 9.11e-19
C39834 a_n4318_39304# a_n4251_39392# 3.13e-19
C39835 a_3626_43646# a_18997_42308# 8.14e-19
C39836 a_10809_44734# SINGLE_ENDED 0.008311f
C39837 a_1239_39587# VDD 0.530104f
C39838 a_13717_47436# a_12465_44636# 0.049141f
C39839 a_14955_47212# a_13507_46334# 2.55e-20
C39840 a_3785_47178# a_n1613_43370# 0.006133f
C39841 a_16327_47482# a_18597_46090# 1.28053f
C39842 a_17591_47464# a_10227_46804# 0.292864f
C39843 a_13487_47204# a_4883_46098# 4.22e-20
C39844 a_16588_47582# a_18143_47464# 4.68e-20
C39845 a_3357_43084# a_5829_43940# 0.00562f
C39846 a_n2661_45010# a_2455_43940# 3.99e-19
C39847 a_n2293_45010# a_1443_43940# 3.99e-19
C39848 a_11322_45546# a_9145_43396# 4.56e-21
C39849 a_626_44172# a_1525_44260# 2.9e-21
C39850 a_10193_42453# a_13667_43396# 5.44e-20
C39851 a_2711_45572# a_17324_43396# 7.1e-20
C39852 a_8746_45002# a_10695_43548# 3.62e-21
C39853 a_n2293_42834# a_2479_44172# 0.021799f
C39854 a_9482_43914# a_9028_43914# 0.092045f
C39855 a_5009_45028# a_3905_42865# 1.03e-19
C39856 a_n2661_43370# a_n809_44244# 5.6e-20
C39857 a_11827_44484# a_20766_44850# 0.004974f
C39858 a_20193_45348# a_20159_44458# 5.71e-19
C39859 a_10440_44484# a_10617_44484# 0.134298f
C39860 a_5883_43914# a_n2661_43922# 0.028328f
C39861 a_21359_45002# a_19279_43940# 8.47e-19
C39862 a_11963_45334# a_10949_43914# 1.06e-20
C39863 a_5742_30871# a_n443_42852# 2.05e-19
C39864 a_15959_42545# a_n357_42282# 9.81e-20
C39865 a_20712_42282# a_13259_45724# 1.03e-19
C39866 a_n2302_38778# a_n2956_38680# 0.038021f
C39867 a_n2860_38778# a_n2956_39304# 8.73e-19
C39868 a_5342_30871# C3_P_btm 8.34e-20
C39869 a_5534_30871# RST_Z 0.031803f
C39870 a_3537_45260# a_5204_45822# 2.3e-20
C39871 a_4574_45260# a_5164_46348# 1.44e-19
C39872 a_413_45260# a_5937_45572# 4.56e-21
C39873 a_10729_43914# a_2063_45854# 0.004795f
C39874 a_16223_45938# a_8049_45260# 0.004651f
C39875 a_2211_45572# a_1609_45822# 8.16e-20
C39876 a_11827_44484# a_14976_45028# 7.51e-20
C39877 a_9241_44734# a_2107_46812# 1.31e-19
C39878 a_n2293_43922# a_n2293_46634# 0.02819f
C39879 a_18911_45144# a_19466_46812# 1.84e-19
C39880 a_4927_45028# a_4185_45028# 0.004584f
C39881 a_n2661_42834# a_n2312_38680# 1.97e-21
C39882 a_18184_42460# a_15227_44166# 3.08e-21
C39883 a_3232_43370# a_3483_46348# 0.220803f
C39884 a_16328_43172# a_4958_30871# 1.29e-20
C39885 a_5342_30871# a_n4064_38528# 0.028644f
C39886 a_n784_42308# a_9223_42460# 1.96e-20
C39887 a_1606_42308# a_7227_42308# 3.31e-20
C39888 a_1755_42282# a_6761_42308# 0.008867f
C39889 a_961_42354# a_5934_30871# 1.72e-20
C39890 a_3318_42354# a_4921_42308# 1.41e-19
C39891 a_13467_32519# C3_N_btm 1.74e-19
C39892 a_4190_30871# C9_N_btm 0.002182f
C39893 a_22545_38993# a_22609_38406# 2.17e-21
C39894 a_22459_39145# a_22705_37990# 7.75e-19
C39895 a_22521_39511# a_22705_38406# 0.004065f
C39896 a_22469_39537# a_22876_39857# 2.68e-19
C39897 a_12891_46348# a_11735_46660# 0.034334f
C39898 a_n2661_46634# a_10150_46912# 0.010702f
C39899 a_n743_46660# a_7411_46660# 5e-20
C39900 a_n1925_46634# a_7577_46660# 0.007837f
C39901 a_2107_46812# a_6540_46812# 5.62e-20
C39902 a_3177_46902# a_3686_47026# 2.6e-19
C39903 a_2609_46660# a_3055_46660# 2.28e-19
C39904 a_11309_47204# a_11813_46116# 0.007374f
C39905 a_n881_46662# a_15009_46634# 0.004074f
C39906 a_n1613_43370# a_3090_45724# 0.039515f
C39907 a_12465_44636# a_14035_46660# 6.36e-21
C39908 a_4883_46098# a_14513_46634# 3.52e-20
C39909 a_16327_47482# a_19123_46287# 0.005309f
C39910 a_16588_47582# a_765_45546# 0.004612f
C39911 a_17591_47464# a_17339_46660# 3.44e-20
C39912 a_11599_46634# a_20841_46902# 9.01e-21
C39913 a_10227_46804# a_15312_46660# 3.7e-20
C39914 a_n237_47217# a_167_45260# 0.280171f
C39915 a_584_46384# a_376_46348# 0.232754f
C39916 a_n1151_42308# a_n1853_46287# 0.024093f
C39917 a_1209_47178# a_1176_45822# 4.3e-19
C39918 a_1239_47204# a_1208_46090# 7.29e-20
C39919 a_n971_45724# a_2698_46116# 0.001385f
C39920 a_3785_47178# a_n2293_46098# 1.6e-20
C39921 a_n1741_47186# a_4185_45028# 4.26e-20
C39922 a_n2109_47186# a_4704_46090# 4.15e-21
C39923 a_949_44458# a_1209_43370# 6.32e-19
C39924 a_1414_42308# a_453_43940# 0.248504f
C39925 a_644_44056# a_895_43940# 0.106452f
C39926 a_742_44458# a_1049_43396# 2.13e-19
C39927 a_18989_43940# a_18797_44260# 9.07e-19
C39928 a_1115_44172# a_2479_44172# 9.15e-20
C39929 a_n2661_43922# a_12495_44260# 2.04e-19
C39930 a_n2661_42834# a_12603_44260# 6.24e-19
C39931 a_n913_45002# a_3935_42891# 5.11e-21
C39932 a_n1059_45260# a_4520_42826# 0.004119f
C39933 a_n2017_45002# a_5111_42852# 1.11e-19
C39934 a_11206_38545# VDD 8.87267f
C39935 a_5343_44458# VDD 0.49245f
C39936 a_19647_42308# RST_Z 4.07e-20
C39937 a_4958_30871# VIN_P 0.025339f
C39938 a_7174_31319# C5_P_btm 3.27e-20
C39939 a_n4209_39590# a_n1838_35608# 2.05e-19
C39940 a_n4064_40160# EN_VIN_BSTR_P 0.187697f
C39941 a_21398_44850# a_20202_43084# 4.42e-20
C39942 a_20980_44850# a_11415_45002# 0.00141f
C39943 a_11341_43940# a_6755_46942# 3.7e-19
C39944 a_n2267_43396# a_n2438_43548# 0.120634f
C39945 a_n97_42460# a_n2293_46634# 0.108602f
C39946 a_3626_43646# a_768_44030# 0.002415f
C39947 a_n2661_43370# a_3316_45546# 0.022024f
C39948 a_11691_44458# a_16375_45002# 1.43e-19
C39949 a_n2293_42834# a_n443_42852# 1.60683f
C39950 a_9159_44484# a_9290_44172# 7.16e-20
C39951 a_6547_43396# a_n1613_43370# 0.154311f
C39952 a_9145_43396# a_12465_44636# 9.6e-20
C39953 a_10695_43548# a_4883_46098# 3.82e-20
C39954 a_10341_43396# a_18597_46090# 0.027979f
C39955 a_12281_43396# a_10227_46804# 6.09e-20
C39956 a_16547_43609# a_12861_44030# 3.22e-19
C39957 a_n1641_43230# a_n2497_47436# 0.001225f
C39958 a_n2472_42826# SMPL_ON_P 3.03e-19
C39959 a_n2956_39768# VDD 0.697168f
C39960 a_n3690_39616# a_n4209_39304# 2.69e-19
C39961 a_n4209_39590# a_n3690_39392# 2.69e-19
C39962 a_n4064_39616# a_n4251_39616# 0.001131f
C39963 a_5934_30871# C0_dummy_P_btm 1.48e-19
C39964 a_6123_31319# C0_N_btm 0.018968f
C39965 a_5932_42308# C5_N_btm 5.59e-19
C39966 a_3090_45724# a_n2293_46098# 0.642755f
C39967 a_15227_44166# a_12741_44636# 0.250453f
C39968 a_19692_46634# a_11415_45002# 0.033537f
C39969 a_n2661_46098# a_n1736_46482# 0.024986f
C39970 a_n2438_43548# a_1337_46116# 0.008585f
C39971 a_5807_45002# a_11387_46482# 2.88e-19
C39972 a_2107_46812# a_1337_46436# 1.09e-19
C39973 a_n743_46660# a_4365_46436# 2.75e-20
C39974 a_4883_46098# a_n357_42282# 4.03e-19
C39975 a_n2312_39304# a_n2472_45546# 0.001998f
C39976 a_n2312_40392# a_n2956_38216# 0.053778f
C39977 en_comp a_15486_42560# 1.51e-21
C39978 a_n913_45002# a_15890_42674# 1.94e-19
C39979 a_n2661_42282# a_7112_43396# 1.53e-19
C39980 a_14539_43914# a_18817_42826# 5.94e-20
C39981 a_n2293_42834# a_n2104_42282# 0.004809f
C39982 a_n356_44636# a_13635_43156# 9.74e-20
C39983 a_1307_43914# a_3823_42558# 6.3e-20
C39984 a_17970_44736# a_18083_42858# 5.77e-21
C39985 a_5891_43370# a_9127_43156# 0.457718f
C39986 a_20640_44752# a_21259_43561# 6.9e-19
C39987 a_20159_44458# a_20301_43646# 3.21e-20
C39988 a_16680_45572# a_16147_45260# 2.09e-19
C39989 a_16855_45546# a_18175_45572# 2.91e-21
C39990 a_5907_45546# a_6431_45366# 9.96e-19
C39991 a_6194_45824# a_6171_45002# 0.006466f
C39992 a_5263_45724# a_5205_44484# 4.99e-21
C39993 a_2711_45572# a_6709_45028# 0.002223f
C39994 a_6229_45572# a_3357_43084# 6.33e-19
C39995 a_6472_45840# a_3232_43370# 0.001072f
C39996 a_7754_38968# RST_Z 9.75e-19
C39997 a_5267_42460# a_4791_45118# 0.138738f
C39998 a_22521_40599# a_22545_38993# 6.99e-20
C39999 a_22469_40625# a_22521_39511# 0.65678f
C40000 CAL_N a_22821_38993# 2.99e-19
C40001 VDAC_N CAL_P 7.22e-21
C40002 a_n4064_37440# EN_VIN_BSTR_P 0.031982f
C40003 a_2998_44172# a_3316_45546# 4.99e-19
C40004 a_1115_44172# a_n443_42852# 4.54e-19
C40005 a_5663_43940# a_n357_42282# 1.55e-19
C40006 a_15868_43402# a_15227_44166# 3.62e-19
C40007 a_n2293_42282# a_n2312_38680# 3.75e-20
C40008 a_2982_43646# a_1823_45246# 0.022597f
C40009 a_4699_43561# a_4185_45028# 0.010947f
C40010 a_19721_31679# a_18194_35068# 1e-19
C40011 a_8349_46414# VDD 0.209819f
C40012 a_5263_45724# a_n971_45724# 1.03e-20
C40013 a_11415_45002# a_20692_30879# 7.79e-19
C40014 a_22591_46660# a_20205_31679# 0.004038f
C40015 a_8016_46348# a_8034_45724# 0.254614f
C40016 a_6419_46155# a_6633_46155# 0.005572f
C40017 a_9823_46155# a_5066_45546# 3.05e-20
C40018 a_19335_46494# a_10809_44734# 7.36e-20
C40019 a_14955_43396# a_15681_43442# 9.54e-19
C40020 a_14021_43940# a_21671_42860# 6.16e-20
C40021 a_n1761_44111# a_196_42282# 2.46e-19
C40022 a_n356_44636# a_18310_42308# 5.53e-19
C40023 a_n1655_43396# a_n4318_38680# 7.29e-20
C40024 a_5063_47570# DATA[2] 7.59e-20
C40025 a_n1545_43230# VDD 1.95e-19
C40026 a_n955_45028# a_n2661_43370# 6.51e-19
C40027 a_21513_45002# a_18494_42460# 8.98e-20
C40028 a_6171_45002# a_6517_45366# 6.95e-19
C40029 a_6431_45366# a_6125_45348# 7.37e-20
C40030 a_5147_45002# a_5009_45028# 0.007368f
C40031 a_4558_45348# a_5093_45028# 0.001257f
C40032 a_20623_45572# a_20193_45348# 4.8e-19
C40033 a_9049_44484# a_9159_44484# 0.031707f
C40034 a_8696_44636# a_10157_44484# 0.004815f
C40035 a_14537_43396# a_16019_45002# 5.14e-20
C40036 a_8162_45546# a_n2661_43922# 3.6e-21
C40037 a_n2946_39866# a_n2442_46660# 0.024649f
C40038 a_n3565_39590# a_n2312_38680# 0.031736f
C40039 a_n2860_39866# a_n2956_39768# 0.001355f
C40040 a_16243_43396# a_n357_42282# 1.3e-19
C40041 a_5111_42852# a_526_44458# 0.265994f
C40042 a_4520_42826# a_n1925_42282# 6.4e-19
C40043 a_2437_43646# a_3315_47570# 8.57e-19
C40044 a_413_45260# a_18479_47436# 2.86e-19
C40045 a_13777_45326# a_4915_47217# 8.78e-22
C40046 a_6171_45002# a_12861_44030# 0.05507f
C40047 a_1423_45028# a_2063_45854# 4.66e-20
C40048 a_16855_45546# a_n743_46660# 0.005475f
C40049 a_16147_45260# a_13747_46662# 0.027471f
C40050 a_18479_45785# a_5807_45002# 0.174313f
C40051 a_17668_45572# a_12549_44172# 5.63e-20
C40052 a_18175_45572# a_13661_43548# 0.029369f
C40053 a_n310_45899# a_n443_42852# 4.25e-19
C40054 a_n97_42460# a_13249_42558# 5.74e-19
C40055 a_12089_42308# a_12895_43230# 4.25e-19
C40056 a_2982_43646# a_5934_30871# 0.178f
C40057 a_3626_43646# a_6123_31319# 0.109715f
C40058 a_12379_42858# a_13635_43156# 0.043475f
C40059 a_12545_42858# a_13113_42826# 0.178024f
C40060 a_12741_44636# EN_OFFSET_CAL 0.230064f
C40061 a_3422_30871# C4_N_btm 1.36e-19
C40062 a_8912_37509# a_11206_38545# 1.26605f
C40063 VDAC_N CAL_N 2.77e-19
C40064 a_12563_42308# VDD 0.254292f
C40065 a_n971_45724# a_n1435_47204# 2.23698f
C40066 a_n1151_42308# a_4915_47217# 0.1374f
C40067 a_2063_45854# a_6491_46660# 9.61e-20
C40068 a_3381_47502# a_n443_46116# 4.13e-20
C40069 a_3785_47178# a_4791_45118# 0.010875f
C40070 a_4223_44672# a_5518_44484# 0.003606f
C40071 a_18479_45785# a_19478_44306# 0.005615f
C40072 a_n2661_43370# a_n2661_42834# 0.306215f
C40073 a_n699_43396# a_5343_44458# 9.51e-20
C40074 a_n2472_45002# a_n3674_39768# 1.13e-19
C40075 a_2274_45254# a_1414_42308# 1.01e-20
C40076 a_n2017_45002# a_7542_44172# 2.92e-21
C40077 a_413_45260# a_2479_44172# 0.008619f
C40078 a_n2293_45010# a_n4318_39768# 1.61e-21
C40079 a_n2661_45010# a_n1644_44306# 7.26e-19
C40080 a_2437_43646# a_2537_44260# 7.55e-20
C40081 a_1576_42282# a_n863_45724# 0.05148f
C40082 a_n327_42558# a_n357_42282# 0.006254f
C40083 a_n784_42308# a_n755_45592# 0.711298f
C40084 a_4880_45572# VDD 0.004682f
C40085 a_4190_30871# RST_Z 0.087843f
C40086 a_14209_32519# EN_VIN_BSTR_N 0.032853f
C40087 a_n2267_44484# a_n2438_43548# 0.120608f
C40088 a_3357_43084# a_11415_45002# 0.053912f
C40089 a_16019_45002# a_3090_45724# 3.78e-20
C40090 a_13556_45296# a_15227_44166# 0.047404f
C40091 a_17970_44736# a_12549_44172# 3.76e-20
C40092 a_742_44458# a_n2293_46634# 2.95e-19
C40093 a_2437_43646# a_12741_44636# 0.023858f
C40094 a_15595_45028# a_14976_45028# 3.96e-19
C40095 a_15415_45028# a_15368_46634# 2.5e-19
C40096 a_8568_45546# a_5066_45546# 0.04527f
C40097 a_2711_45572# a_14180_46482# 3.42e-20
C40098 a_327_44734# a_765_45546# 5.49e-20
C40099 a_n356_44636# a_n1613_43370# 5.31e-19
C40100 a_9313_44734# SMPL_ON_N 2.16e-20
C40101 a_14112_44734# a_10227_46804# 1.24e-19
C40102 a_14673_44172# a_12861_44030# 0.015418f
C40103 a_n809_44244# a_n2497_47436# 0.029871f
C40104 a_n2840_42282# a_n4318_38216# 0.015074f
C40105 a_n3674_38680# a_n2472_42282# 5e-19
C40106 a_17701_42308# a_16522_42674# 7.63e-21
C40107 a_13661_43548# a_n743_46660# 1.74e-19
C40108 a_n881_46662# a_2959_46660# 2.16e-20
C40109 a_n1613_43370# a_3699_46634# 0.344308f
C40110 a_4791_45118# a_3090_45724# 0.206257f
C40111 a_6151_47436# a_12991_46634# 2.17e-19
C40112 a_4915_47217# a_14084_46812# 0.038663f
C40113 a_16327_47482# a_6755_46942# 0.067305f
C40114 a_10227_46804# a_10428_46928# 0.060058f
C40115 a_n1059_45260# a_16409_43396# 4.57e-19
C40116 a_n913_45002# a_16547_43609# 4.63e-21
C40117 a_n2017_45002# a_16977_43638# 6.48e-21
C40118 a_3232_43370# a_10695_43548# 4.03e-21
C40119 a_3537_45260# a_9885_43646# 2e-19
C40120 a_n2293_42834# a_n229_43646# 0.001042f
C40121 a_10193_42453# a_21195_42852# 0.005652f
C40122 a_11967_42832# a_20980_44850# 8.49e-19
C40123 a_19615_44636# a_19789_44512# 0.006584f
C40124 a_1307_43914# a_6765_43638# 2.03e-20
C40125 a_n2661_43370# a_n1352_43396# 3.84e-21
C40126 a_n2661_42834# a_2998_44172# 0.790177f
C40127 a_5708_44484# a_5013_44260# 3.54e-19
C40128 a_n2661_43922# a_2889_44172# 0.001413f
C40129 a_17517_44484# a_17730_32519# 0.00864f
C40130 a_20679_44626# a_18579_44172# 1.41e-20
C40131 a_14539_43914# a_15682_43940# 0.161926f
C40132 a_20692_30879# C6_N_btm 0.080378f
C40133 a_20205_31679# C7_N_btm 1.43e-20
C40134 a_8560_45348# VDD 0.004463f
C40135 a_6123_31319# C10_P_btm 1.34e-19
C40136 a_5932_42308# C5_P_btm 5.59e-19
C40137 a_8423_43396# a_n971_45724# 0.001593f
C40138 a_n2661_43370# a_5066_45546# 4.51e-19
C40139 a_3537_45260# a_3503_45724# 0.00137f
C40140 a_413_45260# a_n443_42852# 0.005091f
C40141 a_327_44734# a_509_45822# 5.3e-20
C40142 a_3232_43370# a_n357_42282# 4.05e-19
C40143 a_11827_44484# a_19900_46494# 1.49e-22
C40144 a_21101_45002# a_21137_46414# 1.79e-19
C40145 a_11691_44458# a_18985_46122# 2.44e-22
C40146 a_6298_44484# a_6165_46155# 2.52e-20
C40147 a_18494_42460# a_10809_44734# 8.81e-22
C40148 a_4223_44672# a_8199_44636# 4.87e-19
C40149 a_9165_43940# a_n1613_43370# 2.36e-20
C40150 a_3052_44056# a_768_44030# 1.06e-19
C40151 a_19615_44636# a_19466_46812# 3.92e-20
C40152 a_13829_44260# a_13661_43548# 0.001195f
C40153 a_5013_44260# a_5257_43370# 0.002385f
C40154 a_20362_44736# a_15227_44166# 4.57e-21
C40155 a_14021_43940# a_5807_45002# 0.001299f
C40156 a_11967_42832# a_19692_46634# 0.032909f
C40157 a_8975_43940# a_3483_46348# 0.016137f
C40158 a_10227_46804# VDD 2.77567f
C40159 a_5932_42308# a_n3420_38528# 0.001859f
C40160 a_18057_42282# a_18548_42308# 0.00278f
C40161 a_4958_30871# a_13258_32519# 0.033151f
C40162 a_5742_30871# a_1736_39587# 7.65e-20
C40163 a_17303_42282# a_19647_42308# 3.68e-19
C40164 a_n743_46660# a_4185_45028# 0.036891f
C40165 a_n2661_46098# a_n1641_46494# 0.035694f
C40166 a_3699_46634# a_n2293_46098# 1.64e-20
C40167 a_2107_46812# a_1823_45246# 0.007836f
C40168 a_1123_46634# a_167_45260# 0.003466f
C40169 a_14976_45028# a_15559_46634# 0.001514f
C40170 a_11735_46660# a_12359_47026# 9.73e-19
C40171 a_11813_46116# a_12156_46660# 0.157972f
C40172 a_10150_46912# a_765_45546# 4.34e-20
C40173 a_12891_46348# a_2324_44458# 0.026746f
C40174 a_12549_44172# a_14840_46494# 9.46e-38
C40175 a_5807_45002# a_11133_46155# 0.00164f
C40176 a_n2661_46634# a_6419_46155# 1.76e-21
C40177 a_n1925_46634# a_4704_46090# 2.8e-20
C40178 a_5342_30871# a_7754_40130# 7.04e-19
C40179 a_16327_47482# a_8049_45260# 0.605463f
C40180 a_n2497_47436# a_3316_45546# 1.34e-19
C40181 a_n237_47217# a_n863_45724# 3.43e-19
C40182 a_n746_45260# a_n452_45724# 3.79e-20
C40183 a_1239_47204# a_n2661_45546# 4.78e-21
C40184 a_n452_47436# a_n1099_45572# 3.76e-20
C40185 a_n2293_42834# a_1793_42852# 1.98e-35
C40186 a_644_44056# a_458_43396# 2.18e-19
C40187 a_2675_43914# a_n97_42460# 1.83e-19
C40188 a_19478_44306# a_14021_43940# 5.41e-20
C40189 a_9313_44734# a_17499_43370# 2.25e-19
C40190 a_20512_43084# a_2982_43646# 0.029475f
C40191 a_n2661_44458# a_3935_42891# 5.85e-22
C40192 a_11341_43940# a_11173_44260# 0.049235f
C40193 a_n967_45348# a_n961_42308# 0.174237f
C40194 a_n1059_45260# a_564_42282# 0.043244f
C40195 a_n2017_45002# a_n1630_35242# 0.111641f
C40196 a_n913_45002# a_n3674_37592# 8.1e-20
C40197 a_453_43940# VDD 0.225569f
C40198 a_11823_42460# a_12016_45572# 1.71e-19
C40199 a_10210_45822# a_10907_45822# 0.013775f
C40200 a_7499_43078# a_8696_44636# 0.155392f
C40201 a_10193_42453# a_16333_45814# 7.72e-20
C40202 C4_N_btm VREF_GND 0.671882f
C40203 C3_N_btm VCM 0.716273f
C40204 C5_N_btm VREF 0.987144f
C40205 C6_N_btm VIN_N 0.391905f
C40206 a_10341_43396# a_6755_46942# 8.9e-20
C40207 a_n2472_42826# a_n2438_43548# 0.026866f
C40208 a_8791_43396# a_3090_45724# 0.00173f
C40209 a_8037_42858# a_768_44030# 4.29e-23
C40210 a_n4318_38680# a_n2956_39768# 0.023624f
C40211 a_7542_44172# a_526_44458# 7.82e-21
C40212 a_11750_44172# a_2324_44458# 4.42e-21
C40213 a_21671_42860# a_13507_46334# 0.001831f
C40214 a_9482_43914# CLK 3.96e-20
C40215 a_17339_46660# VDD 0.555596f
C40216 a_12741_44636# a_22959_46124# 3.35e-19
C40217 a_15227_44166# a_16375_45002# 0.117865f
C40218 a_22959_46660# a_10809_44734# 0.015306f
C40219 a_6165_46155# a_5937_45572# 1.14e-20
C40220 a_11967_42832# a_16877_43172# 0.003239f
C40221 a_18494_42460# a_18548_42308# 0.005603f
C40222 a_7287_43370# a_8147_43396# 2.55e-19
C40223 a_18184_42460# a_19511_42282# 0.058931f
C40224 a_19778_44110# a_19647_42308# 2.28e-21
C40225 a_n2293_43922# a_n1736_42282# 4.89e-19
C40226 a_5891_43370# a_1755_42282# 3.89e-20
C40227 a_10405_44172# a_10518_42984# 2.78e-20
C40228 a_19319_43548# a_19700_43370# 0.006809f
C40229 a_6197_43396# a_6452_43396# 0.06121f
C40230 a_10729_43914# a_10083_42826# 5.47e-19
C40231 a_3815_47204# DATA[2] 0.022461f
C40232 a_n1151_42308# DATA[5] 0.006171f
C40233 a_19963_31679# C4_N_btm 0.001041f
C40234 a_19479_31679# C7_N_btm 1.43e-20
C40235 a_2711_45572# a_16112_44458# 0.183744f
C40236 a_10490_45724# a_n2661_44458# 2.68e-21
C40237 a_413_45260# a_2680_45002# 0.01804f
C40238 a_n913_45002# a_6171_45002# 8.52e-21
C40239 a_n2017_45002# a_5205_44484# 2.49e-20
C40240 a_4905_42826# a_n357_42282# 0.026713f
C40241 a_3080_42308# a_n755_45592# 0.237742f
C40242 a_3539_42460# a_n2661_45546# 0.091495f
C40243 a_13814_43218# a_3090_45724# 2.67e-19
C40244 a_10533_42308# a_n2293_46634# 2.12e-21
C40245 a_3422_30871# C6_P_btm 2.2e-19
C40246 a_17730_32519# EN_VIN_BSTR_N 0.072552f
C40247 a_n906_45572# VDD 2.32e-19
C40248 a_13527_45546# a_12891_46348# 0.002777f
C40249 a_7227_45028# a_n1925_46634# 5.87e-19
C40250 a_10180_45724# a_5807_45002# 6.9e-20
C40251 a_6667_45809# a_n743_46660# 0.001764f
C40252 a_13163_45724# a_12549_44172# 0.172293f
C40253 a_16147_45260# a_11599_46634# 0.065926f
C40254 a_18909_45814# a_12861_44030# 2.11e-19
C40255 a_n2810_45028# SMPL_ON_P 0.039597f
C40256 a_n2109_45247# a_n746_45260# 1.91e-20
C40257 a_n2017_45002# a_n971_45724# 0.048447f
C40258 a_2437_43646# a_3160_47472# 0.003877f
C40259 a_18783_43370# a_18083_42858# 9.54e-20
C40260 a_16664_43396# a_16414_43172# 4.88e-19
C40261 a_15743_43084# a_17701_42308# 1.11e-19
C40262 a_18429_43548# a_18249_42858# 0.001117f
C40263 a_5649_42852# a_7765_42852# 1.28e-20
C40264 a_4361_42308# a_8387_43230# 5.06e-20
C40265 a_743_42282# a_10835_43094# 8.66e-20
C40266 a_n2012_43396# a_n2104_42282# 2.27e-20
C40267 a_n1352_43396# COMP_P 1.02e-19
C40268 a_5829_43940# a_5755_42308# 9.03e-21
C40269 a_11341_43940# a_14456_42282# 4.56e-23
C40270 a_15493_43396# a_15803_42450# 8.19e-21
C40271 a_n4318_39304# a_n3674_37592# 0.024848f
C40272 a_n4318_38680# a_n1545_43230# 2.34e-20
C40273 a_15037_43396# a_5342_30871# 9.74e-22
C40274 a_15227_44166# RST_Z 2.45e-20
C40275 a_12816_46660# CLK 6.39e-21
C40276 a_18834_46812# START 0.001199f
C40277 a_7754_39964# a_7754_38968# 1.48e-20
C40278 a_n4064_37984# a_n4209_37414# 0.027993f
C40279 a_2113_38308# a_3754_38470# 2.91e-19
C40280 a_n3420_37984# a_n3565_37414# 0.032929f
C40281 a_n3690_38304# a_n3690_37440# 0.050585f
C40282 a_n2472_42282# VDD 0.278905f
C40283 a_3232_43370# a_3363_44484# 0.103472f
C40284 a_n913_45002# a_14673_44172# 3.55e-20
C40285 a_21513_45002# a_20640_44752# 1.55e-19
C40286 a_4574_45260# a_n2661_42834# 4.61e-21
C40287 a_3537_45260# a_n2661_43922# 0.058875f
C40288 a_13249_42308# a_10949_43914# 3.22e-19
C40289 a_18911_45144# a_20193_45348# 5.06e-21
C40290 a_19778_44110# a_11691_44458# 0.013164f
C40291 a_16922_45042# a_17969_45144# 0.002405f
C40292 a_17613_45144# a_17801_45144# 7.06e-21
C40293 a_11823_42460# a_14955_43940# 6.42e-21
C40294 a_10193_42453# a_15493_43396# 0.024143f
C40295 a_5837_45028# a_5883_43914# 4.44e-21
C40296 a_n2661_43370# a_n1352_44484# 0.001902f
C40297 a_21005_45260# a_11827_44484# 0.005914f
C40298 a_21101_45002# a_21359_45002# 0.22264f
C40299 a_15486_42560# a_4185_45028# 6.43e-20
C40300 a_20712_42282# a_20202_43084# 0.028679f
C40301 a_n1630_35242# a_526_44458# 9.42e-21
C40302 a_4649_42852# a_n863_45724# 8.36e-21
C40303 a_564_42282# a_n1925_42282# 2.11e-19
C40304 a_7573_43172# a_n357_42282# 9.51e-19
C40305 a_5742_30871# a_8199_44636# 5.25e-20
C40306 a_10723_42308# a_8953_45546# 2.61e-20
C40307 a_18114_32519# SMPL_ON_N 0.02927f
C40308 a_12607_44458# a_12861_44030# 0.020604f
C40309 a_n2661_42834# a_n2497_47436# 0.099608f
C40310 a_n356_44636# a_4791_45118# 0.001203f
C40311 a_6109_44484# a_2063_45854# 1.19e-20
C40312 a_4927_45028# a_5257_43370# 0.003815f
C40313 a_2437_43646# a_13607_46688# 1.22e-21
C40314 a_413_45260# a_10554_47026# 1.94e-20
C40315 a_21363_45546# a_15227_44166# 6.55e-20
C40316 a_20841_45814# a_19466_46812# 1.64e-19
C40317 a_2711_45572# a_13925_46122# 5.04e-19
C40318 a_10193_42453# a_3483_46348# 0.359034f
C40319 a_20273_45572# a_19692_46634# 0.004885f
C40320 a_4361_42308# a_16522_42674# 0.002806f
C40321 a_4190_30871# a_17303_42282# 0.279034f
C40322 a_7765_42852# a_7963_42308# 9.95e-19
C40323 a_8037_42858# a_6123_31319# 5.06e-20
C40324 a_n2293_42282# COMP_P 0.026882f
C40325 a_15743_43084# a_21613_42308# 1.45e-19
C40326 a_7871_42858# a_5934_30871# 0.001545f
C40327 a_12465_44636# a_16285_47570# 1.31e-20
C40328 a_13507_46334# a_5807_45002# 1.64614f
C40329 a_20990_47178# a_13747_46662# 1.78e-20
C40330 a_18479_47436# a_20916_46384# 0.014237f
C40331 a_19386_47436# a_19594_46812# 0.069651f
C40332 a_14955_47212# a_n743_46660# 6.75e-21
C40333 a_19787_47423# a_19321_45002# 0.029499f
C40334 a_n1741_47186# a_5257_43370# 1.22e-19
C40335 a_2063_45854# a_4646_46812# 0.093604f
C40336 a_n443_46116# a_2959_46660# 0.036727f
C40337 a_n971_45724# a_3633_46660# 2.76e-19
C40338 a_949_44458# a_895_43940# 0.002952f
C40339 a_2779_44458# a_2479_44172# 0.001425f
C40340 a_9482_43914# a_13565_43940# 3.82e-19
C40341 a_n699_43396# a_453_43940# 0.006917f
C40342 a_742_44458# a_2675_43914# 2.91e-21
C40343 a_11823_42460# a_5649_42852# 2.49e-19
C40344 a_n2661_43922# a_11541_44484# 0.004005f
C40345 a_1307_43914# a_8487_44056# 4.35e-19
C40346 a_n1059_45260# a_n1557_42282# 0.031252f
C40347 a_2274_45254# VDD 0.256655f
C40348 COMP_P a_22521_40055# 7.41e-20
C40349 a_16237_45028# a_11415_45002# 1.72e-19
C40350 a_19113_45348# a_12741_44636# 0.003982f
C40351 a_14309_45348# a_3483_46348# 2.79e-20
C40352 a_n2065_43946# a_n2438_43548# 0.265458f
C40353 a_n984_44318# a_n2293_46634# 2.17e-21
C40354 a_9313_44734# a_8270_45546# 7.8e-20
C40355 a_5205_44484# a_526_44458# 2.73e-20
C40356 a_2437_43646# a_16375_45002# 2.49e-20
C40357 a_n2293_42834# a_8199_44636# 0.048304f
C40358 a_7639_45394# a_5937_45572# 2.11e-19
C40359 a_15682_43940# a_11453_44696# 1.72e-19
C40360 a_21115_43940# a_18597_46090# 0.015966f
C40361 a_22223_43948# a_18479_47436# 1.31e-20
C40362 a_n1352_43396# a_n2497_47436# 0.061218f
C40363 a_11551_42558# a_12563_42308# 2.06e-19
C40364 a_2351_42308# a_7174_31319# 4.88e-21
C40365 a_n3674_37592# a_n4334_40480# 7.51e-19
C40366 COMP_P a_n3565_39590# 4.08e-21
C40367 a_5342_30871# C6_N_btm 0.012f
C40368 a_5534_30871# C8_N_btm 5.29e-19
C40369 C3_P_btm VIN_P 0.455045f
C40370 C7_P_btm VCM 1.58335f
C40371 C6_P_btm VREF_GND 0.836236f
C40372 RST_Z EN_OFFSET_CAL 0.044122f
C40373 C5_P_btm VREF 0.987144f
C40374 a_19321_45002# a_20107_46660# 0.003274f
C40375 a_19594_46812# a_19551_46910# 0.07027f
C40376 a_8667_46634# a_6755_46942# 0.011524f
C40377 a_10428_46928# a_10467_46802# 0.820079f
C40378 a_10150_46912# a_10623_46897# 7.99e-20
C40379 a_7577_46660# a_6999_46987# 5.54e-20
C40380 a_5257_43370# a_7832_46660# 2.48e-21
C40381 a_13747_46662# a_20273_46660# 1.3e-20
C40382 a_n971_45724# a_526_44458# 0.21769f
C40383 a_n1151_42308# a_10809_44734# 0.334692f
C40384 a_n1435_47204# a_12594_46348# 1.19e-20
C40385 a_12861_44030# a_10903_43370# 0.378457f
C40386 a_13381_47204# a_13351_46090# 7.4e-20
C40387 a_4883_46098# a_3147_46376# 1.86e-19
C40388 a_n913_45002# a_8292_43218# 0.001438f
C40389 a_n2293_42834# a_n1379_43218# 4.33e-19
C40390 a_18494_42460# a_19177_43646# 7.87e-20
C40391 a_19778_44110# a_4190_30871# 5.46e-20
C40392 a_7499_43078# a_9377_42558# 2.82e-19
C40393 a_10193_42453# a_8791_42308# 2.96e-20
C40394 a_16922_45042# a_4361_42308# 0.00825f
C40395 a_11967_42832# a_18533_44260# 0.001389f
C40396 a_18184_42460# a_21259_43561# 5.43e-20
C40397 a_n356_44636# a_8791_43396# 5.34e-22
C40398 a_8975_43940# a_10695_43548# 7.03e-21
C40399 a_n2661_42834# a_1568_43370# 1.03e-19
C40400 a_n2661_43922# a_1049_43396# 2.6e-21
C40401 a_9482_43914# a_5534_30871# 1.74e-21
C40402 a_14815_43914# VDD 0.307386f
C40403 a_n3565_38502# VCM 0.035399f
C40404 a_n3420_38528# VREF 2.43e-19
C40405 a_n4064_38528# VIN_P 0.044919f
C40406 a_2711_45572# a_11962_45724# 0.054424f
C40407 a_5024_45822# a_4880_45572# 6.84e-19
C40408 a_7227_45028# a_7499_43078# 5.28e-22
C40409 a_13887_32519# SMPL_ON_N 0.029238f
C40410 a_n2293_42282# a_n2497_47436# 1.08e-20
C40411 a_18783_43370# a_12549_44172# 2.61e-20
C40412 a_10651_43940# a_3090_45724# 0.014051f
C40413 a_9885_43646# a_n2293_46634# 0.005638f
C40414 a_12603_44260# a_13059_46348# 3.73e-20
C40415 a_4699_43561# a_5257_43370# 2.14e-19
C40416 a_13837_43396# a_13661_43548# 1.48e-20
C40417 a_n97_42460# a_6755_46942# 2.11e-19
C40418 a_949_44458# a_1609_45822# 0.005374f
C40419 a_2779_44458# a_n443_42852# 1.63e-20
C40420 a_8975_43940# a_n357_42282# 1.39e-20
C40421 a_5495_43940# a_3483_46348# 3.25e-20
C40422 a_2437_43646# RST_Z 0.082469f
C40423 a_10467_46802# VDD 0.401016f
C40424 a_7174_31319# C4_N_btm 2.64e-20
C40425 a_13258_32519# C7_N_btm 1.33e-20
C40426 a_n1630_35242# a_n3690_37440# 1.11e-19
C40427 a_5934_30871# a_n4064_37984# 2.14e-19
C40428 a_n3674_37592# a_n2946_37690# 4.03e-21
C40429 COMP_P a_3726_37500# 0.00602f
C40430 a_n1925_46634# a_2957_45546# 1.1e-20
C40431 a_n743_46660# a_997_45618# 2.04e-19
C40432 a_8667_46634# a_8049_45260# 0.00101f
C40433 a_n2438_43548# a_n755_45592# 0.213107f
C40434 a_1123_46634# a_n863_45724# 2.27e-20
C40435 a_n133_46660# a_n357_42282# 1.78e-19
C40436 a_33_46660# a_n1099_45572# 5.76e-21
C40437 a_171_46873# a_310_45028# 1.19e-19
C40438 a_2107_46812# a_n2293_45546# 2.33e-20
C40439 a_19333_46634# a_18819_46122# 0.003156f
C40440 a_15227_44166# a_18985_46122# 0.287996f
C40441 a_14180_46812# a_10903_43370# 7.73e-19
C40442 a_3090_45724# a_6945_45028# 2.98e-19
C40443 a_14084_46812# a_10809_44734# 0.004861f
C40444 a_17737_43940# a_17499_43370# 0.013048f
C40445 a_n97_42460# a_1209_43370# 0.027601f
C40446 a_14021_43940# a_13667_43396# 4.76e-19
C40447 a_21381_43940# a_2982_43646# 0.236232f
C40448 a_15493_43396# a_16137_43396# 0.023247f
C40449 a_11967_42832# a_5342_30871# 0.077151f
C40450 a_104_43370# a_458_43396# 0.07022f
C40451 a_5891_43370# a_9306_43218# 5.41e-19
C40452 a_n2956_37592# a_n3420_39072# 6.43e-20
C40453 a_n1821_43396# VDD 3.05e-20
C40454 a_21188_45572# a_21513_45002# 0.002147f
C40455 a_21363_45546# a_2437_43646# 0.006526f
C40456 a_20107_45572# a_22591_45572# 3.89e-21
C40457 a_15903_45785# a_6171_45002# 0.011492f
C40458 a_3775_45552# a_n2661_43370# 1.33e-21
C40459 a_20273_45572# a_3357_43084# 0.358383f
C40460 a_16137_43396# a_3483_46348# 6.08e-20
C40461 a_12895_43230# a_3090_45724# 0.004563f
C40462 a_n2840_42282# a_n2956_39768# 3.63e-20
C40463 a_n1557_42282# a_n1925_42282# 0.013245f
C40464 a_1241_43940# a_n863_45724# 6.18e-19
C40465 a_1427_43646# a_526_44458# 0.028942f
C40466 a_14358_43442# a_9290_44172# 0.001132f
C40467 a_10341_43396# a_8953_45546# 0.001386f
C40468 a_9803_43646# a_10903_43370# 2.58e-19
C40469 a_6123_31319# a_n2312_40392# 7.4e-21
C40470 a_n2302_40160# SMPL_ON_P 1.79e-19
C40471 a_8034_45724# VDD 0.812726f
C40472 a_6194_45824# a_4883_46098# 9.26e-21
C40473 a_6229_45572# a_6151_47436# 0.002879f
C40474 a_11652_45724# a_11459_47204# 7.77e-21
C40475 a_8697_45822# a_4791_45118# 1.06e-20
C40476 a_8120_45572# a_n1151_42308# 5.11e-19
C40477 a_19900_46494# a_20009_46494# 0.007416f
C40478 a_20075_46420# a_20254_46482# 0.007399f
C40479 a_19335_46494# a_19443_46116# 0.057222f
C40480 a_17021_43396# a_16823_43084# 0.002675f
C40481 a_n2661_42282# a_5379_42460# 0.121051f
C40482 a_2982_43646# a_18249_42858# 6.61e-20
C40483 a_3626_43646# a_18083_42858# 9.29e-20
C40484 a_15743_43084# a_4361_42308# 0.020459f
C40485 a_1568_43370# a_n2293_42282# 3.41e-20
C40486 a_15903_45785# a_14673_44172# 1.01e-20
C40487 a_9482_43914# a_11691_44458# 0.616964f
C40488 a_14537_43396# a_11827_44484# 0.076354f
C40489 a_5093_45028# a_n2661_43370# 0.005328f
C40490 a_2274_45254# a_n699_43396# 1.36e-20
C40491 a_6171_45002# a_n2661_44458# 0.001196f
C40492 a_2680_45002# a_2779_44458# 1.99e-19
C40493 a_2382_45260# a_4223_44672# 5.91e-19
C40494 a_13657_42558# a_13059_46348# 3.57e-21
C40495 a_17303_42282# a_15227_44166# 1.37e-19
C40496 a_n13_43084# a_n443_42852# 0.13203f
C40497 a_2905_42968# a_n357_42282# 0.011153f
C40498 a_3863_42891# a_526_44458# 8.86e-21
C40499 a_5342_30871# a_13259_45724# 2.89e-19
C40500 a_961_42354# a_1138_42852# 2.56e-20
C40501 a_17538_32519# EN_VIN_BSTR_N 0.06758f
C40502 a_n2302_37690# SMPL_ON_P 3.04e-19
C40503 a_16020_45572# a_6755_46942# 0.010518f
C40504 a_2437_43646# a_2609_46660# 9.86e-20
C40505 a_8191_45002# a_768_44030# 1.08e-20
C40506 a_n467_45028# a_n2293_46634# 0.008099f
C40507 a_n2810_45028# a_n2438_43548# 0.009971f
C40508 a_4927_45028# a_5807_45002# 6.39e-19
C40509 a_413_45260# a_n2661_46634# 0.029743f
C40510 a_22780_39857# VDD 2.73e-20
C40511 a_n1352_44484# a_n2497_47436# 0.006874f
C40512 a_n1991_42858# a_n1329_42308# 0.001762f
C40513 a_n1423_42826# COMP_P 3.47e-19
C40514 a_n1853_43023# a_n961_42308# 2.96e-20
C40515 a_n4318_38680# a_n2472_42282# 4.31e-19
C40516 a_12281_43396# a_11633_42558# 4.33e-21
C40517 a_10341_43396# a_14456_42282# 2.53e-20
C40518 a_12895_43230# a_12991_43230# 0.013793f
C40519 a_n3674_39304# a_n4318_38216# 0.043431f
C40520 a_13113_42826# a_13157_43218# 3.69e-19
C40521 a_4361_42308# a_1606_42308# 1.99e-20
C40522 a_2982_43646# a_21125_42558# 3.84e-19
C40523 a_n1736_43218# a_n3674_38680# 3.47e-20
C40524 a_22959_46124# RST_Z 0.001356f
C40525 a_10809_44734# START 0.002613f
C40526 a_16327_47482# a_18780_47178# 5.16e-20
C40527 a_13717_47436# a_21811_47423# 6.87e-20
C40528 a_12861_44030# a_4883_46098# 0.076083f
C40529 a_16588_47582# a_10227_46804# 0.039575f
C40530 a_n2216_39866# VDD 0.004696f
C40531 a_2063_45854# a_9804_47204# 0.249806f
C40532 a_n1151_42308# a_n881_46662# 1.41446f
C40533 a_14311_47204# a_13507_46334# 1.05e-20
C40534 a_n1435_47204# a_12465_44636# 0.002293f
C40535 a_3381_47502# a_n1613_43370# 5.5e-21
C40536 a_4700_47436# a_4842_47570# 0.007833f
C40537 a_n1741_47186# a_5807_45002# 0.029376f
C40538 a_3357_43084# a_5745_43940# 0.003915f
C40539 a_n2661_45010# a_2253_43940# 0.003669f
C40540 a_n2293_45010# a_1241_43940# 0.005122f
C40541 a_16922_45042# a_20397_44484# 3.67e-19
C40542 a_9482_43914# a_8333_44056# 6.18e-20
C40543 a_626_44172# a_1241_44260# 1.9e-19
C40544 a_18494_42460# a_18579_44172# 2.2e-19
C40545 a_2711_45572# a_17499_43370# 2.44e-19
C40546 a_11823_42460# a_8685_43396# 0.057344f
C40547 a_8746_45002# a_9803_43646# 1.37e-20
C40548 a_1307_43914# a_3499_42826# 0.532672f
C40549 a_n2293_42834# a_2127_44172# 3.16e-21
C40550 a_n2661_43370# a_n1549_44318# 8.71e-21
C40551 a_11827_44484# a_20835_44721# 0.009929f
C40552 a_15004_44636# a_9313_44734# 6.27e-21
C40553 a_10334_44484# a_10617_44484# 0.003683f
C40554 a_5883_43914# a_n2661_42834# 0.106812f
C40555 a_8701_44490# a_n2661_43922# 0.00848f
C40556 a_21101_45002# a_19279_43940# 6.46e-20
C40557 a_15803_42450# a_n357_42282# 1.12e-19
C40558 a_20107_42308# a_13259_45724# 1.03e-19
C40559 a_n4064_38528# a_n2956_38680# 0.058755f
C40560 a_5342_30871# C4_P_btm 8.98e-20
C40561 a_5534_30871# C2_P_btm 7.46e-20
C40562 a_3537_45260# a_5164_46348# 0.003403f
C40563 a_4558_45348# a_4704_46090# 6.71e-22
C40564 a_2437_43646# a_18985_46122# 4.38e-21
C40565 a_n913_45002# a_10903_43370# 0.021559f
C40566 en_comp a_9290_44172# 1.1e-20
C40567 a_413_45260# a_8199_44636# 4.56e-21
C40568 a_3357_43084# a_18189_46348# 4.56e-21
C40569 a_10405_44172# a_2063_45854# 0.001338f
C40570 a_3499_42826# a_n443_46116# 4.85e-21
C40571 a_19778_44110# a_15227_44166# 6.82e-20
C40572 a_11827_44484# a_3090_45724# 0.066595f
C40573 a_5691_45260# a_3483_46348# 0.005653f
C40574 a_18587_45118# a_19466_46812# 7.19e-20
C40575 a_5111_44636# a_4185_45028# 3.83e-19
C40576 a_n2661_43922# a_n2293_46634# 0.023539f
C40577 a_n2293_43922# a_n2442_46660# 7.85e-20
C40578 a_10193_42453# a_n357_42282# 0.634772f
C40579 a_16020_45572# a_8049_45260# 0.002165f
C40580 a_1990_45572# a_1609_45822# 0.002458f
C40581 a_16751_45260# a_12741_44636# 0.01378f
C40582 a_3823_42558# a_3905_42558# 0.171361f
C40583 a_2351_42308# a_5932_42308# 4.34e-21
C40584 a_n784_42308# a_8791_42308# 3.86e-20
C40585 a_1606_42308# a_6761_42308# 1.94e-20
C40586 a_1184_42692# a_5934_30871# 8.33e-21
C40587 a_13467_32519# C2_N_btm 0.001797f
C40588 a_4190_30871# C8_N_btm 4.06e-19
C40589 a_22521_39511# a_22609_38406# 0.23688f
C40590 a_22521_40055# a_22705_37990# 0.016815f
C40591 a_22459_39145# a_22609_37990# 0.172129f
C40592 a_22469_39537# a_22780_39857# 1.79e-19
C40593 a_n743_46660# a_5257_43370# 0.036418f
C40594 a_n2661_46634# a_9863_46634# 0.010932f
C40595 a_n1925_46634# a_7715_46873# 0.01948f
C40596 a_2107_46812# a_5732_46660# 0.00317f
C40597 a_2609_46660# a_3686_47026# 1.46e-19
C40598 a_5807_45002# a_7832_46660# 0.001677f
C40599 a_2443_46660# a_3055_46660# 0.001881f
C40600 a_11309_47204# a_11735_46660# 0.003123f
C40601 a_12465_44636# a_13885_46660# 0.006386f
C40602 a_4883_46098# a_14180_46812# 8.02e-20
C40603 a_16763_47508# a_765_45546# 0.005699f
C40604 a_4915_47217# a_12741_44636# 0.031734f
C40605 a_11599_46634# a_20273_46660# 0.003014f
C40606 a_10227_46804# a_14447_46660# 2.5e-20
C40607 a_16327_47482# a_18285_46348# 3.07e-20
C40608 a_13717_47436# a_22000_46634# 3.86e-20
C40609 a_n237_47217# a_2202_46116# 0.049087f
C40610 a_584_46384# a_n1076_46494# 5.23e-20
C40611 a_n1151_42308# a_n2157_46122# 0.027101f
C40612 a_1209_47178# a_1208_46090# 7.67e-19
C40613 a_n971_45724# a_2521_46116# 6.68e-20
C40614 a_n746_45260# a_167_45260# 0.234425f
C40615 a_n2109_47186# a_4419_46090# 3.48e-20
C40616 a_949_44458# a_458_43396# 0.001416f
C40617 a_15433_44458# a_15493_43940# 0.001343f
C40618 a_18287_44626# a_19319_43548# 1.07e-20
C40619 a_1467_44172# a_453_43940# 0.05905f
C40620 a_1115_44172# a_2127_44172# 2.04e-20
C40621 a_17517_44484# a_17973_43940# 4.57e-20
C40622 a_10193_42453# a_18707_42852# 0.003123f
C40623 a_742_44458# a_1209_43370# 1.04e-19
C40624 a_175_44278# a_895_43940# 2.38e-19
C40625 a_18989_43940# a_18533_44260# 3.53e-19
C40626 a_n2661_42834# a_12495_44260# 8.52e-19
C40627 a_n913_45002# a_3681_42891# 1.8e-20
C40628 a_n1059_45260# a_3935_42891# 0.004841f
C40629 a_n2017_45002# a_4520_42826# 5.33e-20
C40630 VDAC_P VDD 5.18919f
C40631 a_4743_44484# VDD 0.266843f
C40632 a_19511_42282# RST_Z 2.38e-20
C40633 a_7174_31319# C6_P_btm 2.51e-19
C40634 a_n2302_37984# a_n2956_38216# 0.041408f
C40635 a_13940_44484# a_3483_46348# 1.24e-19
C40636 a_n2129_43609# a_n2438_43548# 0.068602f
C40637 a_3540_43646# a_768_44030# 0.002561f
C40638 a_n2661_43370# a_3218_45724# 6.79e-20
C40639 a_6197_43396# a_n881_46662# 6.52e-20
C40640 a_5891_43370# a_2324_44458# 7.07e-20
C40641 a_6765_43638# a_n1613_43370# 0.164755f
C40642 a_9803_43646# a_4883_46098# 0.002651f
C40643 a_16243_43396# a_12861_44030# 9.34e-20
C40644 a_n2840_42826# SMPL_ON_P 7.81e-19
C40645 a_n4334_39616# a_n4334_39392# 0.052468f
C40646 a_n3565_39590# a_n4209_39304# 5.4667f
C40647 a_n4209_39590# a_n3565_39304# 0.032081f
C40648 a_n4064_40160# a_n4064_39072# 0.06545f
C40649 a_n3420_39616# a_n3607_39616# 0.001546f
C40650 a_n2840_46634# VDD 0.306342f
C40651 a_5934_30871# C0_P_btm 0.015126f
C40652 a_6123_31319# C0_dummy_N_btm 1.31e-19
C40653 a_5932_42308# C4_N_btm 0.032349f
C40654 a_19692_46634# a_20202_43084# 0.172738f
C40655 a_19466_46812# a_11415_45002# 0.037852f
C40656 a_15227_44166# a_20820_30879# 5.72e-19
C40657 a_16751_46987# a_17829_46910# 2.45e-20
C40658 a_5807_45002# a_10586_45546# 0.001693f
C40659 a_12891_46348# a_12839_46116# 0.038804f
C40660 a_n2661_46098# a_n2956_38680# 0.123968f
C40661 a_n743_46660# a_1337_46116# 0.004248f
C40662 a_9863_46634# a_8199_44636# 2.9e-20
C40663 a_8667_46634# a_8953_45546# 0.002384f
C40664 a_8492_46660# a_5937_45572# 0.002914f
C40665 a_n2312_39304# a_n2661_45546# 0.022905f
C40666 a_n2017_45002# a_15720_42674# 1.72e-19
C40667 en_comp a_15051_42282# 1.64e-19
C40668 a_n913_45002# a_15959_42545# 3.53e-19
C40669 a_n1059_45260# a_15890_42674# 2.22e-20
C40670 a_2382_45260# a_5742_30871# 1.17e-20
C40671 a_5111_44636# a_9803_42558# 2.44e-21
C40672 a_14539_43914# a_18249_42858# 2.08e-19
C40673 a_742_44458# a_3059_42968# 1.47e-19
C40674 a_n356_44636# a_12895_43230# 1.3e-20
C40675 a_n2293_42834# a_n4318_38216# 7.97e-19
C40676 a_11967_42832# a_743_42282# 0.043946f
C40677 a_1307_43914# a_3318_42354# 0.001768f
C40678 a_17767_44458# a_18083_42858# 1.98e-19
C40679 a_16979_44734# a_17333_42852# 4.43e-22
C40680 a_17517_44484# a_22591_43396# 7.11e-20
C40681 a_20159_44458# a_4190_30871# 1.81e-20
C40682 a_5891_43370# a_8387_43230# 0.010767f
C40683 a_16855_45546# a_16147_45260# 1.95e-19
C40684 a_15765_45572# a_18341_45572# 0.001304f
C40685 a_8696_44636# a_16377_45572# 2.13e-20
C40686 a_5907_45546# a_6171_45002# 0.001025f
C40687 a_6194_45824# a_3232_43370# 1.03e-19
C40688 a_2711_45572# a_7229_43940# 0.001392f
C40689 a_n97_42460# a_8953_45546# 0.015611f
C40690 a_20753_42852# a_18479_47436# 2.93e-20
C40691 a_3823_42558# a_4791_45118# 0.005746f
C40692 a_15681_43442# a_13059_46348# 2.56e-21
C40693 a_2998_44172# a_3218_45724# 1.18e-19
C40694 a_644_44056# a_n443_42852# 1.15e-19
C40695 a_5495_43940# a_n357_42282# 1.86e-21
C40696 a_3080_42308# a_3483_46348# 2.72e-21
C40697 a_2896_43646# a_1823_45246# 6.58e-19
C40698 a_22521_40599# a_22521_39511# 0.365591f
C40699 CAL_N a_22545_38993# 0.01247f
C40700 a_n4064_37440# a_n923_35174# 0.002259f
C40701 a_6886_37412# CAL_P 0.002915f
C40702 a_18114_32519# a_18194_35068# 6.3e-20
C40703 a_19721_31679# EN_VIN_BSTR_N 0.005343f
C40704 a_8016_46348# VDD 1.42798f
C40705 a_2711_45572# a_n237_47217# 0.025745f
C40706 a_4099_45572# a_n971_45724# 8.72e-19
C40707 a_6511_45714# a_n1741_47186# 4.36e-21
C40708 a_3775_45552# a_n2497_47436# 4.13e-21
C40709 a_11415_45002# a_20205_31679# 0.070403f
C40710 a_20202_43084# a_20692_30879# 3.23e-19
C40711 a_7920_46348# a_8034_45724# 0.032141f
C40712 a_6419_46155# a_6347_46155# 6.64e-19
C40713 a_9569_46155# a_5066_45546# 2.22e-20
C40714 a_19900_46494# a_21137_46414# 3.02e-20
C40715 a_20075_46420# a_6945_45028# 1.64e-20
C40716 a_19553_46090# a_10809_44734# 5.04e-21
C40717 a_n4064_39072# a_n4064_37440# 0.046264f
C40718 a_15095_43370# a_15681_43442# 3.23e-21
C40719 a_n229_43646# a_n13_43084# 3.17e-20
C40720 a_14021_43940# a_21195_42852# 8.07e-21
C40721 a_n1761_44111# a_n473_42460# 0.110251f
C40722 a_648_43396# a_743_42282# 4.53e-21
C40723 a_17730_32519# a_n1630_35242# 5.92e-20
C40724 a_10341_43396# a_10149_43396# 7.68e-19
C40725 a_13667_43396# a_13943_43396# 0.00119f
C40726 a_3539_42460# a_4361_42308# 0.027414f
C40727 a_14205_43396# a_15781_43660# 9.18e-21
C40728 a_9145_43396# a_16547_43609# 2.43e-21
C40729 a_2982_43646# a_5649_42852# 0.205161f
C40730 a_n356_44636# a_18220_42308# 5.19e-19
C40731 a_n1821_43396# a_n4318_38680# 1.73e-19
C40732 a_4842_47570# DATA[2] 1.24e-19
C40733 a_n1736_43218# VDD 0.082445f
C40734 a_6171_45002# a_6125_45348# 4.58e-19
C40735 a_2382_45260# a_n2293_42834# 0.026697f
C40736 a_4558_45348# a_5009_45028# 0.013349f
C40737 a_8696_44636# a_9838_44484# 0.004732f
C40738 a_14537_43396# a_15595_45028# 5.49e-20
C40739 a_13777_45326# a_1307_43914# 3.69e-21
C40740 a_15037_45618# a_15004_44636# 5.28e-20
C40741 a_n2302_39866# a_n2956_39768# 0.037924f
C40742 a_n3420_39616# a_n2442_46660# 0.00978f
C40743 a_743_42282# a_13259_45724# 0.066992f
C40744 a_3935_42891# a_n1925_42282# 0.010366f
C40745 a_4520_42826# a_526_44458# 0.247914f
C40746 a_16137_43396# a_n357_42282# 1.09442f
C40747 a_10765_43646# a_n443_42852# 6.06e-19
C40748 a_2437_43646# a_3094_47570# 9.06e-19
C40749 a_n913_45002# a_4883_46098# 1.34e-19
C40750 a_413_45260# a_18143_47464# 4.35e-19
C40751 a_13556_45296# a_4915_47217# 0.146395f
C40752 a_3232_43370# a_12861_44030# 2.11e-21
C40753 a_1423_45028# a_584_46384# 1.63e-19
C40754 a_1307_43914# a_n1151_42308# 3.38e-20
C40755 a_16115_45572# a_n743_46660# 0.012735f
C40756 a_2711_45572# a_8270_45546# 0.063301f
C40757 a_8568_45546# a_7577_46660# 1.67e-20
C40758 a_18175_45572# a_5807_45002# 0.004334f
C40759 a_16147_45260# a_13661_43548# 0.002524f
C40760 a_17786_45822# a_13747_46662# 0.005559f
C40761 a_n356_45724# a_1609_45822# 5.07e-20
C40762 a_n23_45546# a_n443_42852# 0.039956f
C40763 a_n755_45592# a_603_45572# 4.44e-20
C40764 a_16137_43396# a_18707_42852# 0.001058f
C40765 a_12089_42308# a_13113_42826# 6.01e-19
C40766 a_5649_42852# a_5837_42852# 0.001623f
C40767 a_n97_42460# a_14456_42282# 0.067807f
C40768 a_2982_43646# a_7963_42308# 8.09e-20
C40769 a_3626_43646# a_7227_42308# 0.004361f
C40770 a_12379_42858# a_12895_43230# 0.109156f
C40771 a_20820_30879# EN_OFFSET_CAL 0.107181f
C40772 a_3422_30871# C3_N_btm 1.1e-19
C40773 a_6886_37412# CAL_N 1.24e-19
C40774 VDAC_N a_11206_38545# 0.15219f
C40775 a_8912_37509# VDAC_P 3.15325f
C40776 a_11633_42558# VDD 0.193501f
C40777 a_n237_47217# a_9313_45822# 0.063143f
C40778 a_n452_47436# a_n1435_47204# 2.2e-19
C40779 a_2063_45854# a_6545_47178# 2.04e-19
C40780 a_3381_47502# a_4791_45118# 3.29e-20
C40781 a_3785_47178# a_4700_47436# 0.090466f
C40782 a_n1151_42308# a_n443_46116# 0.099874f
C40783 a_3815_47204# a_4007_47204# 0.224415f
C40784 a_n699_43396# a_4743_44484# 0.235328f
C40785 a_4223_44672# a_5343_44458# 0.229803f
C40786 a_18479_45785# a_15493_43396# 0.235084f
C40787 a_n2661_44458# a_12607_44458# 1.59e-19
C40788 a_327_44734# a_453_43940# 8.52e-21
C40789 a_413_45260# a_2127_44172# 0.104737f
C40790 a_n2661_45010# a_n3674_39768# 0.001075f
C40791 a_2437_43646# a_2253_44260# 2.98e-19
C40792 a_n784_42308# a_n357_42282# 0.008228f
C40793 a_196_42282# a_n755_45592# 0.090568f
C40794 a_1067_42314# a_n863_45724# 0.289393f
C40795 a_4190_30871# C2_P_btm 9.13e-20
C40796 a_14209_32519# a_11530_34132# 0.004282f
C40797 a_n2129_44697# a_n2438_43548# 0.060059f
C40798 a_n2661_43370# a_7577_46660# 3.63e-21
C40799 a_15595_45028# a_3090_45724# 0.00235f
C40800 a_9482_43914# a_15227_44166# 0.020073f
C40801 a_n452_44636# a_n2293_46634# 3.66e-20
C40802 a_17767_44458# a_12549_44172# 1.63e-20
C40803 a_19479_31679# a_11415_45002# 0.224531f
C40804 a_15415_45028# a_14976_45028# 0.027906f
C40805 a_3357_43084# a_20202_43084# 0.029548f
C40806 a_21513_45002# a_12741_44636# 1.26e-19
C40807 a_2437_43646# a_20820_30879# 0.006482f
C40808 a_8162_45546# a_5066_45546# 0.025437f
C40809 a_6171_45002# a_14035_46660# 3.2e-20
C40810 a_413_45260# a_765_45546# 0.031429f
C40811 a_14033_45822# a_13925_46122# 0.001241f
C40812 a_n1655_44484# a_n1613_43370# 0.003155f
C40813 a_13857_44734# a_10227_46804# 4.26e-19
C40814 a_n2472_43914# SMPL_ON_P 3.53e-19
C40815 a_n1549_44318# a_n2497_47436# 0.018493f
C40816 a_16795_42852# a_17124_42282# 3.59e-19
C40817 a_n2840_42282# a_n2472_42282# 7.52e-19
C40818 a_5534_30871# a_4958_30871# 0.024536f
C40819 a_17701_42308# a_16104_42674# 7.22e-21
C40820 a_7309_42852# a_6123_31319# 9.07e-19
C40821 a_14097_32519# COMP_P 7e-21
C40822 a_5807_45002# a_n743_46660# 0.669712f
C40823 a_n1613_43370# a_2959_46660# 0.187029f
C40824 a_2747_46873# a_3877_44458# 8.98e-21
C40825 a_9313_45822# a_8270_45546# 0.0271f
C40826 a_4915_47217# a_13607_46688# 0.082884f
C40827 a_10227_46804# a_10150_46912# 0.236747f
C40828 a_n2017_45002# a_16409_43396# 1.12e-20
C40829 a_n913_45002# a_16243_43396# 3.59e-20
C40830 a_n1059_45260# a_16547_43609# 0.024317f
C40831 a_3232_43370# a_9803_43646# 2.81e-21
C40832 a_6171_45002# a_9145_43396# 3.37e-21
C40833 a_n2293_42834# a_n1655_43396# 3.89e-19
C40834 a_10193_42453# a_21356_42826# 1.27e-19
C40835 a_n2661_43370# a_n1177_43370# 3.12e-21
C40836 a_11967_42832# a_19789_44512# 5.08e-19
C40837 a_1307_43914# a_6197_43396# 7.34e-20
C40838 a_14539_43914# a_14955_43940# 0.064683f
C40839 a_n2661_42834# a_2889_44172# 0.005688f
C40840 a_626_44172# a_648_43396# 0.04847f
C40841 a_n2661_43922# a_2675_43914# 0.002037f
C40842 a_17517_44484# a_22591_44484# 0.196232f
C40843 a_20766_44850# a_19279_43940# 0.021466f
C40844 a_16112_44458# a_15682_43940# 0.006723f
C40845 a_5932_42308# C6_P_btm 3.73e-19
C40846 a_20205_31679# C6_N_btm 1.26e-20
C40847 a_20692_30879# C5_N_btm 3.17e-19
C40848 a_21005_45260# a_21137_46414# 1.84e-20
C40849 a_19113_45348# a_18985_46122# 6.36e-21
C40850 a_11691_44458# a_18819_46122# 2.75e-19
C40851 a_n2661_44458# a_10903_43370# 4.92e-19
C40852 a_8487_44056# a_n1613_43370# 3.38e-21
C40853 a_14401_32519# SMPL_ON_N 0.029323f
C40854 a_11967_42832# a_19466_46812# 8.14e-20
C40855 a_5244_44056# a_5257_43370# 6.32e-19
C40856 a_2455_43940# a_768_44030# 0.005192f
C40857 a_13565_44260# a_13661_43548# 3.81e-19
C40858 a_16751_45260# a_16375_45002# 0.047561f
C40859 a_3429_45260# a_3503_45724# 2.71e-19
C40860 a_n37_45144# a_n443_42852# 0.137227f
C40861 a_3537_45260# a_3316_45546# 0.078381f
C40862 a_413_45260# a_509_45822# 1.95e-19
C40863 a_10057_43914# a_3483_46348# 0.00873f
C40864 a_17591_47464# VDD 0.421992f
C40865 a_5934_30871# comp_n 1.4e-19
C40866 a_18057_42282# a_18310_42308# 0.011913f
C40867 a_5742_30871# a_1239_39587# 1.45e-19
C40868 a_17303_42282# a_19511_42282# 0.001918f
C40869 a_n743_46660# a_3699_46348# 0.010053f
C40870 a_n2661_46098# a_n1423_46090# 0.021984f
C40871 a_2959_46660# a_n2293_46098# 5.68e-21
C40872 a_2107_46812# a_1138_42852# 1.62e-19
C40873 a_3090_45724# a_15559_46634# 2.45e-20
C40874 a_14976_45028# a_15368_46634# 0.097092f
C40875 a_11735_46660# a_12156_46660# 0.086708f
C40876 a_9863_46634# a_765_45546# 3.07e-20
C40877 a_12549_44172# a_15015_46420# 7.35e-20
C40878 a_5807_45002# a_11189_46129# 0.001199f
C40879 a_n2661_46634# a_6165_46155# 2.58e-20
C40880 a_13661_43548# a_9290_44172# 0.00745f
C40881 a_11309_47204# a_2324_44458# 2.57e-20
C40882 a_6151_47436# a_13259_45724# 1.86e-20
C40883 a_n2497_47436# a_3218_45724# 2.25e-20
C40884 a_n1741_47186# a_n755_45592# 1.26e-21
C40885 a_n2109_47186# a_1848_45724# 5.91e-22
C40886 a_n971_45724# a_n452_45724# 0.03667f
C40887 a_n815_47178# a_n1099_45572# 3.58e-22
C40888 a_n746_45260# a_n863_45724# 0.664707f
C40889 a_n1925_46634# a_4419_46090# 3.01e-19
C40890 a_n2293_42834# a_1709_42852# 2.82e-20
C40891 a_175_44278# a_458_43396# 4.64e-19
C40892 a_895_43940# a_n97_42460# 0.002734f
C40893 a_14673_44172# a_9145_43396# 1.46e-19
C40894 a_15493_43396# a_14021_43940# 0.139192f
C40895 a_9313_44734# a_16759_43396# 8.78e-20
C40896 a_11827_44484# a_12379_42858# 2.49e-21
C40897 a_15367_44484# a_8685_43396# 2.8e-22
C40898 a_n967_45348# a_n1329_42308# 0.033651f
C40899 a_n1059_45260# a_n3674_37592# 1.1e-19
C40900 en_comp a_n961_42308# 6.61e-20
C40901 a_n2017_45002# a_564_42282# 0.013024f
C40902 a_1414_42308# VDD 0.657887f
C40903 a_11823_42460# a_11778_45572# 8.46e-20
C40904 a_8568_45546# a_8696_44636# 4.42e-20
C40905 a_10193_42453# a_15765_45572# 1.09e-19
C40906 C3_N_btm VREF_GND 0.67174f
C40907 C2_N_btm VCM 0.716172f
C40908 C4_N_btm VREF 0.98728f
C40909 C5_N_btm VIN_N 0.502041f
C40910 a_14021_43940# a_3483_46348# 0.066924f
C40911 a_8147_43396# a_3090_45724# 0.002892f
C40912 a_n2840_42826# a_n2438_43548# 2.22e-21
C40913 a_7765_42852# a_768_44030# 1.22e-20
C40914 a_n3674_39304# a_n2956_39768# 0.023853f
C40915 a_10807_43548# a_2324_44458# 1.65e-20
C40916 a_21195_42852# a_13507_46334# 0.005401f
C40917 a_20820_30879# a_22959_46124# 0.00389f
C40918 a_19466_46812# a_13259_45724# 5.7e-20
C40919 a_3483_46348# a_11133_46155# 0.001334f
C40920 a_12741_44636# a_10809_44734# 0.088683f
C40921 a_4185_45028# a_9290_44172# 4.71e-19
C40922 a_7920_46348# a_8016_46348# 0.318386f
C40923 a_5343_44458# a_5742_30871# 9.93e-21
C40924 a_11967_42832# a_16328_43172# 0.001925f
C40925 a_18494_42460# a_18310_42308# 0.001869f
C40926 a_n2293_43922# a_n3674_38216# 0.032717f
C40927 a_5891_43370# a_1606_42308# 5.17e-20
C40928 a_8975_43940# a_8685_42308# 1.95e-22
C40929 a_n2661_42834# a_n4318_37592# 1.57e-19
C40930 a_19319_43548# a_19268_43646# 0.17076f
C40931 a_2982_43646# a_8685_43396# 6.82e-20
C40932 a_6031_43396# a_6655_43762# 9.73e-19
C40933 a_6293_42852# a_6452_43396# 0.157972f
C40934 a_7287_43370# a_7112_43396# 0.234322f
C40935 a_10405_44172# a_10083_42826# 1.98e-19
C40936 a_3785_47178# DATA[2] 0.119025f
C40937 a_4915_47217# RST_Z 5.15e-19
C40938 a_n1151_42308# DATA[4] 8.05e-22
C40939 a_19963_31679# C3_N_btm 0.041776f
C40940 a_19479_31679# C6_N_btm 1.26e-20
C40941 a_12281_43396# VDD 0.341026f
C40942 a_8746_45002# a_n2661_44458# 0.017636f
C40943 a_8696_44636# a_n2661_43370# 0.674122f
C40944 a_2711_45572# a_15004_44636# 5.78e-22
C40945 a_413_45260# a_2382_45260# 0.048205f
C40946 a_n913_45002# a_3232_43370# 6.56e-20
C40947 a_15051_42282# a_13661_43548# 1.21e-20
C40948 a_5742_30871# a_n2956_39768# 7.02e-21
C40949 a_13569_43230# a_3090_45724# 1.94e-19
C40950 a_104_43370# a_n443_42852# 0.003607f
C40951 a_4699_43561# a_n755_45592# 2.57e-21
C40952 a_3080_42308# a_n357_42282# 0.023702f
C40953 a_3626_43646# a_n2661_45546# 0.009175f
C40954 a_3422_30871# C7_P_btm 2.94e-19
C40955 a_n1013_45572# VDD 4.04e-19
C40956 a_11823_42460# a_768_44030# 0.066425f
C40957 a_13163_45724# a_12891_46348# 0.009037f
C40958 a_12791_45546# a_12549_44172# 0.083854f
C40959 a_10053_45546# a_5807_45002# 3.59e-20
C40960 a_6598_45938# a_n1925_46634# 8.63e-21
C40961 a_6511_45714# a_n743_46660# 0.003331f
C40962 a_15903_45785# a_4883_46098# 1.41e-19
C40963 a_17786_45822# a_11599_46634# 2.55e-20
C40964 a_18341_45572# a_12861_44030# 0.026945f
C40965 a_n2293_45010# a_n746_45260# 0.023201f
C40966 a_3357_43084# a_2063_45854# 0.023045f
C40967 a_2437_43646# a_2905_45572# 0.003457f
C40968 a_18429_43548# a_17333_42852# 0.003673f
C40969 a_18525_43370# a_18083_42858# 0.016073f
C40970 a_n1853_43023# a_685_42968# 1.6e-20
C40971 a_15743_43084# a_17595_43084# 7.44e-20
C40972 a_5649_42852# a_7871_42858# 1.53e-20
C40973 a_743_42282# a_10518_42984# 2.81e-20
C40974 a_4361_42308# a_8605_42826# 3.01e-20
C40975 a_5745_43940# a_5755_42308# 5.58e-22
C40976 a_15493_43396# a_15764_42576# 1.23e-21
C40977 a_17538_32519# a_n1630_35242# 4.52e-20
C40978 a_n1076_43230# a_n967_43230# 0.007416f
C40979 a_n901_43156# a_n722_43218# 0.007399f
C40980 a_n1641_43230# a_n1533_42852# 0.057222f
C40981 a_n4318_38680# a_n1736_43218# 4.04e-20
C40982 a_12991_46634# CLK 5.91e-20
C40983 a_17609_46634# START 4.81e-19
C40984 a_n3690_38304# a_n3565_37414# 6.38e-20
C40985 a_n3420_37984# a_n4334_37440# 0.008459f
C40986 a_7754_39632# a_7754_39300# 0.296258f
C40987 a_n3674_38680# VDD 0.503323f
C40988 a_3065_45002# a_n2293_43922# 3.78e-20
C40989 a_n1059_45260# a_14673_44172# 7.92e-21
C40990 a_5111_44636# a_5708_44484# 0.002882f
C40991 a_3537_45260# a_n2661_42834# 0.097192f
C40992 a_10193_42453# a_19328_44172# 4.1e-19
C40993 a_13249_42308# a_10729_43914# 3.94e-20
C40994 a_16922_45042# a_17896_45144# 0.003722f
C40995 a_11823_42460# a_13483_43940# 0.029429f
C40996 a_n2293_42834# a_5343_44458# 0.165923f
C40997 a_n2661_43370# a_n1177_44458# 0.002135f
C40998 a_21005_45260# a_21359_45002# 0.001885f
C40999 a_20567_45036# a_11827_44484# 0.004169f
C41000 a_18911_45144# a_11691_44458# 0.013593f
C41001 a_18587_45118# a_20193_45348# 4.24e-21
C41002 a_20107_42308# a_20202_43084# 0.002968f
C41003 a_15051_42282# a_4185_45028# 4.66e-19
C41004 a_564_42282# a_526_44458# 1.5e-19
C41005 a_n3674_37592# a_n1925_42282# 0.072052f
C41006 a_9803_42558# a_9290_44172# 0.094028f
C41007 a_10533_42308# a_8953_45546# 7.15e-20
C41008 a_2711_45572# a_13759_46122# 2.27e-19
C41009 a_n2661_44458# a_4883_46098# 0.019556f
C41010 a_n998_44484# a_n1151_42308# 7.11e-19
C41011 a_10180_45724# a_3483_46348# 0.047643f
C41012 a_20107_45572# a_19692_46634# 0.001896f
C41013 a_5111_44636# a_5257_43370# 0.22597f
C41014 a_20623_45572# a_15227_44166# 0.002557f
C41015 a_2437_43646# a_12816_46660# 1.78e-20
C41016 a_20273_45572# a_19466_46812# 0.328586f
C41017 a_19700_43370# a_7174_31319# 2.53e-19
C41018 a_15743_43084# a_21887_42336# 3.74e-20
C41019 a_4190_30871# a_4958_30871# 11.510201f
C41020 a_7765_42852# a_6123_31319# 6.64e-19
C41021 a_n2293_42282# a_n4318_37592# 0.004341f
C41022 a_7871_42858# a_7963_42308# 3.99e-19
C41023 a_21259_43561# a_17303_42282# 9.51e-21
C41024 a_n914_42852# a_n4318_38216# 5.63e-21
C41025 a_14311_47204# a_n743_46660# 6.88e-21
C41026 a_18597_46090# a_19594_46812# 6.44e-19
C41027 a_19386_47436# a_19321_45002# 0.086877f
C41028 a_n1435_47204# a_33_46660# 3.84e-20
C41029 a_2063_45854# a_3877_44458# 0.024649f
C41030 a_n971_45724# a_5275_47026# 6.84e-21
C41031 a_n443_46116# a_3177_46902# 0.019328f
C41032 a_2905_45572# a_3686_47026# 1.64e-19
C41033 a_949_44458# a_2479_44172# 3.43e-19
C41034 a_n699_43396# a_1414_42308# 0.104607f
C41035 a_742_44458# a_895_43940# 0.025021f
C41036 a_10193_42453# a_20749_43396# 1.81e-19
C41037 a_1307_43914# a_8415_44056# 5.17e-19
C41038 a_n2661_43922# a_10809_44484# 1.69e-19
C41039 a_3065_45002# a_n97_42460# 0.019675f
C41040 a_n913_45002# a_4905_42826# 0.101072f
C41041 a_n2017_45002# a_n1557_42282# 0.090464f
C41042 a_n4209_38502# a_n2810_45572# 0.066112f
C41043 a_1667_45002# VDD 0.315476f
C41044 COMP_P a_22780_40945# 3.32e-19
C41045 a_20193_45348# a_11415_45002# 0.007211f
C41046 a_13711_45394# a_3483_46348# 0.002278f
C41047 a_n2472_43914# a_n2438_43548# 0.032003f
C41048 a_n809_44244# a_n2293_46634# 5.01e-20
C41049 a_18479_45785# a_n357_42282# 2.83e-19
C41050 a_3537_45260# a_5066_45546# 1.14e-19
C41051 a_2304_45348# a_2324_44458# 1.74e-19
C41052 a_7418_45394# a_5937_45572# 2.23e-19
C41053 a_15493_43396# a_13507_46334# 2.29e-20
C41054 a_20935_43940# a_18597_46090# 0.008467f
C41055 a_11341_43940# a_18479_47436# 0.009284f
C41056 a_15493_43940# a_10227_46804# 0.00594f
C41057 a_n2433_43396# SMPL_ON_P 2.87e-19
C41058 a_n1177_43370# a_n2497_47436# 0.062743f
C41059 a_5742_30871# a_12563_42308# 1.19e-20
C41060 a_2123_42473# a_7174_31319# 4.88e-21
C41061 a_n3674_37592# a_n4315_30879# 7.52e-19
C41062 a_n4318_38216# a_n4064_39616# 0.024304f
C41063 a_11551_42558# a_11633_42558# 0.171361f
C41064 a_n3674_38216# a_n3420_39616# 0.02009f
C41065 a_5342_30871# C5_N_btm 9.85e-20
C41066 a_5534_30871# C7_N_btm 0.060228f
C41067 C4_P_btm VIN_P 0.50261f
C41068 C6_P_btm VREF 1.41944f
C41069 DATA[0] DATA[1] 1.62e-19
C41070 C8_P_btm VCM 2.61094f
C41071 C7_P_btm VREF_GND 1.61142f
C41072 a_3067_47026# a_3090_45724# 1.04e-20
C41073 a_13747_46662# a_20411_46873# 3.16e-20
C41074 a_13661_43548# a_20273_46660# 5.45e-20
C41075 a_10150_46912# a_10467_46802# 0.102355f
C41076 a_7927_46660# a_6755_46942# 0.036549f
C41077 a_19321_45002# a_19551_46910# 0.009214f
C41078 a_7577_46660# a_6682_46987# 3.94e-20
C41079 a_5257_43370# a_6086_46660# 1.63e-19
C41080 a_19594_46812# a_19123_46287# 0.002216f
C41081 a_n881_46662# a_12741_44636# 7.98e-20
C41082 a_13717_47436# a_10903_43370# 0.001667f
C41083 a_13381_47204# a_12594_46348# 3.26e-21
C41084 a_n1435_47204# a_12005_46116# 9.73e-21
C41085 a_13507_46334# a_3483_46348# 1.37e-19
C41086 a_3065_45002# a_3935_43218# 5.01e-19
C41087 a_3537_45260# a_n2293_42282# 0.001815f
C41088 a_n1059_45260# a_8292_43218# 0.002071f
C41089 a_n2293_42834# a_n1545_43230# 8.56e-19
C41090 a_12607_44458# a_9145_43396# 2.06e-20
C41091 a_7499_43078# a_9293_42558# 1.64e-19
C41092 a_10193_42453# a_8685_42308# 3e-20
C41093 a_1423_45028# a_8952_43230# 6.06e-21
C41094 a_8975_43940# a_9803_43646# 8.14e-21
C41095 a_n356_44636# a_8147_43396# 6.99e-22
C41096 a_n2661_43922# a_1209_43370# 1.01e-21
C41097 a_n2661_42834# a_1049_43396# 6.94e-20
C41098 a_14539_43914# a_8685_43396# 5.25e-19
C41099 a_17517_44484# a_20974_43370# 1.2e-20
C41100 a_13556_45296# a_13460_43230# 1.23e-19
C41101 a_10057_43914# a_10695_43548# 0.148476f
C41102 a_18911_45144# a_4190_30871# 1.03e-21
C41103 a_14112_44734# VDD 0.004001f
C41104 a_n3565_38502# VREF_GND 0.001993f
C41105 a_2711_45572# a_11652_45724# 0.013232f
C41106 a_5013_44260# a_3483_46348# 0.002821f
C41107 a_3905_42865# a_4185_45028# 0.09316f
C41108 a_18525_43370# a_12549_44172# 3.14e-20
C41109 a_15493_43940# a_17339_46660# 0.020994f
C41110 a_10555_43940# a_3090_45724# 0.005028f
C41111 a_12495_44260# a_13059_46348# 2e-20
C41112 a_13749_43396# a_13661_43548# 1.53e-20
C41113 a_14955_43396# a_n2293_46634# 0.002132f
C41114 a_949_44458# a_n443_42852# 0.0015f
C41115 a_n2661_43922# a_8049_45260# 2.89e-19
C41116 a_10057_43914# a_n357_42282# 9.91e-20
C41117 a_742_44458# a_1609_45822# 2.73e-20
C41118 a_10428_46928# VDD 0.278873f
C41119 a_13258_32519# C6_N_btm 1.87e-19
C41120 a_7174_31319# C3_N_btm 3.5e-20
C41121 a_n3674_37592# a_n3420_37440# 0.073321f
C41122 a_n1630_35242# a_n3565_37414# 6.25e-19
C41123 a_n784_42308# a_n4064_37440# 0.014901f
C41124 a_n2293_46634# a_3316_45546# 0.067277f
C41125 a_n743_46660# a_n755_45592# 0.020454f
C41126 a_6969_46634# a_5066_45546# 1.41e-19
C41127 a_33_46660# a_380_45546# 1.08e-19
C41128 a_n133_46660# a_310_45028# 8.97e-20
C41129 a_171_46873# a_n1099_45572# 5.56e-21
C41130 a_7927_46660# a_8049_45260# 7.61e-20
C41131 a_n2438_43548# a_n357_42282# 0.026249f
C41132 a_14035_46660# a_10903_43370# 2e-19
C41133 a_765_45546# a_6165_46155# 6.78e-20
C41134 a_15227_44166# a_18819_46122# 0.288885f
C41135 a_15009_46634# a_6945_45028# 5.03e-20
C41136 a_13607_46688# a_10809_44734# 0.002497f
C41137 a_19466_46812# a_18189_46348# 0.001238f
C41138 a_n97_42460# a_458_43396# 0.013064f
C41139 a_11967_42832# a_15279_43071# 0.027468f
C41140 a_n4318_40392# a_n3674_37592# 0.032206f
C41141 a_19721_31679# a_n1630_35242# 1.04e-19
C41142 a_5891_43370# a_9061_43230# 7.06e-20
C41143 a_n2956_37592# a_n3690_39392# 1.91e-20
C41144 a_n2810_45028# a_n3420_39072# 6.67e-21
C41145 en_comp a_n3565_39304# 2.05e-19
C41146 a_n1190_43762# VDD 7.62e-19
C41147 a_20528_45572# a_20719_45572# 4.61e-19
C41148 a_21363_45546# a_21513_45002# 0.06363f
C41149 a_20623_45572# a_2437_43646# 2e-20
C41150 a_20107_45572# a_3357_43084# 0.308463f
C41151 a_15599_45572# a_6171_45002# 0.001026f
C41152 a_7227_45028# a_n2661_43370# 0.026158f
C41153 a_20273_45572# a_19479_31679# 4.39e-20
C41154 a_743_42282# a_20202_43084# 0.135735f
C41155 a_13113_42826# a_3090_45724# 0.003304f
C41156 a_961_42354# a_768_44030# 1.48e-21
C41157 a_5837_43172# a_5257_43370# 3.27e-20
C41158 a_n1557_42282# a_526_44458# 0.31675f
C41159 a_11341_43940# a_n443_42852# 0.51832f
C41160 a_14021_43940# a_n357_42282# 3.16e-19
C41161 a_9145_43396# a_10903_43370# 0.041756f
C41162 a_9885_43646# a_8953_45546# 0.011162f
C41163 a_14579_43548# a_9290_44172# 0.007608f
C41164 a_6765_43638# a_6945_45028# 4.3e-20
C41165 a_5742_30871# a_10227_46804# 6.15e-19
C41166 a_15803_42450# a_12861_44030# 5.43e-20
C41167 a_n3420_39616# w_1575_34946# 0.036508f
C41168 a_n4064_40160# SMPL_ON_P 2.22e-19
C41169 a_5907_45546# a_4883_46098# 2.75e-20
C41170 a_11525_45546# a_11459_47204# 1.91e-21
C41171 a_10193_42453# a_12861_44030# 1.83e-19
C41172 a_19553_46090# a_19443_46116# 0.097745f
C41173 a_10809_44734# a_16375_45002# 6.42e-20
C41174 a_16855_43396# a_16823_43084# 0.005656f
C41175 a_19268_43646# a_19095_43396# 0.032587f
C41176 a_3422_30871# a_17124_42282# 6.32e-20
C41177 a_n2661_42282# a_5267_42460# 2.34e-19
C41178 a_15743_43084# a_13467_32519# 0.02051f
C41179 a_2982_43646# a_17333_42852# 3.68e-20
C41180 a_3626_43646# a_17701_42308# 0.003224f
C41181 a_8685_43396# a_7871_42858# 0.004749f
C41182 a_18783_43370# a_4361_42308# 7.79e-21
C41183 a_17324_43396# a_5649_42852# 1.08e-21
C41184 a_n4209_37414# C1_P_btm 0.043983f
C41185 a_5907_45546# a_5663_43940# 2.08e-20
C41186 a_15599_45572# a_14673_44172# 9.73e-20
C41187 a_13348_45260# a_11691_44458# 2.44e-20
C41188 a_5009_45028# a_n2661_43370# 0.003943f
C41189 a_n2293_42834# a_8560_45348# 3.09e-20
C41190 a_3232_43370# a_n2661_44458# 0.468391f
C41191 a_2382_45260# a_2779_44458# 1.06e-19
C41192 a_n913_45002# a_8975_43940# 4.06e-21
C41193 a_3065_45002# a_742_44458# 2.17e-20
C41194 a_1184_42692# a_1138_42852# 0.00134f
C41195 a_4958_30871# a_15227_44166# 1.39e-20
C41196 a_n1076_43230# a_n443_42852# 0.003517f
C41197 a_1847_42826# a_n755_45592# 0.053279f
C41198 a_8483_43230# a_526_44458# 0.004236f
C41199 a_17538_32519# a_11530_34132# 0.002953f
C41200 a_n4064_37440# SMPL_ON_P 6.21e-20
C41201 a_2437_43646# a_2443_46660# 3.88e-20
C41202 a_n37_45144# a_n2661_46634# 2.93e-21
C41203 a_5111_44636# a_5807_45002# 0.204193f
C41204 a_n955_45028# a_n2293_46634# 4.55e-21
C41205 a_13556_45296# a_n881_46662# 4.04e-20
C41206 a_n2433_44484# SMPL_ON_P 2.73e-19
C41207 a_n1177_44458# a_n2497_47436# 1.74e-19
C41208 a_22469_39537# VDD 0.356405f
C41209 a_743_42282# a_n327_42308# 5.05e-21
C41210 a_14358_43442# a_14113_42308# 7.16e-21
C41211 a_n1991_42858# COMP_P 1.96e-19
C41212 a_n1641_43230# a_n1736_42282# 3.46e-19
C41213 a_12281_43396# a_11551_42558# 0.007065f
C41214 a_14579_43548# a_15051_42282# 0.002402f
C41215 a_n4318_39304# a_n4064_39072# 0.017224f
C41216 a_n4318_38680# a_n3674_38680# 3.04229f
C41217 a_13467_32519# a_1606_42308# 0.002946f
C41218 a_12895_43230# a_12800_43218# 0.049827f
C41219 a_13113_42826# a_12991_43230# 3.16e-19
C41220 a_12379_42858# a_13569_43230# 2.56e-19
C41221 a_10809_44734# RST_Z 0.00392f
C41222 a_6945_45028# SINGLE_ENDED 0.021393f
C41223 a_n2860_39866# VDD 0.004232f
C41224 a_n1151_42308# a_n1613_43370# 1.19311f
C41225 a_16327_47482# a_18479_47436# 0.723416f
C41226 a_13717_47436# a_4883_46098# 2.67e-19
C41227 a_13487_47204# a_13507_46334# 1.68e-19
C41228 a_16763_47508# a_10227_46804# 0.070681f
C41229 a_16588_47582# a_17591_47464# 0.001438f
C41230 a_3160_47472# a_n881_46662# 0.070909f
C41231 a_2063_45854# a_8128_46384# 0.032153f
C41232 a_n2293_45010# a_726_44056# 8.78e-19
C41233 a_8746_45002# a_9145_43396# 1.83e-20
C41234 a_n356_44636# a_7_44811# 0.005265f
C41235 a_18184_42460# a_18579_44172# 0.161593f
C41236 a_2711_45572# a_16759_43396# 6.88e-21
C41237 a_10180_45724# a_10695_43548# 1.07e-21
C41238 a_n2293_42834# a_453_43940# 1.92e-20
C41239 a_18114_32519# a_17517_44484# 0.055077f
C41240 a_11827_44484# a_20679_44626# 0.030022f
C41241 a_11691_44458# a_19615_44636# 0.001633f
C41242 a_20193_45348# a_11967_42832# 0.01602f
C41243 a_13720_44458# a_9313_44734# 1.1e-21
C41244 a_8103_44636# a_n2661_43922# 0.008682f
C41245 a_21359_45002# a_20835_44721# 2.3e-19
C41246 a_21101_45002# a_20766_44850# 0.01337f
C41247 a_21005_45260# a_19279_43940# 4.39e-21
C41248 a_11787_45002# a_10729_43914# 3.79e-21
C41249 a_10951_45334# a_10949_43914# 8.94e-19
C41250 a_10775_45002# a_10807_43548# 1.41e-19
C41251 a_15764_42576# a_n357_42282# 8.52e-20
C41252 a_13258_32519# a_13259_45724# 0.037974f
C41253 a_n4064_38528# a_n2956_39304# 0.001421f
C41254 a_n2946_38778# a_n2956_38680# 0.14863f
C41255 a_5342_30871# C5_P_btm 9.85e-20
C41256 a_5534_30871# C3_P_btm 7.69e-20
C41257 a_4574_45260# a_4704_46090# 1.1e-20
C41258 a_2437_43646# a_18819_46122# 2.62e-20
C41259 a_3537_45260# a_5068_46348# 1.38e-20
C41260 a_n1059_45260# a_10903_43370# 0.028694f
C41261 a_3357_43084# a_17715_44484# 9.87e-21
C41262 a_2537_44260# a_n443_46116# 5.68e-19
C41263 a_7584_44260# a_n1151_42308# 9.64e-20
C41264 a_4558_45348# a_4419_46090# 0.00116f
C41265 a_1307_43914# a_12741_44636# 0.05146f
C41266 a_4927_45028# a_3483_46348# 0.032156f
C41267 a_18911_45144# a_15227_44166# 3.32e-20
C41268 a_n2661_43922# a_n2442_46660# 1.33e-20
C41269 a_5147_45002# a_4185_45028# 5.45e-19
C41270 a_18315_45260# a_19466_46812# 9.44e-20
C41271 a_n2661_42834# a_n2293_46634# 0.025484f
C41272 a_17478_45572# a_8049_45260# 0.010438f
C41273 a_3823_42558# a_3581_42558# 3.68e-20
C41274 a_1755_42282# a_6481_42558# 0.012532f
C41275 a_5534_30871# a_n4064_38528# 0.057361f
C41276 a_5342_30871# a_n3420_38528# 0.028503f
C41277 a_2123_42473# a_5932_42308# 4.34e-21
C41278 a_n784_42308# a_8685_42308# 1.58e-20
C41279 a_1576_42282# a_5934_30871# 2.52e-20
C41280 a_961_42354# a_6123_31319# 1.52e-20
C41281 a_13467_32519# C1_N_btm 0.031032f
C41282 a_4190_30871# C7_N_btm 2.94e-19
C41283 a_22521_39511# CAL_P 0.027034f
C41284 a_22521_40055# a_22609_37990# 0.234448f
C41285 a_22459_39145# a_22705_38406# 6.64e-21
C41286 a_22545_38993# a_22876_39857# 4.42e-19
C41287 a_3080_42308# a_n4064_37440# 1.61e-19
C41288 a_n2661_46634# a_8492_46660# 0.009944f
C41289 a_n1925_46634# a_7411_46660# 0.047823f
C41290 a_2107_46812# a_5907_46634# 0.003718f
C41291 a_5807_45002# a_6086_46660# 1.02e-19
C41292 a_11309_47204# a_11186_47026# 0.004771f
C41293 a_n881_46662# a_13607_46688# 2.29e-20
C41294 a_4883_46098# a_14035_46660# 0.019262f
C41295 a_13507_46334# a_14513_46634# 9.96e-20
C41296 a_18597_46090# a_16388_46812# 0.011997f
C41297 a_16023_47582# a_765_45546# 0.006051f
C41298 a_16327_47482# a_17829_46910# 7.11e-21
C41299 a_10227_46804# a_14226_46660# 4.83e-20
C41300 a_11599_46634# a_20411_46873# 0.00162f
C41301 a_13717_47436# a_21188_46660# 2.12e-21
C41302 a_n2109_47186# a_4185_45028# 1.33e-19
C41303 a_n971_45724# a_167_45260# 1.89e-19
C41304 a_n1151_42308# a_n2293_46098# 0.040266f
C41305 a_n237_47217# a_1823_45246# 0.370766f
C41306 a_584_46384# a_n901_46420# 3.34e-19
C41307 a_n1741_47186# a_3483_46348# 4.84e-20
C41308 a_742_44458# a_458_43396# 4.92e-20
C41309 a_6298_44484# a_n97_42460# 5.4e-19
C41310 a_1467_44172# a_1414_42308# 0.335735f
C41311 a_n984_44318# a_895_43940# 2.65e-20
C41312 a_1115_44172# a_453_43940# 0.150214f
C41313 a_17517_44484# a_17737_43940# 9.06e-20
C41314 a_18248_44752# a_19319_43548# 1.93e-20
C41315 a_14815_43914# a_15493_43940# 8.51e-20
C41316 a_14537_43396# a_16823_43084# 9.22e-21
C41317 a_n2661_42834# a_11816_44260# 1.53e-19
C41318 a_n913_45002# a_2905_42968# 0.009485f
C41319 a_n1059_45260# a_3681_42891# 0.003573f
C41320 a_n2017_45002# a_3935_42891# 4.3e-21
C41321 a_8912_37509# VDD 18.3523f
C41322 a_n699_43396# VDD 0.922998f
C41323 a_7174_31319# C7_P_btm 9.97e-20
C41324 a_n4064_40160# a_n1532_35090# 6.3e-20
C41325 a_n4064_37984# a_n2956_38216# 0.054267f
C41326 a_n3607_38304# a_n2810_45572# 5.7e-20
C41327 a_18579_44172# a_12741_44636# 0.002357f
C41328 a_20596_44850# a_11415_45002# 8.83e-20
C41329 a_n2433_43396# a_n2438_43548# 0.415301f
C41330 a_2982_43646# a_768_44030# 0.0012f
C41331 a_n2661_42282# a_3090_45724# 0.039366f
C41332 a_n2661_43370# a_2957_45546# 3.26e-20
C41333 a_20193_45348# a_13259_45724# 0.014145f
C41334 a_18494_42460# a_20254_46482# 2.45e-20
C41335 a_n2661_43922# a_8953_45546# 0.024071f
C41336 a_6197_43396# a_n1613_43370# 0.03252f
C41337 a_8685_43396# a_11453_44696# 9.12e-22
C41338 a_9145_43396# a_4883_46098# 0.02956f
C41339 a_10341_43396# a_18479_47436# 1.96e-19
C41340 a_16137_43396# a_12861_44030# 3.28e-19
C41341 a_n1991_42858# a_n2497_47436# 9.6e-20
C41342 a_743_42282# a_2063_45854# 1.93e-20
C41343 a_n4209_39590# a_n4334_39392# 3.3e-19
C41344 a_n4334_39616# a_n4209_39304# 3.3e-19
C41345 a_n4315_30879# a_n2302_39072# 6.48e-20
C41346 a_n2302_39866# a_n2216_39866# 0.011479f
C41347 a_n3690_39616# a_n3607_39616# 0.007692f
C41348 a_n4064_40160# a_n2946_39072# 2.04e-20
C41349 a_n3420_39616# a_n4251_39616# 0.0016f
C41350 a_22612_30879# VDD 3.2377f
C41351 a_5934_30871# C1_P_btm 0.011025f
C41352 a_6123_31319# C0_dummy_P_btm 1.31e-19
C41353 a_5932_42308# C3_N_btm 0.121156f
C41354 a_17609_46634# a_12741_44636# 5.71e-21
C41355 a_15227_44166# a_22591_46660# 1.6e-20
C41356 a_19466_46812# a_20202_43084# 2.86e-21
C41357 a_16388_46812# a_19123_46287# 4.8e-20
C41358 a_16434_46987# a_17829_46910# 4.36e-20
C41359 a_16721_46634# a_18285_46348# 2.92e-20
C41360 a_16751_46987# a_765_45546# 1.47e-19
C41361 a_n2661_46098# a_n2956_39304# 0.008823f
C41362 a_19594_46812# a_8049_45260# 9.33e-20
C41363 a_n743_46660# a_835_46155# 4.14e-19
C41364 a_2107_46812# a_739_46482# 5.16e-20
C41365 a_n881_46662# a_16375_45002# 2.62e-19
C41366 a_8667_46634# a_5937_45572# 0.001106f
C41367 a_8492_46660# a_8199_44636# 2.51e-19
C41368 a_16327_47482# a_n443_42852# 2.73e-21
C41369 a_13507_46334# a_n357_42282# 0.001222f
C41370 a_n2312_39304# a_n2810_45572# 0.044713f
C41371 a_n2312_40392# a_n2661_45546# 7.42e-20
C41372 en_comp a_14113_42308# 3.72e-20
C41373 a_n913_45002# a_15803_42450# 8.35e-19
C41374 a_n2017_45002# a_15890_42674# 0.00307f
C41375 a_5111_44636# a_9223_42460# 1.34e-20
C41376 a_n1059_45260# a_15959_42545# 0.002635f
C41377 a_n2661_42282# a_6547_43396# 0.00581f
C41378 a_742_44458# a_2987_42968# 7.44e-19
C41379 a_1307_43914# a_2903_42308# 6.88e-22
C41380 a_14539_43914# a_17333_42852# 0.072085f
C41381 a_n356_44636# a_13113_42826# 5.02e-21
C41382 a_n2293_42834# a_n2472_42282# 0.002489f
C41383 a_22315_44484# a_15743_43084# 2.11e-21
C41384 a_19615_44636# a_4190_30871# 1.28e-21
C41385 a_5891_43370# a_8605_42826# 0.0011f
C41386 a_8375_44464# a_8387_43230# 6.17e-22
C41387 a_22959_43948# VDD 0.297936f
C41388 a_16115_45572# a_16147_45260# 6.95e-19
C41389 a_8696_44636# a_16211_45572# 2.41e-20
C41390 a_5907_45546# a_3232_43370# 0.001196f
C41391 a_6194_45824# a_5691_45260# 1.08e-19
C41392 a_3775_45552# a_3537_45260# 1.46e-19
C41393 a_2711_45572# a_7276_45260# 0.00282f
C41394 a_10193_42453# a_n913_45002# 0.562004f
C41395 a_7499_43078# en_comp 8.68e-21
C41396 a_n97_42460# a_5937_45572# 1.46e-20
C41397 a_18707_42852# a_13507_46334# 6.67e-19
C41398 a_2903_42308# a_n443_46116# 7.96e-21
C41399 a_3318_42354# a_4791_45118# 2.33e-20
C41400 a_4699_43561# a_3483_46348# 2.57e-21
C41401 a_4093_43548# a_4185_45028# 4.24e-20
C41402 a_1987_43646# a_1823_45246# 2.6e-20
C41403 a_8952_43230# a_4646_46812# 3.88e-21
C41404 a_n2293_42282# a_n2293_46634# 7.31e-22
C41405 a_14621_43646# a_13059_46348# 2.44e-20
C41406 a_16823_43084# a_3090_45724# 7.78e-20
C41407 a_2675_43914# a_3316_45546# 4.27e-20
C41408 a_175_44278# a_n443_42852# 0.003303f
C41409 a_5013_44260# a_n357_42282# 2.45e-20
C41410 a_n3674_39768# a_n2956_38216# 0.031697f
C41411 CAL_N a_22521_39511# 0.023597f
C41412 a_22469_40625# a_22459_39145# 0.245891f
C41413 a_n3420_37440# EN_VIN_BSTR_P 0.040234f
C41414 a_22959_45036# RST_Z 0.001356f
C41415 a_18114_32519# EN_VIN_BSTR_N 0.187697f
C41416 a_7920_46348# VDD 0.100184f
C41417 a_1609_45572# a_n237_47217# 2.16e-20
C41418 a_6472_45840# a_n1741_47186# 9.06e-21
C41419 a_2112_39137# a_3754_38470# 2.65e-20
C41420 a_3483_46348# a_10586_45546# 0.099824f
C41421 a_20202_43084# a_20205_31679# 1.27e-19
C41422 a_765_45546# a_n23_45546# 8.66e-20
C41423 a_22365_46825# a_20692_30879# 7.03e-19
C41424 a_9625_46129# a_5066_45546# 1.5e-20
C41425 a_19900_46494# a_20708_46348# 2.56e-19
C41426 a_19335_46494# a_6945_45028# 1.78e-20
C41427 a_18985_46122# a_10809_44734# 9.49e-20
C41428 a_14205_43396# a_15681_43442# 3.24e-20
C41429 a_9145_43396# a_16243_43396# 2.75e-21
C41430 a_2982_43646# a_13678_32519# 2.63e-21
C41431 a_14021_43940# a_21356_42826# 6.95e-20
C41432 a_n1761_44111# a_n961_42308# 0.002207f
C41433 a_3626_43646# a_4361_42308# 5.20633f
C41434 a_12293_43646# a_12281_43396# 0.01129f
C41435 a_13667_43396# a_13837_43396# 0.001675f
C41436 a_n356_44636# a_18214_42558# 5.42e-19
C41437 a_10341_43396# a_9885_43396# 9.63e-20
C41438 a_n1331_43914# COMP_P 5.76e-20
C41439 a_n881_46662# RST_Z 0.351994f
C41440 a_22612_30879# a_22469_39537# 1.3e-19
C41441 a_n4318_38680# VDD 0.417422f
C41442 a_6171_45002# a_5837_45348# 9.51e-21
C41443 a_21513_45002# a_19778_44110# 1.82e-19
C41444 a_3232_43370# a_6125_45348# 0.001449f
C41445 a_n967_45348# a_n2661_43370# 0.016831f
C41446 a_3537_45260# a_5093_45028# 0.009279f
C41447 a_7499_43078# a_10617_44484# 5.41e-19
C41448 a_13556_45296# a_1307_43914# 0.007672f
C41449 a_8696_44636# a_5883_43914# 0.004598f
C41450 a_14537_43396# a_15415_45028# 4.17e-20
C41451 a_20273_45572# a_20193_45348# 5.61e-19
C41452 a_4649_42852# a_1823_45246# 0.042816f
C41453 a_n4064_39616# a_n2956_39768# 0.058734f
C41454 a_n4209_39590# a_n2312_38680# 0.020921f
C41455 a_n3690_39616# a_n2442_46660# 5.77e-19
C41456 a_5934_30871# a_8270_45546# 2.28e-21
C41457 a_10341_43396# a_n443_42852# 0.23026f
C41458 a_3935_42891# a_526_44458# 0.012937f
C41459 a_3681_42891# a_n1925_42282# 9.76e-21
C41460 a_n1059_45260# a_4883_46098# 0.001764f
C41461 a_413_45260# a_10227_46804# 3.82e-19
C41462 a_9482_43914# a_4915_47217# 0.269756f
C41463 a_16333_45814# a_n743_46660# 0.014466f
C41464 a_8162_45546# a_7577_46660# 5.56e-21
C41465 a_16147_45260# a_5807_45002# 3.67e-19
C41466 a_n356_45724# a_n443_42852# 0.056063f
C41467 a_n755_45592# a_509_45572# 1.66e-20
C41468 a_n357_42282# a_603_45572# 7.72e-19
C41469 a_15743_43084# a_18695_43230# 5.34e-19
C41470 a_5649_42852# a_5193_42852# 0.003625f
C41471 a_n97_42460# a_13575_42558# 0.179828f
C41472 a_2982_43646# a_6123_31319# 0.163265f
C41473 a_3626_43646# a_6761_42308# 0.006571f
C41474 a_12379_42858# a_13113_42826# 0.06628f
C41475 a_12089_42308# a_12545_42858# 0.261463f
C41476 a_16759_43396# a_16877_42852# 6.34e-20
C41477 a_11415_45002# CLK 6.94e-20
C41478 a_22591_46660# EN_OFFSET_CAL 0.047938f
C41479 a_3422_30871# C2_N_btm 9.13e-20
C41480 VDAC_N VDAC_P 4.74149f
C41481 a_11551_42558# VDD 0.192086f
C41482 a_n815_47178# a_n1435_47204# 0.003452f
C41483 a_2063_45854# a_6151_47436# 0.448977f
C41484 a_2905_45572# a_4915_47217# 0.001556f
C41485 a_n1741_47186# a_13487_47204# 1.17e-19
C41486 a_n1151_42308# a_4791_45118# 1.16458f
C41487 a_3785_47178# a_4007_47204# 0.106797f
C41488 a_3160_47472# a_n443_46116# 0.018382f
C41489 a_4223_44672# a_4743_44484# 0.043867f
C41490 a_18479_45785# a_19328_44172# 0.003851f
C41491 a_n2661_44458# a_8975_43940# 0.075732f
C41492 a_20193_45348# a_18989_43940# 4.63e-22
C41493 a_413_45260# a_453_43940# 5.59e-20
C41494 a_n913_45002# a_5495_43940# 4.51e-22
C41495 a_n2840_45002# a_n3674_39768# 0.00158f
C41496 a_n1630_35242# a_n863_45724# 3.34e-20
C41497 a_196_42282# a_n357_42282# 0.033292f
C41498 a_n473_42460# a_n755_45592# 0.061354f
C41499 a_5024_45822# VDD 0.004293f
C41500 a_4190_30871# C3_P_btm 1.1e-19
C41501 a_13887_32519# EN_VIN_BSTR_N 0.031746f
C41502 a_n2433_44484# a_n2438_43548# 0.421822f
C41503 a_n2661_43370# a_7715_46873# 3.07e-20
C41504 a_22223_45572# a_11415_45002# 0.021019f
C41505 a_14797_45144# a_14976_45028# 0.137651f
C41506 a_15415_45028# a_3090_45724# 0.009288f
C41507 a_n1352_44484# a_n2293_46634# 2.08e-20
C41508 a_16979_44734# a_12549_44172# 1.34e-19
C41509 a_2437_43646# a_22591_46660# 7.95e-19
C41510 a_19479_31679# a_20202_43084# 9.39e-20
C41511 a_14033_45822# a_13759_46122# 1.75e-20
C41512 a_10544_45572# a_2324_44458# 2.77e-19
C41513 a_n1821_44484# a_n1613_43370# 9.54e-19
C41514 a_13468_44734# a_10227_46804# 7.33e-20
C41515 a_n2840_43914# SMPL_ON_P 9.38e-19
C41516 a_n1331_43914# a_n2497_47436# 0.003514f
C41517 a_n2840_42282# a_n3674_38680# 0.154001f
C41518 a_7309_42852# a_7227_42308# 4.85e-19
C41519 a_22400_42852# COMP_P 0.614467f
C41520 a_4190_30871# a_n4064_38528# 0.031783f
C41521 a_5342_30871# a_15761_42308# 1e-19
C41522 a_768_44030# a_2107_46812# 0.087742f
C41523 a_n881_46662# a_2609_46660# 1.09e-19
C41524 a_n1613_43370# a_3177_46902# 0.209276f
C41525 a_4915_47217# a_12816_46660# 0.006808f
C41526 a_15673_47210# a_6755_46942# 1.86e-19
C41527 a_10227_46804# a_9863_46634# 0.278164f
C41528 a_n913_45002# a_16137_43396# 3.32e-19
C41529 a_n2017_45002# a_16547_43609# 8.08e-20
C41530 a_n1059_45260# a_16243_43396# 0.012252f
C41531 a_3232_43370# a_9145_43396# 1.89e-19
C41532 a_n2293_42834# a_n1821_43396# 7.71e-19
C41533 a_n356_44636# a_n2661_42282# 2.54767f
C41534 a_14539_43914# a_13483_43940# 8.72e-20
C41535 a_11967_42832# a_20596_44850# 2.49e-19
C41536 a_10193_42453# a_20922_43172# 0.059157f
C41537 a_16922_45042# a_19319_43548# 1.84e-20
C41538 a_1307_43914# a_6293_42852# 2.54e-19
C41539 a_n2661_43370# a_n1917_43396# 3.88e-20
C41540 a_n2661_42834# a_2675_43914# 0.024352f
C41541 a_n2661_43922# a_895_43940# 0.002919f
C41542 a_17517_44484# a_22485_44484# 0.110643f
C41543 a_20835_44721# a_19279_43940# 0.036128f
C41544 a_20362_44736# a_18579_44172# 6.86e-20
C41545 a_20205_31679# C5_N_btm 0.00105f
C41546 a_20692_30879# C4_N_btm 5.85e-20
C41547 a_5932_42308# C7_P_btm 0.003981f
C41548 a_1606_42308# VCM 0.152876f
C41549 a_3065_45002# a_3503_45724# 9.76e-20
C41550 a_n143_45144# a_n443_42852# 0.104427f
C41551 a_3429_45260# a_3316_45546# 0.142842f
C41552 a_5111_44636# a_n755_45592# 0.004145f
C41553 a_19113_45348# a_18819_46122# 5.65e-21
C41554 a_21005_45260# a_20708_46348# 1.01e-20
C41555 a_n2661_44458# a_11387_46155# 4.75e-21
C41556 a_8415_44056# a_n1613_43370# 4.2e-21
C41557 a_3457_43396# a_584_46384# 0.120485f
C41558 a_6197_43396# a_4791_45118# 1.47e-19
C41559 a_2253_43940# a_768_44030# 0.004046f
C41560 a_19279_43940# a_3090_45724# 0.046663f
C41561 a_3905_42865# a_5257_43370# 0.106385f
C41562 a_n2293_42834# a_8034_45724# 0.00209f
C41563 a_1307_43914# a_16375_45002# 0.101951f
C41564 a_16588_47582# VDD 0.282243f
C41565 a_18727_42674# a_18214_42558# 0.035505f
C41566 a_18057_42282# a_18220_42308# 0.01135f
C41567 a_5934_30871# a_1736_39043# 5.23e-20
C41568 a_17124_42282# a_7174_31319# 5.22e-20
C41569 a_18907_42674# a_19332_42282# 0.017308f
C41570 a_5534_30871# a_7754_40130# 0.002632f
C41571 a_n1925_46634# a_4185_45028# 2.83e-19
C41572 a_n743_46660# a_3483_46348# 0.050648f
C41573 a_n2661_46098# a_n1991_46122# 0.025798f
C41574 a_1123_46634# a_1823_45246# 1.41e-19
C41575 a_948_46660# a_1138_42852# 4.64e-20
C41576 a_2107_46812# a_1176_45822# 1.38e-19
C41577 a_15009_46634# a_15559_46634# 4.99e-19
C41578 a_3090_45724# a_15368_46634# 0.440843f
C41579 a_6755_46942# a_16388_46812# 0.002525f
C41580 a_12549_44172# a_14275_46494# 4.53e-20
C41581 a_5807_45002# a_9290_44172# 0.00233f
C41582 a_n2661_46634# a_5497_46414# 2.47e-20
C41583 a_4883_46098# a_n1925_42282# 5.4e-19
C41584 a_n2497_47436# a_2957_45546# 2.23e-21
C41585 a_n237_47217# a_n2293_45546# 0.002405f
C41586 a_n2109_47186# a_997_45618# 4.13e-22
C41587 a_n971_45724# a_n863_45724# 0.199707f
C41588 a_327_47204# a_n2661_45546# 5.19e-21
C41589 a_n746_45260# a_n1079_45724# 9.3e-19
C41590 a_2479_44172# a_n97_42460# 0.196935f
C41591 a_19328_44172# a_14021_43940# 1.77e-20
C41592 a_9313_44734# a_16977_43638# 1.9e-20
C41593 a_n2661_44458# a_2905_42968# 1.46e-21
C41594 a_n356_44636# a_16823_43084# 0.003531f
C41595 a_n913_45002# a_n784_42308# 0.005856f
C41596 a_n1059_45260# a_n327_42558# 6.01e-20
C41597 en_comp a_n1329_42308# 5.94e-20
C41598 a_n967_45348# COMP_P 0.00202f
C41599 a_n2017_45002# a_n3674_37592# 0.241068f
C41600 a_n2293_45010# a_n1630_35242# 1.46e-20
C41601 a_1467_44172# VDD 0.391994f
C41602 a_10193_42453# a_15903_45785# 2.18e-20
C41603 a_11823_42460# a_11688_45572# 8.92e-20
C41604 a_11962_45724# a_12016_45572# 0.002378f
C41605 C2_N_btm VREF_GND 0.671742f
C41606 C1_N_btm VCM 0.716121f
C41607 C3_N_btm VREF 0.984942f
C41608 C4_N_btm VIN_N 0.50261f
C41609 a_13829_44260# a_3483_46348# 0.002792f
C41610 a_1443_43940# a_1138_42852# 7.84e-21
C41611 a_7112_43396# a_3090_45724# 0.004584f
C41612 a_7871_42858# a_768_44030# 8.9e-21
C41613 a_n2293_43922# a_n443_42852# 0.021367f
C41614 a_n2661_43922# a_1609_45822# 7.32e-20
C41615 a_21356_42826# a_13507_46334# 1.5e-19
C41616 a_5742_30871# VDAC_P 0.030356f
C41617 a_17609_46634# a_16375_45002# 2.49e-19
C41618 a_20820_30879# a_10809_44734# 0.234047f
C41619 a_3483_46348# a_11189_46129# 0.001012f
C41620 a_12741_44636# a_22223_46124# 1.14e-19
C41621 a_5204_45822# a_5937_45572# 2.47e-19
C41622 a_6419_46155# a_8016_46348# 1.19e-20
C41623 a_11967_42832# a_15785_43172# 0.003242f
C41624 a_18494_42460# a_18220_42308# 7.47e-19
C41625 a_6547_43396# a_7112_43396# 7.99e-20
C41626 a_n2661_42834# a_n1736_42282# 6.4e-21
C41627 a_n2293_43922# a_n2104_42282# 0.009285f
C41628 a_9672_43914# a_10083_42826# 8.52e-20
C41629 a_19319_43548# a_15743_43084# 0.035611f
C41630 a_18533_43940# a_18783_43370# 0.00197f
C41631 a_6031_43396# a_6452_43396# 0.086708f
C41632 a_3381_47502# DATA[2] 1.73e-19
C41633 a_n1151_42308# DATA[3] 5.14e-19
C41634 a_19479_31679# C5_N_btm 1.11e-20
C41635 a_12293_43646# VDD 0.005635f
C41636 a_10193_42453# a_n2661_44458# 3e-19
C41637 a_2711_45572# a_13720_44458# 0.001214f
C41638 a_413_45260# a_2274_45254# 0.002353f
C41639 a_n1059_45260# a_3232_43370# 1.26e-19
C41640 a_743_42282# a_17715_44484# 1.09e-20
C41641 a_13635_43156# a_12741_44636# 1.35e-21
C41642 a_5534_30871# a_11415_45002# 4.51e-21
C41643 a_n97_42460# a_n443_42852# 0.822111f
C41644 a_4235_43370# a_n755_45592# 6.26e-21
C41645 a_4699_43561# a_n357_42282# 1.83e-20
C41646 a_1427_43646# a_n863_45724# 0.006268f
C41647 a_3422_30871# C8_P_btm 4.06e-19
C41648 a_7_45899# VDD 0.001958f
C41649 a_11823_42460# a_12549_44172# 0.624462f
C41650 a_12427_45724# a_768_44030# 1.64e-22
C41651 a_9049_44484# a_5807_45002# 8.47e-20
C41652 a_6667_45809# a_n1925_46634# 1.11e-20
C41653 a_6472_45840# a_n743_46660# 0.006296f
C41654 a_12791_45546# a_12891_46348# 0.012918f
C41655 a_6977_45572# a_n1613_43370# 0.001505f
C41656 a_18479_45785# a_12861_44030# 0.058482f
C41657 a_n913_45002# SMPL_ON_P 1.07e-20
C41658 a_n967_45348# a_n2497_47436# 0.021003f
C41659 a_3357_43084# a_584_46384# 0.060446f
C41660 a_n2472_45002# a_n746_45260# 9.92e-21
C41661 a_n2293_45010# a_n971_45724# 0.549225f
C41662 a_2437_43646# a_2952_47436# 0.007981f
C41663 a_16375_45002# a_19443_46116# 4.21e-20
C41664 a_18429_43548# a_18083_42858# 1.96e-19
C41665 a_n1423_42826# a_n1533_42852# 0.097745f
C41666 a_4361_42308# a_8037_42858# 1.08e-19
C41667 a_743_42282# a_10083_42826# 2.64e-19
C41668 a_10555_44260# a_10533_42308# 3.68e-22
C41669 a_15493_43396# a_15486_42560# 2.06e-19
C41670 a_n3674_39304# a_n1736_43218# 3.4e-21
C41671 a_15743_43084# a_16795_42852# 5.64e-20
C41672 VDAC_Pi a_3754_39134# 0.012307f
C41673 a_2113_38308# VDAC_Ni 0.315941f
C41674 a_n3420_37984# a_n4209_37414# 0.03f
C41675 a_n2840_42282# VDD 0.294987f
C41676 a_5111_44636# a_5608_44484# 0.002582f
C41677 a_n2017_45002# a_14673_44172# 8.16e-21
C41678 a_5147_45002# a_5708_44484# 0.055267f
C41679 a_8953_45002# a_5891_43370# 4.12e-19
C41680 a_3065_45002# a_n2661_43922# 0.023551f
C41681 a_n2661_43370# a_n1917_44484# 0.002293f
C41682 a_17023_45118# a_16981_45144# 7.47e-21
C41683 a_16922_45042# a_17801_45144# 0.005123f
C41684 a_10193_42453# a_18451_43940# 0.20167f
C41685 a_n2293_42834# a_4743_44484# 7.24e-21
C41686 a_18494_42460# a_11827_44484# 0.031498f
C41687 a_18911_45144# a_19113_45348# 0.054737f
C41688 a_21005_45260# a_21101_45002# 0.419086f
C41689 a_18587_45118# a_11691_44458# 3.11e-20
C41690 a_11823_42460# a_12429_44172# 0.018664f
C41691 a_13258_32519# a_20202_43084# 0.685083f
C41692 a_15486_42560# a_3483_46348# 6.47e-22
C41693 a_14113_42308# a_4185_45028# 1.2e-19
C41694 a_6101_43172# a_n357_42282# 0.001097f
C41695 a_9223_42460# a_9290_44172# 2.46e-19
C41696 a_10545_42558# a_8953_45546# 2.8e-20
C41697 CAL_N a_16327_47482# 0.001106f
C41698 a_2711_45572# a_13351_46090# 6.51e-20
C41699 a_5437_45600# a_5204_45822# 5.76e-19
C41700 a_18545_45144# a_11453_44696# 2.11e-20
C41701 a_n1243_44484# a_n1151_42308# 1.58e-19
C41702 a_9313_44734# a_n971_45724# 2.29e-20
C41703 a_10053_45546# a_3483_46348# 0.002243f
C41704 a_7499_43078# a_4185_45028# 2.72e-19
C41705 a_20107_45572# a_19466_46812# 0.283769f
C41706 a_14309_45028# a_768_44030# 3.22e-19
C41707 a_5147_45002# a_5257_43370# 0.836149f
C41708 a_20841_45814# a_15227_44166# 3.03e-19
C41709 a_413_45260# a_10467_46802# 1.23e-20
C41710 a_2437_43646# a_12991_46634# 9.73e-20
C41711 a_3357_43084# a_11901_46660# 5.71e-20
C41712 a_5111_44636# a_5429_46660# 5.34e-20
C41713 a_4361_42308# a_13921_42308# 3.34e-19
C41714 a_15743_43084# a_21335_42336# 3.06e-20
C41715 a_n2293_42282# a_n1736_42282# 4.89e-19
C41716 a_7871_42858# a_6123_31319# 0.010286f
C41717 a_11453_44696# a_768_44030# 0.031665f
C41718 a_10227_46804# a_20916_46384# 0.013668f
C41719 a_18597_46090# a_19321_45002# 0.024487f
C41720 a_19787_47423# a_13747_46662# 1.81e-19
C41721 a_19386_47436# a_19452_47524# 0.006978f
C41722 a_18479_47436# a_20843_47204# 0.021416f
C41723 a_18780_47178# a_19594_46812# 2.12e-19
C41724 a_n1435_47204# a_171_46873# 5.97e-20
C41725 a_9067_47204# a_2107_46812# 1.22e-20
C41726 a_13487_47204# a_n743_46660# 2.02e-20
C41727 a_n2109_47186# a_5257_43370# 0.153164f
C41728 a_n971_45724# a_5072_46660# 4.58e-21
C41729 a_n443_46116# a_2609_46660# 0.349838f
C41730 a_3815_47204# a_3524_46660# 1.6e-20
C41731 a_4007_47204# a_3699_46634# 0.008067f
C41732 a_584_46384# a_3877_44458# 1.42e-20
C41733 a_949_44458# a_2127_44172# 0.006932f
C41734 a_n2661_44458# a_5495_43940# 1.41e-20
C41735 a_n699_43396# a_1467_44172# 0.030347f
C41736 a_4223_44672# a_1414_42308# 2.93e-20
C41737 a_742_44458# a_2479_44172# 0.019563f
C41738 a_11649_44734# a_11541_44484# 5.37e-19
C41739 a_13857_44734# a_14112_44734# 0.005172f
C41740 a_1307_43914# a_7499_43940# 0.005916f
C41741 a_n143_45144# a_n229_43646# 1.73e-21
C41742 a_n913_45002# a_3080_42308# 0.044741f
C41743 a_n1059_45260# a_4905_42826# 0.027099f
C41744 a_327_44734# VDD 0.667364f
C41745 a_22400_42852# a_22705_37990# 1.13e-20
C41746 a_11691_44458# a_11415_45002# 0.047412f
C41747 a_20193_45348# a_20202_43084# 0.116706f
C41748 a_13490_45394# a_3483_46348# 0.001975f
C41749 a_949_44458# a_765_45546# 3.16e-19
C41750 a_n2840_43914# a_n2438_43548# 1.6e-21
C41751 a_n1549_44318# a_n2293_46634# 9.06e-21
C41752 a_8855_44734# a_8270_45546# 1.44e-35
C41753 a_3232_43370# a_n1925_42282# 0.021554f
C41754 a_n2293_42834# a_8016_46348# 6.15e-21
C41755 a_9482_43914# a_10809_44734# 0.001033f
C41756 a_13483_43940# a_11453_44696# 1.03e-20
C41757 a_21115_43940# a_18479_47436# 0.001943f
C41758 a_14021_43940# a_12861_44030# 0.035798f
C41759 a_n2661_43370# a_4419_46090# 0.002591f
C41760 a_n4318_39304# SMPL_ON_P 0.039268f
C41761 a_n1917_43396# a_n2497_47436# 0.012526f
C41762 a_1755_42282# a_7174_31319# 1.94e-20
C41763 a_n4318_37592# a_n4334_39616# 7.61e-20
C41764 COMP_P a_n4209_39590# 0.010869f
C41765 a_5934_30871# a_10149_42308# 4.13e-20
C41766 a_5342_30871# C4_N_btm 8.98e-20
C41767 a_5534_30871# C6_N_btm 0.01116f
C41768 C5_P_btm VIN_P 0.502041f
C41769 C7_P_btm VREF 1.818f
C41770 a_4190_30871# a_7754_40130# 4.95e-20
C41771 C9_P_btm VCM 6.06251f
C41772 C8_P_btm VREF_GND 2.58605f
C41773 a_n1151_42308# a_6945_45028# 0.024325f
C41774 a_13747_46662# a_20107_46660# 2.33e-21
C41775 a_12549_44172# a_18280_46660# 0.03199f
C41776 a_13661_43548# a_20411_46873# 3e-19
C41777 a_n743_46660# a_14513_46634# 2.15e-20
C41778 a_10150_46912# a_10428_46928# 0.118759f
C41779 a_9863_46634# a_10467_46802# 0.043587f
C41780 a_8145_46902# a_6755_46942# 0.02566f
C41781 a_n2293_46634# a_13059_46348# 0.207934f
C41782 a_7577_46660# a_6969_46634# 6.14e-19
C41783 a_5257_43370# a_5841_46660# 5.15e-20
C41784 a_19321_45002# a_19123_46287# 2.27e-20
C41785 a_16750_47204# a_765_45546# 1.34e-19
C41786 a_n1435_47204# a_10903_43370# 1.64e-20
C41787 a_2382_45260# a_4156_43218# 6.43e-19
C41788 a_10193_42453# a_8325_42308# 3.66e-20
C41789 a_7499_43078# a_9803_42558# 0.158876f
C41790 a_5891_43370# a_3626_43646# 0.00315f
C41791 a_1307_43914# a_10991_42826# 1.82e-20
C41792 a_1423_45028# a_9127_43156# 2.04e-20
C41793 a_n2293_42834# a_n1736_43218# 0.005982f
C41794 a_n2661_42834# a_1209_43370# 2.79e-20
C41795 a_10057_43914# a_9803_43646# 0.001251f
C41796 a_17517_44484# a_14401_32519# 8.5e-19
C41797 a_13556_45296# a_13635_43156# 8.03e-21
C41798 a_9482_43914# a_13460_43230# 1.07e-20
C41799 a_8975_43940# a_9145_43396# 1.06e-19
C41800 a_13857_44734# VDD 0.18416f
C41801 a_n4209_38502# VCM 0.035344f
C41802 a_n3565_38502# VREF 0.056031f
C41803 a_n3420_38528# VIN_P 0.053985f
C41804 a_2711_45572# a_11525_45546# 0.0154f
C41805 a_7227_45028# a_8162_45546# 0.003048f
C41806 a_6667_45809# a_7499_43078# 2.77e-21
C41807 a_20835_44721# a_20708_46348# 1.53e-20
C41808 a_5244_44056# a_3483_46348# 2.37e-21
C41809 a_18429_43548# a_12549_44172# 3.26e-20
C41810 a_9801_43940# a_3090_45724# 0.004765f
C41811 a_15095_43370# a_n2293_46634# 3.1e-19
C41812 a_n2661_42834# a_8049_45260# 5.27e-20
C41813 a_10440_44484# a_n357_42282# 1.65e-21
C41814 a_742_44458# a_n443_42852# 0.168627f
C41815 a_10150_46912# VDD 0.284144f
C41816 a_13258_32519# C5_N_btm 1.87e-19
C41817 a_7174_31319# C2_N_btm 1.86e-20
C41818 a_n2293_46634# a_3218_45724# 0.001771f
C41819 a_n1925_46634# a_997_45618# 5.01e-21
C41820 a_n2438_43548# a_310_45028# 2.28e-20
C41821 a_n743_46660# a_n357_42282# 0.03365f
C41822 a_1123_46634# a_n2293_45546# 1.17e-21
C41823 a_n1021_46688# a_n755_45592# 1.15e-20
C41824 a_6755_46942# a_5066_45546# 1.35e-19
C41825 a_n133_46660# a_n1099_45572# 5.35e-21
C41826 a_8145_46902# a_8049_45260# 4.44e-19
C41827 a_15227_44166# a_17957_46116# 0.0045f
C41828 a_18834_46812# a_18819_46122# 3.09e-19
C41829 a_14084_46812# a_6945_45028# 5.12e-21
C41830 a_12816_46660# a_10809_44734# 0.011603f
C41831 a_13885_46660# a_10903_43370# 5.54e-19
C41832 a_n3674_37592# a_n3690_37440# 0.071822f
C41833 a_6123_31319# a_n4064_37984# 1.56e-19
C41834 a_5934_30871# a_n3420_37984# 2.14e-19
C41835 a_15682_43940# a_16759_43396# 0.013707f
C41836 a_n97_42460# a_n229_43646# 0.046961f
C41837 a_n1761_44111# a_685_42968# 5.14e-21
C41838 a_11967_42832# a_5534_30871# 0.017079f
C41839 a_18114_32519# a_n1630_35242# 6.72e-20
C41840 a_n2012_43396# a_n1821_43396# 4.61e-19
C41841 a_18451_43940# a_16137_43396# 2.49e-19
C41842 a_n2956_37592# a_n3565_39304# 0.0261f
C41843 a_n1809_43762# VDD 0.142403f
C41844 a_20841_45814# a_2437_43646# 3.5e-21
C41845 a_18479_45785# a_n913_45002# 1.19e-20
C41846 a_8696_44636# a_3537_45260# 1.04e-19
C41847 a_20107_45572# a_19479_31679# 5.42e-21
C41848 a_20273_45572# a_22223_45572# 1.24e-19
C41849 a_15781_43660# a_4185_45028# 4.43e-21
C41850 a_1184_42692# a_768_44030# 6.5e-19
C41851 a_12545_42858# a_3090_45724# 0.002446f
C41852 a_13565_43940# a_13259_45724# 3.63e-19
C41853 a_766_43646# a_526_44458# 1.14e-19
C41854 a_4905_42826# a_n1925_42282# 8.84e-21
C41855 a_13667_43396# a_9290_44172# 0.136018f
C41856 a_10341_43396# a_8199_44636# 2.94e-19
C41857 a_6197_43396# a_6945_45028# 4.56e-21
C41858 a_11323_42473# a_10227_46804# 4.75e-21
C41859 a_15764_42576# a_12861_44030# 1.78e-19
C41860 a_n4334_40480# SMPL_ON_P 1.83e-19
C41861 a_5066_45546# a_8049_45260# 0.076918f
C41862 a_18985_46122# a_19443_46116# 0.027606f
C41863 a_3499_42826# a_3581_42558# 1.79e-19
C41864 a_n2293_43922# a_1736_39587# 3.88e-21
C41865 a_n2661_42282# a_3823_42558# 1.12e-19
C41866 a_2982_43646# a_18083_42858# 1.03e-19
C41867 a_17499_43370# a_5649_42852# 8.65e-21
C41868 a_18579_44172# a_17303_42282# 8.14e-21
C41869 a_15743_43084# a_19095_43396# 0.012939f
C41870 a_1209_43370# a_n2293_42282# 3.21e-21
C41871 a_133_42852# VDD 0.184203f
C41872 a_13159_45002# a_11691_44458# 1.4e-19
C41873 a_2809_45028# a_n2661_43370# 0.003105f
C41874 a_8696_44636# a_11541_44484# 1.04e-19
C41875 a_n2293_42834# a_8488_45348# 1.54e-20
C41876 a_327_44734# a_n699_43396# 1.13e-20
C41877 a_2382_45260# a_949_44458# 2.24e-19
C41878 a_5691_45260# a_n2661_44458# 2.93e-20
C41879 a_n913_45002# a_10057_43914# 1.12e-19
C41880 a_n1059_45260# a_8975_43940# 5.1e-19
C41881 a_5534_30871# a_13259_45724# 0.032063f
C41882 a_n901_43156# a_n443_42852# 0.367747f
C41883 a_1847_42826# a_n357_42282# 0.037548f
C41884 a_8292_43218# a_526_44458# 0.02177f
C41885 a_19332_42282# a_3090_45724# 1.58e-19
C41886 a_14401_32519# EN_VIN_BSTR_N 0.772414f
C41887 a_n2946_37690# SMPL_ON_P 2.4e-19
C41888 a_15861_45028# a_6755_46942# 0.033041f
C41889 a_n913_45002# a_n2438_43548# 6.79e-21
C41890 a_5147_45002# a_5807_45002# 0.035651f
C41891 a_2437_43646# a_n2661_46098# 0.025093f
C41892 en_comp a_n2312_38680# 5.01e-19
C41893 a_n659_45366# a_n2293_46634# 6.05e-19
C41894 a_9482_43914# a_n881_46662# 1.52e-20
C41895 a_13711_45394# a_12861_44030# 6.53e-20
C41896 a_n1917_44484# a_n2497_47436# 0.011319f
C41897 a_n2661_44458# SMPL_ON_P 0.002144f
C41898 a_22821_38993# VDD 0.431879f
C41899 a_n1076_43230# a_n4318_38216# 2.24e-19
C41900 a_14579_43548# a_14113_42308# 9.55e-20
C41901 a_n1991_42858# a_n4318_37592# 3.9e-19
C41902 a_n1853_43023# COMP_P 5.05e-20
C41903 a_n2157_42858# a_n1329_42308# 1.45e-20
C41904 a_743_42282# a_2351_42308# 0.00729f
C41905 a_12281_43396# a_5742_30871# 9.39e-19
C41906 a_n3674_39304# a_n3674_38680# 0.17962f
C41907 a_12545_42858# a_12991_43230# 2.28e-19
C41908 a_n4318_39304# a_n2946_39072# 4.19e-20
C41909 a_22223_46124# RST_Z 1.13e-19
C41910 a_6945_45028# START 0.029602f
C41911 a_n2302_39866# VDD 0.361509f
C41912 a_2905_45572# a_n881_46662# 0.050468f
C41913 a_3160_47472# a_n1613_43370# 0.043254f
C41914 a_3785_47178# a_5063_47570# 2.94e-19
C41915 a_n1151_42308# a_3411_47243# 2.47e-19
C41916 a_n1435_47204# a_4883_46098# 2.09e-20
C41917 a_16763_47508# a_17591_47464# 0.010417f
C41918 a_13717_47436# a_21496_47436# 6.95e-20
C41919 a_12861_44030# a_13507_46334# 0.315418f
C41920 a_16023_47582# a_10227_46804# 0.036076f
C41921 a_16327_47482# a_18143_47464# 1.35e-19
C41922 a_n443_46116# a_3094_47570# 3.58e-19
C41923 a_n2109_47186# a_5807_45002# 0.003143f
C41924 a_n913_45002# a_14021_43940# 2.81e-19
C41925 a_16922_45042# a_3422_30871# 5.99e-20
C41926 a_1307_43914# a_2253_44260# 7.63e-19
C41927 a_n356_44636# a_n310_44811# 0.006879f
C41928 a_10193_42453# a_9145_43396# 0.02642f
C41929 a_2711_45572# a_16977_43638# 2.53e-20
C41930 a_10180_45724# a_9803_43646# 8.22e-23
C41931 a_10775_45002# a_10949_43914# 1.24e-19
C41932 a_n2293_42834# a_1414_42308# 0.02233f
C41933 a_n2661_43370# a_n1899_43946# 6.55e-21
C41934 a_11827_44484# a_20640_44752# 0.016882f
C41935 a_11691_44458# a_11967_42832# 0.041904f
C41936 a_5883_43914# a_9159_44484# 0.049132f
C41937 a_8103_44636# a_n2661_42834# 6.31e-20
C41938 a_6298_44484# a_n2661_43922# 0.048814f
C41939 a_21359_45002# a_20679_44626# 9.5e-19
C41940 a_10951_45334# a_10729_43914# 2.14e-21
C41941 a_21101_45002# a_20835_44721# 4.69e-19
C41942 a_21005_45260# a_20766_44850# 1.08e-19
C41943 a_20567_45036# a_19279_43940# 1.73e-21
C41944 a_19778_44110# a_18579_44172# 0.268475f
C41945 a_10533_42308# a_n443_42852# 1.11e-21
C41946 a_15486_42560# a_n357_42282# 1.89e-20
C41947 a_19647_42308# a_13259_45724# 1.03e-19
C41948 a_n2946_38778# a_n2956_39304# 0.004064f
C41949 a_n3420_38528# a_n2956_38680# 0.233147f
C41950 a_5342_30871# C6_P_btm 0.012f
C41951 a_5534_30871# C4_P_btm 8.01e-20
C41952 a_15861_45028# a_8049_45260# 0.001507f
C41953 a_3537_45260# a_4704_46090# 4.91e-19
C41954 a_3357_43084# a_17583_46090# 1.42e-21
C41955 a_413_45260# a_8016_46348# 1.13e-21
C41956 a_n2017_45002# a_10903_43370# 0.029479f
C41957 a_3065_45002# a_5164_46348# 1.51e-21
C41958 a_2253_44260# a_n443_46116# 0.0014f
C41959 a_4574_45260# a_4419_46090# 3.99e-20
C41960 a_16019_45002# a_12741_44636# 5.77e-19
C41961 a_5111_44636# a_3483_46348# 0.340106f
C41962 a_18587_45118# a_15227_44166# 0.040339f
C41963 a_18911_45144# a_18834_46812# 1.88e-21
C41964 a_n2661_42834# a_n2442_46660# 7.66e-20
C41965 a_4558_45348# a_4185_45028# 0.059418f
C41966 a_556_44484# a_n2438_43548# 0.011144f
C41967 a_3823_42558# a_3497_42558# 2.37e-20
C41968 a_3318_42354# a_3581_42558# 0.011552f
C41969 a_n784_42308# a_8325_42308# 2.26e-20
C41970 a_1755_42282# a_5932_42308# 0.046344f
C41971 a_1184_42692# a_6123_31319# 7.32e-21
C41972 a_5267_42460# a_5379_42460# 0.156424f
C41973 a_1067_42314# a_5934_30871# 1.02e-20
C41974 a_4190_30871# C6_N_btm 0.005085f
C41975 a_22821_38993# a_22469_39537# 0.039707f
C41976 a_22521_40055# a_22705_38406# 0.010302f
C41977 a_22459_39145# a_22609_38406# 0.12318f
C41978 a_22521_39511# a_22876_39857# 0.011942f
C41979 a_22545_38993# a_22780_39857# 0.003614f
C41980 a_n97_42460# CAL_N 8.11e-21
C41981 a_n1925_46634# a_5257_43370# 0.01497f
C41982 a_n2661_46634# a_8667_46634# 0.007776f
C41983 a_2107_46812# a_5167_46660# 0.002706f
C41984 a_2959_46660# a_3067_47026# 0.057222f
C41985 a_5807_45002# a_5841_46660# 2.18e-20
C41986 a_n881_46662# a_12816_46660# 5.76e-20
C41987 a_13507_46334# a_14180_46812# 3.77e-20
C41988 a_4883_46098# a_13885_46660# 5.17e-20
C41989 a_11599_46634# a_20107_46660# 0.266678f
C41990 a_16327_47482# a_765_45546# 0.043622f
C41991 a_13717_47436# a_21363_46634# 3.19e-20
C41992 a_n1741_47186# a_3147_46376# 1.56e-20
C41993 a_n971_45724# a_2202_46116# 3.09e-20
C41994 a_n237_47217# a_1138_42852# 2.57e-19
C41995 a_3160_47472# a_n2293_46098# 1.31e-19
C41996 a_15433_44458# a_11341_43940# 4.01e-21
C41997 a_644_44056# a_453_43940# 0.077973f
C41998 a_1115_44172# a_1414_42308# 0.134389f
C41999 a_n2661_44458# a_3080_42308# 1.4e-21
C42000 a_n2661_42834# a_11173_44260# 0.002687f
C42001 a_n809_44244# a_895_43940# 1.44e-19
C42002 a_11823_42460# a_14853_42852# 9.4e-19
C42003 a_n1059_45260# a_2905_42968# 0.002465f
C42004 a_n2017_45002# a_3681_42891# 1.04e-20
C42005 a_n913_45002# a_2075_43172# 0.175893f
C42006 VDAC_N VDD 4.61811f
C42007 a_4223_44672# VDD 2.99073f
C42008 a_7174_31319# C8_P_btm 7.53e-20
C42009 a_n2946_37984# a_n2956_38216# 0.150404f
C42010 a_n4318_39304# a_n2438_43548# 9.42e-19
C42011 a_2896_43646# a_768_44030# 0.005068f
C42012 a_2982_43646# a_12549_44172# 5e-19
C42013 a_11691_44458# a_13259_45724# 0.337184f
C42014 a_6031_43396# a_n881_46662# 1.13e-19
C42015 a_n2661_43922# a_5937_45572# 0.048264f
C42016 a_n2661_42834# a_8953_45546# 0.019463f
C42017 a_n2293_43922# a_8199_44636# 6.69e-20
C42018 a_7640_43914# a_2324_44458# 3.17e-20
C42019 a_6293_42852# a_n1613_43370# 0.004944f
C42020 a_n1853_43023# a_n2497_47436# 4.11e-19
C42021 a_743_42282# a_584_46384# 3.35e-20
C42022 a_n4209_39590# a_n4209_39304# 0.045123f
C42023 a_n4315_30879# a_n4064_39072# 0.036792f
C42024 a_n4064_40160# a_n3420_39072# 0.052668f
C42025 a_n3565_39590# a_n3607_39616# 0.001003f
C42026 a_n4064_39616# a_n2216_39866# 0.005567f
C42027 a_21588_30879# VDD 1.78413f
C42028 a_6123_31319# C0_P_btm 0.018968f
C42029 a_5932_42308# C2_N_btm 0.011289f
C42030 a_15227_44166# a_11415_45002# 0.047556f
C42031 a_16388_46812# a_18285_46348# 0.028532f
C42032 a_19692_46634# a_20885_46660# 0.002303f
C42033 a_16721_46634# a_17829_46910# 8.81e-20
C42034 a_19321_45002# a_8049_45260# 0.030309f
C42035 a_768_44030# a_14180_46482# 0.00983f
C42036 a_n743_46660# a_518_46155# 4.76e-19
C42037 a_9863_46634# a_8016_46348# 0.001599f
C42038 a_8667_46634# a_8199_44636# 0.005444f
C42039 a_n2312_39304# a_n2840_45546# 0.003056f
C42040 a_n2312_40392# a_n2810_45572# 0.052551f
C42041 a_n913_45002# a_15764_42576# 5.85e-19
C42042 a_n2017_45002# a_15959_42545# 0.004519f
C42043 a_n1059_45260# a_15803_42450# 0.008866f
C42044 a_10807_43548# a_3626_43646# 0.001709f
C42045 a_n2661_42282# a_6765_43638# 2.44e-19
C42046 a_n2293_42834# a_n3674_38680# 0.010983f
C42047 a_742_44458# a_1793_42852# 0.010622f
C42048 a_14539_43914# a_18083_42858# 0.00221f
C42049 a_n356_44636# a_12545_42858# 4.75e-20
C42050 a_1307_43914# a_2713_42308# 4.75e-19
C42051 a_n699_43396# a_133_42852# 1.03e-19
C42052 a_11967_42832# a_4190_30871# 0.002622f
C42053 a_3422_30871# a_15743_43084# 0.022574f
C42054 a_5891_43370# a_8037_42858# 0.12253f
C42055 a_15493_43940# VDD 1.4617f
C42056 a_16333_45814# a_16147_45260# 1.26e-19
C42057 a_15599_45572# a_18341_45572# 1.38e-21
C42058 a_15765_45572# a_18175_45572# 6.29e-20
C42059 a_8696_44636# a_16842_45938# 1.95e-20
C42060 a_5907_45546# a_5691_45260# 0.001013f
C42061 a_3775_45552# a_3429_45260# 0.001061f
C42062 a_2711_45572# a_5205_44484# 8.29e-19
C42063 a_10193_42453# a_n1059_45260# 0.440111f
C42064 a_2675_43914# a_3218_45724# 6.54e-21
C42065 a_n984_44318# a_n443_42852# 1.59e-20
C42066 a_5244_44056# a_n357_42282# 2.74e-21
C42067 a_3905_42865# a_n755_45592# 4.59e-20
C42068 a_n4318_39768# a_n2956_38216# 0.045702f
C42069 a_n97_42460# a_8199_44636# 0.003284f
C42070 a_2713_42308# a_n443_46116# 1.17e-19
C42071 a_8515_42308# a_n971_45724# 3.09e-19
C42072 a_22521_40599# a_22459_39145# 1.41583f
C42073 a_22469_40625# a_22521_40055# 0.076632f
C42074 a_n2302_37690# a_n1838_35608# 5.27e-19
C42075 a_n3420_37440# a_n923_35174# 0.002091f
C42076 a_6293_42852# a_n2293_46098# 0.001583f
C42077 a_n2293_42282# a_n2442_46660# 5.92e-20
C42078 a_14537_43646# a_13059_46348# 0.003923f
C42079 a_19700_43370# a_19692_46634# 4.58e-19
C42080 a_9127_43156# a_4646_46812# 4.29e-21
C42081 a_22223_45036# RST_Z 1.13e-19
C42082 a_6419_46155# VDD 0.094119f
C42083 a_2711_45572# a_n971_45724# 0.214535f
C42084 a_6194_45824# a_n1741_47186# 3.64e-21
C42085 a_6511_45714# a_n2109_47186# 5.45e-21
C42086 a_n4064_39072# a_n3420_37440# 0.051893f
C42087 a_n3420_39072# a_n4064_37440# 0.047151f
C42088 a_n4064_39616# VDAC_P 0.008251f
C42089 a_12741_44636# a_20254_46482# 3.54e-19
C42090 a_765_45546# a_n356_45724# 3.13e-19
C42091 a_22365_46825# a_20205_31679# 0.002648f
C42092 a_8953_45546# a_5066_45546# 0.191859f
C42093 a_7920_46348# a_8062_46482# 0.007833f
C42094 a_20075_46420# a_20708_46348# 0.017547f
C42095 a_19553_46090# a_6945_45028# 1.78e-21
C42096 a_18819_46122# a_10809_44734# 7.49e-20
C42097 a_2982_43646# a_21855_43396# 2.81e-19
C42098 a_n229_43646# a_n901_43156# 3.1e-19
C42099 a_14021_43940# a_20922_43172# 6.69e-20
C42100 a_13667_43396# a_13749_43396# 0.005781f
C42101 a_14205_43396# a_14621_43646# 2.64e-19
C42102 a_n1761_44111# a_n1329_42308# 7.38e-20
C42103 a_n4318_40392# a_n4064_39072# 2.29e-21
C42104 a_3422_30871# a_1606_42308# 0.022481f
C42105 a_n1899_43946# COMP_P 4.56e-21
C42106 a_n2293_43922# a_13070_42354# 0.002481f
C42107 a_21588_30879# a_22469_39537# 1.05e-19
C42108 a_22612_30879# a_22821_38993# 1.98e-19
C42109 a_n3674_39304# VDD 0.587205f
C42110 a_3537_45260# a_5009_45028# 0.001769f
C42111 a_5691_45260# a_6125_45348# 0.003935f
C42112 en_comp a_n2661_43370# 0.164814f
C42113 a_21188_45572# a_11827_44484# 1.57e-20
C42114 a_8696_44636# a_8701_44490# 0.095858f
C42115 a_14537_43396# a_14797_45144# 0.082443f
C42116 a_9482_43914# a_1307_43914# 0.010221f
C42117 a_20107_45572# a_20193_45348# 8.83e-19
C42118 a_n2946_39866# a_n2956_39768# 0.14868f
C42119 a_n3565_39590# a_n2442_46660# 0.134948f
C42120 a_3681_42891# a_526_44458# 0.002914f
C42121 a_2905_42968# a_n1925_42282# 1.42e-20
C42122 a_4190_30871# a_13259_45724# 0.271537f
C42123 a_9885_43646# a_n443_42852# 0.001927f
C42124 a_n913_45002# a_13507_46334# 0.023897f
C42125 a_n2017_45002# a_4883_46098# 1.86e-19
C42126 a_413_45260# a_17591_47464# 4.35e-19
C42127 a_626_44172# a_584_46384# 0.450256f
C42128 a_1307_43914# a_2905_45572# 1.08e-21
C42129 a_15765_45572# a_n743_46660# 0.026376f
C42130 a_8568_45546# a_7411_46660# 0.001217f
C42131 a_8696_44636# a_n2293_46634# 3.28e-20
C42132 a_16377_45572# a_13661_43548# 1.08e-20
C42133 a_n356_45724# a_509_45822# 2.78e-19
C42134 a_310_45028# a_603_45572# 8.28e-19
C42135 a_1848_45724# a_2307_45899# 6.64e-19
C42136 a_3218_45724# a_2277_45546# 7.5e-20
C42137 a_3316_45546# a_1609_45822# 1.08e-19
C42138 a_n357_42282# a_509_45572# 3.18e-19
C42139 a_15743_43084# a_18504_43218# 2.23e-19
C42140 a_n97_42460# a_13070_42354# 0.02477f
C42141 a_2982_43646# a_7227_42308# 6.66e-20
C42142 a_12379_42858# a_12545_42858# 0.810394f
C42143 a_16977_43638# a_16877_42852# 6.98e-20
C42144 a_11415_45002# EN_OFFSET_CAL 0.14622f
C42145 VDAC_N a_8912_37509# 3.43288f
C42146 a_3422_30871# C1_N_btm 7.67e-20
C42147 a_6886_37412# VDAC_P 0.062773f
C42148 a_5700_37509# a_11206_38545# 4.96e-20
C42149 a_5742_30871# VDD 0.556959f
C42150 a_n1605_47204# a_n1435_47204# 0.110832f
C42151 a_n1741_47186# a_12861_44030# 5.74e-20
C42152 a_n1151_42308# a_4700_47436# 0.01362f
C42153 a_2905_45572# a_n443_46116# 0.14923f
C42154 a_3785_47178# a_3815_47204# 0.270823f
C42155 a_4223_44672# a_n699_43396# 0.217586f
C42156 a_11691_44458# a_18989_43940# 0.066207f
C42157 a_n2661_44458# a_10057_43914# 0.007497f
C42158 a_16147_45260# a_15493_43396# 9.87e-21
C42159 a_413_45260# a_1414_42308# 0.12534f
C42160 a_n913_45002# a_5013_44260# 7.77e-21
C42161 a_n1059_45260# a_5495_43940# 1.76e-21
C42162 a_n2840_45002# a_n4318_39768# 0.002422f
C42163 a_n473_42460# a_n357_42282# 0.179066f
C42164 a_564_42282# a_n863_45724# 1.21e-19
C42165 a_n961_42308# a_n755_45592# 2.27e-20
C42166 a_4190_30871# C4_P_btm 1.36e-19
C42167 a_13887_32519# a_11530_34132# 0.005035f
C42168 VDAC_N a_22612_30879# 0.011363f
C42169 a_16147_45260# a_3483_46348# 6.65e-20
C42170 a_n2661_44458# a_n2438_43548# 0.136664f
C42171 a_n2661_43370# a_7411_46660# 5.29e-21
C42172 a_2437_43646# a_11415_45002# 0.01065f
C42173 a_14797_45144# a_3090_45724# 9.53e-19
C42174 a_n1177_44458# a_n2293_46634# 1.56e-19
C42175 a_14539_43914# a_12549_44172# 0.110516f
C42176 a_14537_43396# a_14976_45028# 0.087031f
C42177 a_20719_45572# a_12741_44636# 3.43e-19
C42178 a_3357_43084# a_20885_46660# 5.68e-19
C42179 a_6977_45572# a_6945_45028# 0.001758f
C42180 a_10306_45572# a_2324_44458# 7.74e-19
C42181 a_9313_44734# a_12465_44636# 2.57e-20
C42182 a_13296_44484# a_12861_44030# 1.28e-19
C42183 a_n1899_43946# a_n2497_47436# 0.040963f
C42184 a_16414_43172# a_16522_42674# 6.05e-20
C42185 a_5342_30871# a_15521_42308# 2.73e-19
C42186 a_5807_45002# a_n1925_46634# 0.933976f
C42187 a_21588_30879# a_22612_30879# 7.53611f
C42188 a_n881_46662# a_2443_46660# 1.1e-19
C42189 a_n1613_43370# a_2609_46660# 0.631348f
C42190 a_3815_47204# a_3090_45724# 6.61e-21
C42191 a_n1151_42308# a_15559_46634# 2.09e-19
C42192 a_4915_47217# a_12991_46634# 0.068619f
C42193 a_6151_47436# a_11901_46660# 2.66e-19
C42194 a_10227_46804# a_8492_46660# 6.27e-21
C42195 a_15811_47375# a_6755_46942# 8.93e-20
C42196 a_5111_44636# a_10695_43548# 6.49e-20
C42197 a_n1059_45260# a_16137_43396# 0.438785f
C42198 a_n2017_45002# a_16243_43396# 9.54e-20
C42199 a_n2293_42834# a_n1190_43762# 8.33e-20
C42200 a_375_42282# a_648_43396# 9.82e-19
C42201 a_13249_42308# a_5342_30871# 7.46e-20
C42202 a_10193_42453# a_19987_42826# 0.164153f
C42203 a_n2661_43370# a_n1699_43638# 7.67e-21
C42204 a_9482_43914# a_9396_43370# 0.011522f
C42205 a_1307_43914# a_6031_43396# 0.002834f
C42206 a_n2661_42834# a_895_43940# 0.095907f
C42207 a_n2661_43922# a_2479_44172# 0.002669f
C42208 a_20159_44458# a_18579_44172# 4.88e-19
C42209 a_17517_44484# a_20512_43084# 0.027951f
C42210 a_20835_44721# a_20766_44850# 0.209641f
C42211 a_20679_44626# a_19279_43940# 0.279785f
C42212 a_15004_44636# a_14955_43940# 2.26e-20
C42213 a_n2293_42834# VDD 0.853754f
C42214 a_20205_31679# C4_N_btm 0.042623f
C42215 a_20692_30879# C3_N_btm 3.19e-20
C42216 a_5932_42308# C8_P_btm 1.4e-19
C42217 a_5934_30871# EN_VIN_BSTR_N 0.073476f
C42218 a_1606_42308# VREF_GND 9e-19
C42219 a_16019_45002# a_16375_45002# 0.032313f
C42220 a_3065_45002# a_3316_45546# 0.141454f
C42221 a_3429_45260# a_3218_45724# 0.001528f
C42222 a_n467_45028# a_n443_42852# 0.007314f
C42223 a_5111_44636# a_n357_42282# 0.033023f
C42224 a_6671_43940# a_n881_46662# 1.87e-19
C42225 a_20567_45036# a_20708_46348# 5.99e-19
C42226 a_11691_44458# a_18189_46348# 6.35e-20
C42227 a_7499_43940# a_n1613_43370# 0.001731f
C42228 a_2813_43396# a_584_46384# 0.00985f
C42229 a_11967_42832# a_15227_44166# 0.132673f
C42230 a_1443_43940# a_768_44030# 0.003817f
C42231 a_15493_43940# a_22612_30879# 1.68e-20
C42232 a_16763_47508# VDD 0.392885f
C42233 a_6123_31319# comp_n 1.63e-19
C42234 a_18057_42282# a_18214_42558# 0.18824f
C42235 a_5934_30871# a_1239_39043# 6.07e-20
C42236 a_33_46660# a_167_45260# 7.22e-22
C42237 a_n743_46660# a_3147_46376# 0.016933f
C42238 a_n2661_46098# a_n1853_46287# 0.019613f
C42239 a_1123_46634# a_1138_42852# 0.00173f
C42240 a_2609_46660# a_n2293_46098# 1.8e-20
C42241 a_948_46660# a_1176_45822# 0.003207f
C42242 a_2107_46812# a_1208_46090# 5e-19
C42243 a_6755_46942# a_13059_46348# 0.239671f
C42244 a_3090_45724# a_14976_45028# 0.730613f
C42245 a_8667_46634# a_765_45546# 1.37e-20
C42246 a_15009_46634# a_15368_46634# 7.72e-19
C42247 a_5807_45002# a_10355_46116# 0.003081f
C42248 a_n2661_46634# a_5204_45822# 1.9e-19
C42249 a_768_44030# a_13925_46122# 0.02161f
C42250 a_12891_46348# a_14275_46494# 4.45e-21
C42251 a_4883_46098# a_526_44458# 0.010154f
C42252 a_12861_44030# a_10586_45546# 9.62e-21
C42253 a_n2497_47436# a_1848_45724# 7.52e-22
C42254 a_n2109_47186# a_n755_45592# 5.59e-21
C42255 a_n971_45724# a_n1079_45724# 0.150623f
C42256 a_n746_45260# a_n2293_45546# 0.404324f
C42257 a_n2293_42834# a_873_42968# 1.97e-20
C42258 a_15433_44458# a_10341_43396# 1.5e-21
C42259 a_18989_43940# a_4190_30871# 1.16e-19
C42260 a_2127_44172# a_n97_42460# 1.47e-19
C42261 a_15493_43940# a_22959_43948# 0.182001f
C42262 a_18451_43940# a_14021_43940# 1.25e-20
C42263 a_9313_44734# a_16409_43396# 6.68e-20
C42264 a_7584_44260# a_7499_43940# 1.48e-19
C42265 a_n1059_45260# a_n784_42308# 0.008929f
C42266 a_n913_45002# a_196_42282# 1.19e-19
C42267 en_comp COMP_P 1.92051f
C42268 a_n2293_45010# a_564_42282# 6.44e-21
C42269 a_n2017_45002# a_n327_42558# 0.005655f
C42270 a_n967_45348# a_n4318_37592# 8.19e-19
C42271 a_1115_44172# VDD 0.165092f
C42272 C1_N_btm VREF_GND 0.673422f
C42273 C0_N_btm VCM 0.717064f
C42274 C2_N_btm VREF 0.987884f
C42275 C3_N_btm VIN_N 0.455045f
C42276 a_11962_45724# a_11778_45572# 5.39e-20
C42277 a_2711_45572# a_19431_45546# 2.71e-21
C42278 a_10193_42453# a_15599_45572# 5.53e-20
C42279 a_11823_42460# a_11136_45572# 5.02e-20
C42280 a_1241_43940# a_1138_42852# 0.006402f
C42281 a_13565_44260# a_3483_46348# 3.95e-19
C42282 a_7287_43370# a_3090_45724# 0.005365f
C42283 a_8685_43396# a_8270_45546# 0.006203f
C42284 a_n1423_42826# a_n2442_46660# 4.46e-21
C42285 a_n2661_43922# a_n443_42852# 0.045456f
C42286 a_10729_43914# a_2324_44458# 2.83e-21
C42287 a_20922_43172# a_13507_46334# 2.68e-20
C42288 a_14097_32519# w_11334_34010# 5.84e-19
C42289 a_11415_45002# a_22959_46124# 0.002009f
C42290 a_13059_46348# a_8049_45260# 0.068978f
C42291 a_15227_44166# a_13259_45724# 0.916975f
C42292 a_3483_46348# a_9290_44172# 0.207611f
C42293 a_12741_44636# a_6945_45028# 0.021699f
C42294 a_22591_46660# a_10809_44734# 0.013929f
C42295 a_7174_31319# a_2113_38308# 8.18e-20
C42296 a_5164_46348# a_5937_45572# 3.66e-19
C42297 a_19808_44306# a_15743_43084# 5.11e-21
C42298 a_5883_43914# a_9293_42558# 2.71e-21
C42299 a_n2293_43922# a_n4318_38216# 5.44e-19
C42300 a_2479_44172# a_3445_43172# 1.16e-19
C42301 a_18184_42460# a_18220_42308# 5.62e-19
C42302 a_11967_42832# a_14635_42282# 0.018349f
C42303 a_19319_43548# a_18783_43370# 9.48e-20
C42304 a_6765_43638# a_7112_43396# 0.051162f
C42305 a_18494_42460# a_18214_42558# 0.012583f
C42306 a_n356_44636# a_5379_42460# 0.038779f
C42307 a_14021_43940# a_17364_32525# 0.007637f
C42308 a_18533_43940# a_18525_43370# 7.52e-19
C42309 a_n1151_42308# DATA[2] 0.01294f
C42310 a_3381_47502# DATA[1] 4.03e-22
C42311 a_2063_45854# CLK 0.271193f
C42312 a_19479_31679# C4_N_btm 9.91e-21
C42313 a_10849_43646# VDD 0.009276f
C42314 a_2711_45572# a_13076_44458# 6.99e-21
C42315 a_15143_45578# a_11691_44458# 3.46e-19
C42316 a_10180_45724# a_n2661_44458# 2.83e-19
C42317 a_413_45260# a_1667_45002# 0.00537f
C42318 a_n2017_45002# a_3232_43370# 1.68e-19
C42319 a_n447_43370# a_n443_42852# 0.002103f
C42320 a_n1557_42282# a_n863_45724# 0.034373f
C42321 a_4235_43370# a_n357_42282# 0.005266f
C42322 a_4093_43548# a_n755_45592# 1.18e-21
C42323 a_2982_43646# a_n2661_45546# 0.007559f
C42324 a_5111_42852# a_1823_45246# 5.16e-20
C42325 a_14113_42308# a_5807_45002# 1.48e-22
C42326 a_1755_42282# a_4646_46812# 1.48e-21
C42327 a_13657_42558# a_13661_43548# 3.59e-20
C42328 a_13157_43218# a_3090_45724# 7.17e-19
C42329 a_3422_30871# C9_P_btm 0.003737f
C42330 a_n310_45899# VDD 0.002211f
C42331 a_12427_45724# a_12549_44172# 0.152925f
C42332 a_7499_43078# a_5807_45002# 6.76e-20
C42333 a_6511_45714# a_n1925_46634# 0.028817f
C42334 a_6194_45824# a_n743_46660# 0.002138f
C42335 a_11823_42460# a_12891_46348# 0.033376f
C42336 a_6469_45572# a_n881_46662# 3.11e-19
C42337 a_6905_45572# a_n1613_43370# 8.54e-19
C42338 a_15037_45618# a_12465_44636# 2.95e-21
C42339 a_15903_45785# a_13507_46334# 7.77e-20
C42340 a_18175_45572# a_12861_44030# 0.031037f
C42341 en_comp a_n2497_47436# 4.47e-20
C42342 a_n2661_45010# a_n746_45260# 0.400342f
C42343 a_2437_43646# a_2553_47502# 0.004656f
C42344 a_16137_43396# a_19987_42826# 2.41e-19
C42345 a_n2267_43396# a_n1329_42308# 8.36e-21
C42346 a_17499_43370# a_17333_42852# 7.75e-20
C42347 a_15743_43084# a_16414_43172# 1.55e-19
C42348 a_5649_42852# a_5755_42852# 0.089078f
C42349 a_4361_42308# a_7765_42852# 3.76e-20
C42350 a_743_42282# a_8952_43230# 3.27e-20
C42351 a_n2129_43609# a_n961_42308# 1.71e-20
C42352 a_15493_43396# a_15051_42282# 3.6e-21
C42353 a_n3674_39304# a_n4318_38680# 2.92578f
C42354 a_n1853_43023# a_133_43172# 6.79e-19
C42355 a_n1991_42858# a_n1533_42852# 0.034619f
C42356 a_n1699_43638# COMP_P 9.19e-20
C42357 a_16292_46812# RST_Z 9.44e-21
C42358 a_22765_42852# VDD 0.006527f
C42359 a_2437_43646# a_11967_42832# 4.65e-20
C42360 a_5147_45002# a_5608_44484# 0.003234f
C42361 a_2382_45260# a_n2293_43922# 5.18e-20
C42362 a_8191_45002# a_5891_43370# 6.65e-19
C42363 a_3065_45002# a_n2661_42834# 0.022516f
C42364 a_2680_45002# a_n2661_43922# 6.61e-20
C42365 a_n2661_43370# a_n1699_44726# 0.001811f
C42366 a_18494_42460# a_21359_45002# 4.97e-21
C42367 a_19778_44110# a_22223_45036# 6.5e-20
C42368 a_10193_42453# a_18326_43940# 0.130866f
C42369 a_n2293_42834# a_n699_43396# 0.00729f
C42370 a_18315_45260# a_11691_44458# 8.2e-21
C42371 a_18184_42460# a_11827_44484# 0.027981f
C42372 a_20567_45036# a_21101_45002# 3.03e-19
C42373 a_18587_45118# a_19113_45348# 2.02e-19
C42374 a_11823_42460# a_11750_44172# 6.71e-20
C42375 a_12427_45724# a_12429_44172# 4.6e-20
C42376 a_19647_42308# a_20202_43084# 6.58e-21
C42377 a_n784_42308# a_n1925_42282# 0.235613f
C42378 a_14635_42282# a_13259_45724# 3.09e-19
C42379 a_9885_42558# a_8953_45546# 0.024699f
C42380 a_10533_42308# a_8199_44636# 4.26e-20
C42381 a_413_45260# a_10428_46928# 1.23e-20
C42382 a_5205_44484# a_6540_46812# 1.12e-21
C42383 a_4558_45348# a_5257_43370# 2.74e-21
C42384 a_5111_44636# a_5263_46660# 5.58e-20
C42385 a_3357_43084# a_11813_46116# 1.83e-20
C42386 a_2711_45572# a_12594_46348# 0.009529f
C42387 a_18450_45144# a_11453_44696# 3.07e-19
C42388 a_20273_45572# a_15227_44166# 2.83e-19
C42389 a_9049_44484# a_3483_46348# 0.117501f
C42390 a_17478_45572# a_17829_46910# 2.26e-21
C42391 a_4361_42308# a_13657_42308# 5.57e-19
C42392 a_7227_42852# a_6123_31319# 0.001591f
C42393 a_16823_43084# a_18057_42282# 2.44e-21
C42394 a_n2293_42282# a_n3674_38216# 0.111055f
C42395 a_15743_43084# a_7174_31319# 3.05e-19
C42396 a_11453_44696# a_12549_44172# 0.066205f
C42397 a_18479_47436# a_19594_46812# 0.108004f
C42398 a_18780_47178# a_19321_45002# 4.23e-20
C42399 a_19386_47436# a_13747_46662# 0.145228f
C42400 a_n1435_47204# a_n133_46660# 2.75e-20
C42401 a_12861_44030# a_n743_46660# 0.100542f
C42402 a_6575_47204# a_2107_46812# 1.07e-19
C42403 a_n971_45724# a_6540_46812# 0.31827f
C42404 a_n443_46116# a_2443_46660# 0.041057f
C42405 a_n1151_42308# a_3067_47026# 7.63e-19
C42406 a_3785_47178# a_3524_46660# 0.002172f
C42407 a_3815_47204# a_3699_46634# 2.44e-19
C42408 a_584_46384# a_3221_46660# 6.04e-20
C42409 a_949_44458# a_453_43940# 0.006129f
C42410 a_2779_44458# a_1414_42308# 5.89e-19
C42411 a_742_44458# a_2127_44172# 0.002775f
C42412 a_n2661_44458# a_5013_44260# 2.48e-20
C42413 a_n699_43396# a_1115_44172# 6.01e-20
C42414 a_11823_42460# a_4361_42308# 0.056415f
C42415 a_1307_43914# a_6671_43940# 0.007083f
C42416 a_13249_42308# a_743_42282# 0.010211f
C42417 a_9482_43914# a_10867_43940# 2.96e-19
C42418 a_18989_43940# a_18753_44484# 4.75e-19
C42419 a_n467_45028# a_n229_43646# 6.99e-21
C42420 a_2382_45260# a_n97_42460# 0.02063f
C42421 a_n913_45002# a_4699_43561# 8.4e-21
C42422 a_n1059_45260# a_3080_42308# 0.025424f
C42423 a_n2017_45002# a_4905_42826# 0.042734f
C42424 a_n2293_45010# a_n1557_42282# 1.08e-20
C42425 a_413_45260# VDD 1.203f
C42426 a_n2661_43370# a_4185_45028# 0.053994f
C42427 a_11827_44484# a_12741_44636# 0.305294f
C42428 a_19113_45348# a_11415_45002# 0.012208f
C42429 a_13105_45348# a_3483_46348# 4.98e-19
C42430 a_2437_43646# a_13259_45724# 3.14e-20
C42431 a_3232_43370# a_526_44458# 0.461444f
C42432 a_n2293_42834# a_7920_46348# 4.35e-20
C42433 a_5837_45028# a_5937_45572# 0.043505f
C42434 a_1423_45028# a_2324_44458# 0.154419f
C42435 a_12429_44172# a_11453_44696# 2.89e-21
C42436 a_18451_43940# a_13507_46334# 2.1e-20
C42437 a_20365_43914# a_18597_46090# 4.85e-21
C42438 a_20935_43940# a_18479_47436# 0.207572f
C42439 a_11341_43940# a_10227_46804# 0.057378f
C42440 a_13829_44260# a_12861_44030# 3.01e-20
C42441 a_n2840_43370# SMPL_ON_P 8.96e-19
C42442 a_n1699_43638# a_n2497_47436# 0.038204f
C42443 a_1606_42308# a_7174_31319# 2.41314f
C42444 a_5742_30871# a_11551_42558# 0.007648f
C42445 a_n4318_38216# a_n3420_39616# 0.023792f
C42446 a_5934_30871# a_9885_42308# 0.001708f
C42447 a_n3674_38680# a_n4064_39616# 0.019915f
C42448 a_5342_30871# C3_N_btm 8.34e-20
C42449 a_5534_30871# C5_N_btm 8.45e-20
C42450 C6_P_btm VIN_P 0.391898f
C42451 C8_P_btm VREF 3.6701f
C42452 C9_P_btm VREF_GND 5.18245f
C42453 C10_P_btm VCM 10.5945f
C42454 SMPL_ON_P a_n1925_42282# 1.26e-19
C42455 a_12549_44172# a_17639_46660# 0.129285f
C42456 a_13661_43548# a_20107_46660# 2.78e-20
C42457 a_n743_46660# a_14180_46812# 4.96e-20
C42458 a_7577_46660# a_6755_46942# 0.035922f
C42459 a_7715_46873# a_6969_46634# 3.3e-19
C42460 a_9863_46634# a_10428_46928# 0.042509f
C42461 a_19321_45002# a_18285_46348# 4.63e-22
C42462 a_13747_46662# a_19551_46910# 0.001463f
C42463 a_5807_45002# a_20411_46873# 1.37e-19
C42464 a_3065_45002# a_n2293_42282# 0.007636f
C42465 a_2382_45260# a_3935_43218# 0.005937f
C42466 a_11691_44458# a_16867_43762# 7.88e-20
C42467 a_7499_43078# a_9223_42460# 0.013802f
C42468 a_1423_45028# a_8387_43230# 4.08e-21
C42469 a_3499_42826# a_n2661_42282# 1.48e-20
C42470 a_9482_43914# a_13635_43156# 3.22e-21
C42471 a_1307_43914# a_10796_42968# 1.45e-20
C42472 a_n2293_42834# a_n4318_38680# 0.007189f
C42473 a_n356_44636# a_7287_43370# 7.66e-21
C42474 a_n2661_42834# a_458_43396# 0.001339f
C42475 a_15004_44636# a_8685_43396# 8.84e-21
C42476 a_10057_43914# a_9145_43396# 0.121499f
C42477 a_13468_44734# VDD 0.004018f
C42478 a_n3565_38216# C2_P_btm 0.040789f
C42479 a_n4209_38502# VREF_GND 0.00199f
C42480 a_2711_45572# a_11322_45546# 0.056109f
C42481 a_6511_45714# a_7499_43078# 1.26e-20
C42482 a_7227_45028# a_7230_45938# 0.170618f
C42483 a_6598_45938# a_8162_45546# 9.36e-20
C42484 a_14205_43396# a_n2293_46634# 0.0055f
C42485 a_17324_43396# a_12549_44172# 6.76e-20
C42486 a_11341_43940# a_17339_46660# 0.023304f
C42487 a_9420_43940# a_3090_45724# 0.00133f
C42488 a_10334_44484# a_n357_42282# 9.23e-21
C42489 a_18579_44172# a_18819_46122# 8.68e-21
C42490 a_13678_32519# SMPL_ON_N 0.029315f
C42491 a_17364_32525# a_13507_46334# 3.3e-20
C42492 a_3905_42865# a_3483_46348# 3.18e-20
C42493 a_2998_44172# a_4185_45028# 0.001414f
C42494 a_20447_31679# a_21589_35634# 3.86e-20
C42495 a_9863_46634# VDD 0.411318f
C42496 a_13258_32519# C4_N_btm 2.18e-19
C42497 a_7174_31319# C1_N_btm 5.34e-20
C42498 a_n2293_46634# a_2957_45546# 0.001699f
C42499 a_n1925_46634# a_n755_45592# 7.2e-20
C42500 a_n743_46660# a_310_45028# 0.143623f
C42501 a_n2438_43548# a_n1099_45572# 7.2e-20
C42502 a_7577_46660# a_8049_45260# 4.87e-20
C42503 a_33_46660# a_n863_45724# 5.8e-20
C42504 a_2107_46812# a_n2661_45546# 9.54e-20
C42505 a_765_45546# a_5204_45822# 1.06e-19
C42506 a_13607_46688# a_6945_45028# 3.26e-20
C42507 a_12991_46634# a_10809_44734# 0.008021f
C42508 a_15227_44166# a_18189_46348# 0.066472f
C42509 a_n3674_37592# a_n3565_37414# 0.129086f
C42510 a_5932_42308# a_2113_38308# 9.09e-20
C42511 a_n1630_35242# a_n4209_37414# 2.12e-19
C42512 a_n784_42308# a_n3420_37440# 0.140549f
C42513 a_15682_43940# a_16977_43638# 0.003291f
C42514 a_18326_43940# a_16137_43396# 3.25e-22
C42515 a_n1352_43396# a_458_43396# 1.68e-20
C42516 a_14021_43940# a_9145_43396# 0.032057f
C42517 a_17517_44484# a_18249_42858# 8.87e-22
C42518 a_11967_42832# a_14543_43071# 0.022161f
C42519 a_19319_43548# a_3626_43646# 4.18e-20
C42520 a_n447_43370# a_n229_43646# 0.08213f
C42521 a_5891_43370# a_7309_42852# 0.071511f
C42522 a_14539_43914# a_14853_42852# 3.54e-21
C42523 a_1307_43914# a_4958_30871# 9.67e-22
C42524 a_n2810_45028# a_n3565_39304# 0.021534f
C42525 en_comp a_n4209_39304# 3.42e-19
C42526 a_n2012_43396# VDD 0.08228f
C42527 a_20623_45572# a_20885_45572# 0.001705f
C42528 a_21188_45572# a_21350_45938# 0.006453f
C42529 a_20107_45572# a_22223_45572# 7.3e-21
C42530 a_6667_45809# a_n2661_43370# 3.11e-20
C42531 a_20273_45572# a_2437_43646# 8.82e-20
C42532 a_4190_30871# a_20202_43084# 4.66e-19
C42533 a_12089_42308# a_3090_45724# 0.002716f
C42534 a_1576_42282# a_768_44030# 6.84e-23
C42535 a_4905_42826# a_526_44458# 0.202895f
C42536 a_3080_42308# a_n1925_42282# 0.897997f
C42537 a_9885_43646# a_8199_44636# 0.007796f
C42538 a_10695_43548# a_9290_44172# 0.011352f
C42539 a_10723_42308# a_10227_46804# 6.28e-21
C42540 a_15486_42560# a_12861_44030# 1.58e-19
C42541 a_n4315_30879# SMPL_ON_P 3.70932f
C42542 a_5527_46155# VDD 2.18e-20
C42543 a_2711_45572# a_12465_44636# 0.027219f
C42544 a_10490_45724# a_11459_47204# 3.69e-22
C42545 a_10193_42453# a_n1435_47204# 9.87e-21
C42546 a_6945_45028# a_16375_45002# 3.78e-20
C42547 a_19553_46090# a_20009_46494# 4.2e-19
C42548 a_19335_46494# a_19597_46482# 0.001705f
C42549 a_9290_44172# a_n357_42282# 0.138435f
C42550 a_18819_46122# a_19443_46116# 9.73e-19
C42551 a_3499_42826# a_3497_42558# 1.79e-19
C42552 a_18783_43370# a_19095_43396# 0.038241f
C42553 a_n2293_43922# a_1239_39587# 1.55e-20
C42554 a_7845_44172# a_7963_42308# 7.62e-22
C42555 a_n2661_42282# a_3318_42354# 1.07e-19
C42556 a_2982_43646# a_17701_42308# 1.83e-19
C42557 a_3626_43646# a_16795_42852# 2.28e-21
C42558 a_15743_43084# a_21487_43396# 1.58e-19
C42559 a_19700_43370# a_743_42282# 0.001969f
C42560 a_458_43396# a_n2293_42282# 1.03e-20
C42561 a_n914_42852# VDD 7.75e-19
C42562 a_13017_45260# a_11691_44458# 1.87e-20
C42563 a_13556_45296# a_11827_44484# 0.05613f
C42564 a_n2293_42834# a_8137_45348# 0.009658f
C42565 a_2448_45028# a_n2661_43370# 2.21e-19
C42566 a_2274_45254# a_949_44458# 3.92e-19
C42567 a_4927_45028# a_n2661_44458# 0.00137f
C42568 a_413_45260# a_n699_43396# 0.100762f
C42569 a_n1059_45260# a_10057_43914# 6.77e-20
C42570 a_2382_45260# a_742_44458# 3.78e-19
C42571 a_14456_42282# a_13059_46348# 0.001136f
C42572 a_685_42968# a_n755_45592# 2.82e-19
C42573 a_791_42968# a_n357_42282# 0.009083f
C42574 a_3935_42891# a_n863_45724# 4.1e-20
C42575 a_7573_43172# a_526_44458# 0.001584f
C42576 a_n1641_43230# a_n443_42852# 8.55e-20
C42577 a_14543_43071# a_13259_45724# 2.13e-20
C42578 COMP_P a_4185_45028# 3.46e-20
C42579 a_1067_42314# a_1138_42852# 3.59e-19
C42580 a_14401_32519# a_11530_34132# 0.004736f
C42581 a_3726_37500# w_1575_34946# 0.007105f
C42582 a_n3420_37440# SMPL_ON_P 0.025729f
C42583 a_15143_45578# a_15227_44166# 0.010748f
C42584 a_11823_42460# a_12359_47026# 5.24e-20
C42585 a_8696_44636# a_6755_46942# 0.04097f
C42586 a_2437_43646# a_1799_45572# 0.002971f
C42587 a_413_45260# a_22612_30879# 0.11791f
C42588 a_n1059_45260# a_n2438_43548# 3.13e-20
C42589 a_n967_45348# a_n2293_46634# 0.007362f
C42590 a_7229_43940# a_768_44030# 0.042486f
C42591 a_n2956_37592# a_n2312_38680# 0.048307f
C42592 a_4558_45348# a_5807_45002# 9.02e-19
C42593 a_n4318_40392# SMPL_ON_P 0.039594f
C42594 a_n1699_44726# a_n2497_47436# 0.012807f
C42595 a_11691_44458# a_2063_45854# 4.35e-20
C42596 a_22545_38993# VDD 0.536989f
C42597 a_n901_43156# a_n4318_38216# 6.06e-21
C42598 a_n1853_43023# a_n4318_37592# 1.26e-19
C42599 a_n1991_42858# a_n1736_42282# 0.0101f
C42600 a_n2157_42858# COMP_P 1.05e-19
C42601 a_12545_42858# a_12800_43218# 0.05936f
C42602 a_n3674_39304# a_n2840_42282# 4.48e-19
C42603 a_743_42282# a_2123_42473# 0.007332f
C42604 a_12281_43396# a_11323_42473# 3.39e-20
C42605 a_2982_43646# a_21613_42308# 0.001693f
C42606 a_3539_42460# a_7174_31319# 4.88e-21
C42607 a_n4318_39304# a_n3420_39072# 0.001411f
C42608 a_10341_42308# a_11136_42852# 0.003f
C42609 a_3080_42308# a_n4315_30879# 5.51e-21
C42610 a_6945_45028# RST_Z 0.022027f
C42611 a_20708_46348# SINGLE_ENDED 9.74e-21
C42612 a_n4064_39616# VDD 1.6861f
C42613 a_2905_45572# a_n1613_43370# 0.044171f
C42614 a_3785_47178# a_4842_47570# 9.52e-19
C42615 a_3160_47472# a_3411_47243# 4.21e-19
C42616 a_n1151_42308# a_3094_47243# 3.77e-19
C42617 a_11599_46634# a_19386_47436# 1.17e-21
C42618 a_16763_47508# a_16588_47582# 0.233657f
C42619 a_13717_47436# a_13507_46334# 3.3e-19
C42620 a_13381_47204# a_4883_46098# 7.29e-21
C42621 a_16327_47482# a_10227_46804# 0.630403f
C42622 a_n237_47217# a_768_44030# 7.54e-19
C42623 a_n1059_45260# a_14021_43940# 0.008971f
C42624 a_413_45260# a_22959_43948# 0.00133f
C42625 a_5343_44458# a_n2293_43922# 2.33e-20
C42626 a_11691_44458# a_19006_44850# 0.005009f
C42627 a_8701_44490# a_9159_44484# 6.03e-19
C42628 a_2711_45572# a_16409_43396# 2.45e-19
C42629 a_n2293_42834# a_1467_44172# 9.22e-22
C42630 a_n2661_43370# a_n1761_44111# 1.12e-20
C42631 a_11827_44484# a_20362_44736# 0.009001f
C42632 a_6298_44484# a_n2661_42834# 0.001263f
C42633 a_5518_44484# a_n2661_43922# 0.011667f
C42634 a_n356_44636# a_n23_44458# 0.220577f
C42635 a_21359_45002# a_20640_44752# 0.013689f
C42636 a_21101_45002# a_20679_44626# 0.001069f
C42637 a_21005_45260# a_20835_44721# 7.06e-20
C42638 a_20567_45036# a_20766_44850# 0.001007f
C42639 a_18494_42460# a_19279_43940# 0.137363f
C42640 a_18911_45144# a_18579_44172# 2.07e-20
C42641 a_10775_45002# a_10729_43914# 1.25e-21
C42642 a_15051_42282# a_n357_42282# 3.44e-19
C42643 a_19511_42282# a_13259_45724# 7.13e-20
C42644 a_n3420_38528# a_n2956_39304# 0.001161f
C42645 a_n3690_38528# a_n2956_38680# 0.015398f
C42646 a_5342_30871# C7_P_btm 5.39e-19
C42647 a_5534_30871# C5_P_btm 8.45e-20
C42648 a_4574_45260# a_4185_45028# 0.006766f
C42649 a_5147_45002# a_3483_46348# 0.363215f
C42650 a_18315_45260# a_15227_44166# 0.272047f
C42651 a_484_44484# a_n2438_43548# 7.2e-20
C42652 a_n2293_43922# a_n2956_39768# 6.42e-20
C42653 a_n2661_43922# a_n2661_46634# 1.58e-19
C42654 a_5205_44484# a_1823_45246# 4.61e-19
C42655 a_8696_44636# a_8049_45260# 0.005215f
C42656 a_7499_43078# a_n755_45592# 0.157526f
C42657 a_21188_45572# a_21137_46414# 1.5e-20
C42658 a_3357_43084# a_15682_46116# 3.34e-20
C42659 a_21363_45546# a_6945_45028# 2.51e-20
C42660 a_2437_43646# a_18189_46348# 3.03e-20
C42661 a_19237_31679# a_13507_46334# 6.88e-20
C42662 a_n2661_42282# a_n1151_42308# 1.58e-19
C42663 a_3537_45260# a_4419_46090# 0.003458f
C42664 a_16751_45260# a_11415_45002# 0.009485f
C42665 a_15595_45028# a_12741_44636# 3.6e-19
C42666 a_n1630_35242# a_5934_30871# 0.039258f
C42667 a_3318_42354# a_3497_42558# 0.010303f
C42668 a_5534_30871# a_n3420_38528# 0.041746f
C42669 a_1606_42308# a_5932_42308# 0.111585f
C42670 a_1755_42282# a_6171_42473# 0.065035f
C42671 a_2713_42308# a_3905_42558# 1.81e-21
C42672 a_1576_42282# a_6123_31319# 2.22e-20
C42673 a_4190_30871# C5_N_btm 1.71e-19
C42674 a_22545_38993# a_22469_39537# 0.049703f
C42675 a_22459_39145# CAL_P 0.005678f
C42676 a_22521_40055# a_22609_38406# 0.1922f
C42677 a_22521_39511# a_22780_39857# 0.01318f
C42678 a_n2661_46634# a_7927_46660# 0.00501f
C42679 a_2107_46812# a_5385_46902# 0.001613f
C42680 a_3177_46902# a_3067_47026# 0.097745f
C42681 a_3699_46634# a_3524_46660# 0.233657f
C42682 a_768_44030# a_8270_45546# 0.03575f
C42683 a_n2661_46098# a_2162_46660# 0.003322f
C42684 a_2959_46660# a_2864_46660# 0.049827f
C42685 a_n1925_46634# a_5429_46660# 4.33e-19
C42686 a_n881_46662# a_12991_46634# 1.56e-19
C42687 a_3080_42308# a_n3420_37440# 7.3e-19
C42688 a_13507_46334# a_14035_46660# 0.027121f
C42689 a_16327_47482# a_17339_46660# 0.058779f
C42690 a_11599_46634# a_19551_46910# 5.02e-19
C42691 a_16241_47178# a_765_45546# 0.004102f
C42692 a_18479_47436# a_16388_46812# 5.74e-20
C42693 a_4915_47217# a_11415_45002# 0.134061f
C42694 a_13717_47436# a_20623_46660# 2.48e-20
C42695 a_n971_45724# a_1823_45246# 0.514159f
C42696 a_327_47204# a_472_46348# 7.59e-19
C42697 a_2905_45572# a_n2293_46098# 0.028964f
C42698 a_n2109_47186# a_3483_46348# 0.03221f
C42699 a_n746_45260# a_1138_42852# 6.98e-20
C42700 a_n237_47217# a_1176_45822# 3.23e-19
C42701 a_5343_44458# a_n97_42460# 3.84e-19
C42702 a_175_44278# a_453_43940# 0.112594f
C42703 a_1115_44172# a_1467_44172# 0.115277f
C42704 a_17061_44734# a_15682_43940# 1.68e-19
C42705 a_14815_43914# a_11341_43940# 0.001047f
C42706 a_n2661_44458# a_4699_43561# 1.98e-20
C42707 a_n2661_42834# a_10555_44260# 0.003997f
C42708 a_644_44056# a_1414_42308# 5.43e-20
C42709 a_n913_45002# a_1847_42826# 0.294312f
C42710 a_n2017_45002# a_2905_42968# 7.95e-20
C42711 a_n967_45348# a_n1533_42852# 0.002483f
C42712 a_6886_37412# VDD 0.235486f
C42713 a_2779_44458# VDD 0.38604f
C42714 a_7174_31319# C9_P_btm 9.33e-20
C42715 a_n4315_30879# a_n1532_35090# 2.87e-19
C42716 a_n3420_37984# a_n2956_38216# 0.208204f
C42717 a_n2302_37984# a_n2810_45572# 0.130495f
C42718 a_n2840_43370# a_n2438_43548# 0.00955f
C42719 a_1987_43646# a_768_44030# 3.01e-19
C42720 a_11827_44484# a_16375_45002# 2.06e-19
C42721 a_6298_44484# a_5066_45546# 7.32e-21
C42722 a_8975_43940# a_526_44458# 3.81e-21
C42723 a_n2661_44458# a_10586_45546# 9.07e-20
C42724 a_n2661_43922# a_8199_44636# 0.04879f
C42725 a_n2661_42834# a_5937_45572# 0.043505f
C42726 a_6109_44484# a_2324_44458# 0.101116f
C42727 a_6031_43396# a_n1613_43370# 0.308901f
C42728 a_10341_43396# a_10227_46804# 0.188948f
C42729 a_n2157_42858# a_n2497_47436# 1.22e-19
C42730 a_n4064_39616# a_n2860_39866# 0.003766f
C42731 a_n4064_40160# a_n3690_39392# 3.42e-19
C42732 a_7174_31319# a_n4209_38502# 5.81e-22
C42733 a_20916_46384# VDD 0.302226f
C42734 a_6123_31319# C1_P_btm 0.011005f
C42735 a_5932_42308# C1_N_btm 0.011049f
C42736 a_15227_44166# a_20202_43084# 0.086371f
C42737 a_16388_46812# a_17829_46910# 1.39e-19
C42738 a_16721_46634# a_765_45546# 0.002907f
C42739 a_19692_46634# a_20719_46660# 0.004558f
C42740 a_5807_45002# a_10044_46482# 5.69e-19
C42741 a_n743_46660# a_3873_46454# 2.25e-19
C42742 a_8492_46660# a_8016_46348# 7.47e-19
C42743 a_4646_46812# a_2324_44458# 0.023652f
C42744 a_n913_45002# a_15486_42560# 2.61e-19
C42745 a_n2017_45002# a_15803_42450# 0.005056f
C42746 a_5111_44636# a_8685_42308# 3.87e-21
C42747 a_n1059_45260# a_15764_42576# 4.65e-19
C42748 a_742_44458# a_1709_42852# 0.001488f
C42749 a_n2661_42282# a_6197_43396# 0.033187f
C42750 a_9165_43940# a_9420_43940# 0.005172f
C42751 a_14539_43914# a_17701_42308# 0.039977f
C42752 a_n356_44636# a_12089_42308# 5.58e-20
C42753 a_5891_43370# a_7765_42852# 0.168516f
C42754 a_8375_44464# a_8037_42858# 4.44e-20
C42755 a_22223_43948# VDD 0.254313f
C42756 a_15765_45572# a_16147_45260# 0.005068f
C42757 a_16680_45572# a_16842_45938# 0.006453f
C42758 a_16115_45572# a_16377_45572# 0.001705f
C42759 a_4099_45572# a_3232_43370# 2.19e-22
C42760 a_3775_45552# a_3065_45002# 3.53e-20
C42761 a_10193_42453# a_n2017_45002# 0.081859f
C42762 a_2711_45572# a_6431_45366# 0.001609f
C42763 a_10341_43396# a_17339_46660# 0.023552f
C42764 a_19268_43646# a_19692_46634# 5.49e-20
C42765 a_8387_43230# a_4646_46812# 4.44e-20
C42766 a_3600_43914# a_n755_45592# 7.02e-21
C42767 a_n809_44244# a_n443_42852# 1.06e-19
C42768 a_3905_42865# a_n357_42282# 0.059842f
C42769 a_22400_42852# a_18597_46090# 2.28e-21
C42770 a_5934_30871# a_n971_45724# 7.07e-19
C42771 CAL_N a_22459_39145# 0.014789f
C42772 a_22521_40599# a_22521_40055# 0.086402f
C42773 a_22469_40625# a_22780_40945# 4.21e-20
C42774 a_n3565_37414# EN_VIN_BSTR_P 0.069167f
C42775 a_4338_37500# CAL_P 0.00316f
C42776 a_6031_43396# a_n2293_46098# 1.36e-21
C42777 a_4093_43548# a_3483_46348# 4.56e-21
C42778 a_6165_46155# VDD 0.204296f
C42779 a_5937_45572# a_5066_45546# 0.419426f
C42780 a_20075_46420# a_19900_46494# 0.233657f
C42781 a_18985_46122# a_6945_45028# 1.4e-20
C42782 a_n3565_39304# a_n2302_37690# 4.02e-19
C42783 a_2112_39137# VDAC_Ni 0.018166f
C42784 a_n1917_43396# a_n1533_42852# 1.04e-19
C42785 a_14579_43548# a_15681_43442# 9.87e-22
C42786 a_2982_43646# a_4361_42308# 0.545077f
C42787 a_14021_43940# a_19987_42826# 1.06e-19
C42788 a_n2293_43922# a_12563_42308# 0.015547f
C42789 a_9313_44734# a_15890_42674# 1.49e-20
C42790 a_14358_43442# a_14621_43646# 0.011552f
C42791 a_14205_43396# a_14537_43646# 3.88e-19
C42792 a_n1761_44111# COMP_P 2.35e-19
C42793 a_n356_44636# a_18907_42674# 2.06e-20
C42794 a_n1809_43762# a_n3674_39304# 9.24e-22
C42795 a_n2012_43396# a_n4318_38680# 1.79e-19
C42796 a_8685_43396# a_16759_43396# 1.34e-19
C42797 a_3315_47570# DATA[2] 9.25e-20
C42798 a_21588_30879# a_22821_38993# 1.81e-19
C42799 a_n13_43084# VDD 0.260551f
C42800 a_3065_45002# a_5093_45028# 1.41e-21
C42801 a_n2956_37592# a_n2661_43370# 0.044152f
C42802 a_5691_45260# a_5837_45348# 0.013377f
C42803 a_20731_45938# a_21005_45260# 2.73e-20
C42804 a_21363_45546# a_11827_44484# 1.3e-22
C42805 a_21188_45572# a_21359_45002# 4.16e-19
C42806 a_10490_45724# a_9313_44734# 4.22e-21
C42807 a_14180_45002# a_14797_45144# 0.070624f
C42808 a_2711_45572# a_16241_44734# 0.03035f
C42809 a_8696_44636# a_8103_44636# 1.41e-19
C42810 a_13556_45296# a_15595_45028# 1.42e-20
C42811 a_13348_45260# a_1307_43914# 3.41e-21
C42812 a_4743_43172# a_4185_45028# 5.73e-19
C42813 a_n3420_39616# a_n2956_39768# 0.233256f
C42814 a_n4334_39616# a_n2442_46660# 6.16e-20
C42815 a_14955_43396# a_n443_42852# 0.076467f
C42816 a_2905_42968# a_526_44458# 0.007721f
C42817 a_15567_42826# a_2324_44458# 7.25e-19
C42818 a_15903_45785# a_n743_46660# 2.48e-19
C42819 a_6598_45938# a_6969_46634# 6.03e-19
C42820 a_8162_45546# a_7411_46660# 4.69e-20
C42821 a_16842_45938# a_13747_46662# 3.67e-19
C42822 a_7227_45028# a_6755_46942# 2.07e-20
C42823 a_16211_45572# a_13661_43548# 6.84e-20
C42824 a_2437_43646# a_2747_46873# 0.003933f
C42825 a_n1059_45260# a_13507_46334# 3.96e-20
C42826 a_413_45260# a_16588_47582# 8.28e-20
C42827 a_9482_43914# a_4791_45118# 6.76e-20
C42828 a_501_45348# a_584_46384# 1.78e-19
C42829 a_1848_45724# a_1990_45899# 0.005572f
C42830 a_310_45028# a_509_45572# 1.27e-19
C42831 a_n1099_45572# a_603_45572# 3.32e-19
C42832 a_n755_45592# a_n310_45572# 0.001154f
C42833 a_3539_42460# a_5932_42308# 4.34e-21
C42834 a_n97_42460# a_12563_42308# 0.001953f
C42835 a_2982_43646# a_6761_42308# 3.92e-20
C42836 a_10341_42308# a_12545_42858# 9.44e-20
C42837 a_12379_42858# a_12089_42308# 0.16885f
C42838 a_20202_43084# EN_OFFSET_CAL 0.001606f
C42839 a_6886_37412# a_8912_37509# 0.339465f
C42840 a_3422_30871# C0_N_btm 6.53e-20
C42841 a_5700_37509# VDAC_P 0.081094f
C42842 a_4338_37500# CAL_N 0.052373f
C42843 a_5088_37509# a_11206_38545# 0.005271f
C42844 a_n237_47217# a_9067_47204# 0.0235f
C42845 SMPL_ON_P a_n1435_47204# 0.082028f
C42846 a_2063_45854# a_5129_47502# 9.87e-20
C42847 a_n1741_47186# a_13717_47436# 6.56e-20
C42848 a_11323_42473# VDD 0.205172f
C42849 a_n1151_42308# a_4007_47204# 0.015013f
C42850 a_3381_47502# a_3815_47204# 0.021997f
C42851 a_2905_45572# a_4791_45118# 0.001355f
C42852 a_2952_47436# a_n443_46116# 9.06e-19
C42853 a_18175_45572# a_18451_43940# 6.66e-21
C42854 a_16751_45260# a_11967_42832# 1.76e-21
C42855 a_2779_44458# a_n699_43396# 0.025176f
C42856 a_n2661_44458# a_10440_44484# 0.005733f
C42857 a_11691_44458# a_18374_44850# 0.02267f
C42858 a_19113_45348# a_18989_43940# 3.13e-19
C42859 a_n1059_45260# a_5013_44260# 2e-20
C42860 a_n2017_45002# a_5495_43940# 8.92e-22
C42861 a_n913_45002# a_5244_44056# 1.75e-21
C42862 a_n961_42308# a_n357_42282# 7.65e-19
C42863 a_n1329_42308# a_n755_45592# 2.67e-21
C42864 a_4190_30871# C5_P_btm 1.71e-19
C42865 VDAC_N a_21588_30879# 0.006893f
C42866 a_n2661_43370# a_5257_43370# 0.027779f
C42867 a_n2661_44458# a_n743_46660# 8.9e-21
C42868 a_2437_43646# a_20202_43084# 0.129143f
C42869 a_13017_45260# a_15227_44166# 5.47e-20
C42870 a_21513_45002# a_11415_45002# 0.050445f
C42871 a_n4318_40392# a_n2438_43548# 0.001259f
C42872 a_16112_44458# a_12549_44172# 1.91e-20
C42873 a_14537_43396# a_3090_45724# 0.530123f
C42874 a_14539_43914# a_12891_46348# 3.29e-20
C42875 a_7227_45028# a_8049_45260# 3.6e-19
C42876 a_10193_42453# a_526_44458# 1.72e-19
C42877 a_3357_43084# a_20719_46660# 0.001371f
C42878 a_8696_44636# a_8953_45546# 0.022578f
C42879 a_14033_45822# a_12594_46348# 0.001526f
C42880 a_6905_45572# a_6945_45028# 7.62e-19
C42881 a_10216_45572# a_2324_44458# 9.53e-19
C42882 a_n1809_44850# a_n1613_43370# 0.012196f
C42883 a_n2293_43922# a_10227_46804# 1.57e-19
C42884 a_11967_42832# a_4915_47217# 1.34e-21
C42885 a_n1761_44111# a_n2497_47436# 0.045728f
C42886 a_n4318_38680# a_n4064_39616# 0.021342f
C42887 a_4190_30871# a_n3420_38528# 0.031855f
C42888 a_n1741_47186# a_14035_46660# 2.61e-20
C42889 a_3785_47178# a_3090_45724# 4.4e-22
C42890 a_n1151_42308# a_15368_46634# 2.09e-19
C42891 a_20916_46384# a_22612_30879# 3.3e-20
C42892 a_n881_46662# a_n2661_46098# 0.096736f
C42893 a_9313_45822# a_8654_47026# 4.81e-20
C42894 a_4915_47217# a_12251_46660# 2.85e-19
C42895 a_9067_47204# a_8270_45546# 9.93e-19
C42896 a_6151_47436# a_11813_46116# 8.68e-20
C42897 a_15507_47210# a_6755_46942# 2.7e-19
C42898 a_10227_46804# a_8667_46634# 6.04e-20
C42899 a_n1613_43370# a_2443_46660# 0.917984f
C42900 a_n2017_45002# a_16137_43396# 0.63011f
C42901 a_5111_44636# a_9803_43646# 0.118936f
C42902 a_n2293_42834# a_n1809_43762# 0.001769f
C42903 a_375_42282# a_548_43396# 6.62e-19
C42904 a_19006_44850# a_18753_44484# 4.61e-19
C42905 a_10193_42453# a_19164_43230# 0.003383f
C42906 a_n2661_43370# a_n2267_43396# 0.001687f
C42907 a_n2661_42834# a_2479_44172# 0.027713f
C42908 a_n2661_43922# a_2127_44172# 0.007786f
C42909 a_19615_44636# a_18579_44172# 0.158449f
C42910 a_20640_44752# a_19279_43940# 0.22152f
C42911 a_20679_44626# a_20766_44850# 0.052825f
C42912 a_20692_30879# C2_N_btm 1.93e-20
C42913 a_5932_42308# C9_P_btm 9.33e-20
C42914 a_5934_30871# a_11530_34132# 8.66e-19
C42915 a_1241_43940# a_768_44030# 0.003504f
C42916 a_15493_43940# a_21588_30879# 1.53e-20
C42917 a_16751_45260# a_13259_45724# 1.84e-20
C42918 a_2382_45260# a_3503_45724# 3.72e-20
C42919 a_3065_45002# a_3218_45724# 0.002508f
C42920 a_5147_45002# a_n357_42282# 1.06e-21
C42921 a_2680_45002# a_3316_45546# 0.050127f
C42922 a_16237_45028# a_15682_46116# 3.39e-20
C42923 a_n2661_44458# a_11189_46129# 2.93e-21
C42924 a_5518_44484# a_5164_46348# 7.19e-19
C42925 a_11691_44458# a_17715_44484# 0.036149f
C42926 a_19113_45348# a_18189_46348# 2.31e-19
C42927 a_6671_43940# a_n1613_43370# 0.03314f
C42928 a_n97_42460# a_10227_46804# 0.18445f
C42929 a_6031_43396# a_4791_45118# 4.86e-20
C42930 a_1512_43396# a_n443_46116# 0.010064f
C42931 a_2437_43396# a_584_46384# 8.66e-20
C42932 a_10157_44484# a_3483_46348# 2.51e-21
C42933 a_5883_43914# a_4185_45028# 4.3e-21
C42934 a_16023_47582# VDD 0.201413f
C42935 a_6123_31319# a_1736_39043# 6.11e-20
C42936 a_18727_42674# a_18907_42674# 0.185422f
C42937 a_n1925_46634# a_3483_46348# 4.03e-19
C42938 a_n743_46660# a_2804_46116# 0.012952f
C42939 a_n2661_46098# a_n2157_46122# 0.227082f
C42940 a_2443_46660# a_n2293_46098# 1.88e-20
C42941 a_1123_46634# a_1176_45822# 0.001261f
C42942 a_948_46660# a_1208_46090# 3.04e-19
C42943 a_2107_46812# a_805_46414# 1.28e-19
C42944 a_15009_46634# a_14976_45028# 0.071873f
C42945 a_12549_44172# a_13925_46122# 5.78e-20
C42946 a_768_44030# a_13759_46122# 0.024686f
C42947 a_5807_45002# a_9823_46155# 0.005199f
C42948 a_n2661_46634# a_5164_46348# 1.31e-19
C42949 a_9804_47204# a_2324_44458# 1.14e-19
C42950 a_4915_47217# a_13259_45724# 0.04489f
C42951 a_n971_45724# a_n2293_45546# 0.097168f
C42952 a_n815_47178# a_n863_45724# 2.42e-20
C42953 a_n1741_47186# a_n1099_45572# 2.08e-20
C42954 a_n809_44244# a_n229_43646# 0.001748f
C42955 a_453_43940# a_n97_42460# 2.8e-19
C42956 a_14815_43914# a_10341_43396# 8.2e-20
C42957 a_n699_43396# a_n13_43084# 0.001012f
C42958 a_9313_44734# a_16547_43609# 0.010576f
C42959 a_3422_30871# a_3626_43646# 1.22e-19
C42960 a_10193_42453# a_21973_42336# 3.78e-21
C42961 a_14539_43914# a_4361_42308# 2.29e-20
C42962 a_3357_43084# a_1755_42282# 4.76e-20
C42963 a_n967_45348# a_n1736_42282# 0.001893f
C42964 a_n913_45002# a_n473_42460# 7.7e-21
C42965 a_n1059_45260# a_196_42282# 4.1e-19
C42966 a_n2017_45002# a_n784_42308# 0.0226f
C42967 en_comp a_n4318_37592# 0.03345f
C42968 a_n2956_37592# COMP_P 1.39e-21
C42969 a_644_44056# VDD 0.147321f
C42970 a_11652_45724# a_11778_45572# 0.001094f
C42971 a_11962_45724# a_11688_45572# 2.07e-20
C42972 a_11525_45546# a_12016_45572# 0.00278f
C42973 C0_N_btm VREF_GND 0.350401f
C42974 C0_dummy_N_btm VCM 0.311452f
C42975 C1_N_btm VREF 0.98698f
C42976 C2_N_btm VIN_N 0.502408f
C42977 a_6547_43396# a_3090_45724# 0.003527f
C42978 a_n97_42460# a_17339_46660# 0.001432f
C42979 a_5755_42852# a_768_44030# 2.35e-21
C42980 a_n2661_42834# a_n443_42852# 0.076984f
C42981 a_18005_44484# a_16375_45002# 8.14e-20
C42982 a_10796_42968# a_n1613_43370# 1.91e-20
C42983 a_19987_42826# a_13507_46334# 6.44e-20
C42984 a_16751_46987# VDD 8.63e-19
C42985 a_12741_44636# a_21137_46414# 2.81e-21
C42986 a_3483_46348# a_10355_46116# 1.51e-21
C42987 a_11415_45002# a_10809_44734# 0.140489f
C42988 a_5742_30871# VDAC_N 0.008249f
C42989 a_n2293_43922# a_n2472_42282# 1.85e-19
C42990 a_n2661_43922# a_n4318_38216# 5.64e-19
C42991 a_3539_42460# a_4181_43396# 3.38e-21
C42992 a_16922_45042# a_20712_42282# 2.62e-20
C42993 a_18494_42460# a_19332_42282# 0.040916f
C42994 a_18184_42460# a_18214_42558# 0.056496f
C42995 a_11967_42832# a_13291_42460# 0.015813f
C42996 a_n356_44636# a_5267_42460# 1.4e-19
C42997 a_n2661_42834# a_n2104_42282# 3.95e-21
C42998 a_14021_43940# a_22959_43396# 0.191956f
C42999 a_6197_43396# a_7112_43396# 0.118423f
C43000 a_2479_44172# a_n2293_42282# 0.059476f
C43001 a_9672_43914# a_9127_43156# 0.001066f
C43002 a_9028_43914# a_8952_43230# 6.18e-20
C43003 a_3160_47472# DATA[2] 5.43e-20
C43004 a_n1151_42308# DATA[1] 0.009539f
C43005 a_10765_43646# VDD 0.00801f
C43006 a_14495_45572# a_11691_44458# 2.65e-20
C43007 a_413_45260# a_327_44734# 0.195096f
C43008 a_n37_45144# a_1667_45002# 1.12e-20
C43009 a_n913_45002# a_5111_44636# 0.070773f
C43010 a_12991_43230# a_3090_45724# 0.001405f
C43011 a_n1352_43396# a_n443_42852# 2.4e-19
C43012 a_4093_43548# a_n357_42282# 0.002194f
C43013 a_7174_31319# a_n2312_39304# 4.73e-21
C43014 a_22775_42308# SMPL_ON_N 9.64e-21
C43015 a_4520_42826# a_1823_45246# 0.053569f
C43016 a_3422_30871# C10_P_btm 0.002966f
C43017 a_n23_45546# VDD 0.150941f
C43018 a_11652_45724# a_768_44030# 4.54e-22
C43019 a_11962_45724# a_12549_44172# 0.034917f
C43020 a_8568_45546# a_5807_45002# 7.37e-22
C43021 a_6472_45840# a_n1925_46634# 9.08e-19
C43022 a_5907_45546# a_n743_46660# 0.002962f
C43023 a_12427_45724# a_12891_46348# 1.55e-19
C43024 a_15599_45572# a_13507_46334# 4.46e-20
C43025 a_16020_45572# a_10227_46804# 3.37e-19
C43026 a_16147_45260# a_12861_44030# 3.97e-19
C43027 a_n2956_37592# a_n2497_47436# 1.14e-20
C43028 a_n2017_45002# SMPL_ON_P 1.46e-21
C43029 a_n2661_45010# a_n971_45724# 0.017233f
C43030 a_2437_43646# a_2063_45854# 0.392331f
C43031 a_16137_43396# a_19164_43230# 9.01e-19
C43032 a_n1699_43638# a_n4318_37592# 9.74e-21
C43033 a_n1917_43396# a_n1736_42282# 7.84e-20
C43034 a_n2267_43396# COMP_P 8.07e-20
C43035 a_17324_43396# a_17701_42308# 0.00643f
C43036 a_17499_43370# a_18083_42858# 0.003663f
C43037 a_15743_43084# a_15567_42826# 0.215954f
C43038 a_5649_42852# a_5111_42852# 0.110096f
C43039 a_4361_42308# a_7871_42858# 6.79e-20
C43040 a_743_42282# a_9127_43156# 2.23e-19
C43041 a_n1641_43230# a_n1379_43218# 0.001705f
C43042 a_n1423_42826# a_n967_43230# 4.2e-19
C43043 a_15559_46634# RST_Z 1.85e-21
C43044 a_11901_46660# CLK 6.62e-20
C43045 a_7754_39964# a_7754_39300# 3.86e-20
C43046 a_20753_42852# VDD 0.193909f
C43047 a_21513_45002# a_11967_42832# 5.76e-19
C43048 a_6171_45002# a_9313_44734# 2.05e-20
C43049 a_2382_45260# a_n2661_43922# 0.026472f
C43050 a_20731_45938# a_20835_44721# 8.44e-21
C43051 a_8191_45002# a_8375_44464# 9.04e-19
C43052 a_2680_45002# a_n2661_42834# 6.24e-21
C43053 a_21188_45572# a_19279_43940# 3.06e-19
C43054 a_11823_42460# a_10807_43548# 4.89e-19
C43055 a_10193_42453# a_18079_43940# 0.076581f
C43056 a_n2293_42834# a_4223_44672# 0.015649f
C43057 a_5837_45028# a_5518_44484# 1.43e-19
C43058 a_n2661_43370# a_n2267_44484# 0.007573f
C43059 a_18494_42460# a_21101_45002# 1.76e-20
C43060 a_19778_44110# a_11827_44484# 0.029054f
C43061 a_17719_45144# a_11691_44458# 2.64e-20
C43062 a_20567_45036# a_21005_45260# 0.015494f
C43063 a_19511_42282# a_20202_43084# 0.082529f
C43064 a_13291_42460# a_13259_45724# 0.089962f
C43065 a_n2293_42282# a_n443_42852# 4.9e-19
C43066 a_n784_42308# a_526_44458# 0.011818f
C43067 a_196_42282# a_n1925_42282# 2.11e-19
C43068 a_8685_42308# a_9290_44172# 1.4e-21
C43069 a_9377_42558# a_8953_45546# 0.007183f
C43070 a_20107_45572# a_15227_44166# 1.29e-19
C43071 a_17478_45572# a_765_45546# 0.00712f
C43072 a_n2661_43370# a_5807_45002# 0.018021f
C43073 a_2809_45028# a_n2293_46634# 4.98e-19
C43074 a_13490_45067# a_768_44030# 2.87e-19
C43075 a_14033_45572# a_13059_46348# 2.71e-20
C43076 a_3357_43084# a_11735_46660# 5.8e-20
C43077 a_413_45260# a_10150_46912# 9.34e-21
C43078 a_2711_45572# a_12005_46116# 6.25e-20
C43079 a_4880_45572# a_5204_45822# 0.046074f
C43080 a_7499_43078# a_3483_46348# 0.207714f
C43081 a_4361_42308# a_11897_42308# 3.73e-19
C43082 a_15743_43084# a_20712_42282# 4.16e-20
C43083 a_743_42282# a_17124_42282# 0.007228f
C43084 a_16823_43084# a_17531_42308# 1.38e-20
C43085 a_7227_42852# a_7227_42308# 3.59e-19
C43086 a_n2293_42282# a_n2104_42282# 0.058363f
C43087 a_19700_43370# a_13258_32519# 1.55e-20
C43088 a_11453_44696# a_12891_46348# 0.029995f
C43089 a_12465_44636# a_16119_47582# 5.64e-20
C43090 a_18597_46090# a_13747_46662# 0.391702f
C43091 a_18479_47436# a_19321_45002# 0.262984f
C43092 a_10227_46804# a_20843_47204# 0.02328f
C43093 a_19386_47436# a_13661_43548# 1.13e-19
C43094 a_n1435_47204# a_n2438_43548# 1.05e-19
C43095 a_7903_47542# a_2107_46812# 1.01e-20
C43096 a_13717_47436# a_n743_46660# 7.97e-20
C43097 a_n237_47217# a_5167_46660# 2.88e-21
C43098 a_n971_45724# a_5732_46660# 0.004372f
C43099 a_3160_47472# a_3067_47026# 0.002863f
C43100 a_3785_47178# a_3699_46634# 0.001286f
C43101 a_n443_46116# a_n2661_46098# 0.198865f
C43102 a_584_46384# a_3055_46660# 1.4e-19
C43103 a_949_44458# a_1414_42308# 0.009641f
C43104 a_742_44458# a_453_43940# 0.001956f
C43105 a_n2661_44458# a_5244_44056# 1.12e-20
C43106 a_n699_43396# a_644_44056# 1.32e-19
C43107 a_1307_43914# a_5829_43940# 0.016223f
C43108 a_9313_44734# a_14673_44172# 6.42e-20
C43109 a_18374_44850# a_18753_44484# 3.16e-19
C43110 a_2274_45254# a_n97_42460# 6.35e-21
C43111 a_n913_45002# a_4235_43370# 9.46e-20
C43112 a_n1059_45260# a_4699_43561# 1.87e-20
C43113 a_n2017_45002# a_3080_42308# 0.034898f
C43114 a_n37_45144# VDD 0.138f
C43115 a_22400_42852# a_22705_38406# 2.84e-20
C43116 a_n2661_43370# a_3699_46348# 5.24e-21
C43117 a_21359_45002# a_12741_44636# 4.18e-19
C43118 a_11915_45394# a_3483_46348# 0.002345f
C43119 a_22959_45036# a_11415_45002# 0.001254f
C43120 a_18374_44850# a_15227_44166# 4.22e-19
C43121 a_7845_44172# a_768_44030# 0.004571f
C43122 a_n1899_43946# a_n2293_46634# 5.11e-21
C43123 a_n356_44636# a_3090_45724# 5.97e-22
C43124 a_5093_45028# a_5937_45572# 9.15e-20
C43125 a_11750_44172# a_11453_44696# 1.03e-20
C43126 a_20623_43914# a_18479_47436# 0.012705f
C43127 a_n2267_43396# a_n2497_47436# 0.222725f
C43128 a_11323_42473# a_11551_42558# 0.062483f
C43129 a_n3674_38216# a_n4334_39616# 9.11e-20
C43130 a_5342_30871# C2_N_btm 7.86e-20
C43131 a_5534_30871# C4_N_btm 8.01e-20
C43132 C9_P_btm VREF 7.369471f
C43133 C7_P_btm VIN_P 1.52449f
C43134 C10_P_btm VREF_GND 10.3207f
C43135 a_n746_45260# a_739_46482# 1.28e-19
C43136 a_n2497_47436# a_1337_46116# 8.17e-21
C43137 a_n1741_47186# a_n1925_42282# 3.03e-20
C43138 a_n743_46660# a_14035_46660# 0.007691f
C43139 a_13747_46662# a_19123_46287# 0.191545f
C43140 a_13661_43548# a_19551_46910# 6.46e-20
C43141 a_8667_46634# a_10467_46802# 2.84e-21
C43142 a_7411_46660# a_6969_46634# 0.033891f
C43143 a_7715_46873# a_6755_46942# 0.089466f
C43144 a_9863_46634# a_10150_46912# 0.233657f
C43145 a_8492_46660# a_10428_46928# 8.55e-21
C43146 a_12549_44172# a_16655_46660# 1.26e-19
C43147 a_n881_46662# a_11415_45002# 0.017774f
C43148 a_n1435_47204# a_11133_46155# 2.19e-21
C43149 a_11459_47204# a_10903_43370# 1.51e-21
C43150 a_12861_44030# a_9290_44172# 0.09212f
C43151 a_6545_47178# a_2324_44458# 2.07e-20
C43152 a_2382_45260# a_3445_43172# 1.08e-19
C43153 a_n2661_42834# a_n229_43646# 0.001251f
C43154 a_n2293_42834# a_n3674_39304# 1.76e-19
C43155 a_16922_45042# a_20556_43646# 0.00844f
C43156 a_7499_43078# a_8791_42308# 0.001313f
C43157 a_5891_43370# a_2982_43646# 5.95e-19
C43158 a_1307_43914# a_10835_43094# 3.58e-20
C43159 a_10334_44484# a_9803_43646# 5.26e-20
C43160 a_n356_44636# a_6547_43396# 9.65e-22
C43161 a_13720_44458# a_8685_43396# 1.78e-22
C43162 a_10440_44484# a_9145_43396# 2.03e-20
C43163 a_13213_44734# VDD 0.184239f
C43164 a_n3565_38216# C3_P_btm 0.001023f
C43165 a_n4209_38502# VREF 0.059621f
C43166 a_n3565_38502# VIN_P 0.029053f
C43167 a_2711_45572# a_10490_45724# 0.036939f
C43168 a_6472_45840# a_7499_43078# 2.82e-21
C43169 a_6667_45809# a_8162_45546# 1.87e-19
C43170 a_3539_42460# a_4646_46812# 1.05e-20
C43171 a_14358_43442# a_n2293_46634# 0.008808f
C43172 a_17499_43370# a_12549_44172# 1.62e-19
C43173 a_9165_43940# a_3090_45724# 0.006052f
C43174 a_14621_43646# a_13661_43548# 1.53e-19
C43175 a_9159_44484# a_8049_45260# 1.3e-21
C43176 a_11967_42832# a_10809_44734# 7.41e-21
C43177 a_20447_31679# a_19864_35138# 1.11e-20
C43178 a_8492_46660# VDD 0.273866f
C43179 a_n4064_38528# a_n3565_38216# 0.028041f
C43180 a_13258_32519# C3_N_btm 2.18e-19
C43181 a_7174_31319# C0_N_btm 0.050478f
C43182 a_n3674_37592# a_n4334_37440# 0.050036f
C43183 a_6123_31319# a_n3420_37984# 0.00363f
C43184 a_n1630_35242# a_8530_39574# 7.09e-20
C43185 a_22400_42852# a_22469_40625# 0.954861f
C43186 a_n2293_46634# a_1848_45724# 0.002657f
C43187 a_n743_46660# a_n1099_45572# 0.108295f
C43188 a_8667_46634# a_8034_45724# 0.001019f
C43189 a_n1925_46634# a_n357_42282# 5.15e-20
C43190 a_15227_44166# a_17715_44484# 0.385336f
C43191 a_12816_46660# a_6945_45028# 3.52e-20
C43192 a_12251_46660# a_10809_44734# 0.023146f
C43193 a_765_45546# a_5164_46348# 6.42e-20
C43194 a_15682_43940# a_16409_43396# 0.007432f
C43195 a_18079_43940# a_16137_43396# 1.32e-20
C43196 a_n1352_43396# a_n229_43646# 2.37e-19
C43197 a_5891_43370# a_5837_42852# 0.010625f
C43198 a_15493_43396# a_15781_43660# 0.047833f
C43199 a_11967_42832# a_13460_43230# 0.038517f
C43200 a_11341_43940# a_12281_43396# 0.002178f
C43201 en_comp a_1343_38525# 0.038003f
C43202 a_n2956_37592# a_n4209_39304# 0.102982f
C43203 a_104_43370# VDD 0.252393f
C43204 a_20841_45814# a_20885_45572# 3.69e-19
C43205 a_20623_45572# a_20719_45572# 0.013793f
C43206 a_18479_45785# a_n2017_45002# 8.68e-20
C43207 a_20107_45572# a_2437_43646# 3.54e-19
C43208 a_15037_45618# a_6171_45002# 6.48e-20
C43209 a_7227_45028# a_7735_45067# 1.1e-19
C43210 a_6511_45714# a_n2661_43370# 6.25e-20
C43211 a_20273_45572# a_21513_45002# 2.44e-19
C43212 a_21259_43561# a_20202_43084# 1.84e-19
C43213 a_16823_43084# a_12741_44636# 0.00226f
C43214 a_12379_42858# a_3090_45724# 0.00513f
C43215 a_4699_43561# a_n1925_42282# 5.23e-20
C43216 a_3080_42308# a_526_44458# 0.041925f
C43217 a_9803_43646# a_9290_44172# 0.010228f
C43218 a_6031_43396# a_6945_45028# 3.75e-20
C43219 a_10341_43396# a_8016_46348# 0.00203f
C43220 a_5932_42308# a_n2312_39304# 4.36e-21
C43221 a_10533_42308# a_10227_46804# 0.001306f
C43222 a_15051_42282# a_12861_44030# 4e-21
C43223 a_5210_46155# VDD 6.34e-20
C43224 a_13904_45546# a_6151_47436# 3.01e-22
C43225 a_18985_46122# a_20009_46494# 2.36e-20
C43226 a_19553_46090# a_19597_46482# 3.69e-19
C43227 a_10809_44734# a_13259_45724# 1.7e-19
C43228 a_5066_45546# a_6633_46155# 0.001122f
C43229 a_7845_44172# a_6123_31319# 1.02e-21
C43230 a_n2661_42282# a_2903_42308# 2.11e-19
C43231 a_2982_43646# a_17595_43084# 3.45e-20
C43232 a_19268_43646# a_743_42282# 7.11e-21
C43233 a_15743_43084# a_20556_43646# 2.78e-21
C43234 a_17324_43396# a_4361_42308# 8.49e-21
C43235 a_15037_45618# a_14673_44172# 1.11e-21
C43236 a_11963_45334# a_11691_44458# 1.33e-19
C43237 a_9482_43914# a_11827_44484# 0.031913f
C43238 a_117_45144# a_n2661_43370# 4.07e-19
C43239 a_8696_44636# a_15463_44811# 3.4e-19
C43240 a_n37_45144# a_n699_43396# 4.14e-19
C43241 a_1667_45002# a_949_44458# 0.008156f
C43242 a_5111_44636# a_n2661_44458# 0.048314f
C43243 a_n913_45002# a_10334_44484# 2.34e-21
C43244 a_n1059_45260# a_10440_44484# 7.97e-22
C43245 a_n2017_45002# a_10057_43914# 5.16e-20
C43246 a_13575_42558# a_13059_46348# 3.09e-21
C43247 a_13460_43230# a_13259_45724# 0.015281f
C43248 a_685_42968# a_n357_42282# 0.004355f
C43249 a_3681_42891# a_n863_45724# 4.05e-19
C43250 a_7309_43172# a_526_44458# 0.003264f
C43251 a_n1423_42826# a_n443_42852# 1.28e-19
C43252 a_421_43172# a_n755_45592# 1.37e-20
C43253 a_n3690_37440# SMPL_ON_P 1.8e-19
C43254 a_16680_45572# a_6755_46942# 9.94e-21
C43255 a_n913_45002# a_n1021_46688# 2.23e-21
C43256 a_n2017_45002# a_n2438_43548# 0.29197f
C43257 a_413_45260# a_21588_30879# 0.041669f
C43258 a_n967_45348# a_n2442_46660# 1.82e-19
C43259 en_comp a_n2293_46634# 0.00109f
C43260 a_n2810_45028# a_n2312_38680# 0.044149f
C43261 a_n2840_44458# SMPL_ON_P 8.99e-19
C43262 a_n2267_44484# a_n2497_47436# 0.025633f
C43263 a_22521_39511# VDD 0.910209f
C43264 a_13105_45348# a_12861_44030# 3.05e-19
C43265 a_n1641_43230# a_n4318_38216# 6.62e-19
C43266 a_n2157_42858# a_n4318_37592# 1.43e-19
C43267 a_n1853_43023# a_n1736_42282# 0.004594f
C43268 a_10922_42852# a_11136_42852# 0.097745f
C43269 a_12089_42308# a_12800_43218# 0.15794f
C43270 a_743_42282# a_1755_42282# 0.058846f
C43271 a_14205_43396# a_14456_42282# 1.85e-20
C43272 a_3626_43646# a_7174_31319# 0.022247f
C43273 a_12379_42858# a_12991_43230# 3.82e-19
C43274 a_14209_32519# a_n784_42308# 0.004411f
C43275 a_n4318_39304# a_n3690_39392# 8.45e-19
C43276 a_n746_45260# a_768_44030# 0.005354f
C43277 a_2952_47436# a_n1613_43370# 2.81e-19
C43278 a_2905_45572# a_3411_47243# 0.005614f
C43279 a_n1151_42308# a_5063_47570# 1.74e-19
C43280 a_n1435_47204# a_13507_46334# 1.53e-21
C43281 a_11599_46634# a_18597_46090# 0.191253f
C43282 a_13717_47436# a_21177_47436# 6.95e-20
C43283 a_11459_47204# a_4883_46098# 2.08e-20
C43284 a_16241_47178# a_10227_46804# 0.022072f
C43285 a_16327_47482# a_17591_47464# 0.339529f
C43286 a_16023_47582# a_16588_47582# 7.99e-20
C43287 a_15673_47210# a_18143_47464# 3.18e-20
C43288 a_n2946_39866# VDD 0.393552f
C43289 a_n2293_43922# VDAC_P 6.46e-20
C43290 a_n2017_45002# a_14021_43940# 1.77e-19
C43291 a_413_45260# a_15493_43940# 0.013529f
C43292 a_11691_44458# a_18588_44850# 0.00186f
C43293 a_1307_43914# a_1241_44260# 7.06e-19
C43294 a_2711_45572# a_16547_43609# 4.49e-19
C43295 a_n2293_42834# a_1115_44172# 9.47e-21
C43296 a_5883_43914# a_5708_44484# 2.58e-19
C43297 a_11827_44484# a_20159_44458# 0.012941f
C43298 a_7499_43078# a_10695_43548# 0.124597f
C43299 a_5518_44484# a_n2661_42834# 1.65e-20
C43300 a_5343_44458# a_n2661_43922# 0.094786f
C43301 a_21101_45002# a_20640_44752# 4.25e-19
C43302 a_21005_45260# a_20679_44626# 2.52e-20
C43303 a_18184_42460# a_19279_43940# 0.132218f
C43304 a_18587_45118# a_18579_44172# 8.05e-19
C43305 a_10775_45002# a_10405_44172# 1.45e-20
C43306 a_14113_42308# a_n357_42282# 5.29e-20
C43307 a_n3565_38502# a_n2956_38680# 0.302523f
C43308 a_16223_45938# VDD 0.132317f
C43309 a_5342_30871# C8_P_btm 0.093874f
C43310 a_5534_30871# C6_P_btm 0.01116f
C43311 a_1307_43914# a_11415_45002# 0.001965f
C43312 a_15415_45028# a_12741_44636# 1.4e-19
C43313 a_3537_45260# a_4185_45028# 1.06643f
C43314 a_4558_45348# a_3483_46348# 0.068916f
C43315 a_17719_45144# a_15227_44166# 0.187414f
C43316 a_5883_43914# a_5257_43370# 0.019234f
C43317 a_5891_43370# a_2107_46812# 1.37e-20
C43318 a_n2661_43922# a_n2956_39768# 1.22e-20
C43319 a_16922_45042# a_19692_46634# 0.055961f
C43320 a_n2661_42834# a_n2661_46634# 1.68e-20
C43321 a_16680_45572# a_8049_45260# 0.005473f
C43322 a_7499_43078# a_n357_42282# 0.259858f
C43323 a_11967_42832# a_n881_46662# 9.73e-21
C43324 a_3357_43084# a_2324_44458# 0.216574f
C43325 a_21363_45546# a_21137_46414# 0.001589f
C43326 a_20623_45572# a_6945_45028# 5.77e-19
C43327 a_n913_45002# a_9290_44172# 0.632534f
C43328 a_2437_43646# a_17715_44484# 3.38e-20
C43329 a_1606_42308# a_6171_42473# 1.34e-20
C43330 a_1755_42282# a_5755_42308# 4.89e-19
C43331 a_1067_42314# a_6123_31319# 9e-21
C43332 a_564_42282# a_5934_30871# 2.52e-20
C43333 a_4190_30871# C4_N_btm 1.36e-19
C43334 a_22545_38993# a_22821_38993# 0.235701f
C43335 a_22521_39511# a_22469_39537# 1.02751f
C43336 a_22521_40055# CAL_P 0.001469f
C43337 a_13747_46662# a_6755_46942# 0.316914f
C43338 a_n2661_46634# a_8145_46902# 0.008097f
C43339 a_2107_46812# a_4817_46660# 0.002361f
C43340 a_2609_46660# a_3067_47026# 0.027317f
C43341 a_2959_46660# a_3524_46660# 7.99e-20
C43342 a_n2661_46098# a_1302_46660# 2.6e-19
C43343 a_n1925_46634# a_5263_46660# 8.56e-19
C43344 a_13507_46334# a_13885_46660# 5.84e-20
C43345 a_11599_46634# a_19123_46287# 0.024241f
C43346 a_15673_47210# a_765_45546# 0.028544f
C43347 a_15811_47375# a_17829_46910# 2.1e-20
C43348 a_13717_47436# a_20841_46902# 1.67e-20
C43349 a_n2497_47436# a_3699_46348# 6.3e-22
C43350 a_n2109_47186# a_3147_46376# 5.93e-20
C43351 a_n1741_47186# a_2698_46116# 9.05e-21
C43352 a_n971_45724# a_1138_42852# 1.34e-20
C43353 a_327_47204# a_376_46348# 1.5e-19
C43354 a_n237_47217# a_1208_46090# 0.003284f
C43355 a_n746_45260# a_1176_45822# 3.33e-20
C43356 a_4743_44484# a_n97_42460# 1.46e-20
C43357 a_n984_44318# a_453_43940# 3.53e-20
C43358 a_16241_44734# a_15682_43940# 2.85e-19
C43359 a_n699_43396# a_104_43370# 0.21575f
C43360 a_18479_45785# a_19164_43230# 0.001979f
C43361 a_175_44278# a_1414_42308# 1.49e-20
C43362 a_n2661_42834# a_9895_44260# 2.38e-19
C43363 a_n913_45002# a_791_42968# 0.054288f
C43364 a_n1059_45260# a_1847_42826# 0.038913f
C43365 a_5700_37509# VDD 1.0734f
C43366 a_949_44458# VDD 1.2275f
C43367 a_7174_31319# C10_P_btm 1.34e-19
C43368 a_n4315_30879# a_n1386_35608# 1.11e-19
C43369 a_n3690_38304# a_n2956_38216# 0.016795f
C43370 a_n4064_37984# a_n2810_45572# 0.094405f
C43371 a_18579_44172# a_11415_45002# 2.58e-23
C43372 a_19279_43940# a_12741_44636# 6.8e-19
C43373 a_3737_43940# a_3877_44458# 1.04e-19
C43374 a_1891_43646# a_768_44030# 5.62e-19
C43375 a_n2661_43370# a_n755_45592# 0.036276f
C43376 a_10057_43914# a_526_44458# 3.21e-19
C43377 a_n2661_42834# a_8199_44636# 0.032396f
C43378 a_9313_44734# a_10903_43370# 0.030402f
C43379 a_9159_44484# a_8953_45546# 0.004058f
C43380 a_5826_44734# a_2324_44458# 9.11e-19
C43381 a_5649_42852# a_n971_45724# 7.13e-21
C43382 a_n4064_39616# a_n2302_39866# 0.239588f
C43383 a_n4315_30879# a_n3420_39072# 0.036979f
C43384 a_n4064_40160# a_n3565_39304# 0.028096f
C43385 a_n4334_39616# a_n4251_39616# 0.007692f
C43386 a_n2946_39866# a_n2860_39866# 0.011479f
C43387 a_n4209_39590# a_n3607_39616# 0.002294f
C43388 a_16750_47204# VDD 6.26e-19
C43389 a_5932_42308# C0_N_btm 0.015561f
C43390 a_17609_46634# a_11415_45002# 5.34e-21
C43391 a_16388_46812# a_765_45546# 0.164902f
C43392 a_16721_46634# a_17339_46660# 0.005637f
C43393 a_15227_44166# a_22365_46825# 3.68e-20
C43394 a_12549_44172# a_12638_46436# 3.01e-19
C43395 a_13747_46662# a_8049_45260# 0.208778f
C43396 a_n2438_43548# a_526_44458# 0.107408f
C43397 a_n743_46660# a_n1925_42282# 0.010043f
C43398 a_12891_46348# a_14180_46482# 1.22e-21
C43399 a_5807_45002# a_9823_46482# 2.88e-19
C43400 a_7927_46660# a_8349_46414# 0.01072f
C43401 a_7577_46660# a_5937_45572# 2.93e-19
C43402 a_8667_46634# a_8016_46348# 1.13e-19
C43403 a_3877_44458# a_2324_44458# 0.153319f
C43404 a_n881_46662# a_13259_45724# 0.507296f
C43405 a_n2017_45002# a_15764_42576# 0.014981f
C43406 a_n1059_45260# a_15486_42560# 2.84e-20
C43407 a_n913_45002# a_15051_42282# 0.003302f
C43408 a_5111_44636# a_8325_42308# 6.44e-22
C43409 a_n2661_42834# a_n1379_43218# 1.92e-19
C43410 a_742_44458# a_945_42968# 4.68e-20
C43411 a_14539_43914# a_17595_43084# 0.141972f
C43412 a_n356_44636# a_12379_42858# 8.61e-20
C43413 a_n2661_42282# a_6293_42852# 0.16527f
C43414 a_5891_43370# a_7871_42858# 0.051552f
C43415 a_11341_43940# VDD 1.23655f
C43416 a_15599_45572# a_18175_45572# 4.17e-21
C43417 a_16115_45572# a_16211_45572# 0.013793f
C43418 a_16333_45814# a_16377_45572# 3.69e-19
C43419 a_15903_45785# a_16147_45260# 0.003162f
C43420 a_15765_45572# a_17786_45822# 1.13e-19
C43421 a_5907_45546# a_5111_44636# 0.01337f
C43422 a_5263_45724# a_4927_45028# 0.001784f
C43423 a_2711_45572# a_6171_45002# 0.457554f
C43424 a_3260_45572# a_413_45260# 4.87e-19
C43425 a_1427_43646# a_1138_42852# 7.47e-20
C43426 a_15743_43084# a_19692_46634# 5.26e-19
C43427 a_8605_42826# a_4646_46812# 9.01e-21
C43428 a_2998_44172# a_n755_45592# 5.92e-21
C43429 a_n3674_39768# a_n2810_45572# 0.023119f
C43430 CAL_N a_22521_40055# 6.29e-19
C43431 a_22521_40599# a_22780_40945# 0.009658f
C43432 a_3726_37500# CAL_P 0.102027f
C43433 a_5497_46414# VDD 0.200657f
C43434 a_6194_45824# a_n2109_47186# 1.26e-19
C43435 a_n3420_39616# VDAC_P 0.005053f
C43436 a_13059_46348# a_n443_42852# 0.09278f
C43437 a_8199_44636# a_5066_45546# 0.178583f
C43438 a_18819_46122# a_6945_45028# 4.66e-20
C43439 a_19335_46494# a_19900_46494# 7.99e-20
C43440 a_18985_46122# a_21137_46414# 5.31e-20
C43441 a_18189_46348# a_10809_44734# 8.9e-20
C43442 a_n3565_39304# a_n4064_37440# 0.028266f
C43443 a_n4064_39072# a_n3565_37414# 0.031386f
C43444 a_n3420_39072# a_n3420_37440# 0.052876f
C43445 a_n1761_44111# a_n4318_37592# 1.64e-20
C43446 a_n1899_43946# a_n1736_42282# 5.43e-21
C43447 a_2982_43646# a_13467_32519# 0.006898f
C43448 a_14021_43940# a_19164_43230# 1.26e-20
C43449 a_9313_44734# a_15959_42545# 6.1e-20
C43450 a_14358_43442# a_14537_43646# 0.010303f
C43451 a_14579_43548# a_14621_43646# 8.44e-19
C43452 a_10341_43396# a_12281_43396# 0.012652f
C43453 a_9145_43396# a_13837_43396# 4.66e-20
C43454 a_n97_42460# a_n1736_43218# 7.3e-22
C43455 a_n356_44636# a_18727_42674# 2.05e-20
C43456 a_n4318_40392# a_n3420_39072# 7.42e-22
C43457 a_3080_42308# a_14209_32519# 0.001913f
C43458 a_n2012_43396# a_n3674_39304# 8.64e-20
C43459 a_3094_47570# DATA[2] 6.24e-20
C43460 a_3315_47570# DATA[1] 1.79e-21
C43461 a_22612_30879# a_22521_39511# 9.02e-20
C43462 a_n1076_43230# VDD 0.292942f
C43463 a_n2810_45028# a_n2661_43370# 0.002593f
C43464 a_3065_45002# a_5009_45028# 6.35e-21
C43465 a_21188_45572# a_21101_45002# 3.83e-19
C43466 a_20731_45938# a_20567_45036# 1.28e-19
C43467 a_8953_45002# a_1423_45028# 0.011739f
C43468 a_21363_45546# a_21359_45002# 0.01738f
C43469 a_20623_45572# a_11827_44484# 1.21e-20
C43470 a_18953_45572# a_11691_44458# 2.11e-20
C43471 a_8746_45002# a_9313_44734# 2.85e-19
C43472 a_2711_45572# a_14673_44172# 0.04263f
C43473 a_9482_43914# a_15595_45028# 0.0011f
C43474 a_13556_45296# a_15415_45028# 1.78e-20
C43475 a_14180_45002# a_14537_43396# 0.143922f
C43476 a_n2302_40160# a_n2312_38680# 4.94e-19
C43477 a_n3690_39616# a_n2956_39768# 0.015398f
C43478 a_n4209_39590# a_n2442_46660# 0.095025f
C43479 a_15095_43370# a_n443_42852# 0.006819f
C43480 a_15781_43660# a_n357_42282# 6.97e-20
C43481 a_2075_43172# a_526_44458# 0.227071f
C43482 a_1847_42826# a_n1925_42282# 2.13e-20
C43483 a_15599_45572# a_n743_46660# 0.022482f
C43484 a_18596_45572# a_12549_44172# 1.55e-20
C43485 a_6667_45809# a_6969_46634# 1.42e-19
C43486 a_6598_45938# a_6755_46942# 2.16e-20
C43487 a_2437_43646# a_2487_47570# 0.001086f
C43488 a_n2017_45002# a_13507_46334# 5.63e-19
C43489 a_413_45260# a_16763_47508# 3.7e-19
C43490 en_comp a_18597_46090# 3.29e-20
C43491 a_13017_45260# a_4915_47217# 0.002063f
C43492 a_6171_45002# a_9313_45822# 1.31e-19
C43493 a_375_42282# a_584_46384# 0.480677f
C43494 a_3602_45348# a_n971_45724# 0.003621f
C43495 a_n755_45592# a_2307_45899# 9.75e-21
C43496 a_n1099_45572# a_509_45572# 0.001017f
C43497 a_380_45546# a_603_45572# 0.011458f
C43498 a_16137_43396# a_17749_42852# 0.001147f
C43499 a_3080_42308# a_4169_42308# 0.001081f
C43500 a_n13_43084# a_133_42852# 0.171361f
C43501 a_n97_42460# a_11633_42558# 0.011546f
C43502 a_3626_43646# a_5932_42308# 0.062334f
C43503 a_10341_42308# a_12089_42308# 0.003265f
C43504 a_18525_43370# a_18504_43218# 6.38e-19
C43505 a_22365_46825# EN_OFFSET_CAL 0.195393f
C43506 a_5088_37509# VDAC_P 1.15441f
C43507 a_3726_37500# CAL_N 0.036205f
C43508 a_4338_37500# a_11206_38545# 0.072616f
C43509 a_6886_37412# VDAC_N 0.067053f
C43510 a_5700_37509# a_8912_37509# 15.051701f
C43511 a_3422_30871# C0_dummy_N_btm 1.28e-20
C43512 a_10723_42308# VDD 0.223902f
C43513 a_n1741_47186# a_n1435_47204# 0.047534f
C43514 a_n237_47217# a_6575_47204# 0.0275f
C43515 a_2063_45854# a_4915_47217# 0.055521f
C43516 a_2905_45572# a_4700_47436# 4.48e-20
C43517 a_n1151_42308# a_3815_47204# 0.01223f
C43518 a_3381_47502# a_3785_47178# 0.00589f
C43519 a_2553_47502# a_n443_46116# 1.33e-19
C43520 a_1307_43914# a_11967_42832# 0.031135f
C43521 a_949_44458# a_n699_43396# 1.66e-19
C43522 a_n2661_44458# a_10334_44484# 0.009408f
C43523 a_11691_44458# a_18443_44721# 0.042634f
C43524 a_13249_42308# a_13565_43940# 0.048533f
C43525 a_327_44734# a_644_44056# 1.79e-19
C43526 a_n913_45002# a_3905_42865# 5e-19
C43527 a_n2017_45002# a_5013_44260# 1.47e-20
C43528 a_n1059_45260# a_5244_44056# 4.98e-21
C43529 a_n1329_42308# a_n357_42282# 7.05e-20
C43530 a_n1630_35242# a_n2956_38216# 4.4e-19
C43531 COMP_P a_n755_45592# 1.75e-21
C43532 a_16823_43084# RST_Z 5.98e-22
C43533 a_4190_30871# C6_P_btm 0.005085f
C43534 a_13678_32519# EN_VIN_BSTR_N 0.031779f
C43535 a_21513_45002# a_20202_43084# 0.13666f
C43536 a_n2840_44458# a_n2438_43548# 0.00955f
C43537 a_13720_44458# a_768_44030# 0.178939f
C43538 a_15004_44636# a_12549_44172# 3.69e-20
C43539 a_5883_43914# a_5807_45002# 0.002403f
C43540 a_20885_45572# a_11415_45002# 4.28e-19
C43541 a_10180_45724# a_526_44458# 4e-22
C43542 a_6598_45938# a_8049_45260# 2.14e-19
C43543 a_2437_43646# a_22365_46825# 0.001459f
C43544 a_15143_45578# a_10809_44734# 1.76e-21
C43545 a_8696_44636# a_5937_45572# 0.041815f
C43546 a_9159_45572# a_2324_44458# 0.003342f
C43547 a_n2012_44484# a_n1613_43370# 2.46e-19
C43548 a_9313_44734# a_4883_46098# 0.015767f
C43549 a_n2661_43922# a_10227_46804# 0.041913f
C43550 a_n2065_43946# a_n2497_47436# 0.036632f
C43551 a_n3674_39304# a_n4064_39616# 0.020873f
C43552 a_n1151_42308# a_14976_45028# 1.72e-19
C43553 a_13661_43548# a_n2293_46634# 0.055067f
C43554 a_20916_46384# a_21588_30879# 5.25e-19
C43555 a_4915_47217# a_12469_46902# 5.76e-19
C43556 a_6575_47204# a_8270_45546# 9.19e-20
C43557 a_6151_47436# a_11735_46660# 1.81e-19
C43558 a_11599_46634# a_6755_46942# 0.321942f
C43559 a_4883_46098# a_5072_46660# 7.49e-20
C43560 a_n1613_43370# a_n2661_46098# 1.40554f
C43561 a_n881_46662# a_1799_45572# 0.028083f
C43562 a_5111_44636# a_9145_43396# 0.057312f
C43563 a_n2293_42834# a_n2012_43396# 0.001738f
C43564 a_10193_42453# a_19339_43156# 0.003128f
C43565 a_1307_43914# a_648_43396# 6.76e-20
C43566 a_n2661_43370# a_n2129_43609# 3.94e-19
C43567 a_n2661_42834# a_2127_44172# 0.019594f
C43568 a_3363_44484# a_3600_43914# 4.63e-19
C43569 a_n2661_43922# a_453_43940# 0.006118f
C43570 a_20640_44752# a_20766_44850# 0.17072f
C43571 a_20362_44736# a_19279_43940# 0.039759f
C43572 a_20679_44626# a_20835_44721# 0.105995f
C43573 a_11967_42832# a_18579_44172# 0.158329f
C43574 a_13249_42308# a_5534_30871# 0.215947f
C43575 a_13720_44458# a_13483_43940# 0.001108f
C43576 a_20692_30879# C1_N_btm 1.3e-20
C43577 a_5932_42308# C10_P_btm 1.34e-19
C43578 a_6123_31319# EN_VIN_BSTR_N 0.050716f
C43579 a_1606_42308# VIN_N 0.014401f
C43580 a_9838_44484# a_3483_46348# 0.014242f
C43581 a_20679_44626# a_3090_45724# 5.62e-22
C43582 a_1307_43914# a_13259_45724# 0.023098f
C43583 a_2382_45260# a_3316_45546# 0.052075f
C43584 a_3065_45002# a_2957_45546# 4.26e-19
C43585 a_n659_45366# a_n443_42852# 1.08e-19
C43586 a_11827_44484# a_18819_46122# 1.7e-21
C43587 a_18494_42460# a_19900_46494# 0.001134f
C43588 a_11691_44458# a_17583_46090# 3.92e-21
C43589 a_n2661_44458# a_9290_44172# 0.027487f
C43590 a_5343_44458# a_5164_46348# 3.87e-20
C43591 a_8685_43396# a_n971_45724# 0.079658f
C43592 a_7287_43370# a_n1151_42308# 2.15e-20
C43593 a_16327_47482# VDD 2.81451f
C43594 a_4958_30871# a_18220_42308# 6.64e-20
C43595 a_6123_31319# a_1239_39043# 6.84e-20
C43596 a_17303_42282# a_18214_42558# 7.99e-21
C43597 a_n743_46660# a_2698_46116# 0.013101f
C43598 a_n2661_46098# a_n2293_46098# 0.063852f
C43599 a_n1925_46634# a_3147_46376# 1.66e-19
C43600 a_n2438_43548# a_2521_46116# 5.14e-19
C43601 a_1123_46634# a_1208_46090# 0.0037f
C43602 a_n133_46660# a_167_45260# 5.4e-22
C43603 a_n2293_46634# a_4185_45028# 0.027799f
C43604 a_2107_46812# a_472_46348# 2.45e-19
C43605 a_15009_46634# a_3090_45724# 0.154981f
C43606 a_8145_46902# a_765_45546# 1.38e-20
C43607 a_6755_46942# a_13693_46688# 0.001956f
C43608 a_768_44030# a_13351_46090# 1.3e-19
C43609 a_12549_44172# a_13759_46122# 5.27e-19
C43610 a_5807_45002# a_9569_46155# 2.47e-19
C43611 a_n2661_46634# a_5068_46348# 3.78e-20
C43612 a_12891_46348# a_13925_46122# 2.71e-21
C43613 a_8128_46384# a_2324_44458# 2.07e-20
C43614 a_n881_46662# a_18189_46348# 2.07e-20
C43615 a_11599_46634# a_8049_45260# 0.14064f
C43616 a_4915_47217# a_14383_46116# 9.48e-19
C43617 a_n1435_47204# a_10586_45546# 4.56e-21
C43618 a_n237_47217# a_n2661_45546# 0.038356f
C43619 a_n2497_47436# a_n755_45592# 0.45034f
C43620 a_n815_47178# a_n1079_45724# 7.01e-21
C43621 a_n971_45724# a_n2956_38216# 1.71e-19
C43622 a_15433_44458# a_14955_43396# 1.98e-19
C43623 a_1414_42308# a_n97_42460# 0.196768f
C43624 a_18079_43940# a_14021_43940# 4.92e-20
C43625 a_11341_43940# a_22959_43948# 4.69e-19
C43626 a_22223_43948# a_15493_43940# 0.051823f
C43627 a_9313_44734# a_16243_43396# 1.87e-19
C43628 a_n699_43396# a_n1076_43230# 0.001631f
C43629 a_n2293_43922# a_12281_43396# 0.147288f
C43630 a_14955_43940# a_15301_44260# 0.013377f
C43631 a_6756_44260# a_6671_43940# 1.48e-19
C43632 a_18989_43940# a_19177_43646# 1.57e-19
C43633 a_18443_44721# a_4190_30871# 3.98e-20
C43634 a_n2293_42834# a_n914_42852# 1.34e-19
C43635 a_n913_45002# a_n961_42308# 9.71e-19
C43636 a_n1059_45260# a_n473_42460# 8.15e-19
C43637 en_comp a_n1736_42282# 6.61e-20
C43638 a_n2017_45002# a_196_42282# 0.010023f
C43639 a_n2956_37592# a_n4318_37592# 0.023082f
C43640 a_n967_45348# a_n3674_38216# 3.49e-20
C43641 a_n2810_45028# COMP_P 1.61e-21
C43642 a_175_44278# VDD 0.20887f
C43643 a_11652_45724# a_11688_45572# 0.001673f
C43644 a_11525_45546# a_11778_45572# 0.011913f
C43645 C0_dummy_P_btm VCM 0.311452f
C43646 C0_N_btm VREF 0.443884f
C43647 C1_N_btm VIN_N 0.39234f
C43648 a_5829_43940# a_n2293_46098# 0.05512f
C43649 a_6765_43638# a_3090_45724# 0.002105f
C43650 a_5111_42852# a_768_44030# 3.09e-21
C43651 a_n1853_43023# a_n2442_46660# 2.67e-21
C43652 a_18579_44172# a_13259_45724# 5.71e-20
C43653 a_5013_44260# a_526_44458# 3.48e-20
C43654 a_9672_43914# a_2324_44458# 1.42e-19
C43655 a_10835_43094# a_n1613_43370# 7.12e-22
C43656 a_19164_43230# a_13507_46334# 1.15e-20
C43657 a_16434_46987# VDD 0.001765f
C43658 a_5742_30871# a_6886_37412# 3.23e-19
C43659 a_17609_46634# a_13259_45724# 9.09e-19
C43660 a_20202_43084# a_10809_44734# 0.014133f
C43661 a_11415_45002# a_22223_46124# 0.011454f
C43662 a_3483_46348# a_9823_46155# 2.75e-19
C43663 a_n2293_43922# a_n3674_38680# 2.31e-20
C43664 a_6293_42852# a_7112_43396# 5.47e-21
C43665 a_3626_43646# a_4181_43396# 2.16e-20
C43666 a_18184_42460# a_19332_42282# 0.042769f
C43667 a_18494_42460# a_18907_42674# 0.11494f
C43668 a_n97_42460# a_12281_43396# 6.17e-19
C43669 a_5883_43914# a_9223_42460# 2.74e-20
C43670 a_n356_44636# a_3823_42558# 1.46e-19
C43671 a_3539_42460# a_3457_43396# 2.02e-20
C43672 a_9028_43914# a_9127_43156# 9.19e-20
C43673 a_n2661_42834# a_n4318_38216# 0.023647f
C43674 a_14021_43940# a_14209_32519# 0.042544f
C43675 a_6031_43396# a_8147_43396# 3.33e-21
C43676 a_6765_43638# a_6547_43396# 0.209641f
C43677 a_6197_43396# a_7287_43370# 0.041762f
C43678 a_2905_45572# DATA[2] 5.19e-19
C43679 a_n1151_42308# DATA[0] 0.088597f
C43680 a_3160_47472# DATA[1] 8.03e-22
C43681 a_2063_45854# DATA[5] 0.001488f
C43682 a_19479_31679# C2_N_btm 0.001057f
C43683 a_10341_43396# VDD 0.401264f
C43684 a_6511_45714# a_5883_43914# 1.33e-21
C43685 a_13249_42308# a_11691_44458# 0.017891f
C43686 a_7227_45028# a_6298_44484# 0.003074f
C43687 a_2711_45572# a_12607_44458# 8.18e-21
C43688 a_9049_44484# a_n2661_44458# 0.015549f
C43689 a_n1059_45260# a_5111_44636# 0.038143f
C43690 a_3935_42891# a_1823_45246# 0.002482f
C43691 a_12800_43218# a_3090_45724# 0.002125f
C43692 a_1568_43370# a_n755_45592# 7.31e-20
C43693 a_n1177_43370# a_n443_42852# 1.95e-19
C43694 a_743_42282# a_2324_44458# 8.04e-21
C43695 a_7174_31319# a_n2312_40392# 6.67e-21
C43696 a_n356_45724# VDD 0.719282f
C43697 a_11525_45546# a_768_44030# 1.76e-21
C43698 a_3775_45552# a_n2661_46634# 1.47e-21
C43699 a_5263_45724# a_n743_46660# 7.27e-19
C43700 a_11962_45724# a_12891_46348# 0.001251f
C43701 a_11652_45724# a_12549_44172# 6.46e-20
C43702 a_15143_45578# a_n881_46662# 0.069805f
C43703 a_15037_45618# a_4883_46098# 7.22e-21
C43704 a_17478_45572# a_10227_46804# 8.9e-22
C43705 a_n2810_45028# a_n2497_47436# 9.88e-21
C43706 a_2437_43646# a_584_46384# 0.302508f
C43707 a_16137_43396# a_19339_43156# 2.87e-19
C43708 a_15682_43940# a_15890_42674# 1.13e-19
C43709 a_n1699_43638# a_n1736_42282# 7.33e-20
C43710 a_n2433_43396# a_n1329_42308# 3.94e-21
C43711 a_17324_43396# a_17595_43084# 6.75e-20
C43712 a_n2157_42858# a_n1533_42852# 9.73e-19
C43713 a_17499_43370# a_17701_42308# 8.78e-19
C43714 a_743_42282# a_8387_43230# 6e-20
C43715 a_15743_43084# a_5342_30871# 0.006894f
C43716 a_n2129_43609# COMP_P 2.54e-20
C43717 a_n1641_43230# a_n1545_43230# 0.013793f
C43718 a_n1423_42826# a_n1379_43218# 3.69e-19
C43719 a_n1991_42858# a_n967_43230# 2.36e-20
C43720 a_n1853_43023# a_n722_43218# 0.001894f
C43721 a_n1076_43230# a_n4318_38680# 1.6e-20
C43722 a_15368_46634# RST_Z 3.47e-20
C43723 a_11813_46116# CLK 2.07e-20
C43724 a_20356_42852# VDD 7.06e-19
C43725 a_3537_45260# a_5708_44484# 3.43e-20
C43726 a_2382_45260# a_n2661_42834# 0.055134f
C43727 a_3232_43370# a_9313_44734# 0.11426f
C43728 a_2274_45254# a_n2661_43922# 5.45e-20
C43729 a_21363_45546# a_19279_43940# 1.63e-19
C43730 a_18494_42460# a_21005_45260# 1.23e-20
C43731 a_19778_44110# a_21359_45002# 6.57e-19
C43732 a_10193_42453# a_17973_43940# 0.084505f
C43733 a_n2293_42834# a_2779_44458# 7.79e-21
C43734 a_n2661_43370# a_n2129_44697# 0.014856f
C43735 a_18184_42460# a_21101_45002# 2.52e-36
C43736 a_16922_45042# a_16237_45028# 3.82e-19
C43737 a_18911_45144# a_11827_44484# 4.77e-20
C43738 a_17613_45144# a_11691_44458# 5.83e-21
C43739 a_11823_42460# a_10949_43914# 0.002042f
C43740 a_n473_42460# a_n1925_42282# 1.12e-19
C43741 a_9885_42558# a_8199_44636# 0.009365f
C43742 a_8325_42308# a_9290_44172# 1.58e-20
C43743 a_9293_42558# a_8953_45546# 0.007436f
C43744 a_8568_45546# a_3483_46348# 0.137016f
C43745 a_17478_45572# a_17339_46660# 2.92e-22
C43746 a_15861_45028# a_765_45546# 0.004302f
C43747 a_19418_45938# a_19466_46812# 2.93e-19
C43748 a_2304_45348# a_2107_46812# 9.3e-21
C43749 a_2437_43646# a_11901_46660# 9.19e-20
C43750 a_413_45260# a_9863_46634# 1.44e-20
C43751 a_3537_45260# a_5257_43370# 0.001934f
C43752 a_7227_45028# a_5937_45572# 0.064518f
C43753 a_2711_45572# a_10903_43370# 0.213719f
C43754 a_4808_45572# a_5204_45822# 7.79e-20
C43755 a_n23_44458# a_n1151_42308# 0.101137f
C43756 a_4361_42308# a_11633_42308# 9.01e-19
C43757 a_5342_30871# a_1606_42308# 0.023615f
C43758 a_743_42282# a_16522_42674# 0.003239f
C43759 a_12800_43218# a_12991_43230# 4.61e-19
C43760 a_15743_43084# a_20107_42308# 1.94e-20
C43761 a_16823_43084# a_17303_42282# 3.24e-21
C43762 a_7227_42852# a_6761_42308# 4.22e-19
C43763 a_n2293_42282# a_n4318_38216# 0.004948f
C43764 a_19700_43370# a_19647_42308# 4.12e-19
C43765 a_2747_46873# a_n881_46662# 5.46e-20
C43766 a_12465_44636# a_15928_47570# 5.23e-20
C43767 a_11453_44696# a_11309_47204# 2.71e-19
C43768 a_10227_46804# a_19594_46812# 0.01518f
C43769 a_19386_47436# a_5807_45002# 2.36e-21
C43770 a_18597_46090# a_13661_43548# 0.266647f
C43771 a_18143_47464# a_19321_45002# 2.46e-20
C43772 a_18780_47178# a_13747_46662# 0.028845f
C43773 a_16588_47582# a_16750_47204# 0.006453f
C43774 a_18479_47436# a_19452_47524# 5.84e-19
C43775 a_n1435_47204# a_n743_46660# 2.75e-20
C43776 a_n971_45724# a_5907_46634# 3.23e-19
C43777 a_n443_46116# a_1799_45572# 0.081828f
C43778 a_n1151_42308# a_3524_46660# 4.19e-20
C43779 a_2905_45572# a_3067_47026# 1.43e-19
C43780 a_n2109_47186# a_5894_47026# 1.64e-19
C43781 a_949_44458# a_1467_44172# 0.004991f
C43782 a_18989_43940# a_18579_44172# 0.035827f
C43783 a_n2661_44458# a_3905_42865# 2.18e-19
C43784 a_n699_43396# a_175_44278# 0.001042f
C43785 a_742_44458# a_1414_42308# 0.052151f
C43786 a_18443_44721# a_18753_44484# 0.013793f
C43787 a_18374_44850# a_18681_44484# 3.69e-19
C43788 a_1307_43914# a_5745_43940# 0.001752f
C43789 a_n1059_45260# a_4235_43370# 0.003711f
C43790 a_n2017_45002# a_4699_43561# 1.2e-20
C43791 a_n913_45002# a_4093_43548# 4.03e-21
C43792 a_3357_43084# a_3539_42460# 0.001767f
C43793 a_n143_45144# VDD 0.092f
C43794 a_22400_42852# a_22609_38406# 1.37e-20
C43795 a_n2661_43370# a_3483_46348# 0.953959f
C43796 a_22223_45036# a_11415_45002# 0.011148f
C43797 a_21101_45002# a_12741_44636# 7.11e-19
C43798 a_18443_44721# a_15227_44166# 0.002052f
C43799 a_7542_44172# a_768_44030# 0.005732f
C43800 a_n1761_44111# a_n2293_46634# 4.77e-21
C43801 a_8696_44636# a_n443_42852# 8.12e-20
C43802 a_5111_44636# a_n1925_42282# 5.66e-21
C43803 a_5009_45028# a_5937_45572# 6.92e-20
C43804 a_13017_45260# a_10809_44734# 1.77e-20
C43805 a_14955_43940# a_12465_44636# 6.55e-20
C43806 a_19862_44208# a_18597_46090# 0.536021f
C43807 a_n2129_43609# a_n2497_47436# 0.216536f
C43808 a_10533_42308# a_11633_42558# 9.27e-21
C43809 a_11323_42473# a_5742_30871# 0.198522f
C43810 COMP_P a_n2302_40160# 4e-20
C43811 a_n3674_38680# a_n3420_39616# 0.020072f
C43812 a_5342_30871# C1_N_btm 9.04e-20
C43813 a_5534_30871# C3_N_btm 7.69e-20
C43814 C10_P_btm VREF 14.773f
C43815 C8_P_btm VIN_P 0.907642f
C43816 a_n746_45260# a_518_46482# 7.09e-19
C43817 a_n1741_47186# a_526_44458# 3.03e-20
C43818 a_2063_45854# a_10809_44734# 0.169005f
C43819 a_13747_46662# a_18285_46348# 1.64e-19
C43820 a_n2661_46634# a_13059_46348# 1.84e-19
C43821 a_13661_43548# a_19123_46287# 0.073049f
C43822 a_n743_46660# a_13885_46660# 1.96e-21
C43823 a_8492_46660# a_10150_46912# 0.00213f
C43824 a_7411_46660# a_6755_46942# 0.265786f
C43825 a_2959_46660# a_3090_45724# 4.18e-19
C43826 a_5807_45002# a_19551_46910# 1.7e-20
C43827 a_5257_43370# a_6969_46634# 6.29e-21
C43828 a_8667_46634# a_10428_46928# 6.23e-20
C43829 a_12549_44172# a_16434_46660# 2.11e-19
C43830 a_n1435_47204# a_11189_46129# 9.06e-22
C43831 a_6151_47436# a_2324_44458# 0.002957f
C43832 a_11459_47204# a_11387_46155# 1.29e-20
C43833 a_18597_46090# a_4185_45028# 1.12e-19
C43834 a_2382_45260# a_n2293_42282# 0.080755f
C43835 a_n2661_42834# a_n1655_43396# 2.44e-19
C43836 a_17730_32519# a_14021_43940# 9.75e-19
C43837 a_16922_45042# a_743_42282# 0.120316f
C43838 a_7499_43078# a_8685_42308# 7.11e-19
C43839 a_1423_45028# a_8037_42858# 1.11e-21
C43840 a_1307_43914# a_10518_42984# 3.51e-21
C43841 a_n2293_42834# a_n13_43084# 0.007462f
C43842 a_n2661_43370# a_n2840_42826# 3.35e-19
C43843 a_10334_44484# a_9145_43396# 1.97e-20
C43844 a_10157_44484# a_9803_43646# 0.001011f
C43845 a_n2293_43922# VDD 0.735248f
C43846 a_n3565_38216# C4_P_btm 9.91e-21
C43847 a_2711_45572# a_8746_45002# 0.010166f
C43848 a_6511_45714# a_8162_45546# 0.004311f
C43849 a_6598_45938# a_6812_45938# 0.097745f
C43850 a_6667_45809# a_7230_45938# 0.049827f
C43851 a_6472_45840# a_8568_45546# 3.47e-20
C43852 a_2998_44172# a_3483_46348# 2.54e-20
C43853 a_3626_43646# a_4646_46812# 4.2e-20
C43854 a_14579_43548# a_n2293_46634# 0.035629f
C43855 a_16759_43396# a_12549_44172# 1.5e-19
C43856 a_14537_43646# a_13661_43548# 1.89e-19
C43857 a_10341_43396# a_22612_30879# 1.26e-21
C43858 a_n2661_43922# a_8034_45724# 6.46e-21
C43859 a_5883_43914# a_n755_45592# 1.16e-19
C43860 a_14209_32519# a_13507_46334# 0.008866f
C43861 a_19963_31679# a_21589_35634# 1.55e-20
C43862 a_8667_46634# VDD 0.39254f
C43863 a_n4064_38528# a_n4334_38304# 0.001145f
C43864 a_n2302_38778# a_n4209_38216# 0.001254f
C43865 a_n2946_38778# a_n3565_38216# 0.001251f
C43866 a_1177_38525# a_2684_37794# 3.29e-20
C43867 a_7174_31319# C0_dummy_N_btm 0.029132f
C43868 a_13258_32519# C2_N_btm 2.75e-19
C43869 a_22400_42852# a_22521_40599# 0.133947f
C43870 a_n3674_37592# a_n4209_37414# 0.044977f
C43871 a_n1630_35242# a_7754_38470# 4.78e-20
C43872 a_n4318_37592# a_n2860_37690# 1.77e-20
C43873 a_7927_46660# a_8034_45724# 9e-20
C43874 a_n2293_46634# a_997_45618# 0.002767f
C43875 a_n1925_46634# a_310_45028# 5.87e-20
C43876 a_n743_46660# a_380_45546# 0.010247f
C43877 a_n1021_46688# a_n1099_45572# 2.81e-21
C43878 a_7411_46660# a_8049_45260# 5.59e-20
C43879 a_1123_46634# a_n2661_45546# 4.02e-20
C43880 a_n133_46660# a_n863_45724# 1.41e-19
C43881 a_n2438_43548# a_n452_45724# 3.99e-20
C43882 a_15227_44166# a_17583_46090# 4.28e-21
C43883 a_765_45546# a_5068_46348# 3.71e-21
C43884 a_12991_46634# a_6945_45028# 1.08e-19
C43885 a_12469_46902# a_10809_44734# 0.014309f
C43886 a_17609_46634# a_18189_46348# 1.41e-19
C43887 a_15682_43940# a_16547_43609# 0.008948f
C43888 a_7499_43940# a_7112_43396# 0.001375f
C43889 a_15493_43396# a_15681_43442# 0.029338f
C43890 a_11967_42832# a_13635_43156# 0.053949f
C43891 a_14539_43914# a_18695_43230# 1.08e-19
C43892 a_13565_44260# a_9145_43396# 2.31e-20
C43893 a_15301_44260# a_8685_43396# 1.7e-20
C43894 a_11341_43940# a_12293_43646# 8.32e-19
C43895 a_n2810_45028# a_n4209_39304# 0.021684f
C43896 a_n97_42460# VDD 3.61113f
C43897 a_20841_45814# a_20719_45572# 3.16e-19
C43898 a_16147_45260# a_n1059_45260# 5.91e-21
C43899 a_20107_45572# a_21513_45002# 8.78e-20
C43900 a_7227_45028# a_7418_45067# 4e-19
C43901 a_10907_45822# a_9482_43914# 3.21e-20
C43902 a_6472_45840# a_n2661_43370# 5.95e-20
C43903 a_10341_42308# a_3090_45724# 0.002812f
C43904 a_4235_43370# a_n1925_42282# 0.199349f
C43905 a_4699_43561# a_526_44458# 1.19e-19
C43906 a_9145_43396# a_9290_44172# 0.103991f
C43907 a_9885_43646# a_8016_46348# 0.001881f
C43908 a_5932_42308# a_n2312_40392# 6.05e-21
C43909 a_14113_42308# a_12861_44030# 1.46e-20
C43910 a_2711_45572# a_4883_46098# 0.041245f
C43911 a_14495_45572# a_4915_47217# 0.001776f
C43912 a_13527_45546# a_6151_47436# 4.69e-21
C43913 a_10193_42453# a_11459_47204# 3.13e-19
C43914 a_8746_45002# a_9313_45822# 5.46e-20
C43915 a_6229_45572# a_4791_45118# 1.28e-19
C43916 a_18819_46122# a_20009_46494# 2.56e-19
C43917 a_5066_45546# a_6347_46155# 7.61e-19
C43918 a_7542_44172# a_6123_31319# 8.34e-21
C43919 a_n2661_42282# a_2713_42308# 1.2e-19
C43920 a_2982_43646# a_16795_42852# 1.51e-20
C43921 a_3626_43646# a_15567_42826# 2.41e-20
C43922 a_19700_43370# a_4190_30871# 0.046581f
C43923 a_15743_43084# a_743_42282# 0.029529f
C43924 a_17499_43370# a_4361_42308# 6.03e-20
C43925 a_104_43370# a_133_42852# 8.41e-20
C43926 en_comp a_22469_40625# 0.021539f
C43927 a_16751_45260# a_17719_45144# 3.82e-19
C43928 a_11787_45002# a_11691_44458# 1.53e-19
C43929 a_13348_45260# a_11827_44484# 3.7e-22
C43930 a_5263_45724# a_5244_44056# 5.95e-21
C43931 a_45_45144# a_n2661_43370# 4.17e-19
C43932 a_8696_44636# a_15146_44811# 1.39e-19
C43933 a_5147_45002# a_n2661_44458# 0.024256f
C43934 a_327_44734# a_949_44458# 0.003334f
C43935 a_413_45260# a_2779_44458# 0.024142f
C43936 a_1667_45002# a_742_44458# 0.002122f
C43937 a_13635_43156# a_13259_45724# 0.017822f
C43938 a_2905_42968# a_n863_45724# 0.269475f
C43939 a_133_43172# a_n755_45592# 0.002433f
C43940 a_n1991_42858# a_n443_42852# 1.6e-19
C43941 a_421_43172# a_n357_42282# 2.38e-19
C43942 a_6101_43172# a_526_44458# 6.27e-21
C43943 a_n3565_37414# SMPL_ON_P 0.016441f
C43944 a_16855_45546# a_6755_46942# 3.44e-19
C43945 a_13249_42308# a_15227_44166# 2.89e-20
C43946 a_413_45260# a_20916_46384# 6.71e-20
C43947 a_n2109_45247# a_n2438_43548# 0.007532f
C43948 a_n1059_45260# a_n1021_46688# 3.15e-21
C43949 a_n913_45002# a_n1925_46634# 1.36e-21
C43950 a_5205_44484# a_768_44030# 0.033081f
C43951 a_3537_45260# a_5807_45002# 0.005102f
C43952 en_comp a_n2442_46660# 0.02478f
C43953 a_n2956_37592# a_n2293_46634# 4.76e-19
C43954 a_8953_45002# a_9804_47204# 0.003283f
C43955 a_n2129_44697# a_n2497_47436# 0.019202f
C43956 a_22780_40081# VDD 2.4e-19
C43957 a_3626_43646# a_20712_42282# 3.92e-19
C43958 a_n1423_42826# a_n4318_38216# 3.57e-19
C43959 a_9145_43396# a_15051_42282# 0.001238f
C43960 a_2982_43646# a_21335_42336# 0.009024f
C43961 a_n2472_42826# a_n4318_37592# 2.65e-20
C43962 a_n2157_42858# a_n1736_42282# 0.001064f
C43963 a_12379_42858# a_12800_43218# 0.089677f
C43964 a_n1991_42858# a_n2104_42282# 2.18e-19
C43965 a_743_42282# a_1606_42308# 0.088097f
C43966 a_14358_43442# a_14456_42282# 1.03e-20
C43967 a_10341_43396# a_11551_42558# 3.11e-22
C43968 a_10991_42826# a_11136_42852# 0.057222f
C43969 a_10765_43646# a_5742_30871# 3.49e-20
C43970 a_n4318_39304# a_n3565_39304# 3.96e-19
C43971 a_15682_46116# CLK 2.6e-19
C43972 a_20708_46348# RST_Z 5.4e-22
C43973 a_19900_46494# START 3.05e-20
C43974 a_n3420_39616# VDD 0.568506f
C43975 a_n971_45724# a_768_44030# 0.069358f
C43976 a_2063_45854# a_n881_46662# 0.612456f
C43977 a_2553_47502# a_n1613_43370# 3.57e-20
C43978 a_2905_45572# a_3094_47243# 0.006879f
C43979 a_2952_47436# a_3411_47243# 6.64e-19
C43980 a_16327_47482# a_16588_47582# 0.276601f
C43981 a_13717_47436# a_20990_47178# 9.85e-20
C43982 a_9313_45822# a_4883_46098# 0.026043f
C43983 a_13381_47204# a_13507_46334# 0.001369f
C43984 a_15673_47210# a_10227_46804# 0.02634f
C43985 a_11599_46634# a_18780_47178# 3.49e-19
C43986 a_n443_46116# a_2747_46873# 0.047485f
C43987 a_8953_45002# a_10405_44172# 1.1e-20
C43988 a_6171_45002# a_15682_43940# 5.04e-19
C43989 a_11691_44458# a_17325_44484# 0.0017f
C43990 a_2711_45572# a_16243_43396# 2.11e-19
C43991 a_7499_43078# a_9803_43646# 0.001386f
C43992 a_18315_45260# a_18579_44172# 1.04e-20
C43993 a_n2293_42834# a_644_44056# 1.25e-20
C43994 a_n2661_43370# a_n2472_43914# 0.00608f
C43995 a_11827_44484# a_19615_44636# 0.006593f
C43996 a_8975_43940# a_9313_44734# 0.391938f
C43997 a_6298_44484# a_9159_44484# 6.91e-21
C43998 a_5343_44458# a_n2661_42834# 0.038788f
C43999 a_4743_44484# a_n2661_43922# 0.008142f
C44000 a_21005_45260# a_20640_44752# 4.55e-20
C44001 a_20567_45036# a_20679_44626# 0.006083f
C44002 a_19778_44110# a_19279_43940# 0.020911f
C44003 a_n3565_38502# a_n2956_39304# 0.001812f
C44004 a_16020_45572# VDD 0.077625f
C44005 a_5534_30871# C7_P_btm 0.060228f
C44006 a_5342_30871# C9_P_btm 5.28e-19
C44007 a_16019_45002# a_11415_45002# 0.007819f
C44008 a_14797_45144# a_12741_44636# 1.29e-20
C44009 a_3537_45260# a_3699_46348# 3.5e-21
C44010 a_16922_45042# a_19466_46812# 0.030378f
C44011 a_4574_45260# a_3483_46348# 0.022358f
C44012 a_17613_45144# a_15227_44166# 0.048772f
C44013 a_6298_44484# a_7715_46873# 3.13e-20
C44014 a_17517_44484# a_12549_44172# 0.019389f
C44015 a_18494_42460# a_3090_45724# 1.58e-20
C44016 a_n2661_42834# a_n2956_39768# 7.06e-20
C44017 a_3429_45260# a_4185_45028# 0.004974f
C44018 a_11691_44458# a_11813_46116# 1.05e-21
C44019 a_16855_45546# a_8049_45260# 0.004398f
C44020 a_20528_45572# a_20075_46420# 5.63e-19
C44021 a_2437_43646# a_17583_46090# 9.89e-22
C44022 a_3357_43084# a_14840_46494# 2.67e-21
C44023 a_413_45260# a_6165_46155# 9.78e-21
C44024 a_n1059_45260# a_9290_44172# 0.092471f
C44025 a_20841_45814# a_6945_45028# 4.67e-19
C44026 a_17730_32519# a_13507_46334# 1.98e-20
C44027 a_n1630_35242# a_6123_31319# 0.036823f
C44028 a_16245_42852# a_15890_42674# 0.001613f
C44029 a_1606_42308# a_5755_42308# 3.31e-20
C44030 a_4190_30871# C3_N_btm 1.1e-19
C44031 a_22521_39511# a_22821_38993# 0.112629f
C44032 a_22521_40055# a_22876_39857# 4.84e-19
C44033 a_22780_40081# a_22469_39537# 1.28e-20
C44034 a_n2661_46634# a_7577_46660# 0.047111f
C44035 a_5807_45002# a_6969_46634# 0.003601f
C44036 a_2107_46812# a_4955_46873# 0.031068f
C44037 a_2443_46660# a_3067_47026# 9.73e-19
C44038 a_2609_46660# a_2864_46660# 0.055869f
C44039 a_13661_43548# a_6755_46942# 0.088986f
C44040 a_n2293_46634# a_5257_43370# 0.061974f
C44041 a_3177_46902# a_3524_46660# 0.051162f
C44042 a_n2661_46098# a_1057_46660# 1.99e-19
C44043 a_11599_46634# a_18285_46348# 0.030958f
C44044 a_10227_46804# a_16388_46812# 8.39e-20
C44045 a_15811_47375# a_765_45546# 0.035109f
C44046 a_13717_47436# a_20273_46660# 2.45e-21
C44047 a_n2497_47436# a_3483_46348# 4.12e-20
C44048 a_n1741_47186# a_2521_46116# 1.08e-20
C44049 a_n971_45724# a_1176_45822# 1.67e-19
C44050 a_2553_47502# a_n2293_46098# 4.34e-23
C44051 a_584_46384# a_n1853_46287# 4.85e-21
C44052 a_n237_47217# a_805_46414# 1.4e-19
C44053 a_n746_45260# a_1208_46090# 3.58e-20
C44054 a_n785_47204# a_376_46348# 1.57e-19
C44055 a_n699_43396# a_n97_42460# 0.152094f
C44056 a_644_44056# a_1115_44172# 0.013441f
C44057 a_14673_44172# a_15682_43940# 0.001963f
C44058 a_n2661_43370# a_10695_43548# 6.82e-21
C44059 a_13249_42308# a_14635_42282# 1.46e-19
C44060 a_n2661_44458# a_4093_43548# 3.38e-20
C44061 a_18479_45785# a_19339_43156# 0.001029f
C44062 a_n2661_42834# a_9801_44260# 2.25e-19
C44063 a_n1059_45260# a_791_42968# 0.122941f
C44064 a_n913_45002# a_685_42968# 0.015577f
C44065 a_n2017_45002# a_1847_42826# 0.017915f
C44066 a_n967_45348# a_n967_43230# 3.59e-19
C44067 a_5088_37509# VDD 1.15925f
C44068 a_742_44458# VDD 1.3845f
C44069 a_19332_42282# RST_Z 4.07e-20
C44070 a_n4315_30879# a_n1838_35608# 2.23e-19
C44071 a_n2946_37984# a_n2810_45572# 0.020842f
C44072 a_n2267_43396# a_n2293_46634# 7.31e-22
C44073 a_n2661_43370# a_n357_42282# 0.034578f
C44074 a_5343_44458# a_5066_45546# 1.18e-21
C44075 a_n2661_43922# a_8016_46348# 0.02895f
C44076 a_9159_44484# a_5937_45572# 0.040512f
C44077 a_5289_44734# a_2324_44458# 0.001168f
C44078 a_8685_43396# a_12465_44636# 5.48e-20
C44079 a_15781_43660# a_12861_44030# 0.025765f
C44080 a_14955_43396# a_10227_46804# 0.035123f
C44081 a_n4209_39590# a_n4251_39616# 0.00226f
C44082 a_n2946_39866# a_n2302_39866# 6.68e-19
C44083 a_n4064_40160# a_n4334_39392# 0.013157f
C44084 a_n3420_39616# a_n2860_39866# 0.002301f
C44085 a_20843_47204# VDD 0.188032f
C44086 a_5932_42308# C0_dummy_N_btm 1.2e-19
C44087 a_14976_45028# a_12741_44636# 3.06e-19
C44088 a_13059_46348# a_765_45546# 4.68e-19
C44089 a_16388_46812# a_17339_46660# 0.24887f
C44090 a_19692_46634# a_19636_46660# 3.77e-19
C44091 a_7577_46660# a_8199_44636# 1.99e-19
C44092 a_7715_46873# a_5937_45572# 1.65e-20
C44093 a_7927_46660# a_8016_46348# 8.96e-19
C44094 a_8145_46902# a_8349_46414# 7.84e-19
C44095 a_n881_46662# a_14383_46116# 1.43e-19
C44096 a_13661_43548# a_8049_45260# 0.032643f
C44097 a_n743_46660# a_526_44458# 0.020498f
C44098 a_12891_46348# a_12638_46436# 0.13727f
C44099 a_12549_44172# a_12379_46436# 3.71e-19
C44100 en_comp a_14456_42282# 8.68e-21
C44101 a_n2017_45002# a_15486_42560# 0.005473f
C44102 a_n1059_45260# a_15051_42282# 6.54e-19
C44103 a_n913_45002# a_14113_42308# 0.029759f
C44104 a_n2661_42834# a_n1545_43230# 3.82e-19
C44105 a_19789_44512# a_15743_43084# 2.77e-21
C44106 a_742_44458# a_873_42968# 7.93e-21
C44107 a_n2293_43922# a_n4318_38680# 2.08e-19
C44108 a_14539_43914# a_16795_42852# 0.037061f
C44109 a_n356_44636# a_10341_42308# 1.92e-20
C44110 a_5891_43370# a_7227_42852# 0.129383f
C44111 a_17517_44484# a_21855_43396# 3.12e-22
C44112 a_n2661_42282# a_6031_43396# 0.036698f
C44113 a_21115_43940# VDD 0.145936f
C44114 a_15599_45572# a_16147_45260# 7.22e-19
C44115 a_16333_45814# a_16211_45572# 3.16e-19
C44116 a_5263_45724# a_5111_44636# 0.00615f
C44117 a_3775_45552# a_2382_45260# 2.04e-19
C44118 a_2711_45572# a_3232_43370# 0.002535f
C44119 a_7499_43078# a_n913_45002# 0.548687f
C44120 a_n1557_42282# a_1138_42852# 0.009215f
C44121 a_n2293_42282# a_n2956_39768# 5.23e-20
C44122 a_8037_42858# a_4646_46812# 0.001539f
C44123 a_18783_43370# a_19692_46634# 1.14e-20
C44124 a_n4318_39768# a_n2810_45572# 0.023737f
C44125 a_2998_44172# a_n357_42282# 4.93e-20
C44126 a_n4064_37984# VCM 0.011087f
C44127 a_n4209_37414# EN_VIN_BSTR_P 0.007584f
C44128 a_n3565_37414# a_n1532_35090# 7.27e-20
C44129 a_7754_38470# a_11530_34132# 7.75e-19
C44130 a_5204_45822# VDD 0.359177f
C44131 a_5907_45546# a_n2109_47186# 8.91e-19
C44132 a_n4209_39304# a_n2302_37690# 3.3e-19
C44133 a_n3565_39304# a_n2946_37690# 2.71e-19
C44134 a_n4064_39072# a_n4334_37440# 3.19e-19
C44135 a_4185_45028# a_8049_45260# 0.014062f
C44136 a_8349_46414# a_5066_45546# 0.005369f
C44137 a_18819_46122# a_21137_46414# 2.71e-21
C44138 a_17715_44484# a_10809_44734# 1.44e-19
C44139 a_19553_46090# a_19900_46494# 0.051162f
C44140 a_18985_46122# a_20708_46348# 2.48e-19
C44141 a_n2065_43946# a_n4318_37592# 2.96e-22
C44142 a_n1761_44111# a_n1736_42282# 3.18e-19
C44143 a_8333_44056# a_8495_42852# 5.85e-22
C44144 a_n2267_43396# a_n1533_42852# 4.05e-20
C44145 a_3539_42460# a_743_42282# 0.054149f
C44146 a_n2293_43922# a_11551_42558# 1.93e-19
C44147 a_9313_44734# a_15803_42450# 8.69e-20
C44148 a_n356_44636# a_18057_42282# 0.087032f
C44149 a_14579_43548# a_14537_43646# 0.001675f
C44150 a_8685_43396# a_16409_43396# 6.54e-20
C44151 a_9145_43396# a_13749_43396# 3.66e-19
C44152 a_3094_47570# DATA[1] 2.62e-21
C44153 a_21588_30879# a_22521_39511# 7.63e-20
C44154 a_n901_43156# VDD 0.475947f
C44155 a_5147_45002# a_6125_45348# 1.1e-19
C44156 a_5111_44636# a_5837_45348# 0.001223f
C44157 a_3065_45002# a_2809_45028# 0.006555f
C44158 a_4927_45028# a_5365_45348# 0.013015f
C44159 a_8191_45002# a_1423_45028# 1.9e-20
C44160 a_n745_45366# a_n2661_43370# 0.005292f
C44161 a_18787_45572# a_11691_44458# 1.34e-19
C44162 a_13777_45326# a_14537_43396# 4.1e-19
C44163 a_9482_43914# a_15415_45028# 0.002812f
C44164 a_13556_45296# a_14797_45144# 2.59e-20
C44165 a_10193_42453# a_9313_44734# 0.078654f
C44166 a_n4064_40160# a_n2312_38680# 8.3e-19
C44167 a_n3565_39590# a_n2956_39768# 0.302561f
C44168 a_n2216_40160# a_n2442_46660# 0.001258f
C44169 a_14205_43396# a_n443_42852# 0.118229f
C44170 a_15681_43442# a_n357_42282# 3.86e-20
C44171 a_1847_42826# a_526_44458# 0.154735f
C44172 a_6511_45714# a_6969_46634# 7.16e-20
C44173 a_6667_45809# a_6755_46942# 1.38e-20
C44174 a_7230_45938# a_5257_43370# 6.16e-21
C44175 a_8696_44636# a_n2661_46634# 2.14e-19
C44176 a_16842_45938# a_5807_45002# 1.8e-19
C44177 a_2437_43646# a_2266_47570# 0.001239f
C44178 a_20447_31679# SMPL_ON_N 0.029368f
C44179 a_413_45260# a_16023_47582# 1.6e-19
C44180 a_3232_43370# a_9313_45822# 1.83e-20
C44181 a_1307_43914# a_2063_45854# 0.005774f
C44182 a_3495_45348# a_n971_45724# 0.005013f
C44183 a_6125_45348# a_n2109_47186# 3.53e-19
C44184 a_n1099_45572# a_n89_45572# 9.15e-19
C44185 a_n755_45592# a_1990_45899# 9.01e-21
C44186 a_380_45546# a_509_45572# 0.010132f
C44187 a_n356_45724# a_7_45899# 0.005265f
C44188 a_1848_45724# a_1609_45822# 0.042695f
C44189 a_16137_43396# a_17665_42852# 0.001078f
C44190 a_3080_42308# a_3905_42308# 8.29e-20
C44191 a_10922_42852# a_12089_42308# 8.07e-21
C44192 a_n97_42460# a_11551_42558# 0.095523f
C44193 a_3626_43646# a_6171_42473# 0.003703f
C44194 a_10341_42308# a_12379_42858# 2.14e-19
C44195 a_n1076_43230# a_133_42852# 1.24e-19
C44196 a_18429_43548# a_18504_43218# 1.16e-19
C44197 a_21076_30879# SINGLE_ENDED 1.21e-19
C44198 a_4338_37500# VDAC_P 0.037246f
C44199 a_3726_37500# a_11206_38545# 0.11542f
C44200 a_5700_37509# VDAC_N 1.09421f
C44201 a_5088_37509# a_8912_37509# 16.1906f
C44202 a_3422_30871# C0_dummy_P_btm 1.28e-20
C44203 a_10533_42308# VDD 0.216201f
C44204 a_3160_47472# a_3815_47204# 1.5e-19
C44205 a_n1151_42308# a_3785_47178# 0.029415f
C44206 a_2905_45572# a_4007_47204# 0.001036f
C44207 a_2063_45854# a_n443_46116# 0.177177f
C44208 a_n1741_47186# a_13381_47204# 4.11e-19
C44209 a_n1920_47178# a_n1435_47204# 0.001089f
C44210 a_n237_47217# a_7903_47542# 0.086772f
C44211 a_16019_45002# a_11967_42832# 8.44e-20
C44212 a_11691_44458# a_18287_44626# 0.032949f
C44213 a_n2661_44458# a_10157_44484# 0.00786f
C44214 a_742_44458# a_n699_43396# 0.047576f
C44215 a_18479_45785# a_17973_43940# 2.56e-22
C44216 a_18494_42460# a_n356_44636# 0.003788f
C44217 a_327_44734# a_175_44278# 0.001132f
C44218 a_n1059_45260# a_3905_42865# 0.01898f
C44219 a_n2017_45002# a_5244_44056# 3.28e-21
C44220 a_n784_42308# a_n863_45724# 0.358682f
C44221 COMP_P a_n357_42282# 3.45e-20
C44222 a_3733_45822# VDD 5.25e-19
C44223 a_4190_30871# C7_P_btm 2.94e-19
C44224 a_13678_32519# a_11530_34132# 0.002459f
C44225 a_n2267_44484# a_n2293_46634# 2.41e-19
C44226 a_13556_45296# a_14976_45028# 0.003018f
C44227 a_13076_44458# a_768_44030# 0.132449f
C44228 a_13720_44458# a_12549_44172# 7.87e-20
C44229 a_9482_43914# a_15368_46634# 3.52e-20
C44230 a_20719_45572# a_11415_45002# 7.75e-19
C44231 a_4880_45572# a_5066_45546# 0.04794f
C44232 a_6667_45809# a_8049_45260# 2.79e-19
C44233 a_14033_45822# a_10903_43370# 0.040019f
C44234 a_8696_44636# a_8199_44636# 0.265919f
C44235 a_n2661_42834# a_10227_46804# 0.024624f
C44236 a_n4318_38680# a_n3420_39616# 0.02534f
C44237 a_5342_30871# a_16104_42674# 4.45e-20
C44238 a_n1151_42308# a_3090_45724# 0.003613f
C44239 a_5807_45002# a_n2293_46634# 9.62e-19
C44240 a_4915_47217# a_11901_46660# 0.004227f
C44241 a_6575_47204# a_8189_46660# 1.95e-20
C44242 a_11599_46634# a_10249_46116# 7.84e-19
C44243 a_14955_47212# a_6755_46942# 4.64e-19
C44244 a_4883_46098# a_6540_46812# 2.72e-20
C44245 a_n1613_43370# a_1799_45572# 0.008733f
C44246 a_n913_45002# a_15781_43660# 8.25e-21
C44247 a_11967_42832# a_18245_44484# 1.94e-19
C44248 a_20362_44736# a_20766_44850# 0.051162f
C44249 a_n356_44636# a_3499_42826# 1.72e-20
C44250 a_n2293_42834# a_104_43370# 0.003003f
C44251 a_n2661_43370# a_n2433_43396# 0.021188f
C44252 a_10193_42453# a_18599_43230# 0.003065f
C44253 a_n2661_42834# a_453_43940# 0.04708f
C44254 a_n2661_43922# a_1414_42308# 0.010195f
C44255 a_20640_44752# a_20835_44721# 0.20669f
C44256 a_20159_44458# a_19279_43940# 0.06519f
C44257 a_20692_30879# C0_N_btm 9.35e-21
C44258 a_6123_31319# a_11530_34132# 0.001062f
C44259 a_5934_30871# EN_VIN_BSTR_P 0.075302f
C44260 a_1606_42308# VIN_P 0.014401f
C44261 a_22469_40625# a_4185_45028# 1.54e-20
C44262 a_5883_43914# a_3483_46348# 5.92e-19
C44263 a_17325_44484# a_15227_44166# 0.001944f
C44264 a_10949_43914# a_2107_46812# 8.95e-21
C44265 a_16019_45002# a_13259_45724# 1.86e-19
C44266 a_2382_45260# a_3218_45724# 5.5e-20
C44267 a_2680_45002# a_2957_45546# 4.36e-19
C44268 a_3537_45260# a_n755_45592# 0.025346f
C44269 a_n967_45348# a_n443_42852# 3.13e-19
C44270 a_2274_45254# a_3316_45546# 8.04e-21
C44271 a_19778_44110# a_20708_46348# 4.6e-21
C44272 a_11691_44458# a_15682_46116# 1.87e-21
C44273 a_18184_42460# a_19900_46494# 4.45e-21
C44274 a_18494_42460# a_20075_46420# 2.66e-19
C44275 a_5343_44458# a_5068_46348# 1.11e-21
C44276 a_17538_32519# a_13507_46334# 8.21e-20
C44277 a_16241_47178# VDD 0.208959f
C44278 a_18057_42282# a_18727_42674# 0.003581f
C44279 a_17303_42282# a_19332_42282# 3.68e-19
C44280 a_n743_46660# a_2521_46116# 0.013075f
C44281 a_n1925_46634# a_2804_46116# 3.92e-20
C44282 a_948_46660# a_472_46348# 7.34e-19
C44283 a_n2661_46098# a_n2472_46090# 0.094589f
C44284 a_n2438_43548# a_167_45260# 0.050543f
C44285 a_1799_45572# a_n2293_46098# 0.014011f
C44286 a_2107_46812# a_376_46348# 7.16e-20
C44287 a_7577_46660# a_765_45546# 0.002481f
C44288 a_6755_46942# a_14543_46987# 4.62e-19
C44289 a_12891_46348# a_13759_46122# 2.87e-20
C44290 a_5807_45002# a_9625_46129# 0.001468f
C44291 a_n2661_46634# a_4704_46090# 1.84e-20
C44292 a_12549_44172# a_13351_46090# 0.014836f
C44293 a_768_44030# a_12594_46348# 0.001137f
C44294 a_n881_46662# a_17715_44484# 0.014166f
C44295 a_14955_47212# a_8049_45260# 1.17e-21
C44296 a_n746_45260# a_n2661_45546# 0.022378f
C44297 a_n2497_47436# a_n357_42282# 0.046314f
C44298 a_n971_45724# a_n2472_45546# 7.36e-20
C44299 a_n2109_47186# a_n1099_45572# 1.08e-20
C44300 a_15433_44458# a_15095_43370# 1.02e-20
C44301 a_18287_44626# a_4190_30871# 4.63e-21
C44302 a_1467_44172# a_n97_42460# 0.190191f
C44303 a_17973_43940# a_14021_43940# 4.61e-20
C44304 a_11341_43940# a_15493_43940# 0.216602f
C44305 a_3422_30871# a_2982_43646# 0.140944f
C44306 a_n699_43396# a_n901_43156# 6.3e-20
C44307 a_n2661_44458# a_685_42968# 1.08e-21
C44308 a_11827_44484# a_10835_43094# 8.97e-20
C44309 a_9313_44734# a_16137_43396# 0.044229f
C44310 a_11823_42460# a_7174_31319# 9.76e-21
C44311 a_14955_43940# a_15037_44260# 0.003935f
C44312 a_n2661_42282# a_6671_43940# 0.002068f
C44313 a_n2661_43922# a_12281_43396# 2.21e-20
C44314 a_n2293_42834# a_4156_43218# 6.26e-20
C44315 a_n2017_45002# a_n473_42460# 0.017082f
C44316 a_n2956_37592# a_n1736_42282# 8.96e-21
C44317 en_comp a_n3674_38216# 0.026738f
C44318 a_n2810_45028# a_n4318_37592# 0.023097f
C44319 a_n1059_45260# a_n961_42308# 3.29e-21
C44320 a_n967_45348# a_n2104_42282# 4.03e-19
C44321 a_n984_44318# VDD 0.281427f
C44322 a_10490_45724# a_12016_45572# 0.003469f
C44323 a_11525_45546# a_11688_45572# 0.011381f
C44324 C0_P_btm VCM 0.717283f
C44325 C0_N_btm VIN_N 0.529671f
C44326 a_5745_43940# a_n2293_46098# 0.019006f
C44327 a_6197_43396# a_3090_45724# 0.010809f
C44328 a_n2157_42858# a_n2442_46660# 5.35e-21
C44329 a_n1423_42826# a_n2956_39768# 3.32e-21
C44330 a_5244_44056# a_526_44458# 4.69e-21
C44331 a_3905_42865# a_n1925_42282# 0.023709f
C44332 a_18245_44484# a_13259_45724# 1.46e-19
C44333 a_9028_43914# a_2324_44458# 4.61e-20
C44334 a_19339_43156# a_13507_46334# 4.77e-21
C44335 a_10951_45334# CLK 0.005907f
C44336 a_16721_46634# VDD 0.186443f
C44337 a_4419_46090# a_5937_45572# 8.29e-20
C44338 a_22365_46825# a_10809_44734# 0.010841f
C44339 a_12741_44636# a_19900_46494# 0.005543f
C44340 a_3483_46348# a_9569_46155# 1.05e-19
C44341 a_11415_45002# a_6945_45028# 0.002828f
C44342 a_20202_43084# a_22223_46124# 1.62e-19
C44343 a_3090_45724# a_19240_46482# 2.23e-19
C44344 a_14976_45028# a_16375_45002# 1.01e-20
C44345 a_n2661_42834# a_n2472_42282# 2.95e-19
C44346 a_16922_45042# a_13258_32519# 4.48e-20
C44347 a_6293_42852# a_7287_43370# 1.04e-20
C44348 a_11967_42832# a_13814_43218# 0.001842f
C44349 a_3626_43646# a_3457_43396# 0.067226f
C44350 a_18494_42460# a_18727_42674# 0.031761f
C44351 a_18184_42460# a_18907_42674# 0.071964f
C44352 a_n356_44636# a_3318_42354# 1.4e-19
C44353 a_14021_43940# a_22591_43396# 0.057848f
C44354 a_6197_43396# a_6547_43396# 0.216095f
C44355 a_6031_43396# a_7112_43396# 0.101963f
C44356 a_2952_47436# DATA[2] 2.12e-19
C44357 a_2905_45572# DATA[1] 1.91e-21
C44358 a_n1151_42308# CLK_DATA 1.24e-21
C44359 a_2063_45854# DATA[4] 3.07e-19
C44360 a_19479_31679# C1_N_btm 0.043983f
C44361 a_9885_43646# VDD 0.190473f
C44362 a_13904_45546# a_11691_44458# 4.03e-21
C44363 a_6598_45938# a_6298_44484# 0.001025f
C44364 a_7499_43078# a_n2661_44458# 0.059442f
C44365 a_2711_45572# a_8975_43940# 6.21e-21
C44366 a_6472_45840# a_5883_43914# 3.93e-22
C44367 a_n37_45144# a_413_45260# 0.021944f
C44368 a_n1059_45260# a_5147_45002# 2.48e-21
C44369 a_n2017_45002# a_5111_44636# 0.024598f
C44370 a_3681_42891# a_1823_45246# 2.81e-20
C44371 a_12089_42308# a_12741_44636# 6.17e-22
C44372 a_9223_42460# a_n2293_46634# 1.9e-20
C44373 a_1568_43370# a_n357_42282# 0.036942f
C44374 a_3080_42308# a_n863_45724# 0.001926f
C44375 a_n1557_42282# a_n2956_38216# 1.25e-20
C44376 a_1049_43396# a_n755_45592# 8.22e-21
C44377 a_22465_38105# a_13507_46334# 9.82e-20
C44378 a_3503_45724# VDD 0.129733f
C44379 a_11322_45546# a_768_44030# 6.14e-20
C44380 a_5907_45546# a_n1925_46634# 6.84e-21
C44381 a_4099_45572# a_n743_46660# 1.05e-19
C44382 a_11525_45546# a_12549_44172# 7.96e-19
C44383 a_7227_45028# a_n2661_46634# 3.38e-20
C44384 a_14495_45572# a_n881_46662# 0.170589f
C44385 a_n2293_45010# SMPL_ON_P 4.92e-20
C44386 a_2437_43646# a_2124_47436# 0.025048f
C44387 a_17478_45572# a_17591_47464# 1.31e-20
C44388 a_15861_45028# a_10227_46804# 0.002162f
C44389 a_16375_45002# a_18051_46116# 0.038793f
C44390 a_14976_45028# RST_Z 2.6e-20
C44391 a_15682_43940# a_15959_42545# 2.38e-19
C44392 a_n2433_43396# COMP_P 0.001151f
C44393 a_16409_43396# a_17333_42852# 1.86e-19
C44394 a_17499_43370# a_17595_43084# 0.002317f
C44395 a_4361_42308# a_5755_42852# 2.34e-20
C44396 a_743_42282# a_8605_42826# 5.66e-20
C44397 a_17324_43396# a_16795_42852# 1.3e-19
C44398 a_n2267_43396# a_n1736_42282# 3.76e-21
C44399 a_16137_43396# a_18599_43230# 0.005055f
C44400 a_n1641_43230# a_n1736_43218# 0.049827f
C44401 a_n1423_42826# a_n1545_43230# 3.16e-19
C44402 a_n1853_43023# a_n967_43230# 8.59e-19
C44403 a_n901_43156# a_n4318_38680# 7.68e-22
C44404 a_15743_43084# a_15279_43071# 1.83e-19
C44405 a_11341_43940# a_5742_30871# 0.0019f
C44406 a_11735_46660# CLK 6.72e-20
C44407 VDAC_Pi a_3754_39466# 0.308867f
C44408 a_20256_42852# VDD 0.001626f
C44409 a_7705_45326# a_7640_43914# 5.79e-20
C44410 a_3232_43370# a_9241_44734# 8.2e-19
C44411 a_20731_45938# a_20640_44752# 2.23e-21
C44412 a_7229_43940# a_5891_43370# 1.39e-19
C44413 a_2274_45254# a_n2661_42834# 1.64e-20
C44414 a_20623_45572# a_19279_43940# 7.39e-21
C44415 a_16501_45348# a_16237_45028# 3.62e-19
C44416 a_11823_42460# a_10729_43914# 8.14e-20
C44417 a_16922_45042# a_20193_45348# 0.328274f
C44418 a_10193_42453# a_17737_43940# 0.02461f
C44419 a_11652_45724# a_11750_44172# 6.11e-20
C44420 a_n2293_42834# a_949_44458# 4.61e-20
C44421 a_5093_45028# a_5343_44458# 4.13e-19
C44422 a_n2661_43370# a_n2433_44484# 0.018595f
C44423 a_18494_42460# a_20567_45036# 5.4e-19
C44424 a_19778_44110# a_21101_45002# 0.008451f
C44425 a_18587_45118# a_11827_44484# 5.85e-20
C44426 a_17023_45118# a_11691_44458# 0.00304f
C44427 a_12427_45724# a_10949_43914# 3.38e-21
C44428 a_14456_42282# a_4185_45028# 1.64e-19
C44429 a_n961_42308# a_n1925_42282# 2.27e-19
C44430 a_13814_43218# a_13259_45724# 5.53e-19
C44431 a_9803_42558# a_8953_45546# 0.031932f
C44432 a_9377_42558# a_8199_44636# 0.001018f
C44433 a_8162_45546# a_3483_46348# 0.009853f
C44434 a_8696_44636# a_765_45546# 0.001141f
C44435 a_15861_45028# a_17339_46660# 5.36e-22
C44436 a_13490_45067# a_12891_46348# 0.00125f
C44437 a_2232_45348# a_2107_46812# 1.12e-19
C44438 a_6171_45002# a_5732_46660# 1.44e-19
C44439 a_8191_45002# a_4646_46812# 7.69e-21
C44440 a_2437_43646# a_11813_46116# 7.51e-20
C44441 a_7227_45028# a_8199_44636# 3.82e-20
C44442 a_6598_45938# a_5937_45572# 2.01e-19
C44443 a_2711_45572# a_11387_46155# 4.02e-20
C44444 a_5024_45822# a_5204_45822# 1.6e-19
C44445 a_19721_31679# a_13507_46334# 8.21e-20
C44446 a_8975_43940# a_9313_45822# 3.56e-20
C44447 a_n356_44636# a_n1151_42308# 0.093166f
C44448 a_700_44734# a_584_46384# 5.41e-19
C44449 a_4361_42308# a_10149_42308# 6.19e-19
C44450 a_743_42282# a_16104_42674# 0.002282f
C44451 a_4190_30871# a_17124_42282# 7.43e-20
C44452 a_5649_42852# a_15890_42674# 5.19e-20
C44453 a_n2293_42282# a_n2472_42282# 0.163758f
C44454 a_15743_43084# a_13258_32519# 1.74e-19
C44455 a_16823_43084# a_4958_30871# 5.65e-19
C44456 a_19700_43370# a_19511_42282# 6.2e-21
C44457 a_2747_46873# a_n1613_43370# 0.03071f
C44458 a_12465_44636# a_768_44030# 0.120859f
C44459 a_10227_46804# a_19321_45002# 0.111029f
C44460 a_18597_46090# a_5807_45002# 0.005073f
C44461 a_18780_47178# a_13661_43548# 0.153988f
C44462 a_18479_47436# a_13747_46662# 0.083389f
C44463 a_13381_47204# a_n743_46660# 1.37e-20
C44464 a_n237_47217# a_4817_46660# 6.61e-20
C44465 a_n971_45724# a_5167_46660# 3.91e-20
C44466 a_n1151_42308# a_3699_46634# 1.12e-19
C44467 a_3381_47502# a_2959_46660# 0.005389f
C44468 a_3160_47472# a_3524_46660# 1.52e-20
C44469 a_584_46384# a_2162_46660# 0.001394f
C44470 a_949_44458# a_1115_44172# 0.016355f
C44471 a_18374_44850# a_18579_44172# 7.6e-20
C44472 a_n699_43396# a_n984_44318# 2.34e-20
C44473 a_742_44458# a_1467_44172# 0.018499f
C44474 a_13213_44734# a_13468_44734# 0.005172f
C44475 a_18443_44721# a_18681_44484# 0.001705f
C44476 a_9482_43914# a_9801_43940# 8.96e-19
C44477 a_1307_43914# a_5326_44056# 0.001893f
C44478 a_n913_45002# a_1756_43548# 3.6e-21
C44479 a_n2017_45002# a_4235_43370# 2.25e-19
C44480 a_n1059_45260# a_4093_43548# 0.001865f
C44481 a_327_44734# a_n97_42460# 2.31e-20
C44482 a_3357_43084# a_3626_43646# 0.018539f
C44483 a_n467_45028# VDD 0.385804f
C44484 a_n2661_43370# a_3147_46376# 9.13e-21
C44485 a_11827_44484# a_11415_45002# 0.169126f
C44486 a_11361_45348# a_3483_46348# 5.71e-19
C44487 a_21005_45260# a_12741_44636# 0.001247f
C44488 a_18287_44626# a_15227_44166# 5.33e-20
C44489 a_5891_43370# a_8270_45546# 0.052984f
C44490 a_7281_43914# a_768_44030# 0.006034f
C44491 a_n2065_43946# a_n2293_46634# 2.74e-19
C44492 a_5111_44636# a_526_44458# 0.338508f
C44493 a_5147_45002# a_n1925_42282# 9.69e-37
C44494 a_11963_45334# a_10809_44734# 4.58e-19
C44495 a_1307_43914# a_17715_44484# 3.38e-21
C44496 a_n822_43940# a_n1613_43370# 2.39e-19
C44497 a_10949_43914# a_11453_44696# 7.02e-20
C44498 a_13483_43940# a_12465_44636# 3.64e-19
C44499 a_n2433_43396# a_n2497_47436# 0.173242f
C44500 a_15493_43940# a_16327_47482# 0.04211f
C44501 a_961_42354# a_7174_31319# 4.84e-21
C44502 a_10533_42308# a_11551_42558# 2.25e-19
C44503 a_10723_42308# a_5742_30871# 0.185564f
C44504 a_1606_42308# a_13258_32519# 0.001369f
C44505 a_n4318_38216# a_n4334_39616# 1.11e-19
C44506 a_5342_30871# C0_N_btm 8.41e-20
C44507 a_5534_30871# C2_N_btm 7.46e-20
C44508 C9_P_btm VIN_P 1.82823f
C44509 a_n1435_47204# a_9290_44172# 6.71e-22
C44510 a_6151_47436# a_14840_46494# 4.06e-20
C44511 a_n2109_47186# a_n1925_42282# 2.07e-20
C44512 a_4883_46098# a_1823_45246# 0.00603f
C44513 a_2747_46873# a_n2293_46098# 3.99e-20
C44514 a_19321_45002# a_17339_46660# 1.05e-20
C44515 a_5257_43370# a_6755_46942# 8.35e-20
C44516 a_6540_46812# a_6682_46660# 0.007833f
C44517 a_8492_46660# a_9863_46634# 5.2e-20
C44518 a_8667_46634# a_10150_46912# 5.2e-20
C44519 a_13661_43548# a_18285_46348# 0.049064f
C44520 a_5807_45002# a_19123_46287# 0.006772f
C44521 a_n2661_42834# a_n1821_43396# 4.8e-19
C44522 a_10193_42453# a_8515_42308# 1.05e-20
C44523 a_16922_45042# a_20301_43646# 0.00515f
C44524 a_3499_42826# a_3820_44260# 5.31e-19
C44525 a_2711_45572# a_15803_42450# 1.02e-20
C44526 a_7499_43078# a_8325_42308# 2.16e-19
C44527 a_9482_43914# a_12545_42858# 1.33e-20
C44528 a_20193_45348# a_15743_43084# 0.060559f
C44529 a_1307_43914# a_10083_42826# 4.67e-20
C44530 a_1423_45028# a_7765_42852# 5.7e-21
C44531 a_n2293_42834# a_n1076_43230# 0.01241f
C44532 a_11691_44458# a_19268_43646# 1.97e-21
C44533 a_n356_44636# a_6197_43396# 1.09e-20
C44534 a_10157_44484# a_9145_43396# 4.85e-21
C44535 a_9838_44484# a_9803_43646# 7.04e-22
C44536 a_n2661_43922# VDD 0.611934f
C44537 a_n4209_38216# C3_P_btm 0.041776f
C44538 a_n3565_38216# C5_P_btm 1.11e-20
C44539 a_n4209_38502# VIN_P 0.028945f
C44540 a_2711_45572# a_10193_42453# 0.218272f
C44541 a_6511_45714# a_7230_45938# 0.088127f
C44542 a_3775_45552# a_4880_45572# 1.54e-21
C44543 a_6667_45809# a_6812_45938# 0.057222f
C44544 a_6472_45840# a_8162_45546# 3.95e-19
C44545 a_5663_43940# a_1823_45246# 5.36e-19
C44546 a_3626_43646# a_3877_44458# 1.07e-19
C44547 a_16977_43638# a_12549_44172# 3.73e-20
C44548 a_13667_43396# a_n2293_46634# 0.011502f
C44549 a_n2661_42834# a_8034_45724# 5.76e-21
C44550 a_5883_43914# a_n357_42282# 1.93e-19
C44551 a_18579_44172# a_17715_44484# 2.18e-19
C44552 a_13467_32519# SMPL_ON_N 0.029246f
C44553 a_22591_43396# a_13507_46334# 0.011335f
C44554 a_19963_31679# a_19864_35138# 1.38e-21
C44555 a_20447_31679# a_18194_35068# 9.11e-20
C44556 a_7927_46660# VDD 0.187888f
C44557 a_n4064_38528# a_n4209_38216# 0.028013f
C44558 a_n3420_38528# a_n3565_38216# 0.035254f
C44559 a_7174_31319# C0_dummy_P_btm 0.029132f
C44560 a_13258_32519# C1_N_btm 0.001902f
C44561 a_22400_42852# CAL_N 0.001609f
C44562 a_22959_46660# a_21076_30879# 0.165603f
C44563 a_n1925_46634# a_n1099_45572# 0.001556f
C44564 a_n743_46660# a_n452_45724# 0.070244f
C44565 a_n2293_46634# a_n755_45592# 0.094759f
C44566 a_n2438_43548# a_n863_45724# 0.07341f
C44567 a_15227_44166# a_15682_46116# 1.07e-20
C44568 a_765_45546# a_4704_46090# 7.8e-21
C44569 a_17609_46634# a_17715_44484# 0.001359f
C44570 a_11901_46660# a_10809_44734# 0.048084f
C44571 a_15682_43940# a_16243_43396# 0.013782f
C44572 a_17737_43940# a_16137_43396# 2.97e-21
C44573 a_7499_43940# a_7287_43370# 8.47e-19
C44574 a_15493_43940# a_10341_43396# 0.051273f
C44575 a_11967_42832# a_12895_43230# 0.035759f
C44576 a_14539_43914# a_18504_43218# 1.37e-19
C44577 a_n447_43370# VDD 0.204801f
C44578 a_20841_45814# a_21350_45938# 2.6e-19
C44579 a_9159_45572# a_8953_45002# 0.001432f
C44580 a_2711_45572# a_14309_45348# 0.002115f
C44581 a_6194_45824# a_n2661_43370# 0.002009f
C44582 a_20273_45572# a_20719_45572# 2.28e-19
C44583 a_564_42282# a_768_44030# 4.13e-22
C44584 a_10922_42852# a_3090_45724# 0.002693f
C44585 a_7309_42852# a_4646_46812# 1.16e-20
C44586 a_4235_43370# a_526_44458# 0.032501f
C44587 a_4093_43548# a_n1925_42282# 0.018682f
C44588 a_5934_30871# a_4883_46098# 0.005052f
C44589 a_13249_42308# a_4915_47217# 0.161597f
C44590 a_13163_45724# a_6151_47436# 1.73e-21
C44591 a_11682_45822# a_2063_45854# 3.96e-19
C44592 a_19900_46494# a_16375_45002# 9.97e-21
C44593 a_19335_46494# a_19431_46494# 0.013793f
C44594 a_6945_45028# a_13259_45724# 7.64e-20
C44595 a_5066_45546# a_8034_45724# 0.242476f
C44596 a_3626_43646# a_5342_30871# 0.08847f
C44597 a_n97_42460# a_133_42852# 0.012177f
C44598 a_18783_43370# a_743_42282# 1.15e-20
C44599 a_19700_43370# a_21259_43561# 8.8e-21
C44600 a_19268_43646# a_4190_30871# 0.035721f
C44601 a_15743_43084# a_20301_43646# 1.96e-20
C44602 a_16759_43396# a_4361_42308# 7.84e-21
C44603 en_comp a_22521_40599# 0.021604f
C44604 a_13159_45002# a_11827_44484# 9.25e-21
C44605 a_8696_44636# a_15433_44458# 0.001482f
C44606 a_18479_45785# a_9313_44734# 5.83e-19
C44607 a_4558_45348# a_n2661_44458# 0.001813f
C44608 a_327_44734# a_742_44458# 0.005551f
C44609 a_413_45260# a_949_44458# 0.018785f
C44610 a_n467_45028# a_n699_43396# 7.07e-21
C44611 a_2075_43172# a_n863_45724# 2.8e-19
C44612 a_n1853_43023# a_n443_42852# 0.141267f
C44613 a_133_43172# a_n357_42282# 0.001058f
C44614 a_12895_43230# a_13259_45724# 6.21e-19
C44615 a_n4334_37440# SMPL_ON_P 4.8e-20
C44616 a_16115_45572# a_6755_46942# 0.004389f
C44617 a_7227_45028# a_765_45546# 2.27e-20
C44618 a_n2293_45010# a_n2438_43548# 0.033143f
C44619 a_n2956_37592# a_n2442_46660# 0.049818f
C44620 a_n2810_45028# a_n2293_46634# 0.004774f
C44621 a_n2433_44484# a_n2497_47436# 0.027254f
C44622 a_22459_39145# VDD 0.682253f
C44623 a_n1991_42858# a_n4318_38216# 4.7e-19
C44624 a_14579_43548# a_14456_42282# 5.92e-19
C44625 a_n2840_42826# a_n4318_37592# 2.65e-20
C44626 a_n2157_42858# a_n3674_38216# 3.67e-19
C44627 a_n1853_43023# a_n2104_42282# 2.35e-20
C44628 a_10341_42308# a_12800_43218# 5.31e-21
C44629 a_12089_42308# a_11554_42852# 8.72e-21
C44630 a_3626_43646# a_20107_42308# 0.001705f
C44631 a_n4318_39304# a_n4334_39392# 0.081919f
C44632 a_10796_42968# a_11136_42852# 0.027606f
C44633 a_13887_32519# a_n784_42308# 0.00652f
C44634 a_10341_43396# a_5742_30871# 3.28e-19
C44635 a_2982_43646# a_7174_31319# 0.081795f
C44636 a_2324_44458# CLK 0.035116f
C44637 a_n3690_39616# VDD 0.358567f
C44638 a_3422_30871# a_n4064_37984# 0.031408f
C44639 a_n2293_43922# VDAC_N 6.46e-20
C44640 a_584_46384# a_n881_46662# 0.286501f
C44641 a_2063_45854# a_n1613_43370# 0.04116f
C44642 a_2952_47436# a_3094_47243# 0.005572f
C44643 a_16327_47482# a_16763_47508# 0.338544f
C44644 a_13717_47436# a_20894_47436# 6.95e-20
C44645 a_15811_47375# a_10227_46804# 0.019973f
C44646 a_11599_46634# a_18479_47436# 0.005025f
C44647 a_16241_47178# a_16588_47582# 0.051162f
C44648 a_15673_47210# a_17591_47464# 1.51e-19
C44649 a_3785_47178# a_3315_47570# 2.31e-21
C44650 a_n1151_42308# a_2583_47243# 1.83e-19
C44651 a_8953_45002# a_9672_43914# 0.00114f
C44652 a_2711_45572# a_16137_43396# 1.42e-19
C44653 a_11691_44458# a_17061_44484# 0.005038f
C44654 a_n2661_43370# a_n2840_43914# 0.008144f
C44655 a_10057_43914# a_9313_44734# 0.139382f
C44656 a_18494_42460# a_20679_44626# 1.25e-20
C44657 a_11827_44484# a_11967_42832# 0.095859f
C44658 a_7499_43078# a_9145_43396# 0.040441f
C44659 a_4743_44484# a_n2661_42834# 9.88e-20
C44660 a_n699_43396# a_n2661_43922# 0.053529f
C44661 a_20567_45036# a_20640_44752# 0.003077f
C44662 a_18911_45144# a_19279_43940# 3.2e-20
C44663 a_n4209_38502# a_n2956_38680# 0.235751f
C44664 a_21076_30879# C10_N_btm 9.75e-19
C44665 a_17478_45572# VDD 0.411207f
C44666 a_5342_30871# C10_P_btm 2.16e-19
C44667 a_5534_30871# C8_P_btm 5.29e-19
C44668 a_15595_45028# a_11415_45002# 0.003773f
C44669 a_14537_43396# a_12741_44636# 0.094691f
C44670 a_3232_43370# a_1823_45246# 0.344002f
C44671 a_3429_45260# a_3699_46348# 7.23e-21
C44672 a_3537_45260# a_3483_46348# 0.605469f
C44673 a_3065_45002# a_4185_45028# 0.060303f
C44674 a_17023_45118# a_15227_44166# 2.94e-19
C44675 a_18184_42460# a_3090_45724# 2.47e-20
C44676 a_15463_44811# a_13661_43548# 1.29e-19
C44677 a_16115_45572# a_8049_45260# 0.004258f
C44678 a_20273_45572# a_6945_45028# 2.17e-19
C44679 a_20841_45814# a_21137_46414# 2.76e-19
C44680 a_20623_45572# a_20708_46348# 9.36e-19
C44681 a_2437_43646# a_15682_46116# 4.97e-20
C44682 a_3357_43084# a_15015_46420# 6.88e-21
C44683 a_n2017_45002# a_9290_44172# 0.089856f
C44684 a_16877_42852# a_15803_42450# 1.15e-19
C44685 a_n784_42308# a_8515_42308# 1.56e-20
C44686 a_3318_42354# a_3823_42558# 1e-19
C44687 a_961_42354# a_5932_42308# 4.31e-21
C44688 a_564_42282# a_6123_31319# 2.22e-20
C44689 a_4190_30871# C2_N_btm 9.13e-20
C44690 a_22521_39511# a_22545_38993# 0.27533f
C44691 a_22459_39145# a_22469_39537# 0.351623f
C44692 a_22521_40055# a_22780_39857# 3.15e-19
C44693 a_n2661_46634# a_7715_46873# 0.007284f
C44694 a_5807_45002# a_6755_46942# 1.47519f
C44695 a_2107_46812# a_4651_46660# 0.003567f
C44696 a_2609_46660# a_3524_46660# 0.118759f
C44697 a_2443_46660# a_2864_46660# 0.090164f
C44698 a_n1925_46634# a_3878_46660# 3.71e-19
C44699 a_n881_46662# a_11901_46660# 1.99e-19
C44700 a_10227_46804# a_13059_46348# 0.656528f
C44701 a_16588_47582# a_16721_46634# 0.001918f
C44702 a_15507_47210# a_765_45546# 0.00763f
C44703 a_17591_47464# a_16388_46812# 2.32e-20
C44704 a_15811_47375# a_17339_46660# 8.97e-20
C44705 a_13717_47436# a_20411_46873# 1.46e-20
C44706 a_n2497_47436# a_3147_46376# 7.92e-21
C44707 a_n1741_47186# a_167_45260# 4.69e-20
C44708 a_n237_47217# a_472_46348# 3.2e-19
C44709 a_n2109_47186# a_2698_46116# 5.63e-21
C44710 a_n785_47204# a_n1076_46494# 9.42e-21
C44711 a_2063_45854# a_n2293_46098# 0.994164f
C44712 a_n746_45260# a_805_46414# 1.34e-19
C44713 a_13249_42308# a_13291_42460# 0.068754f
C44714 a_n699_43396# a_n447_43370# 0.040315f
C44715 a_n2661_43370# a_9803_43646# 6.41e-22
C44716 a_9313_44734# a_14021_43940# 0.014591f
C44717 a_4223_44672# a_n97_42460# 1.53e-19
C44718 a_n1761_44111# a_895_43940# 7.07e-21
C44719 a_n2661_42834# a_9248_44260# 1.02e-20
C44720 a_n1059_45260# a_685_42968# 0.103646f
C44721 a_n967_45348# a_n1379_43218# 3.56e-19
C44722 a_4338_37500# VDD 0.525635f
C44723 a_n452_44636# VDD 0.112149f
C44724 a_18907_42674# RST_Z 1.72e-20
C44725 a_n3420_37984# a_n2810_45572# 6.34e-19
C44726 a_n1557_42282# a_768_44030# 1.25e-19
C44727 a_n4318_39304# a_n2312_38680# 0.023234f
C44728 a_10807_43548# a_8270_45546# 9.25e-21
C44729 a_n2129_43609# a_n2293_46634# 4.29e-21
C44730 a_11827_44484# a_13259_45724# 0.062801f
C44731 a_n2661_43370# a_310_45028# 0.027265f
C44732 a_9159_44484# a_8199_44636# 4.07e-19
C44733 a_n2661_42834# a_8016_46348# 0.041785f
C44734 a_5205_44734# a_2324_44458# 5.38e-19
C44735 a_15681_43442# a_12861_44030# 0.137136f
C44736 a_15095_43370# a_10227_46804# 0.264777f
C44737 a_n2946_39866# a_n4064_39616# 0.053228f
C44738 a_n4064_40160# a_n4209_39304# 0.04848f
C44739 a_n3420_39616# a_n2302_39866# 1.28e-19
C44740 a_n4315_30879# a_n3565_39304# 0.048127f
C44741 a_19594_46812# VDD 0.349555f
C44742 a_5932_42308# C0_dummy_P_btm 1.2e-19
C44743 a_15559_46634# a_11415_45002# 1.37e-20
C44744 a_3090_45724# a_12741_44636# 0.093609f
C44745 a_7715_46873# a_8199_44636# 2.07e-21
C44746 a_7577_46660# a_8349_46414# 0.001417f
C44747 a_7411_46660# a_5937_45572# 2.28e-21
C44748 a_7927_46660# a_7920_46348# 3.44e-19
C44749 a_n1925_46634# a_n1925_42282# 1.31e-19
C44750 a_n2438_43548# a_1431_46436# 4.38e-20
C44751 a_12891_46348# a_12379_46436# 0.006296f
C44752 a_n743_46660# a_2981_46116# 0.003499f
C44753 a_5807_45002# a_8049_45260# 1.37423f
C44754 a_19692_46634# a_18900_46660# 5.55e-20
C44755 en_comp a_13575_42558# 4.34e-21
C44756 a_n2017_45002# a_15051_42282# 0.006558f
C44757 a_n1059_45260# a_14113_42308# 4.15e-19
C44758 a_n2661_42834# a_n1736_43218# 5.14e-19
C44759 a_n2293_43922# a_n3674_39304# 1.03e-19
C44760 a_n356_44636# a_10922_42852# 2.27e-20
C44761 a_1307_43914# a_2351_42308# 0.00376f
C44762 a_14539_43914# a_16414_43172# 2.71e-20
C44763 a_15493_43940# a_n97_42460# 0.009021f
C44764 a_7640_43914# a_7871_42858# 3.94e-21
C44765 a_14021_43940# a_20974_43370# 0.893848f
C44766 a_5891_43370# a_5755_42852# 0.160849f
C44767 a_20935_43940# VDD 0.184334f
C44768 a_16333_45814# a_16842_45938# 2.6e-19
C44769 a_15765_45572# a_16211_45572# 2.28e-19
C44770 a_5263_45724# a_5147_45002# 5.54e-20
C44771 a_2711_45572# a_5691_45260# 0.004189f
C44772 a_7499_43078# a_n1059_45260# 0.277353f
C44773 a_n4064_37984# VREF_GND 0.047292f
C44774 a_4905_42826# a_1823_45246# 0.110836f
C44775 a_7765_42852# a_4646_46812# 0.122773f
C44776 a_15868_43402# a_3090_45724# 2.14e-21
C44777 a_2889_44172# a_n357_42282# 4.18e-22
C44778 a_n1899_43946# a_n443_42852# 2.87e-20
C44779 a_n4318_39768# a_n2840_45546# 7.96e-20
C44780 a_2351_42308# a_n443_46116# 2.33e-20
C44781 a_5164_46348# VDD 0.717083f
C44782 a_5263_45724# a_n2109_47186# 9.21e-19
C44783 a_n3565_39590# VDAC_P 0.003547f
C44784 a_2684_37794# VDAC_Pi 0.133177f
C44785 a_n3565_39304# a_n3420_37440# 0.032339f
C44786 a_n4209_39304# a_n4064_37440# 0.029715f
C44787 a_n4064_39072# a_n4209_37414# 0.030589f
C44788 a_n3420_39072# a_n3565_37414# 0.031846f
C44789 a_8016_46348# a_5066_45546# 0.054471f
C44790 a_9290_44172# a_526_44458# 0.200352f
C44791 a_6419_46155# a_6640_46482# 0.007833f
C44792 a_18819_46122# a_20708_46348# 2.33e-20
C44793 a_18985_46122# a_19900_46494# 0.118759f
C44794 a_17583_46090# a_10809_44734# 2.89e-21
C44795 a_18189_46348# a_6945_45028# 4.84e-20
C44796 a_n2065_43946# a_n1736_42282# 3.49e-22
C44797 a_104_43370# a_n13_43084# 7.16e-19
C44798 a_2982_43646# a_21487_43396# 0.169809f
C44799 a_14021_43940# a_18599_43230# 5.88e-20
C44800 a_9313_44734# a_15764_42576# 3.58e-20
C44801 a_n2293_43922# a_5742_30871# 0.098838f
C44802 a_n356_44636# a_17531_42308# 0.030778f
C44803 a_3626_43646# a_743_42282# 0.147999f
C44804 a_10341_43396# a_10849_43646# 1.08e-20
C44805 a_8685_43396# a_16547_43609# 7.59e-20
C44806 a_n1761_44111# a_n3674_38216# 5.92e-21
C44807 a_22612_30879# a_22459_39145# 7.31e-20
C44808 a_n1641_43230# VDD 0.203991f
C44809 a_5147_45002# a_5837_45348# 2.22e-19
C44810 a_5111_44636# a_5365_45348# 0.001271f
C44811 a_2680_45002# a_2809_45028# 0.062574f
C44812 a_4927_45028# a_5105_45348# 0.007617f
C44813 a_7705_45326# a_1423_45028# 2.06e-22
C44814 a_n913_45002# a_n2661_43370# 0.031604f
C44815 a_20623_45572# a_21101_45002# 0.00299f
C44816 a_10180_45724# a_9313_44734# 6.72e-20
C44817 a_11963_45334# a_1307_43914# 1.89e-20
C44818 a_13556_45296# a_14537_43396# 0.590856f
C44819 a_13777_45326# a_14180_45002# 0.002746f
C44820 a_9482_43914# a_14797_45144# 0.003056f
C44821 a_n4334_40480# a_n2312_38680# 3.37e-19
C44822 a_14358_43442# a_n443_42852# 0.037176f
C44823 a_791_42968# a_526_44458# 7.15e-19
C44824 a_685_42968# a_n1925_42282# 1.12e-20
C44825 a_6812_45938# a_5257_43370# 3.92e-20
C44826 a_6472_45840# a_6969_46634# 2.28e-19
C44827 a_6511_45714# a_6755_46942# 2.73e-20
C44828 a_19431_45546# a_12549_44172# 1.86e-19
C44829 a_413_45260# a_16327_47482# 2.72e-19
C44830 a_8953_45002# a_6151_47436# 4.09e-20
C44831 a_14180_45002# a_n1151_42308# 1.97e-20
C44832 a_1307_43914# a_584_46384# 0.314947f
C44833 a_2903_45348# a_n971_45724# 0.004883f
C44834 a_5837_45348# a_n2109_47186# 8.23e-19
C44835 a_n1099_45572# a_n310_45572# 2.46e-19
C44836 a_n863_45724# a_603_45572# 3.59e-21
C44837 a_n356_45724# a_n310_45899# 0.006879f
C44838 a_1848_45724# a_n443_42852# 5.35e-20
C44839 a_n755_45592# a_2277_45546# 0.065177f
C44840 a_10796_42968# a_12545_42858# 0.002859f
C44841 a_10991_42826# a_12089_42308# 3.42e-21
C44842 a_16137_43396# a_16877_42852# 0.010276f
C44843 a_15743_43084# a_15785_43172# 3.98e-19
C44844 a_n1076_43230# a_n914_42852# 0.006453f
C44845 a_n97_42460# a_5742_30871# 0.259664f
C44846 a_2982_43646# a_5932_42308# 0.073161f
C44847 a_3626_43646# a_5755_42308# 0.003368f
C44848 a_16243_43396# a_16245_42852# 5.04e-20
C44849 a_6031_43396# a_5379_42460# 1.01e-19
C44850 a_3726_37500# VDAC_P 0.059581f
C44851 a_5700_37509# a_6886_37412# 0.13762f
C44852 a_5088_37509# VDAC_N 0.420254f
C44853 a_4338_37500# a_8912_37509# 0.331796f
C44854 a_3422_30871# C0_P_btm 6.53e-20
C44855 a_10545_42558# VDD 0.004307f
C44856 a_3160_47472# a_3785_47178# 2.34e-19
C44857 a_2063_45854# a_4791_45118# 0.039758f
C44858 a_2905_45572# a_3815_47204# 0.00535f
C44859 a_n1151_42308# a_3381_47502# 0.051194f
C44860 a_584_46384# a_n443_46116# 0.496286f
C44861 a_n2109_47186# a_n1435_47204# 0.041807f
C44862 a_n1741_47186# a_11459_47204# 0.015445f
C44863 a_n237_47217# a_7227_47204# 0.013654f
C44864 a_n971_45724# a_6575_47204# 0.01923f
C44865 a_11691_44458# a_18248_44752# 0.040333f
C44866 a_n452_44636# a_n699_43396# 1.94e-21
C44867 a_n2661_44458# a_9838_44484# 0.006567f
C44868 a_11827_44484# a_18989_43940# 0.054716f
C44869 a_n2293_42834# a_n2293_43922# 0.031735f
C44870 a_949_44458# a_2779_44458# 5.8e-19
C44871 a_18184_42460# a_n356_44636# 0.05602f
C44872 a_16147_45260# a_18079_43940# 2.34e-19
C44873 a_413_45260# a_175_44278# 1.05e-19
C44874 a_n2017_45002# a_3905_42865# 5.53e-19
C44875 a_n913_45002# a_2998_44172# 1.35e-20
C44876 a_196_42282# a_n863_45724# 1.25e-19
C44877 a_n3674_37592# a_n2956_38216# 0.025763f
C44878 a_n4318_37592# a_n357_42282# 4.71e-21
C44879 a_3638_45822# VDD 2.13e-19
C44880 a_4190_30871# C8_P_btm 4.06e-19
C44881 a_13076_44458# a_12549_44172# 5.14e-20
C44882 a_8560_45348# a_7577_46660# 3.58e-21
C44883 a_14180_45002# a_14084_46812# 1.82e-22
C44884 a_13720_44458# a_12891_46348# 8.1e-19
C44885 a_9482_43914# a_14976_45028# 6.03e-19
C44886 a_n2661_44458# a_n2312_38680# 1.97e-21
C44887 a_n2129_44697# a_n2293_46634# 5.68e-19
C44888 a_13556_45296# a_3090_45724# 0.032207f
C44889 a_12883_44458# a_768_44030# 6.59e-19
C44890 a_21350_45938# a_11415_45002# 8.06e-20
C44891 a_6511_45714# a_8049_45260# 0.001936f
C44892 a_15143_45578# a_6945_45028# 1.11e-21
C44893 a_12016_45572# a_10903_43370# 3.71e-20
C44894 a_9313_44734# a_13507_46334# 0.145766f
C44895 a_n3674_39304# a_n3420_39616# 0.152699f
C44896 a_5342_30871# a_13921_42308# 8.71e-20
C44897 a_5837_42852# a_5932_42308# 4.77e-19
C44898 a_n1151_42308# a_15009_46634# 8.05e-19
C44899 a_14311_47204# a_6755_46942# 1.38e-20
C44900 a_11599_46634# a_10554_47026# 7.33e-21
C44901 a_4915_47217# a_11813_46116# 1.35e-19
C44902 a_6575_47204# a_8023_46660# 1.23e-19
C44903 a_9313_45822# a_8035_47026# 1.13e-19
C44904 a_6151_47436# a_10768_47026# 8.29e-20
C44905 a_4883_46098# a_5732_46660# 3.05e-22
C44906 a_n1613_43370# a_645_46660# 0.001903f
C44907 a_n881_46662# a_479_46660# 3.54e-19
C44908 a_20843_47204# a_21588_30879# 1e-19
C44909 a_n1059_45260# a_15781_43660# 4.06e-20
C44910 a_18114_32519# a_14021_43940# 2.66e-19
C44911 a_11967_42832# a_18005_44484# 2.11e-19
C44912 a_11823_42460# a_15567_42826# 3.26e-19
C44913 a_20362_44736# a_20835_44721# 7.99e-20
C44914 a_n2293_42834# a_n97_42460# 0.17628f
C44915 a_n2661_43370# a_n4318_39304# 0.00535f
C44916 a_10193_42453# a_18817_42826# 0.002321f
C44917 a_13249_42308# a_13460_43230# 0.014543f
C44918 a_5891_43370# a_7845_44172# 0.119969f
C44919 a_18588_44850# a_18579_44172# 9.38e-20
C44920 a_n2661_42834# a_1414_42308# 0.081864f
C44921 a_n2661_43922# a_1467_44172# 0.002845f
C44922 a_19615_44636# a_19279_43940# 1.59e-19
C44923 a_20640_44752# a_20679_44626# 0.582607f
C44924 a_5837_45028# VDD 0.191549f
C44925 a_5934_30871# a_n923_35174# 0.009397f
C44926 a_22521_40599# a_4185_45028# 3.39e-20
C44927 a_8701_44490# a_3483_46348# 1.31e-20
C44928 a_14815_43914# a_13059_46348# 0.004368f
C44929 a_20362_44736# a_3090_45724# 1.21e-21
C44930 a_15301_44260# a_12549_44172# 4.3e-19
C44931 a_15493_43396# a_n2293_46634# 4.09e-19
C44932 a_15595_45028# a_13259_45724# 2.25e-19
C44933 a_14537_43396# a_16375_45002# 3.44e-20
C44934 a_2382_45260# a_2957_45546# 2.8e-21
C44935 a_3429_45260# a_n755_45592# 2.78e-19
C44936 a_n37_45144# a_n23_45546# 0.001445f
C44937 a_3537_45260# a_n357_42282# 0.200175f
C44938 a_19778_44110# a_19900_46494# 9.85e-21
C44939 a_11691_44458# a_2324_44458# 0.045025f
C44940 a_18184_42460# a_20075_46420# 1.99e-20
C44941 a_4223_44672# a_5204_45822# 5.85e-20
C44942 a_11827_44484# a_18189_46348# 1.03e-19
C44943 a_20974_43370# a_13507_46334# 0.017855f
C44944 a_15673_47210# VDD 0.569224f
C44945 a_17303_42282# a_18907_42674# 1.62e-19
C44946 a_n743_46660# a_167_45260# 0.045398f
C44947 a_n1925_46634# a_2698_46116# 8.92e-20
C44948 a_n2661_46098# a_n2840_46090# 0.170439f
C44949 a_1123_46634# a_472_46348# 0.001483f
C44950 a_33_46660# a_1176_45822# 5.48e-19
C44951 a_383_46660# a_805_46414# 0.01072f
C44952 a_n2293_46634# a_3483_46348# 0.157275f
C44953 a_14084_46812# a_15009_46634# 4.66e-19
C44954 a_7715_46873# a_765_45546# 0.001838f
C44955 a_12891_46348# a_13351_46090# 0.019821f
C44956 a_5807_45002# a_8953_45546# 0.00249f
C44957 a_12549_44172# a_12594_46348# 0.031894f
C44958 a_n881_46662# a_17583_46090# 0.003148f
C44959 a_n2312_39304# a_n2956_38680# 0.048558f
C44960 a_14311_47204# a_8049_45260# 4.71e-21
C44961 a_11459_47204# a_10586_45546# 1.75e-22
C44962 a_n971_45724# a_n2661_45546# 0.083094f
C44963 a_n2497_47436# a_310_45028# 4.48e-20
C44964 a_n2661_46634# a_4419_46090# 1.65e-19
C44965 a_18248_44752# a_4190_30871# 2.51e-20
C44966 a_1115_44172# a_n97_42460# 1.16e-19
C44967 a_11341_43940# a_22223_43948# 0.175191f
C44968 a_14673_44172# a_8685_43396# 9.41e-20
C44969 a_21115_43940# a_15493_43940# 0.0516f
C44970 a_17737_43940# a_14021_43940# 2.4e-20
C44971 a_n2661_42282# a_5829_43940# 0.002389f
C44972 a_10193_42453# a_21421_42336# 1.05e-20
C44973 a_n2293_42834# a_3935_43218# 9.69e-20
C44974 en_comp a_n2104_42282# 0.002636f
C44975 a_n2017_45002# a_n961_42308# 0.012655f
C44976 a_n2810_45028# a_n1736_42282# 9.69e-21
C44977 a_n2956_37592# a_n3674_38216# 0.023192f
C44978 a_n967_45348# a_n4318_38216# 3e-20
C44979 a_n913_45002# COMP_P 1.4e-20
C44980 a_n809_44244# VDD 0.47719f
C44981 C0_P_btm VREF_GND 0.350485f
C44982 C1_P_btm VCM 0.716121f
C44983 a_2711_45572# a_18479_45785# 0.032371f
C44984 a_10490_45724# a_11778_45572# 0.004273f
C44985 a_11525_45546# a_11136_45572# 1.53e-19
C44986 C0_dummy_N_btm VIN_N 0.544204f
C44987 a_6293_42852# a_3090_45724# 0.003062f
C44988 a_3935_42891# a_768_44030# 2.15e-21
C44989 a_3905_42865# a_526_44458# 0.321601f
C44990 a_3600_43914# a_n1925_42282# 2.11e-19
C44991 a_18005_44484# a_13259_45724# 3.54e-19
C44992 a_12429_44172# a_12594_46348# 5.47e-22
C44993 a_10083_42826# a_n1613_43370# 1.52e-19
C44994 a_21195_42852# a_18597_46090# 0.01512f
C44995 a_18599_43230# a_13507_46334# 0.00421f
C44996 a_10775_45002# CLK 0.058141f
C44997 a_16388_46812# VDD 0.797417f
C44998 a_7174_31319# a_n4064_37984# 0.003259f
C44999 a_20885_46660# a_10809_44734# 3.49e-19
C45000 a_22365_46825# a_22223_46124# 0.011912f
C45001 a_12741_44636# a_20075_46420# 0.027561f
C45002 a_20202_43084# a_6945_45028# 0.02248f
C45003 a_3483_46348# a_9625_46129# 0.038063f
C45004 a_11415_45002# a_21137_46414# 6.03e-22
C45005 a_15559_46634# a_13259_45724# 9.61e-21
C45006 a_3090_45724# a_16375_45002# 0.026416f
C45007 a_5883_43914# a_8685_42308# 1.31e-20
C45008 a_1414_42308# a_n2293_42282# 1.08e-20
C45009 a_2982_43646# a_4181_43396# 1.27e-20
C45010 a_11967_42832# a_13569_43230# 8.29e-19
C45011 a_14021_43940# a_13887_32519# 0.020984f
C45012 a_6293_42852# a_6547_43396# 3.12e-19
C45013 a_18184_42460# a_18727_42674# 0.044914f
C45014 a_18494_42460# a_18057_42282# 0.085802f
C45015 a_n356_44636# a_2903_42308# 2.77e-19
C45016 a_n2661_42834# a_n3674_38680# 0.03399f
C45017 a_6031_43396# a_7287_43370# 0.042271f
C45018 a_6197_43396# a_6765_43638# 0.17072f
C45019 a_8333_44056# a_8387_43230# 7.4e-22
C45020 a_2553_47502# DATA[2] 2.89e-20
C45021 a_2952_47436# DATA[1] 7.06e-21
C45022 a_14955_43396# VDD 0.401358f
C45023 a_13527_45546# a_11691_44458# 2.01e-21
C45024 a_8568_45546# a_n2661_44458# 4.32e-21
C45025 a_6667_45809# a_6298_44484# 0.001371f
C45026 a_8696_44636# a_8560_45348# 6.21e-19
C45027 a_2711_45572# a_10057_43914# 7.42e-20
C45028 a_6194_45824# a_5883_43914# 1.36e-19
C45029 a_n2017_45002# a_5147_45002# 4.93e-22
C45030 a_n467_45028# a_327_44734# 6.38e-20
C45031 a_n2661_45010# a_3232_43370# 3.31e-19
C45032 a_14456_42282# a_5807_45002# 3.82e-19
C45033 a_13575_42558# a_13661_43548# 1.71e-20
C45034 a_11554_42852# a_3090_45724# 0.001994f
C45035 a_1049_43396# a_n357_42282# 0.001179f
C45036 a_5649_42852# a_10903_43370# 9.98e-20
C45037 a_17678_43396# a_17715_44484# 5.41e-20
C45038 a_3316_45546# VDD 0.428912f
C45039 a_6598_45938# a_n2661_46634# 2.77e-21
C45040 a_11322_45546# a_12549_44172# 0.001723f
C45041 a_13249_42308# a_n881_46662# 9.77e-19
C45042 a_n913_45002# a_n2497_47436# 0.019337f
C45043 a_n2472_45002# SMPL_ON_P 1.75e-19
C45044 a_2437_43646# a_1431_47204# 0.001971f
C45045 a_8696_44636# a_10227_46804# 0.089585f
C45046 a_15037_45618# a_13507_46334# 1.52e-20
C45047 a_18243_46436# a_18051_46116# 6.96e-20
C45048 a_19240_46482# a_19431_46494# 4.61e-19
C45049 a_15682_43940# a_15803_42450# 4.66e-19
C45050 a_n2433_43396# a_n4318_37592# 2.5e-20
C45051 a_n1076_43230# a_n13_43084# 3.14e-19
C45052 a_4361_42308# a_5111_42852# 5.5e-20
C45053 a_743_42282# a_8037_42858# 5.74e-20
C45054 a_n2129_43609# a_n1736_42282# 1.65e-20
C45055 a_n1991_42858# a_n1545_43230# 2.28e-19
C45056 a_n2157_42858# a_n967_43230# 2.56e-19
C45057 a_n1853_43023# a_n1379_43218# 0.002143f
C45058 a_n1641_43230# a_n4318_38680# 4.97e-20
C45059 a_16547_43609# a_17333_42852# 2.75e-20
C45060 a_14401_32519# a_n784_42308# 0.003982f
C45061 a_11341_43940# a_11323_42473# 2.29e-19
C45062 a_16137_43396# a_18817_42826# 8.32e-19
C45063 a_11186_47026# CLK 6.21e-21
C45064 a_3090_45724# RST_Z 1.8e-20
C45065 a_19326_42852# VDD 4.6e-19
C45066 a_6709_45028# a_7640_43914# 8.38e-19
C45067 a_3232_43370# a_8855_44734# 0.001723f
C45068 a_3537_45260# a_3363_44484# 9.26e-20
C45069 a_327_44734# a_n2661_43922# 0.005571f
C45070 a_21188_45572# a_20679_44626# 3.17e-20
C45071 a_20623_45572# a_20766_44850# 1.55e-20
C45072 a_18315_45260# a_11827_44484# 9.63e-19
C45073 a_18184_42460# a_20567_45036# 9.9e-21
C45074 a_16405_45348# a_16237_45028# 8.13e-19
C45075 a_11322_45546# a_12429_44172# 5.73e-21
C45076 a_11525_45546# a_11750_44172# 1.43e-21
C45077 a_n2293_42834# a_742_44458# 0.039916f
C45078 a_n2661_43370# a_n2661_44458# 1.0558f
C45079 a_10193_42453# a_15682_43940# 0.003859f
C45080 a_19778_44110# a_21005_45260# 0.135527f
C45081 a_16922_45042# a_11691_44458# 0.428229f
C45082 a_2711_45572# a_14021_43940# 0.029672f
C45083 a_13575_42558# a_4185_45028# 8.71e-20
C45084 a_n1329_42308# a_n1925_42282# 5.81e-19
C45085 a_13569_43230# a_13259_45724# 1.73e-19
C45086 a_9223_42460# a_8953_45546# 0.166987f
C45087 a_9885_42558# a_8016_46348# 5.79e-20
C45088 a_10907_45822# a_11415_45002# 0.050963f
C45089 a_8696_44636# a_17339_46660# 6.71e-19
C45090 a_1423_45028# a_2107_46812# 0.022467f
C45091 a_7705_45326# a_4646_46812# 0.003014f
C45092 a_3232_43370# a_5732_46660# 2.77e-21
C45093 a_2437_43646# a_11735_46660# 6.77e-20
C45094 a_413_45260# a_8667_46634# 2.03e-20
C45095 a_6171_45002# a_5907_46634# 1.1e-20
C45096 a_17613_45144# a_n881_46662# 0.001826f
C45097 a_6667_45809# a_5937_45572# 0.002606f
C45098 a_2711_45572# a_11133_46155# 1.16e-20
C45099 a_18114_32519# a_13507_46334# 0.001272f
C45100 a_n1655_44484# a_n1151_42308# 1.11e-19
C45101 a_4361_42308# a_9885_42308# 0.001144f
C45102 a_17021_43396# a_4958_30871# 5.45e-20
C45103 a_5534_30871# a_1606_42308# 0.030581f
C45104 a_15743_43084# a_19647_42308# 7.14e-19
C45105 a_5649_42852# a_15959_42545# 1.03e-19
C45106 a_19268_43646# a_19511_42282# 1.08e-19
C45107 a_20692_30879# a_21589_35634# 4.41e-20
C45108 a_12465_44636# a_12549_44172# 0.093222f
C45109 a_2747_46873# a_3411_47243# 6.35e-21
C45110 a_16327_47482# a_20916_46384# 3.47e-19
C45111 a_11599_46634# a_n2661_46634# 0.067552f
C45112 a_18780_47178# a_5807_45002# 1.88e-20
C45113 a_18479_47436# a_13661_43548# 0.024025f
C45114 a_17591_47464# a_19321_45002# 6.33e-21
C45115 a_18143_47464# a_13747_46662# 3.2e-19
C45116 a_11459_47204# a_n743_46660# 3.96e-21
C45117 a_6491_46660# a_2107_46812# 7.39e-21
C45118 a_n1435_47204# a_n1925_46634# 1.17e-19
C45119 a_n237_47217# a_4955_46873# 0.032268f
C45120 a_n971_45724# a_5385_46902# 5.88e-20
C45121 a_3160_47472# a_3699_46634# 7.39e-19
C45122 a_3381_47502# a_3177_46902# 2.56e-19
C45123 a_n1151_42308# a_2959_46660# 3.22e-19
C45124 a_2905_45572# a_3524_46660# 0.011982f
C45125 a_584_46384# a_1302_46660# 5.41e-21
C45126 a_n443_46116# a_479_46660# 1.72e-19
C45127 a_18443_44721# a_18579_44172# 5.4e-19
C45128 a_n2661_44458# a_2998_44172# 2.23e-19
C45129 a_n699_43396# a_n809_44244# 1.25e-19
C45130 a_18374_44850# a_18245_44484# 4.2e-19
C45131 a_18248_44752# a_18753_44484# 2.28e-19
C45132 a_742_44458# a_1115_44172# 0.001155f
C45133 a_1307_43914# a_5025_43940# 0.003108f
C45134 a_n37_45144# a_104_43370# 2.79e-21
C45135 a_n913_45002# a_1568_43370# 0.098659f
C45136 a_n1059_45260# a_1756_43548# 6.3e-22
C45137 a_n2017_45002# a_4093_43548# 5.54e-21
C45138 a_n967_45348# a_n1655_43396# 2.02e-19
C45139 a_413_45260# a_n97_42460# 1.07e-21
C45140 a_3357_43084# a_3540_43646# 0.001122f
C45141 a_n2302_39072# a_n2956_38216# 3.61e-19
C45142 a_n955_45028# VDD 0.004233f
C45143 a_n2661_43370# a_2804_46116# 1.16e-20
C45144 a_20567_45036# a_12741_44636# 0.007778f
C45145 a_21359_45002# a_11415_45002# 0.015551f
C45146 a_11827_44484# a_20202_43084# 0.032881f
C45147 a_8704_45028# a_3483_46348# 7.47e-19
C45148 a_18248_44752# a_15227_44166# 0.001323f
C45149 a_8375_44464# a_8270_45546# 1.34e-20
C45150 a_6453_43914# a_768_44030# 0.006009f
C45151 a_4558_45348# a_n1925_42282# 0.001226f
C45152 a_16751_45260# a_15682_46116# 3.1e-20
C45153 a_11787_45002# a_10809_44734# 0.007368f
C45154 a_10729_43914# a_11453_44696# 5.66e-20
C45155 a_12429_44172# a_12465_44636# 0.003194f
C45156 a_5326_44056# a_4791_45118# 1.55e-19
C45157 a_n4318_39304# a_n2497_47436# 3.31e-20
C45158 a_15493_43396# a_18597_46090# 1.64e-21
C45159 a_19862_44208# a_18479_47436# 0.138185f
C45160 a_1184_42692# a_7174_31319# 6.06e-21
C45161 a_10533_42308# a_5742_30871# 0.020913f
C45162 a_10723_42308# a_11323_42473# 0.008191f
C45163 a_n4318_37592# a_n4064_40160# 0.079413f
C45164 a_5534_30871# C1_N_btm 1.06e-19
C45165 a_5342_30871# C0_dummy_N_btm 1.91e-20
C45166 a_21589_35634# VIN_N 0.029423f
C45167 C10_P_btm VIN_P 3.66034f
C45168 START SINGLE_ENDED 0.002177f
C45169 a_11459_47204# a_11189_46129# 7.59e-19
C45170 a_n2109_47186# a_526_44458# 4.75e-20
C45171 a_2063_45854# a_6945_45028# 0.074119f
C45172 a_2609_46660# a_3090_45724# 2.67e-20
C45173 a_13747_46662# a_765_45546# 7.33e-19
C45174 a_5807_45002# a_18285_46348# 0.006196f
C45175 a_n2661_42834# a_n1190_43762# 1.25e-19
C45176 a_2711_45572# a_15764_42576# 1.23e-20
C45177 a_10193_42453# a_5934_30871# 6.18e-20
C45178 a_16922_45042# a_4190_30871# 0.353708f
C45179 a_n2293_43922# a_n2012_43396# 0.011692f
C45180 a_1307_43914# a_8952_43230# 1.54e-20
C45181 a_1423_45028# a_7871_42858# 3.55e-21
C45182 a_n2293_42834# a_n901_43156# 0.021108f
C45183 a_19113_45348# a_19268_43646# 1.84e-21
C45184 a_11691_44458# a_15743_43084# 3.24e-19
C45185 a_n356_44636# a_6293_42852# 2.26e-20
C45186 a_22485_44484# a_14021_43940# 1.69e-19
C45187 a_9838_44484# a_9145_43396# 2.26e-22
C45188 a_n2661_42834# VDD 1.00348f
C45189 a_n4209_38216# C4_P_btm 0.001041f
C45190 a_n3565_38216# C6_P_btm 1.26e-20
C45191 a_2711_45572# a_10180_45724# 0.01318f
C45192 a_6472_45840# a_7230_45938# 0.05936f
C45193 a_6511_45714# a_6812_45938# 9.73e-19
C45194 a_6598_45938# a_6428_45938# 2.6e-19
C45195 a_5495_43940# a_1823_45246# 0.001058f
C45196 a_2982_43646# a_4646_46812# 2.9e-20
C45197 a_10695_43548# a_n2293_46634# 0.007256f
C45198 a_16409_43396# a_12549_44172# 3.09e-19
C45199 a_7499_43940# a_3090_45724# 0.025901f
C45200 a_n699_43396# a_3316_45546# 1.1e-20
C45201 a_8103_44636# a_n755_45592# 4.46e-21
C45202 a_20362_44736# a_20075_46420# 4.79e-20
C45203 a_20159_44458# a_19900_46494# 7.47e-21
C45204 a_13887_32519# a_13507_46334# 0.08088f
C45205 a_20447_31679# EN_VIN_BSTR_N 0.002888f
C45206 a_8145_46902# VDD 0.199702f
C45207 a_n4064_38528# a_n3607_38528# 7.1e-19
C45208 a_n3420_38528# a_n4334_38304# 0.014479f
C45209 a_n2946_38778# a_n4209_38216# 5.32e-20
C45210 a_n3690_38528# a_n3565_38216# 7.97e-20
C45211 a_13258_32519# C0_N_btm 0.033333f
C45212 a_7174_31319# C0_P_btm 0.050478f
C45213 a_12741_44636# a_21076_30879# 0.00607f
C45214 a_n2293_46634# a_n357_42282# 0.034749f
C45215 a_n2661_46634# a_1848_45724# 2.19e-20
C45216 a_n743_46660# a_n863_45724# 0.007504f
C45217 a_n133_46660# a_n2293_45546# 1.48e-22
C45218 a_7577_46660# a_8034_45724# 1.64e-20
C45219 a_13661_43548# a_n443_42852# 0.045364f
C45220 a_3090_45724# a_18985_46122# 1.47e-19
C45221 a_15227_44166# a_2324_44458# 0.190521f
C45222 a_17609_46634# a_17583_46090# 0.008733f
C45223 a_11813_46116# a_10809_44734# 0.001353f
C45224 a_n4318_37592# a_n4064_37440# 0.04779f
C45225 a_n1630_35242# a_3754_38470# 9.47e-20
C45226 a_5932_42308# a_n4064_37984# 0.003117f
C45227 a_765_45546# a_4419_46090# 8e-20
C45228 a_15682_43940# a_16137_43396# 0.004591f
C45229 a_7542_44172# a_4361_42308# 2.2e-21
C45230 a_17517_44484# a_17595_43084# 1.18e-21
C45231 a_11967_42832# a_13113_42826# 0.021992f
C45232 a_n1352_43396# a_n1190_43762# 0.006453f
C45233 a_n1917_43396# a_n1655_43396# 0.001705f
C45234 a_14539_43914# a_17141_43172# 0.00164f
C45235 a_22223_43948# a_10341_43396# 0.002507f
C45236 en_comp a_1736_39587# 8.86e-19
C45237 a_n1352_43396# VDD 0.288329f
C45238 a_11682_45822# a_11963_45334# 2.91e-20
C45239 a_5907_45546# a_n2661_43370# 0.007276f
C45240 a_13249_42308# a_1307_43914# 0.056917f
C45241 a_20273_45572# a_21350_45938# 1.46e-19
C45242 a_5837_42852# a_4646_46812# 1.26e-20
C45243 a_10991_42826# a_3090_45724# 0.004747f
C45244 a_4093_43548# a_526_44458# 0.107158f
C45245 a_8685_43396# a_10903_43370# 0.031035f
C45246 a_n356_44636# RST_Z 2.99e-19
C45247 a_5066_45546# VDD 1.34058f
C45248 a_2711_45572# a_13507_46334# 9.2e-19
C45249 a_13904_45546# a_4915_47217# 0.013453f
C45250 a_11280_45822# a_2063_45854# 0.009384f
C45251 a_8953_45546# a_n755_45592# 3.44e-19
C45252 a_19553_46090# a_19431_46494# 3.16e-19
C45253 a_19335_46494# a_19240_46482# 0.049827f
C45254 a_4185_45028# a_n443_42852# 0.027973f
C45255 a_11967_42832# a_18214_42558# 8.49e-19
C45256 a_7281_43914# a_7227_42308# 1.21e-20
C45257 a_2982_43646# a_15567_42826# 2.67e-20
C45258 a_3499_42826# a_3318_42354# 4.85e-19
C45259 a_18525_43370# a_743_42282# 5.58e-21
C45260 a_16243_43396# a_5649_42852# 8.11e-21
C45261 a_15743_43084# a_4190_30871# 0.290729f
C45262 a_9396_43370# a_8952_43230# 6.44e-19
C45263 a_16977_43638# a_4361_42308# 4.56e-21
C45264 a_n2661_46098# DATA[1] 9e-20
C45265 a_n2293_42282# VDD 0.464485f
C45266 en_comp CAL_N 0.024527f
C45267 a_13017_45260# a_11827_44484# 2.91e-21
C45268 a_16751_45260# a_17023_45118# 0.13675f
C45269 a_8696_44636# a_14815_43914# 0.002482f
C45270 a_10193_42453# a_20512_43084# 0.086337f
C45271 a_6125_45348# a_n2661_43370# 8.72e-19
C45272 a_4574_45260# a_n2661_44458# 6.04e-19
C45273 a_413_45260# a_742_44458# 0.001341f
C45274 a_327_44734# a_n452_44636# 5.28e-19
C45275 a_n913_45002# a_5883_43914# 1.2e-19
C45276 a_n784_42308# a_1823_45246# 6e-20
C45277 a_n2157_42858# a_n443_42852# 8.79e-20
C45278 a_1847_42826# a_n863_45724# 0.216819f
C45279 a_4520_42826# a_n2661_45546# 2.03e-19
C45280 a_5457_43172# a_526_44458# 7.33e-19
C45281 a_13113_42826# a_13259_45724# 1.98e-19
C45282 a_n4209_37414# SMPL_ON_P 8.3e-19
C45283 a_6598_45938# a_765_45546# 2.98e-21
C45284 a_16333_45814# a_6755_46942# 0.001253f
C45285 a_n2472_45002# a_n2438_43548# 0.023014f
C45286 a_n745_45366# a_n2293_46634# 0.006631f
C45287 a_6171_45002# a_768_44030# 0.027851f
C45288 a_n2810_45028# a_n2442_46660# 0.045466f
C45289 a_8191_45002# a_8128_46384# 2.38e-19
C45290 a_11827_44484# a_2063_45854# 8.5e-20
C45291 a_n2661_44458# a_n2497_47436# 0.138848f
C45292 a_22521_40055# VDD 1.04757f
C45293 a_19335_46494# START 6.85e-21
C45294 a_14840_46494# CLK 5.5e-21
C45295 a_n1853_43023# a_n4318_38216# 8.05e-19
C45296 a_n2157_42858# a_n2104_42282# 0.011248f
C45297 a_10835_43094# a_11136_42852# 9.73e-19
C45298 a_12379_42858# a_11554_42852# 2.33e-21
C45299 a_3626_43646# a_13258_32519# 0.006214f
C45300 a_2982_43646# a_20712_42282# 0.003556f
C45301 a_n4318_39304# a_n4209_39304# 0.135369f
C45302 a_4190_30871# a_1606_42308# 0.018892f
C45303 a_9145_43396# a_13657_42558# 4.78e-19
C45304 a_17364_32525# COMP_P 9.77e-21
C45305 a_20075_46420# RST_Z 3.65e-21
C45306 a_n3565_39590# VDD 1.26658f
C45307 a_584_46384# a_n1613_43370# 0.085833f
C45308 a_16327_47482# a_16023_47582# 0.159305f
C45309 a_15507_47210# a_10227_46804# 0.23187f
C45310 a_15673_47210# a_16588_47582# 0.125324f
C45311 a_9863_47436# a_4883_46098# 9.51e-21
C45312 a_3785_47178# a_3094_47570# 1.78e-21
C45313 a_n1151_42308# a_2266_47243# 2.81e-19
C45314 a_13717_47436# a_19787_47423# 6.87e-20
C45315 a_8953_45002# a_9028_43914# 0.001179f
C45316 a_6171_45002# a_13483_43940# 2.43e-21
C45317 a_7499_43078# a_8423_43396# 4.14e-19
C45318 a_11691_44458# a_16789_44484# 3.16e-19
C45319 a_18494_42460# a_20640_44752# 1.1e-19
C45320 a_5343_44458# a_9159_44484# 2.67e-20
C45321 a_11827_44484# a_19006_44850# 0.002956f
C45322 a_n2293_42834# a_n984_44318# 1.22e-19
C45323 a_18184_42460# a_20679_44626# 7.45e-21
C45324 a_19778_44110# a_20835_44721# 8.16e-19
C45325 a_10440_44484# a_9313_44734# 0.027369f
C45326 a_n699_43396# a_n2661_42834# 0.131393f
C45327 a_4223_44672# a_n2661_43922# 0.059715f
C45328 a_21359_45002# a_11967_42832# 1.28e-19
C45329 a_20567_45036# a_20362_44736# 6.75e-19
C45330 a_15861_45028# VDD 0.690795f
C45331 a_21076_30879# C9_N_btm 0.001137f
C45332 a_5534_30871# C9_P_btm 7.29e-20
C45333 a_15415_45028# a_11415_45002# 0.0035f
C45334 a_3065_45002# a_3699_46348# 3.29e-21
C45335 a_3429_45260# a_3483_46348# 4.53e-19
C45336 a_17613_45144# a_17609_46634# 4.03e-21
C45337 a_3537_45260# a_3147_46376# 1.82e-19
C45338 a_16922_45042# a_15227_44166# 0.533576f
C45339 a_15433_44458# a_13747_46662# 1.47e-21
C45340 a_3363_44484# a_n2293_46634# 0.001146f
C45341 a_14673_44172# a_768_44030# 2.39e-20
C45342 a_19778_44110# a_3090_45724# 9.48e-19
C45343 a_5343_44458# a_7715_46873# 2.03e-20
C45344 a_16333_45814# a_8049_45260# 0.002964f
C45345 a_8696_44636# a_8034_45724# 9.58e-21
C45346 a_20273_45572# a_21137_46414# 0.002347f
C45347 a_20107_45572# a_6945_45028# 1.37e-19
C45348 a_3357_43084# a_14275_46494# 4.55e-22
C45349 a_413_45260# a_5204_45822# 4.29e-21
C45350 a_2437_43646# a_2324_44458# 0.011046f
C45351 a_20841_45814# a_20708_46348# 1.63e-19
C45352 en_comp a_8199_44636# 4.34e-21
C45353 a_22485_44484# a_13507_46334# 0.008777f
C45354 a_16245_42852# a_15803_42450# 4.81e-19
C45355 a_1755_42282# a_4921_42308# 0.002752f
C45356 a_n784_42308# a_5934_30871# 0.142087f
C45357 a_1184_42692# a_5932_42308# 4.31e-21
C45358 a_4190_30871# C1_N_btm 7.67e-20
C45359 a_22459_39145# a_22821_38993# 0.013073f
C45360 a_22521_40055# a_22469_39537# 0.037283f
C45361 a_5807_45002# a_10249_46116# 0.041839f
C45362 a_n2661_46634# a_7411_46660# 0.023716f
C45363 a_2107_46812# a_4646_46812# 0.03082f
C45364 a_3177_46902# a_2959_46660# 0.209641f
C45365 a_2609_46660# a_3699_46634# 0.042415f
C45366 a_2443_46660# a_3524_46660# 0.102325f
C45367 a_n2661_46098# a_2864_46660# 7.93e-22
C45368 a_n1925_46634# a_3633_46660# 2.55e-19
C45369 a_n881_46662# a_11813_46116# 8.63e-20
C45370 a_16588_47582# a_16388_46812# 3.64e-19
C45371 a_11599_46634# a_765_45546# 0.332797f
C45372 a_16763_47508# a_16721_46634# 0.005734f
C45373 a_10227_46804# a_15227_46910# 0.00877f
C45374 a_13717_47436# a_20107_46660# 1.28e-20
C45375 a_n2497_47436# a_2804_46116# 8.29e-22
C45376 a_n1741_47186# a_2202_46116# 6.06e-23
C45377 a_584_46384# a_n2293_46098# 0.039917f
C45378 a_n746_45260# a_472_46348# 0.002816f
C45379 a_n2109_47186# a_2521_46116# 1.58e-20
C45380 a_n237_47217# a_376_46348# 2.21e-19
C45381 a_2779_44458# a_n97_42460# 1.5e-20
C45382 a_175_44278# a_644_44056# 0.00101f
C45383 a_n699_43396# a_n1352_43396# 0.003121f
C45384 a_n2661_43370# a_9145_43396# 1.28e-20
C45385 a_n2017_45002# a_685_42968# 9.17e-20
C45386 a_n967_45348# a_n1545_43230# 5.71e-19
C45387 a_3726_37500# VDD 0.341303f
C45388 a_n1352_44484# VDD 0.276725f
C45389 a_18727_42674# RST_Z 3.5e-20
C45390 a_n3690_38304# a_n2810_45572# 4.13e-19
C45391 a_19279_43940# a_11415_45002# 0.003698f
C45392 a_15493_43396# a_6755_46942# 8.69e-20
C45393 a_n2661_43370# a_n1099_45572# 2.12e-19
C45394 a_10157_44484# a_526_44458# 4.13e-20
C45395 a_4181_44734# a_2324_44458# 3.09e-19
C45396 a_5708_44484# a_5937_45572# 5.12e-19
C45397 a_4361_42308# a_n971_45724# 6.67e-20
C45398 a_14621_43646# a_12861_44030# 1.73e-20
C45399 a_14205_43396# a_10227_46804# 0.422372f
C45400 a_8685_43396# a_4883_46098# 0.011038f
C45401 a_n3420_39616# a_n4064_39616# 6.66063f
C45402 a_n3565_39590# a_n2860_39866# 2.96e-19
C45403 a_7174_31319# comp_n 1.92e-19
C45404 a_19321_45002# VDD 1.01574f
C45405 a_5932_42308# C0_P_btm 0.015561f
C45406 a_22165_42308# CAL_N 8.8e-21
C45407 a_22959_47212# a_20692_30879# 1.9e-19
C45408 a_18597_46090# a_n357_42282# 0.250702f
C45409 a_8145_46902# a_7920_46348# 8.72e-19
C45410 a_7577_46660# a_8016_46348# 0.003484f
C45411 a_7411_46660# a_8199_44636# 1.09e-20
C45412 a_5257_43370# a_5937_45572# 0.262028f
C45413 a_n2438_43548# a_1337_46436# 0.001827f
C45414 a_n743_46660# a_1431_46436# 0.004109f
C45415 a_n2312_38680# a_n1925_42282# 4.88e-20
C45416 a_n1925_46634# a_526_44458# 1.65e-19
C45417 a_19692_46634# a_18280_46660# 2.23e-20
C45418 a_19333_46634# a_19636_46660# 0.001377f
C45419 a_13059_46348# a_15312_46660# 3.94e-19
C45420 a_6755_46942# a_3483_46348# 0.014154f
C45421 a_15368_46634# a_11415_45002# 0.001587f
C45422 a_n2017_45002# a_14113_42308# 0.006853f
C45423 en_comp a_13070_42354# 4.34e-21
C45424 a_5205_44484# a_6761_42308# 1.57e-19
C45425 a_17517_44484# a_13467_32519# 2.74e-21
C45426 a_1307_43914# a_2123_42473# 0.001341f
C45427 a_n356_44636# a_10991_42826# 4.8e-20
C45428 a_11967_42832# a_16823_43084# 0.093759f
C45429 a_14539_43914# a_15567_42826# 1.35e-20
C45430 a_n2293_43922# a_n13_43084# 4.46e-21
C45431 a_n2661_42834# a_n4318_38680# 0.102282f
C45432 a_14021_43940# a_14401_32519# 0.059818f
C45433 a_18579_44172# a_19700_43370# 0.175511f
C45434 a_n699_43396# a_n2293_42282# 5.03e-21
C45435 a_7640_43914# a_7227_42852# 1.75e-20
C45436 a_20623_43914# VDD 0.258478f
C45437 a_15765_45572# a_16842_45938# 1.46e-19
C45438 a_7499_43078# a_n2017_45002# 0.065458f
C45439 a_2711_45572# a_4927_45028# 0.006854f
C45440 a_n3420_37984# VCM 0.014539f
C45441 a_3080_42308# a_1823_45246# 0.049986f
C45442 a_15743_43084# a_15227_44166# 0.513622f
C45443 a_7871_42858# a_4646_46812# 0.26422f
C45444 a_1414_42308# a_3218_45724# 3.53e-21
C45445 a_2675_43914# a_n357_42282# 1.8e-19
C45446 a_15493_43396# a_8049_45260# 6.61e-22
C45447 a_n1761_44111# a_n443_42852# 0.007283f
C45448 a_895_43940# a_n755_45592# 8.1e-20
C45449 a_7754_39632# RST_Z 0.030938f
C45450 a_n4064_37984# VREF 3.68e-19
C45451 a_20753_42852# a_16327_47482# 0.00568f
C45452 a_n4209_37414# a_n1532_35090# 8.48e-20
C45453 a_n3565_37414# a_n1838_35608# 1.2e-19
C45454 a_5068_46348# VDD 0.085085f
C45455 a_2711_45572# a_n1741_47186# 6.27e-20
C45456 a_4099_45572# a_n2109_47186# 8.98e-22
C45457 a_3483_46348# a_8049_45260# 0.012066f
C45458 a_765_45546# a_1848_45724# 2.79e-19
C45459 a_7920_46348# a_5066_45546# 0.04093f
C45460 a_18985_46122# a_20075_46420# 0.042415f
C45461 a_18819_46122# a_19900_46494# 0.102355f
C45462 a_19553_46090# a_19335_46494# 0.209641f
C45463 a_17715_44484# a_6945_45028# 8.4e-20
C45464 a_15682_46116# a_10809_44734# 4.63e-19
C45465 a_1736_39043# VDAC_Ni 5.86e-19
C45466 a_n3565_39304# a_n3690_37440# 2.75e-19
C45467 a_n4209_39304# a_n2946_37690# 2.26e-19
C45468 a_n3420_39072# a_n4334_37440# 2.36e-19
C45469 a_n3565_38216# a_n2216_37984# 0.003076f
C45470 a_n2433_43396# a_n1533_42852# 1.07e-19
C45471 a_n97_42460# a_n13_43084# 0.13246f
C45472 a_8685_43396# a_16243_43396# 3.52e-19
C45473 a_2982_43646# a_20556_43646# 8.33e-20
C45474 a_n2293_43922# a_11323_42473# 3.54e-20
C45475 a_9313_44734# a_15486_42560# 8.95e-20
C45476 a_n356_44636# a_17303_42282# 0.10316f
C45477 a_10341_43396# a_10765_43646# 7.4e-20
C45478 a_4905_42826# a_5649_42852# 0.003104f
C45479 a_n1761_44111# a_n2104_42282# 1.67e-20
C45480 a_19237_31679# COMP_P 1.7e-20
C45481 a_n1352_43396# a_n4318_38680# 2.18e-20
C45482 a_2747_46873# DATA[2] 5.46e-20
C45483 a_7_47243# DATA[0] 0.001094f
C45484 a_22612_30879# a_22521_40055# 4.85e-20
C45485 a_21588_30879# a_22459_39145# 6.4e-20
C45486 a_n1423_42826# VDD 0.211036f
C45487 a_20623_45572# a_21005_45260# 0.002863f
C45488 a_n1059_45260# a_n2661_43370# 0.03635f
C45489 a_6709_45028# a_1423_45028# 2.16e-20
C45490 a_20841_45814# a_21101_45002# 0.001934f
C45491 a_n467_45028# a_n2293_42834# 8.59e-21
C45492 a_2382_45260# a_2809_45028# 0.034331f
C45493 a_5147_45002# a_5365_45348# 0.001577f
C45494 a_4558_45348# a_5837_45348# 5.43e-21
C45495 a_3232_43370# a_3602_45348# 7.02e-20
C45496 a_10053_45546# a_9313_44734# 5.63e-20
C45497 a_9482_43914# a_14537_43396# 0.040878f
C45498 a_11787_45002# a_1307_43914# 1.91e-21
C45499 a_20107_45572# a_11827_44484# 2.61e-21
C45500 a_20273_45572# a_21359_45002# 5.74e-20
C45501 a_12800_43218# a_12741_44636# 3.89e-21
C45502 a_n4315_30879# a_n2312_38680# 0.024522f
C45503 a_n2302_40160# a_n2442_46660# 0.017419f
C45504 a_n4209_39590# a_n2956_39768# 0.334714f
C45505 a_14579_43548# a_n443_42852# 0.04846f
C45506 a_685_42968# a_526_44458# 1.6e-19
C45507 a_16823_43084# a_13259_45724# 0.017563f
C45508 a_15037_45618# a_n743_46660# 3.95e-20
C45509 a_6472_45840# a_6755_46942# 1.91e-20
C45510 a_19963_31679# SMPL_ON_N 0.029334f
C45511 a_413_45260# a_16241_47178# 8.41e-20
C45512 a_13777_45326# a_n1151_42308# 2.49e-21
C45513 a_2809_45348# a_n971_45724# 0.00154f
C45514 a_n863_45724# a_509_45572# 3.95e-21
C45515 a_n755_45592# a_1609_45822# 0.12055f
C45516 a_n356_45724# a_n23_45546# 0.360492f
C45517 a_997_45618# a_n443_42852# 0.093108f
C45518 a_16137_43396# a_16245_42852# 0.016079f
C45519 a_3080_42308# a_5934_30871# 1.27306f
C45520 a_n97_42460# a_11323_42473# 0.003208f
C45521 a_2982_43646# a_6171_42473# 8.09e-20
C45522 a_10796_42968# a_12089_42308# 1.05e-19
C45523 a_10922_42852# a_10341_42308# 0.053077f
C45524 a_10835_43094# a_12545_42858# 3.81e-19
C45525 a_12741_44636# SINGLE_ENDED 1.02e-19
C45526 a_21076_30879# RST_Z 0.052228f
C45527 a_5088_37509# a_6886_37412# 0.136505f
C45528 a_4338_37500# VDAC_N 0.046178f
C45529 a_3726_37500# a_8912_37509# 0.267651f
C45530 a_3422_30871# C1_P_btm 7.67e-20
C45531 a_9885_42558# VDD 0.18767f
C45532 a_3160_47472# a_3381_47502# 0.099936f
C45533 a_2124_47436# a_n443_46116# 6.88e-22
C45534 a_2905_45572# a_3785_47178# 0.013619f
C45535 a_n2288_47178# a_n1435_47204# 2.38e-19
C45536 a_n1741_47186# a_9313_45822# 0.102019f
C45537 a_n971_45724# a_7903_47542# 7.01e-19
C45538 a_n237_47217# a_6851_47204# 8.46e-19
C45539 a_n2661_44458# a_5883_43914# 0.010478f
C45540 a_742_44458# a_2779_44458# 2.48e-21
C45541 a_11691_44458# a_17970_44736# 0.040435f
C45542 a_11827_44484# a_18374_44850# 0.004504f
C45543 a_16147_45260# a_17973_43940# 1.63e-19
C45544 a_10193_42453# a_21381_43940# 1.29e-19
C45545 a_n2293_42834# a_n2661_43922# 0.03113f
C45546 a_n37_45144# a_175_44278# 8.37e-20
C45547 a_n913_45002# a_2889_44172# 6.01e-22
C45548 a_n1059_45260# a_2998_44172# 3.88e-20
C45549 a_n1736_42282# a_n357_42282# 2.32e-20
C45550 a_n1630_35242# a_n2810_45572# 5.26e-19
C45551 a_3775_45552# VDD 0.089667f
C45552 a_13467_32519# EN_VIN_BSTR_N 0.031982f
C45553 a_4190_30871# C9_P_btm 0.002182f
C45554 a_14127_45572# a_3483_46348# 1.22e-19
C45555 a_13076_44458# a_12891_46348# 0.182315f
C45556 a_9482_43914# a_3090_45724# 0.029795f
C45557 a_n2433_44484# a_n2293_46634# 7.85e-20
C45558 a_12607_44458# a_768_44030# 0.215512f
C45559 a_12883_44458# a_12549_44172# 7.5e-19
C45560 a_n4318_40392# a_n2312_38680# 0.023897f
C45561 a_20528_45572# a_12741_44636# 0.006514f
C45562 a_6298_44484# a_5807_45002# 1.01e-19
C45563 a_21350_45938# a_20202_43084# 1.43e-19
C45564 a_19610_45572# a_11415_45002# 5.19e-19
C45565 a_2711_45572# a_10586_45546# 0.295169f
C45566 a_7227_45028# a_8034_45724# 2.26e-19
C45567 a_7499_43078# a_526_44458# 0.2203f
C45568 a_6472_45840# a_8049_45260# 4.08e-19
C45569 a_5024_45822# a_5066_45546# 3.47e-19
C45570 a_413_45260# a_16721_46634# 6.74e-22
C45571 a_13904_45546# a_10809_44734# 9.68e-22
C45572 a_8696_44636# a_8016_46348# 0.031525f
C45573 a_11778_45572# a_10903_43370# 3.1e-20
C45574 a_15433_44458# a_11599_46634# 1.57e-21
C45575 a_14635_42282# a_1606_42308# 1.94e-20
C45576 a_n3674_39304# a_n3690_39616# 4.64e-19
C45577 a_5342_30871# a_13657_42308# 1.2e-20
C45578 a_5193_42852# a_5932_42308# 8.62e-21
C45579 a_n1151_42308# a_14084_46812# 0.063788f
C45580 a_2905_45572# a_3090_45724# 0.006554f
C45581 a_n237_47217# a_10425_46660# 2.5e-20
C45582 a_4883_46098# a_5907_46634# 5.32e-21
C45583 a_11599_46634# a_10623_46897# 3.51e-20
C45584 a_4915_47217# a_11735_46660# 3.49e-19
C45585 a_13487_47204# a_6755_46942# 1.18e-19
C45586 a_6151_47436# a_8846_46660# 0.002879f
C45587 a_2747_46873# a_3067_47026# 4.09e-19
C45588 a_n1613_43370# a_479_46660# 1.79e-19
C45589 a_9804_47204# a_2107_46812# 0.033493f
C45590 a_20843_47204# a_20916_46384# 8.16e-20
C45591 a_3232_43370# a_8685_43396# 8.91e-20
C45592 a_3537_45260# a_9803_43646# 2.53e-19
C45593 a_n2017_45002# a_15781_43660# 2.42e-20
C45594 a_11823_42460# a_5342_30871# 0.044603f
C45595 a_n2293_42834# a_n447_43370# 0.006668f
C45596 a_n2661_43370# a_n2840_43370# 0.172532f
C45597 a_10193_42453# a_18249_42858# 0.038446f
C45598 a_13249_42308# a_13635_43156# 0.004017f
C45599 a_5891_43370# a_7542_44172# 0.002369f
C45600 a_n2661_42834# a_1467_44172# 0.028215f
C45601 a_n2661_43922# a_1115_44172# 0.004853f
C45602 a_17517_44484# a_22315_44484# 0.063928f
C45603 a_20362_44736# a_20679_44626# 0.102355f
C45604 a_11967_42832# a_19279_43940# 0.070262f
C45605 a_12883_44458# a_12429_44172# 8.45e-19
C45606 a_5093_45028# VDD 0.168437f
C45607 a_5934_30871# a_n1532_35090# 1.62e-19
C45608 a_6123_31319# EN_VIN_BSTR_P 0.052187f
C45609 CAL_N a_4185_45028# 0.002972f
C45610 a_8103_44636# a_3483_46348# 0.00166f
C45611 a_15037_44260# a_12549_44172# 4.91e-19
C45612 a_15415_45028# a_13259_45724# 1.67e-19
C45613 a_n2661_43370# a_n1925_42282# 0.027962f
C45614 a_3065_45002# a_n755_45592# 0.027852f
C45615 a_n143_45144# a_n23_45546# 0.004979f
C45616 a_n37_45144# a_n356_45724# 0.001109f
C45617 a_413_45260# a_3503_45724# 7.76e-19
C45618 a_11691_44458# a_14840_46494# 2.41e-21
C45619 a_19778_44110# a_20075_46420# 1.42e-20
C45620 a_4223_44672# a_5164_46348# 2.5e-21
C45621 a_4743_44484# a_4704_46090# 4.57e-21
C45622 a_11827_44484# a_17715_44484# 0.037803f
C45623 a_14401_32519# a_13507_46334# 0.001279f
C45624 a_15811_47375# VDD 0.979053f
C45625 a_4958_30871# a_18907_42674# 2.39e-20
C45626 a_5932_42308# comp_n 2.3e-19
C45627 a_17303_42282# a_18727_42674# 3.04e-19
C45628 a_17531_42308# a_18057_42282# 0.00822f
C45629 a_n2661_46634# a_4185_45028# 1.65e-19
C45630 a_n2293_46634# a_3147_46376# 1.96e-19
C45631 a_n743_46660# a_2202_46116# 0.012092f
C45632 a_601_46902# a_805_46414# 7.84e-19
C45633 a_n1925_46634# a_2521_46116# 8.92e-20
C45634 a_383_46660# a_472_46348# 8.96e-19
C45635 a_n2438_43548# a_1823_45246# 0.002972f
C45636 a_171_46873# a_1176_45822# 5.65e-20
C45637 a_6755_46942# a_14513_46634# 0.036712f
C45638 a_7411_46660# a_765_45546# 0.003093f
C45639 a_768_44030# a_10903_43370# 0.082359f
C45640 a_12891_46348# a_12594_46348# 0.088156f
C45641 a_5807_45002# a_5937_45572# 0.038681f
C45642 a_n881_46662# a_15682_46116# 7.66e-19
C45643 a_n2312_40392# a_n2956_38680# 0.052782f
C45644 a_n2312_39304# a_n2956_39304# 6.38528f
C45645 a_13487_47204# a_8049_45260# 1.12e-20
C45646 a_9313_45822# a_10586_45546# 6.08e-20
C45647 a_n2497_47436# a_n1099_45572# 0.004833f
C45648 SMPL_ON_P a_n2293_45546# 8.05e-20
C45649 a_10193_42453# a_21125_42558# 8.15e-20
C45650 a_644_44056# a_n97_42460# 1.26e-20
C45651 a_14815_43914# a_14205_43396# 1.84e-19
C45652 a_15682_43940# a_14021_43940# 5.96e-19
C45653 a_20935_43940# a_15493_43940# 0.037795f
C45654 a_175_44278# a_104_43370# 1.89e-21
C45655 a_n2661_42282# a_5745_43940# 9.04e-20
C45656 a_742_44458# a_n13_43084# 4.27e-21
C45657 a_n2293_42834# a_3445_43172# 7.71e-20
C45658 a_n2017_45002# a_n1329_42308# 0.018315f
C45659 a_n2956_37592# a_n2104_42282# 8.96e-21
C45660 a_20447_31679# a_n1630_35242# 1.81e-19
C45661 a_n2810_45028# a_n3674_38216# 0.023217f
C45662 en_comp a_n4318_38216# 0.064646f
C45663 a_n1549_44318# VDD 0.200608f
C45664 C1_P_btm VREF_GND 0.673422f
C45665 a_10193_42453# a_12016_45572# 0.001841f
C45666 a_10490_45724# a_11688_45572# 0.003828f
C45667 a_2711_45572# a_18175_45572# 1.3e-21
C45668 a_11322_45546# a_11136_45572# 0.044092f
C45669 C0_P_btm VREF 0.443926f
C45670 a_5025_43940# a_n2293_46098# 0.002209f
C45671 a_6031_43396# a_3090_45724# 0.00482f
C45672 a_2982_43646# a_19692_46634# 0.003269f
C45673 a_3681_42891# a_768_44030# 1.91e-20
C45674 a_n1853_43023# a_n2956_39768# 1.99e-21
C45675 a_2998_44172# a_n1925_42282# 0.02835f
C45676 a_3600_43914# a_526_44458# 9.66e-19
C45677 a_13483_43940# a_10903_43370# 1.22e-19
C45678 a_8952_43230# a_n1613_43370# 0.213002f
C45679 a_18817_42826# a_13507_46334# 0.001318f
C45680 a_8953_45002# CLK 0.310391f
C45681 a_13059_46348# VDD 0.955445f
C45682 a_20719_46660# a_10809_44734# 6.1e-19
C45683 a_20202_43084# a_21137_46414# 0.006423f
C45684 a_4185_45028# a_8199_44636# 1.24e-19
C45685 a_3483_46348# a_8953_45546# 0.133493f
C45686 a_12741_44636# a_19335_46494# 1.88e-20
C45687 a_11415_45002# a_20708_46348# 5.4e-21
C45688 a_6755_46942# a_n357_42282# 3.13e-20
C45689 a_5257_43370# a_n443_42852# 0.016836f
C45690 a_15368_46634# a_13259_45724# 0.0178f
C45691 a_2553_47502# DATA[1] 5.06e-21
C45692 a_16922_45042# a_19511_42282# 2.37e-20
C45693 a_6293_42852# a_6765_43638# 2.33e-20
C45694 a_2982_43646# a_3457_43396# 0.074308f
C45695 a_18494_42460# a_17531_42308# 1.14e-19
C45696 a_18184_42460# a_18057_42282# 0.19301f
C45697 a_n356_44636# a_2713_42308# 1.57e-19
C45698 a_n2661_42834# a_n2840_42282# 0.001339f
C45699 a_14021_43940# a_22223_43396# 0.028989f
C45700 a_6031_43396# a_6547_43396# 0.105995f
C45701 a_9028_43914# a_8037_42858# 1.46e-19
C45702 a_8333_44056# a_8605_42826# 6.56e-22
C45703 a_15095_43370# VDD 0.169652f
C45704 a_8162_45546# a_n2661_44458# 1.47e-20
C45705 a_14495_45572# a_11827_44484# 1.5e-20
C45706 a_6511_45714# a_6298_44484# 0.001903f
C45707 a_5907_45546# a_5883_43914# 1.52e-20
C45708 a_3775_45552# a_n699_43396# 2.51e-21
C45709 a_n143_45144# a_n37_45144# 0.13675f
C45710 a_n913_45002# a_3537_45260# 0.148413f
C45711 a_n467_45028# a_413_45260# 2.64e-19
C45712 a_15890_42674# a_12549_44172# 5.15e-21
C45713 a_11301_43218# a_3090_45724# 0.001286f
C45714 a_458_43396# a_n755_45592# 0.001112f
C45715 a_1209_43370# a_n357_42282# 1.52e-19
C45716 a_4235_43370# a_n863_45724# 1.09e-20
C45717 a_n2267_43396# a_n443_42852# 9.52e-20
C45718 a_3218_45724# VDD 0.133843f
C45719 a_6667_45809# a_n2661_46634# 5.79e-21
C45720 a_4099_45572# a_n1925_46634# 2.99e-20
C45721 a_2711_45572# a_n743_46660# 0.525746f
C45722 a_8746_45002# a_768_44030# 0.001081f
C45723 a_10490_45724# a_12549_44172# 0.00731f
C45724 a_11322_45546# a_12891_46348# 1.18e-20
C45725 a_11525_45546# a_11309_47204# 0.004008f
C45726 a_13904_45546# a_n881_46662# 9.09e-19
C45727 a_n2661_45010# SMPL_ON_P 0.006065f
C45728 a_n1059_45260# a_n2497_47436# 0.073215f
C45729 a_2437_43646# a_1239_47204# 4.55e-19
C45730 a_16680_45572# a_10227_46804# 2.11e-19
C45731 a_16223_45938# a_16327_47482# 0.016725f
C45732 a_18147_46436# a_18051_46116# 1.26e-19
C45733 a_15682_43940# a_15764_42576# 3.53e-20
C45734 a_n2129_43609# a_n3674_38216# 1.65e-20
C45735 a_n2267_43396# a_n2104_42282# 4.83e-20
C45736 a_16759_43396# a_16795_42852# 9.47e-19
C45737 a_16243_43396# a_17333_42852# 4.48e-19
C45738 a_n901_43156# a_n13_43084# 0.014329f
C45739 a_n1991_42858# a_n1736_43218# 0.064178f
C45740 a_4361_42308# a_4520_42826# 6.25e-20
C45741 a_743_42282# a_7765_42852# 8.69e-20
C45742 a_16137_43396# a_18249_42858# 0.021561f
C45743 a_n2433_43396# a_n1736_42282# 5.66e-21
C45744 a_n4318_39304# a_n4318_37592# 0.023243f
C45745 a_n1853_43023# a_n1545_43230# 0.004472f
C45746 a_n1423_42826# a_n4318_38680# 1.78e-20
C45747 a_n1641_43230# a_n3674_39304# 1.48e-21
C45748 a_10768_47026# CLK 0.005946f
C45749 a_11735_46660# DATA[5] 4.37e-19
C45750 a_15009_46634# RST_Z 8.66e-21
C45751 a_7754_39964# a_7754_39632# 0.296522f
C45752 a_14097_32519# VDD 0.284675f
C45753 a_20841_45814# a_20766_44850# 3.35e-20
C45754 a_20623_45572# a_20835_44721# 3.31e-20
C45755 a_21188_45572# a_20640_44752# 1.97e-20
C45756 a_21363_45546# a_20679_44626# 3.09e-22
C45757 a_327_44734# a_n2661_42834# 0.001646f
C45758 a_413_45260# a_n2661_43922# 0.031184f
C45759 a_7229_43940# a_7640_43914# 0.177622f
C45760 a_5205_44484# a_5891_43370# 7.79e-20
C45761 a_5111_44636# a_9313_44734# 6.57e-20
C45762 a_3232_43370# a_8783_44734# 0.001081f
C45763 a_18479_45785# a_20512_43084# 2.57e-19
C45764 a_n2661_43370# a_n4318_40392# 0.005935f
C45765 a_16922_45042# a_19113_45348# 0.002269f
C45766 a_16321_45348# a_16237_45028# 9.85e-19
C45767 a_10490_45724# a_12429_44172# 8.84e-22
C45768 a_11322_45546# a_11750_44172# 5.99e-21
C45769 a_19778_44110# a_20567_45036# 0.044967f
C45770 a_17719_45144# a_11827_44484# 2.79e-20
C45771 a_18184_42460# a_18494_42460# 1.31047f
C45772 a_13070_42354# a_4185_45028# 8.35e-20
C45773 COMP_P a_n1925_42282# 0.071512f
C45774 a_3059_42968# a_n357_42282# 7.39e-19
C45775 a_9803_42558# a_8199_44636# 0.036259f
C45776 a_8791_42308# a_8953_45546# 0.006945f
C45777 a_16680_45572# a_17339_46660# 2.93e-21
C45778 a_17668_45572# a_15227_44166# 2.59e-20
C45779 a_6709_45028# a_4646_46812# 0.031325f
C45780 a_5691_45260# a_5732_46660# 9.85e-21
C45781 a_413_45260# a_7927_46660# 1.45e-20
C45782 a_3232_43370# a_5907_46634# 1.41e-20
C45783 a_17023_45118# a_n881_46662# 2.61e-20
C45784 a_6511_45714# a_5937_45572# 9.66e-19
C45785 a_2711_45572# a_11189_46129# 0.011492f
C45786 a_6667_45809# a_8199_44636# 4.59e-21
C45787 a_5891_43370# a_n971_45724# 0.084717f
C45788 a_n1821_44484# a_n1151_42308# 1.76e-19
C45789 a_7640_43914# a_n237_47217# 4.56e-21
C45790 a_4880_45572# a_4419_46090# 0.032829f
C45791 a_20205_31679# a_21589_35634# 3.35e-20
C45792 a_20692_30879# a_19864_35138# 1.26e-20
C45793 a_16855_43396# a_4958_30871# 1.08e-19
C45794 a_15743_43084# a_19511_42282# 1.59e-20
C45795 a_5649_42852# a_15803_42450# 2.29e-19
C45796 a_n2293_42282# a_n2840_42282# 2.81e-19
C45797 a_12465_44636# a_12891_46348# 0.033919f
C45798 a_2747_46873# a_3094_47243# 9.52e-20
C45799 a_4883_46098# a_768_44030# 0.045313f
C45800 a_10227_46804# a_13747_46662# 0.16398f
C45801 a_18479_47436# a_5807_45002# 2.73e-19
C45802 a_18143_47464# a_13661_43548# 0.011802f
C45803 a_16327_47482# a_16750_47204# 3.03e-19
C45804 a_6545_47178# a_2107_46812# 0.028617f
C45805 a_9313_45822# a_n743_46660# 0.029372f
C45806 a_12861_44030# a_n2293_46634# 6.64e-19
C45807 a_n971_45724# a_4817_46660# 1.65e-19
C45808 a_n237_47217# a_4651_46660# 7.27e-20
C45809 a_n1741_47186# a_6540_46812# 7e-21
C45810 a_3160_47472# a_2959_46660# 0.00952f
C45811 a_3381_47502# a_2609_46660# 0.00165f
C45812 a_n1151_42308# a_3177_46902# 0.006126f
C45813 a_n2109_47186# a_5275_47026# 0.001536f
C45814 a_584_46384# a_1057_46660# 6.68e-21
C45815 a_2905_45572# a_3699_46634# 0.00292f
C45816 a_742_44458# a_644_44056# 7.77e-19
C45817 a_18287_44626# a_18579_44172# 0.107662f
C45818 a_11823_42460# a_743_42282# 0.147603f
C45819 a_10193_42453# a_5649_42852# 0.003188f
C45820 a_9482_43914# a_9165_43940# 0.002619f
C45821 a_18989_43940# a_19279_43940# 0.053948f
C45822 a_1307_43914# a_3992_43940# 0.005165f
C45823 a_n1059_45260# a_1568_43370# 0.011697f
C45824 a_3357_43084# a_2982_43646# 0.01988f
C45825 a_n967_45348# a_n1821_43396# 3.3e-19
C45826 a_n659_45366# VDD 2.89e-19
C45827 a_14097_32519# a_22469_39537# 1.25e-20
C45828 a_n2661_43370# a_2698_46116# 1.36e-20
C45829 a_18494_42460# a_12741_44636# 0.114105f
C45830 a_21101_45002# a_11415_45002# 0.018873f
C45831 a_21359_45002# a_20202_43084# 0.008822f
C45832 a_7735_45067# a_3483_46348# 2.41e-19
C45833 a_17970_44736# a_15227_44166# 0.002254f
C45834 a_5663_43940# a_768_44030# 0.011502f
C45835 a_7640_43914# a_8270_45546# 2.57e-20
C45836 a_4558_45348# a_526_44458# 7.28e-20
C45837 a_4574_45260# a_n1925_42282# 3.52e-19
C45838 a_1307_43914# a_15682_46116# 0.001505f
C45839 a_10951_45334# a_10809_44734# 0.015679f
C45840 a_n1441_43940# a_n1613_43370# 0.012196f
C45841 a_11341_43940# a_16327_47482# 0.063063f
C45842 a_10533_42308# a_11323_42473# 0.002638f
C45843 a_1576_42282# a_7174_31319# 9.76e-21
C45844 a_n4318_37592# a_n4334_40480# 7.27e-20
C45845 COMP_P a_n4315_30879# 3.39e-19
C45846 a_n3674_38680# a_n4334_39616# 1.39e-19
C45847 a_5534_30871# C0_N_btm 8.49e-20
C45848 a_5342_30871# C0_dummy_P_btm 1.91e-20
C45849 a_19864_35138# VIN_N 0.367112f
C45850 RST_Z SINGLE_ENDED 0.0318f
C45851 EN_VIN_BSTR_N VCM 0.927905f
C45852 a_9313_45822# a_11189_46129# 1.48e-22
C45853 a_n1435_47204# a_9823_46155# 4.27e-21
C45854 a_4915_47217# a_2324_44458# 0.022906f
C45855 a_n2497_47436# a_n1925_42282# 0.004955f
C45856 a_n971_45724# a_n722_46482# 1.89e-19
C45857 a_n2312_39304# a_n1991_46122# 0.00213f
C45858 a_5807_45002# a_17829_46910# 3.44e-20
C45859 a_2443_46660# a_3090_45724# 2.52e-20
C45860 a_8667_46634# a_8492_46660# 0.233657f
C45861 a_13661_43548# a_765_45546# 1.39e-19
C45862 a_13747_46662# a_17339_46660# 0.015626f
C45863 a_3357_43084# a_5837_42852# 2.16e-20
C45864 a_n2661_42834# a_n1809_43762# 0.003072f
C45865 a_20512_43084# a_14021_43940# 0.030282f
C45866 a_1307_43914# a_9127_43156# 5.14e-20
C45867 a_n2293_42834# a_n1641_43230# 0.014975f
C45868 a_16922_45042# a_21259_43561# 0.108631f
C45869 a_17517_44484# a_19319_43548# 3.23e-20
C45870 a_11691_44458# a_18783_43370# 7.32e-20
C45871 a_n356_44636# a_6031_43396# 1.37e-20
C45872 a_n2293_43922# a_104_43370# 1.18e-21
C45873 a_9482_43914# a_12379_42858# 3.35e-19
C45874 a_8975_43940# a_8685_43396# 2.13e-20
C45875 a_5883_43914# a_9145_43396# 0.004333f
C45876 a_11649_44734# VDD 0.003396f
C45877 a_n4209_38216# C5_P_btm 1.11e-20
C45878 a_n3565_38216# C7_P_btm 1.43e-20
C45879 a_2711_45572# a_10053_45546# 0.018932f
C45880 a_6472_45840# a_6812_45938# 0.027606f
C45881 a_5013_44260# a_1823_45246# 0.001797f
C45882 a_9803_43646# a_n2293_46634# 0.01299f
C45883 a_16547_43609# a_12549_44172# 4.68e-19
C45884 a_6671_43940# a_3090_45724# 0.00493f
C45885 a_n699_43396# a_3218_45724# 1.28e-20
C45886 a_20159_44458# a_20075_46420# 1.46e-19
C45887 a_22223_43396# a_13507_46334# 0.006729f
C45888 a_20749_43396# a_18597_46090# 0.005121f
C45889 a_19963_31679# a_18194_35068# 1.2e-19
C45890 a_19479_31679# a_21589_35634# 7.02e-21
C45891 a_7577_46660# VDD 0.249866f
C45892 a_n4064_38528# a_n4251_38528# 0.001077f
C45893 a_n3420_38528# a_n4209_38216# 0.050044f
C45894 a_n3565_38502# a_n3565_38216# 0.0433f
C45895 a_7174_31319# C1_P_btm 5.34e-20
C45896 a_n784_42308# a_8530_39574# 1.98e-19
C45897 a_n4318_37592# a_n2946_37690# 3.13e-20
C45898 a_12741_44636# a_22959_46660# 0.17409f
C45899 a_20820_30879# a_21076_30879# 8.6867f
C45900 a_765_45546# a_4185_45028# 7.51e-20
C45901 a_n2661_46634# a_997_45618# 3.38e-22
C45902 a_n2293_46634# a_310_45028# 0.020873f
C45903 a_n2438_43548# a_n2293_45546# 0.051617f
C45904 a_n1021_46688# a_n863_45724# 5e-21
C45905 a_33_46660# a_n2661_45546# 4.08e-20
C45906 a_5807_45002# a_n443_42852# 1.54e-19
C45907 a_7715_46873# a_8034_45724# 9.01e-19
C45908 a_n743_46660# a_n1079_45724# 1.23e-19
C45909 a_3090_45724# a_18819_46122# 2.43e-19
C45910 a_12359_47026# a_12594_46348# 1.26e-19
C45911 a_11901_46660# a_6945_45028# 1.36e-19
C45912 a_11735_46660# a_10809_44734# 0.030929f
C45913 a_n97_42460# a_104_43370# 0.027998f
C45914 a_15493_43940# a_14955_43396# 0.013181f
C45915 a_11967_42832# a_12545_42858# 0.028062f
C45916 a_n1917_43396# a_n1821_43396# 0.013793f
C45917 a_n1699_43638# a_n1655_43396# 3.69e-19
C45918 a_14539_43914# a_16877_43172# 9.62e-19
C45919 a_11341_43940# a_10341_43396# 0.289072f
C45920 en_comp a_1239_39587# 0.003125f
C45921 a_n1177_43370# VDD 0.354704f
C45922 a_11778_45572# a_3232_43370# 1.29e-19
C45923 a_20623_45572# a_20731_45938# 0.057222f
C45924 a_11682_45822# a_11787_45002# 4.49e-20
C45925 a_5263_45724# a_n2661_43370# 8.75e-19
C45926 a_10796_42968# a_3090_45724# 0.004117f
C45927 a_14097_32519# a_22612_30879# 0.059759f
C45928 a_1756_43548# a_526_44458# 0.01292f
C45929 a_1568_43370# a_n1925_42282# 1.62e-21
C45930 a_6452_43396# a_2324_44458# 1.62e-20
C45931 a_10053_45546# a_9313_45822# 4.44e-20
C45932 a_11823_42460# a_6151_47436# 4.56e-21
C45933 a_10907_45822# a_2063_45854# 0.22153f
C45934 a_19335_46494# a_16375_45002# 4.62e-20
C45935 a_18985_46122# a_19431_46494# 2.28e-19
C45936 a_17957_46116# a_18051_46116# 0.062574f
C45937 a_8953_45546# a_n357_42282# 0.054106f
C45938 a_8791_43396# a_8952_43230# 6.83e-19
C45939 a_9396_43370# a_9127_43156# 0.00282f
C45940 a_16409_43396# a_4361_42308# 2.27e-20
C45941 a_18783_43370# a_4190_30871# 0.044615f
C45942 a_15743_43084# a_21259_43561# 6.3e-20
C45943 a_2982_43646# a_5342_30871# 0.178973f
C45944 a_16137_43396# a_5649_42852# 5.5e-20
C45945 a_19268_43646# a_19177_43646# 0.001446f
C45946 a_3626_43646# a_5534_30871# 0.082646f
C45947 a_n2661_46098# DATA[0] 4.59e-20
C45948 a_1799_45572# DATA[1] 0.004719f
C45949 a_22959_42860# VDD 0.30747f
C45950 en_comp a_11206_38545# 0.002407f
C45951 a_16751_45260# a_16922_45042# 0.12103f
C45952 a_11963_45334# a_11827_44484# 3.47e-20
C45953 a_2711_45572# a_5244_44056# 3.02e-22
C45954 a_1307_43914# a_17023_45118# 9.26e-21
C45955 a_8696_44636# a_14112_44734# 8.58e-19
C45956 a_5837_45348# a_n2661_43370# 4.55e-19
C45957 a_3537_45260# a_n2661_44458# 0.056342f
C45958 a_327_44734# a_n1352_44484# 5.64e-20
C45959 a_n1059_45260# a_5883_43914# 1.35e-19
C45960 a_n784_42308# a_1138_42852# 3.74e-20
C45961 a_791_42968# a_n863_45724# 0.338631f
C45962 a_3935_42891# a_n2661_45546# 1.6e-19
C45963 a_12545_42858# a_13259_45724# 3.09e-19
C45964 a_5193_43172# a_526_44458# 3.3e-19
C45965 a_15143_45578# a_15368_46634# 0.105334f
C45966 a_11682_45822# a_11813_46116# 2.39e-19
C45967 a_15765_45572# a_6755_46942# 0.026052f
C45968 a_6171_45002# a_12549_44172# 0.029809f
C45969 a_n2661_45010# a_n2438_43548# 0.220364f
C45970 a_413_45260# a_19594_46812# 4.71e-20
C45971 a_n913_45002# a_n2293_46634# 0.024406f
C45972 a_3232_43370# a_768_44030# 0.224083f
C45973 a_n2017_45002# a_n2312_38680# 8.38e-22
C45974 a_3357_43084# a_2107_46812# 0.033995f
C45975 en_comp a_n2956_39768# 0.003442f
C45976 a_22780_40945# VDD 1.38e-19
C45977 a_n2157_42858# a_n4318_38216# 0.001336f
C45978 a_10341_42308# a_11554_42852# 0.170124f
C45979 a_743_42282# a_961_42354# 0.016854f
C45980 a_3626_43646# a_19647_42308# 0.170024f
C45981 a_2982_43646# a_20107_42308# 0.003276f
C45982 a_10922_42852# a_10752_42852# 2.6e-19
C45983 a_5649_42852# a_n784_42308# 0.043382f
C45984 a_n1991_42858# a_n3674_38680# 1.73e-20
C45985 a_19553_46090# START 1.2e-21
C45986 a_15015_46420# CLK 7.59e-21
C45987 a_19335_46494# RST_Z 1.49e-21
C45988 a_n4334_39616# VDD 0.385881f
C45989 a_3422_30871# a_n3420_37984# 0.031681f
C45990 a_1431_47204# a_n881_46662# 3.11e-20
C45991 a_2124_47436# a_n1613_43370# 2.83e-20
C45992 a_9067_47204# a_4883_46098# 1.74e-20
C45993 a_11599_46634# a_10227_46804# 0.60865f
C45994 a_16241_47178# a_16023_47582# 0.209641f
C45995 a_15507_47210# a_17591_47464# 1.96e-21
C45996 a_15673_47210# a_16763_47508# 0.042509f
C45997 a_n1151_42308# a_3315_47570# 0.003697f
C45998 a_4007_47204# a_2747_46873# 3.71e-20
C45999 a_12861_44030# a_18597_46090# 0.045766f
C46000 a_13717_47436# a_19386_47436# 8e-20
C46001 a_21101_45002# a_11967_42832# 1.52e-19
C46002 a_n1809_44850# a_n356_44636# 5.9e-21
C46003 a_2779_44458# a_n2661_43922# 0.013114f
C46004 a_4223_44672# a_n2661_42834# 0.031905f
C46005 a_5518_44484# a_5708_44484# 0.045837f
C46006 a_10334_44484# a_9313_44734# 0.018652f
C46007 a_18494_42460# a_20362_44736# 0.004144f
C46008 a_20567_45036# a_20159_44458# 0.001074f
C46009 a_19778_44110# a_20679_44626# 5.45e-21
C46010 a_n2293_42834# a_n809_44244# 0.001759f
C46011 a_10193_42453# a_8685_43396# 0.024858f
C46012 a_n2661_44458# a_11541_44484# 0.053139f
C46013 a_7499_43078# a_8317_43396# 3.9e-19
C46014 a_5105_45348# a_3905_42865# 3.58e-20
C46015 a_19256_45572# a_19319_43548# 8.54e-21
C46016 a_11691_44458# a_16335_44484# 2.35e-19
C46017 a_11827_44484# a_18588_44850# 4.54e-19
C46018 a_6171_45002# a_12429_44172# 1.87e-21
C46019 a_9223_42460# a_n443_42852# 1.18e-20
C46020 a_14456_42282# a_n357_42282# 7.69e-20
C46021 a_19332_42282# a_13259_45724# 1.03e-19
C46022 a_8696_44636# VDD 1.12228f
C46023 a_21076_30879# C8_N_btm 0.384801f
C46024 a_5534_30871# C10_P_btm 1.08e-19
C46025 a_14797_45144# a_11415_45002# 0.021281f
C46026 a_13777_45326# a_12741_44636# 4.48e-20
C46027 a_5518_44484# a_5257_43370# 0.095452f
C46028 a_3429_45260# a_3147_46376# 1.69e-19
C46029 a_3065_45002# a_3483_46348# 0.001025f
C46030 a_18911_45144# a_3090_45724# 0.190188f
C46031 a_15433_44458# a_13661_43548# 0.038412f
C46032 a_14673_44172# a_12549_44172# 0.024138f
C46033 a_2382_45260# a_4185_45028# 0.008734f
C46034 a_15765_45572# a_8049_45260# 0.012841f
C46035 a_3260_45572# a_3316_45546# 4.85e-19
C46036 a_20273_45572# a_20708_46348# 4.47e-20
C46037 a_20107_45572# a_21137_46414# 0.002164f
C46038 a_2437_43646# a_14840_46494# 1.19e-36
C46039 a_20512_43084# a_13507_46334# 0.497215f
C46040 a_196_42282# a_5934_30871# 3.42e-20
C46041 a_2713_42308# a_3823_42558# 6.62e-20
C46042 a_2903_42308# a_3318_42354# 0.003549f
C46043 a_1606_42308# a_4921_42308# 4.1e-20
C46044 a_n784_42308# a_7963_42308# 1.56e-20
C46045 a_1576_42282# a_5932_42308# 8.68e-21
C46046 a_4190_30871# C0_N_btm 6.53e-20
C46047 a_22521_40055# a_22821_38993# 0.131339f
C46048 a_22459_39145# a_22545_38993# 0.121283f
C46049 a_22780_40081# a_22521_39511# 1.39e-19
C46050 a_n2661_46634# a_5257_43370# 0.005264f
C46051 a_5807_45002# a_10554_47026# 0.003779f
C46052 a_2107_46812# a_3877_44458# 0.070722f
C46053 a_n743_46660# a_6540_46812# 7.69e-21
C46054 a_2443_46660# a_3699_46634# 0.043475f
C46055 a_2609_46660# a_2959_46660# 0.216095f
C46056 a_1799_45572# a_2864_46660# 3.88e-20
C46057 a_n881_46662# a_11735_46660# 1.34e-19
C46058 a_11453_44696# a_19692_46634# 0.05834f
C46059 a_11599_46634# a_17339_46660# 0.131185f
C46060 a_14955_47212# a_765_45546# 0.004861f
C46061 a_16763_47508# a_16388_46812# 5.51e-19
C46062 a_10227_46804# a_13693_46688# 0.002261f
C46063 a_16327_47482# a_16434_46987# 0.00105f
C46064 a_12861_44030# a_19123_46287# 0.002675f
C46065 a_n2497_47436# a_2698_46116# 1.45e-22
C46066 a_n2109_47186# a_167_45260# 4.41e-20
C46067 a_n1741_47186# a_1823_45246# 8.12e-20
C46068 a_n971_45724# a_472_46348# 5.63e-20
C46069 a_n746_45260# a_376_46348# 0.010981f
C46070 a_949_44458# a_n97_42460# 1.25e-19
C46071 a_n699_43396# a_n1177_43370# 0.060973f
C46072 a_742_44458# a_104_43370# 5.46e-21
C46073 a_n1899_43946# a_453_43940# 7e-20
C46074 a_n2293_43922# a_11341_43940# 0.026007f
C46075 a_13249_42308# a_13814_43218# 1.82e-19
C46076 a_n2293_45010# a_791_42968# 3.6e-20
C46077 a_n913_45002# a_n1533_42852# 4.76e-20
C46078 a_n967_45348# a_n1736_43218# 0.001166f
C46079 a_n3607_37440# VDD 2.79e-20
C46080 a_n1177_44458# VDD 0.347966f
C46081 a_18057_42282# RST_Z 1.94e-20
C46082 a_19279_43940# a_20202_43084# 0.020761f
C46083 a_20766_44850# a_11415_45002# 0.001727f
C46084 a_4905_42826# a_768_44030# 4.03e-20
C46085 a_4223_44672# a_5066_45546# 2.22e-20
C46086 a_n2661_43370# a_380_45546# 4.07e-20
C46087 a_9838_44484# a_526_44458# 1.68e-22
C46088 a_117_45144# a_n443_42852# 6.39e-19
C46089 a_9313_44734# a_9290_44172# 0.140741f
C46090 a_n998_43396# a_n1613_43370# 0.001965f
C46091 a_14537_43646# a_12861_44030# 1.95e-20
C46092 a_14358_43442# a_10227_46804# 0.019948f
C46093 a_10341_43396# a_16327_47482# 0.159266f
C46094 a_n3420_39616# a_n2946_39866# 0.236674f
C46095 a_n3690_39616# a_n4064_39616# 0.085414f
C46096 a_n3565_39590# a_n2302_39866# 0.044102f
C46097 a_7174_31319# a_1736_39043# 7.24e-20
C46098 a_n4209_39590# a_n2216_39866# 0.001361f
C46099 a_n4315_30879# a_n4209_39304# 0.032541f
C46100 a_n4064_40160# a_n3607_39616# 5.58e-20
C46101 a_5932_42308# C1_P_btm 0.011049f
C46102 a_7577_46660# a_7920_46348# 5.66e-19
C46103 a_7411_46660# a_8349_46414# 0.001959f
C46104 a_7715_46873# a_8016_46348# 0.009008f
C46105 a_5807_45002# a_6633_46155# 1.37e-19
C46106 a_n743_46660# a_1337_46436# 0.004605f
C46107 a_171_46873# a_518_46482# 9.21e-19
C46108 a_15227_44166# a_19636_46660# 6.47e-19
C46109 a_19692_46634# a_17639_46660# 2.07e-22
C46110 a_15227_46910# a_15312_46660# 1.48e-19
C46111 a_10249_46116# a_3483_46348# 1.46e-20
C46112 a_14976_45028# a_11415_45002# 0.039578f
C46113 a_18579_44172# a_19268_43646# 6.28e-19
C46114 a_n2661_42834# a_n3674_39304# 0.038671f
C46115 a_11341_43940# a_n97_42460# 1.85e-19
C46116 a_1307_43914# a_1755_42282# 1.63e-19
C46117 a_n2293_43922# a_n1076_43230# 1.7e-20
C46118 a_n356_44636# a_10796_42968# 4.72e-20
C46119 a_14539_43914# a_5342_30871# 2.82e-20
C46120 a_14021_43940# a_21381_43940# 0.022437f
C46121 a_5111_44636# a_8515_42308# 5.49e-21
C46122 en_comp a_12563_42308# 8.68e-21
C46123 a_n2017_45002# a_13657_42558# 0.0086f
C46124 a_3537_45260# a_8325_42308# 3.11e-21
C46125 a_20365_43914# VDD 0.261299f
C46126 a_15599_45572# a_16211_45572# 3.82e-19
C46127 a_2711_45572# a_5111_44636# 0.00298f
C46128 a_n3420_37984# VREF_GND 0.047887f
C46129 a_4699_43561# a_1823_45246# 0.003517f
C46130 a_7227_42852# a_4646_46812# 0.032378f
C46131 a_n2065_43946# a_n443_42852# 5.59e-21
C46132 a_1414_42308# a_2957_45546# 9.39e-21
C46133 a_2479_44172# a_n755_45592# 1.32e-20
C46134 a_3905_42865# a_n863_45724# 1.11e-19
C46135 a_895_43940# a_n357_42282# 0.008143f
C46136 a_8495_42852# a_n1613_43370# 0.012196f
C46137 a_20356_42852# a_16327_47482# 7.6e-21
C46138 a_1755_42282# a_n443_46116# 3.6e-20
C46139 a_n4209_37414# a_n1386_35608# 6.24e-22
C46140 a_18494_42460# RST_Z 5.9e-20
C46141 a_4704_46090# VDD 0.225404f
C46142 a_n4209_39590# VDAC_P 0.006893f
C46143 a_765_45546# a_997_45618# 0.026457f
C46144 a_6419_46155# a_5066_45546# 0.038923f
C46145 a_5164_46348# a_5527_46155# 0.005527f
C46146 a_5204_45822# a_5210_46155# 8.95e-19
C46147 a_18819_46122# a_20075_46420# 0.043567f
C46148 a_18985_46122# a_19335_46494# 0.210876f
C46149 a_17583_46090# a_6945_45028# 6.47e-21
C46150 a_2324_44458# a_10809_44734# 0.026995f
C46151 a_n3565_39304# a_n3565_37414# 0.029571f
C46152 a_n4209_39304# a_n3420_37440# 0.033347f
C46153 a_n3420_39072# a_n4209_37414# 0.030579f
C46154 a_n3565_38216# a_n2860_37984# 0.001043f
C46155 C9_N_btm C10_N_btm 53.3168f
C46156 a_n2065_43946# a_n2104_42282# 2.12e-21
C46157 a_8685_43396# a_16137_43396# 0.003201f
C46158 a_2982_43646# a_743_42282# 0.047135f
C46159 a_n97_42460# a_n1076_43230# 4.69e-19
C46160 a_14021_43940# a_18249_42858# 4.16e-20
C46161 a_n2293_43922# a_10723_42308# 8.6e-20
C46162 a_9313_44734# a_15051_42282# 2.49e-19
C46163 a_n356_44636# a_4958_30871# 0.46356f
C46164 a_3626_43646# a_4190_30871# 0.070713f
C46165 a_9145_43396# a_14621_43646# 0.00367f
C46166 a_n310_47243# DATA[0] 0.002781f
C46167 a_2747_46873# DATA[1] 3.15e-21
C46168 a_21588_30879# a_22521_40055# 3.72e-20
C46169 a_n1991_42858# VDD 0.575656f
C46170 a_9482_43914# a_14180_45002# 0.022677f
C46171 a_13556_45296# a_13777_45326# 0.101558f
C46172 a_10951_45334# a_1307_43914# 3.62e-21
C46173 a_9049_44484# a_9313_44734# 0.034936f
C46174 a_13017_45260# a_15415_45028# 5.39e-21
C46175 a_13348_45260# a_14537_43396# 3.8e-20
C46176 a_n2017_45002# a_n2661_43370# 0.038361f
C46177 a_7229_43940# a_1423_45028# 0.024468f
C46178 a_20623_45572# a_20567_45036# 0.001339f
C46179 a_20841_45814# a_21005_45260# 3.92e-20
C46180 a_2382_45260# a_2448_45028# 0.009378f
C46181 a_4558_45348# a_5365_45348# 7.9e-20
C46182 a_5147_45002# a_5105_45348# 2.26e-21
C46183 a_20273_45572# a_21101_45002# 0.014321f
C46184 a_n4064_40160# a_n2442_46660# 0.006941f
C46185 a_13667_43396# a_n443_42852# 0.035517f
C46186 a_421_43172# a_526_44458# 3.36e-20
C46187 a_9159_45572# a_2107_46812# 6.31e-20
C46188 a_3357_43084# a_11453_44696# 0.020072f
C46189 a_413_45260# a_15673_47210# 2.52e-19
C46190 en_comp a_10227_46804# 2.31e-20
C46191 a_n913_45002# a_18597_46090# 0.126328f
C46192 a_6709_45028# a_6545_47178# 1.46e-20
C46193 a_1423_45028# a_n237_47217# 5.23e-20
C46194 a_2304_45348# a_n971_45724# 0.00123f
C46195 a_n863_45724# a_n89_45572# 8.15e-19
C46196 a_n452_45724# a_n310_45572# 0.007833f
C46197 a_n755_45592# a_n443_42852# 0.469263f
C46198 a_16137_43396# a_15953_42852# 2.65e-19
C46199 a_10991_42826# a_10341_42308# 0.035667f
C46200 a_10835_43094# a_12089_42308# 2.32e-19
C46201 a_10796_42968# a_12379_42858# 3.81e-19
C46202 a_3539_42460# a_4921_42308# 3.77e-19
C46203 a_2982_43646# a_5755_42308# 2.01e-19
C46204 a_n97_42460# a_10723_42308# 7.44e-19
C46205 a_22959_46660# RST_Z 0.001115f
C46206 a_4338_37500# a_6886_37412# 1.95816f
C46207 a_3726_37500# VDAC_N 0.06247f
C46208 a_5088_37509# a_5700_37509# 1.48771f
C46209 a_9377_42558# VDD 0.007808f
C46210 a_2952_47436# a_3785_47178# 6.47e-19
C46211 a_2063_45854# a_4007_47204# 3.64e-20
C46212 a_2905_45572# a_3381_47502# 0.208262f
C46213 a_3160_47472# a_n1151_42308# 0.357683f
C46214 a_n2497_47436# a_n1435_47204# 0.010029f
C46215 a_n1741_47186# a_11031_47542# 0.00728f
C46216 a_n237_47217# a_6491_46660# 0.002119f
C46217 a_n971_45724# a_7227_47204# 0.009537f
C46218 a_742_44458# a_949_44458# 0.185221f
C46219 a_16237_45028# a_14539_43914# 1.93e-19
C46220 a_n2661_44458# a_8701_44490# 0.00716f
C46221 a_11691_44458# a_17767_44458# 0.060949f
C46222 a_11827_44484# a_18443_44721# 0.007717f
C46223 a_16147_45260# a_17737_43940# 8.05e-21
C46224 a_n2293_42834# a_n2661_42834# 0.202366f
C46225 a_15861_45028# a_15493_43940# 4.14e-20
C46226 a_n913_45002# a_2675_43914# 2.72e-20
C46227 a_n1059_45260# a_2889_44172# 4.48e-22
C46228 a_n2017_45002# a_2998_44172# 2.57e-20
C46229 a_7227_45028# VDD 0.501104f
C46230 a_13467_32519# a_11530_34132# 0.002259f
C46231 a_4190_30871# C10_P_btm 0.446355f
C46232 a_14033_45572# a_3483_46348# 0.003201f
C46233 a_12607_44458# a_12549_44172# 0.033279f
C46234 a_12883_44458# a_12891_46348# 0.018059f
C46235 a_8560_45348# a_7411_46660# 2.42e-21
C46236 a_5518_44484# a_5807_45002# 7.14e-20
C46237 a_13777_45326# a_13607_46688# 2.78e-21
C46238 a_1423_45028# a_8270_45546# 0.023554f
C46239 a_8975_43940# a_768_44030# 0.124155f
C46240 a_n2661_44458# a_n2293_46634# 0.029279f
C46241 a_19365_45572# a_11415_45002# 1.55e-19
C46242 a_6194_45824# a_8049_45260# 4.11e-20
C46243 a_413_45260# a_16388_46812# 4.56e-20
C46244 a_13527_45546# a_10809_44734# 3.56e-21
C46245 a_11688_45572# a_10903_43370# 2.55e-20
C46246 a_10617_44484# a_10227_46804# 0.006757f
C46247 a_5837_42852# a_5755_42308# 4.85e-19
C46248 a_13291_42460# a_1606_42308# 1.35e-20
C46249 a_n4318_38680# a_n4334_39616# 1.78e-19
C46250 a_17701_42308# a_15890_42674# 2.84e-21
C46251 a_7573_43172# a_6123_31319# 2.33e-20
C46252 a_5534_30871# a_13921_42308# 5.65e-20
C46253 a_12861_44030# a_6755_46942# 0.376009f
C46254 a_6151_47436# a_8601_46660# 6.03e-19
C46255 a_2952_47436# a_3090_45724# 8.88e-21
C46256 a_n1151_42308# a_13607_46688# 0.005534f
C46257 a_n237_47217# a_10185_46660# 7.66e-20
C46258 a_n1741_47186# a_12347_46660# 2.12e-19
C46259 a_4883_46098# a_5167_46660# 1.64e-20
C46260 a_11599_46634# a_10467_46802# 0.261176f
C46261 a_10227_46804# a_7411_46660# 2.95e-22
C46262 a_2747_46873# a_2864_46660# 0.174836f
C46263 a_n1613_43370# a_1110_47026# 6.37e-19
C46264 a_n881_46662# a_n935_46688# 8.8e-19
C46265 a_8128_46384# a_2107_46812# 0.028382f
C46266 a_5807_45002# a_n2661_46634# 0.087532f
C46267 a_12607_44458# a_12429_44172# 4.52e-19
C46268 a_11967_42832# a_20766_44850# 0.042853f
C46269 a_20159_44458# a_20679_44626# 0.043567f
C46270 a_20362_44736# a_20640_44752# 0.118759f
C46271 a_17517_44484# a_3422_30871# 0.073987f
C46272 a_n2661_43922# a_644_44056# 1.23e-19
C46273 a_7640_43914# a_7845_44172# 0.021949f
C46274 a_n2661_42834# a_1115_44172# 0.011443f
C46275 a_5891_43370# a_7281_43914# 4.34e-19
C46276 a_n2293_42834# a_n1352_43396# 0.006475f
C46277 a_11823_42460# a_15279_43071# 0.010476f
C46278 a_10193_42453# a_17333_42852# 0.032471f
C46279 a_13249_42308# a_12895_43230# 0.002542f
C46280 a_18479_45785# a_5649_42852# 4.56e-21
C46281 a_3537_45260# a_9145_43396# 0.002981f
C46282 a_n2017_45002# a_15681_43442# 1.9e-21
C46283 a_5111_44636# a_7466_43396# 0.002133f
C46284 a_5009_45028# VDD 0.151712f
C46285 a_6123_31319# a_n923_35174# 0.008058f
C46286 a_6298_44484# a_3483_46348# 0.017162f
C46287 a_5343_44458# a_4185_45028# 5.81e-20
C46288 a_15682_43940# a_n743_46660# 0.001683f
C46289 a_15493_43940# a_19321_45002# 0.050579f
C46290 a_9672_43914# a_2107_46812# 0.079349f
C46291 a_14761_44260# a_12549_44172# 1.08e-19
C46292 a_14797_45144# a_13259_45724# 0.092924f
C46293 a_n2661_43370# a_526_44458# 0.054473f
C46294 a_n2293_42834# a_5066_45546# 3.17e-20
C46295 a_n143_45144# a_n356_45724# 3.1e-21
C46296 a_3065_45002# a_n357_42282# 0.023226f
C46297 a_413_45260# a_3316_45546# 0.110075f
C46298 a_2680_45002# a_n755_45592# 5.6e-20
C46299 a_n967_45348# a_n1013_45572# 2.46e-19
C46300 a_11827_44484# a_17583_46090# 6.39e-21
C46301 a_19778_44110# a_19335_46494# 4.32e-19
C46302 a_11691_44458# a_15015_46420# 4.75e-21
C46303 a_4223_44672# a_5068_46348# 1.13e-20
C46304 a_21381_43940# a_13507_46334# 5.15e-20
C46305 a_n97_42460# a_16327_47482# 0.113034f
C46306 a_4743_44484# a_4419_46090# 8.99e-21
C46307 a_15507_47210# VDD 0.441662f
C46308 a_17303_42282# a_18057_42282# 7.14e-19
C46309 a_5932_42308# a_1736_39043# 8.72e-20
C46310 a_4958_30871# a_18727_42674# 2.08e-20
C46311 a_5742_30871# a_n3565_39590# 7.02e-21
C46312 a_n2293_46634# a_2804_46116# 1.38e-20
C46313 a_n743_46660# a_1823_45246# 0.04372f
C46314 a_n1925_46634# a_167_45260# 3.51e-19
C46315 a_n2438_43548# a_1138_42852# 0.646257f
C46316 a_383_46660# a_376_46348# 3.44e-19
C46317 a_n133_46660# a_1176_45822# 3.41e-19
C46318 a_33_46660# a_805_46414# 0.001417f
C46319 a_5257_43370# a_765_45546# 0.002074f
C46320 a_6755_46942# a_14180_46812# 0.063843f
C46321 a_13607_46688# a_14084_46812# 0.014875f
C46322 a_5807_45002# a_8199_44636# 0.001797f
C46323 a_12549_44172# a_10903_43370# 0.792848f
C46324 a_12891_46348# a_12005_46116# 0.001509f
C46325 a_n881_46662# a_2324_44458# 0.085939f
C46326 a_n2312_40392# a_n2956_39304# 0.052343f
C46327 a_5342_30871# a_n4064_37984# 0.028465f
C46328 a_4915_47217# a_12839_46116# 2.59e-20
C46329 a_12861_44030# a_8049_45260# 0.109405f
C46330 a_n2497_47436# a_380_45546# 9.69e-22
C46331 a_n815_47178# a_n2661_45546# 4.98e-21
C46332 SMPL_ON_P a_n2956_38216# 0.0385f
C46333 a_14955_43940# a_14021_43940# 1.99e-20
C46334 a_20623_43914# a_15493_43940# 0.040969f
C46335 a_21115_43940# a_11341_43940# 0.008031f
C46336 a_14539_43914# a_743_42282# 3.58e-20
C46337 a_175_44278# a_n97_42460# 2.88e-20
C46338 a_n2293_42834# a_n2293_42282# 0.018879f
C46339 a_n2293_43922# a_10341_43396# 0.022718f
C46340 en_comp a_n2472_42282# 0.018838f
C46341 a_n2017_45002# COMP_P 0.012669f
C46342 a_n2810_45028# a_n2104_42282# 9.69e-21
C46343 a_n2956_37592# a_n4318_38216# 0.023067f
C46344 a_n1331_43914# VDD 0.203823f
C46345 a_2711_45572# a_16147_45260# 0.028186f
C46346 a_10193_42453# a_11778_45572# 0.004713f
C46347 a_10490_45724# a_11136_45572# 0.048799f
C46348 C0_dummy_P_btm VIN_P 0.544204f
C46349 C1_P_btm VREF 0.98698f
C46350 a_2905_42968# a_768_44030# 4.25e-19
C46351 a_n2157_42858# a_n2956_39768# 3.98e-21
C46352 a_3626_43646# a_15227_44166# 1.37e-19
C46353 a_2998_44172# a_526_44458# 0.028337f
C46354 a_12429_44172# a_10903_43370# 0.116356f
C46355 a_9127_43156# a_n1613_43370# 0.267842f
C46356 a_11136_42852# a_2063_45854# 2.55e-20
C46357 a_20922_43172# a_18597_46090# 0.021228f
C46358 a_18249_42858# a_13507_46334# 5.85e-19
C46359 a_15227_46910# VDD 0.229766f
C46360 a_7174_31319# a_n3420_37984# 7.78e-20
C46361 a_5742_30871# a_3726_37500# 0.001929f
C46362 a_5204_45822# a_5497_46414# 0.099282f
C46363 a_5164_46348# a_6165_46155# 3.3e-19
C46364 a_21350_47026# a_10809_44734# 1.68e-19
C46365 a_20202_43084# a_20708_46348# 0.001267f
C46366 a_3483_46348# a_5937_45572# 0.767636f
C46367 a_11415_45002# a_19900_46494# 1.14e-20
C46368 a_765_45546# a_1337_46116# 0.011452f
C46369 a_14180_46812# a_8049_45260# 1.24e-21
C46370 a_14976_45028# a_13259_45724# 0.018965f
C46371 a_8333_44056# a_8037_42858# 2.79e-21
C46372 a_6031_43396# a_6765_43638# 0.053479f
C46373 a_6293_42852# a_6197_43396# 0.213423f
C46374 a_14021_43940# a_5649_42852# 0.005268f
C46375 a_n97_42460# a_10341_43396# 0.917198f
C46376 a_18494_42460# a_17303_42282# 6.74e-19
C46377 a_18184_42460# a_17531_42308# 0.001442f
C46378 a_2982_43646# a_2813_43396# 0.096538f
C46379 a_11967_42832# a_13157_43218# 0.002086f
C46380 a_n1151_42308# RST_Z 0.004602f
C46381 a_2063_45854# DATA[1] 8.67e-20
C46382 a_14205_43396# VDD 0.311811f
C46383 a_13249_42308# a_11827_44484# 0.029876f
C46384 a_6472_45840# a_6298_44484# 0.002101f
C46385 a_n1059_45260# a_3537_45260# 0.162323f
C46386 a_n955_45028# a_413_45260# 1.19e-20
C46387 a_1847_42826# a_1823_45246# 1.28e-20
C46388 a_15959_42545# a_12549_44172# 2.73e-19
C46389 a_11229_43218# a_3090_45724# 7.17e-19
C46390 a_458_43396# a_n357_42282# 0.016095f
C46391 a_4093_43548# a_n863_45724# 9.16e-21
C46392 a_n1557_42282# a_n2810_45572# 1.35e-20
C46393 a_n229_43646# a_n755_45592# 0.049717f
C46394 a_n2129_43609# a_n443_42852# 1.4e-19
C46395 a_16823_43084# a_17715_44484# 4.72e-20
C46396 a_3422_30871# EN_VIN_BSTR_N 0.182769f
C46397 a_2957_45546# VDD 0.192471f
C46398 a_10193_42453# a_768_44030# 0.030504f
C46399 a_6511_45714# a_n2661_46634# 1.3e-20
C46400 a_6428_45938# a_5807_45002# 3.09e-19
C46401 a_1260_45572# a_n2438_43548# 0.001032f
C46402 a_11322_45546# a_11309_47204# 2.89e-19
C46403 a_13527_45546# a_n881_46662# 1.35e-19
C46404 a_n2017_45002# a_n2497_47436# 0.125552f
C46405 a_2437_43646# a_1209_47178# 0.025116f
C46406 a_n2840_45002# SMPL_ON_P 7.52e-19
C46407 a_16020_45572# a_16327_47482# 0.001041f
C46408 a_16375_45002# a_19240_46482# 3.8e-20
C46409 a_n2129_43609# a_n2104_42282# 1.48e-19
C46410 a_n2433_43396# a_n3674_38216# 8.11e-21
C46411 a_16977_43638# a_16795_42852# 7.5e-19
C46412 a_n901_43156# a_n1076_43230# 0.234322f
C46413 a_n1853_43023# a_n1736_43218# 0.183149f
C46414 a_743_42282# a_7871_42858# 9.63e-20
C46415 a_16137_43396# a_17333_42852# 0.01487f
C46416 a_3626_43646# a_14635_42282# 0.002593f
C46417 a_n1991_42858# a_n4318_38680# 5.47e-19
C46418 a_n2157_42858# a_n1545_43230# 3.82e-19
C46419 a_14084_46812# RST_Z 2.99e-19
C46420 a_22400_42852# VDD 0.829052f
C46421 a_11652_45724# a_10729_43914# 5.99e-20
C46422 a_20107_45572# a_19279_43940# 1.81e-19
C46423 a_17613_45144# a_11827_44484# 9.36e-21
C46424 a_19778_44110# a_18494_42460# 0.04586f
C46425 a_n2661_43370# a_n2840_44458# 0.011391f
C46426 a_5093_45028# a_4223_44672# 4.9e-19
C46427 a_10490_45724# a_11750_44172# 1.05e-21
C46428 a_10193_42453# a_13483_43940# 2.57e-19
C46429 a_8704_45028# a_n2661_44458# 1.59e-19
C46430 a_20841_45814# a_20835_44721# 0.001113f
C46431 a_20623_45572# a_20679_44626# 6.43e-21
C46432 a_21363_45546# a_20640_44752# 9.91e-23
C46433 a_n37_45144# a_n2661_43922# 4.45e-20
C46434 a_413_45260# a_n2661_42834# 0.023284f
C46435 a_20528_45572# a_20159_44458# 2.85e-20
C46436 a_7229_43940# a_6109_44484# 5.71e-20
C46437 a_3232_43370# a_8333_44734# 8.77e-20
C46438 a_7276_45260# a_7640_43914# 1.59e-19
C46439 a_12563_42308# a_4185_45028# 1.64e-19
C46440 a_n4318_37592# a_n1925_42282# 0.024213f
C46441 a_2987_42968# a_n357_42282# 4.17e-19
C46442 a_8685_42308# a_8953_45546# 0.250058f
C46443 a_9223_42460# a_8199_44636# 0.065156f
C46444 a_5437_45600# a_3483_46348# 9.84e-20
C46445 a_7229_43940# a_4646_46812# 0.104864f
C46446 a_413_45260# a_8145_46902# 2.46e-21
C46447 a_16922_45042# a_n881_46662# 4.59e-20
C46448 a_6511_45714# a_8199_44636# 1.7e-19
C46449 a_6472_45840# a_5937_45572# 0.001997f
C46450 a_2711_45572# a_9290_44172# 0.030631f
C46451 a_16237_45028# a_11453_44696# 0.008411f
C46452 a_8375_44464# a_n971_45724# 0.007671f
C46453 a_6109_44484# a_n237_47217# 4.56e-21
C46454 a_4808_45572# a_4419_46090# 0.004093f
C46455 a_5755_42852# a_5932_42308# 0.012644f
C46456 a_5649_42852# a_15764_42576# 1.57e-19
C46457 a_4361_42308# a_15890_42674# 0.004318f
C46458 a_20205_31679# a_19864_35138# 9.62e-21
C46459 a_16375_45002# START 1.03e-19
C46460 a_4883_46098# a_12549_44172# 0.021771f
C46461 a_10227_46804# a_13661_43548# 0.072131f
C46462 a_17591_47464# a_13747_46662# 1.16e-19
C46463 a_16241_47178# a_16750_47204# 2.6e-19
C46464 a_18143_47464# a_5807_45002# 1.77e-19
C46465 a_6151_47436# a_2107_46812# 0.019997f
C46466 a_n971_45724# a_4955_46873# 4.2e-20
C46467 a_n237_47217# a_4646_46812# 0.020773f
C46468 a_n1151_42308# a_2609_46660# 3.74e-19
C46469 a_3381_47502# a_2443_46660# 8.51e-19
C46470 a_2905_45572# a_2959_46660# 0.005466f
C46471 a_3160_47472# a_3177_46902# 0.009123f
C46472 a_2063_45854# a_2864_46660# 0.002177f
C46473 a_18248_44752# a_18579_44172# 0.001274f
C46474 a_n2661_44458# a_2675_43914# 9.03e-20
C46475 a_1307_43914# a_3737_43940# 0.058797f
C46476 a_18287_44626# a_18245_44484# 2.56e-19
C46477 a_n143_45144# a_n97_42460# 1.93e-21
C46478 a_n913_45002# a_1209_43370# 7.74e-20
C46479 a_n2017_45002# a_1568_43370# 4.02e-19
C46480 a_2437_43646# a_3626_43646# 6e-20
C46481 a_n967_45348# a_n1190_43762# 1.32e-19
C46482 a_3357_43084# a_2896_43646# 2.67e-19
C46483 a_n967_45348# VDD 0.556063f
C46484 a_22400_42852# a_22469_39537# 0.019601f
C46485 a_21005_45260# a_11415_45002# 0.01592f
C46486 a_18184_42460# a_12741_44636# 0.041879f
C46487 a_21101_45002# a_20202_43084# 4.9e-19
C46488 a_7418_45067# a_3483_46348# 3.85e-19
C46489 a_17767_44458# a_15227_44166# 0.023473f
C46490 a_5495_43940# a_768_44030# 0.017815f
C46491 a_11691_44458# a_18900_46660# 6.04e-20
C46492 a_4574_45260# a_526_44458# 6.77e-19
C46493 a_3537_45260# a_n1925_42282# 0.055426f
C46494 a_16019_45002# a_15682_46116# 5.53e-19
C46495 a_10775_45002# a_10809_44734# 0.022389f
C46496 a_1307_43914# a_2324_44458# 0.129761f
C46497 a_n630_44306# a_n1613_43370# 0.003389f
C46498 a_7499_43940# a_n1151_42308# 4.39e-20
C46499 a_21115_43940# a_16327_47482# 2.26e-21
C46500 a_10533_42308# a_10723_42308# 0.23663f
C46501 a_1067_42314# a_7174_31319# 4.88e-21
C46502 a_n3674_38216# a_n4064_40160# 0.02459f
C46503 a_5342_30871# C0_P_btm 8.41e-20
C46504 a_5534_30871# C0_dummy_N_btm 2.22e-20
C46505 RST_Z START 0.033428f
C46506 a_19120_35138# VIN_N 0.001664f
C46507 EN_VIN_BSTR_N VREF_GND 0.85739f
C46508 a_9313_45822# a_9290_44172# 4.81e-22
C46509 a_11031_47542# a_11189_46129# 8.25e-21
C46510 a_n1435_47204# a_9569_46155# 2.34e-20
C46511 a_n2497_47436# a_526_44458# 0.06857f
C46512 a_n443_46116# a_2324_44458# 0.055032f
C46513 a_10227_46804# a_4185_45028# 3.04e-19
C46514 a_n2312_39304# a_n1853_46287# 3.91e-19
C46515 a_7927_46660# a_8492_46660# 7.99e-20
C46516 a_5807_45002# a_765_45546# 0.103324f
C46517 a_13661_43548# a_17339_46660# 0.599051f
C46518 a_4646_46812# a_8270_45546# 1.8e-19
C46519 a_10057_43914# a_8685_43396# 0.007406f
C46520 a_n2661_43922# a_104_43370# 7.49e-21
C46521 a_11691_44458# a_18525_43370# 1.92e-20
C46522 a_11827_44484# a_19700_43370# 4.41e-21
C46523 a_n2293_42834# a_n1423_42826# 0.011631f
C46524 a_n2293_43922# a_n97_42460# 0.136247f
C46525 a_1307_43914# a_8387_43230# 3.33e-20
C46526 a_n356_44636# a_1512_43396# 5.7e-20
C46527 a_n2661_42834# a_n2012_43396# 0.001847f
C46528 a_9159_44484# VDD 0.004886f
C46529 a_n4209_38216# C6_P_btm 1.26e-20
C46530 a_n3565_38216# C8_P_btm 1.65e-20
C46531 a_2711_45572# a_9049_44484# 0.025215f
C46532 a_5244_44056# a_1823_45246# 5.63e-19
C46533 a_16243_43396# a_12549_44172# 0.001317f
C46534 a_5829_43940# a_3090_45724# 0.003937f
C46535 a_9145_43396# a_n2293_46634# 0.238561f
C46536 a_15493_43940# a_13059_46348# 1.93e-19
C46537 a_n2661_44458# a_2277_45546# 1.47e-21
C46538 a_6298_44484# a_n357_42282# 3.34e-19
C46539 a_n2129_44697# a_n443_42852# 8.3e-20
C46540 a_n699_43396# a_2957_45546# 2.21e-19
C46541 a_11967_42832# a_19900_46494# 2.43e-21
C46542 a_5649_42852# a_13507_46334# 0.136078f
C46543 a_19479_31679# a_19864_35138# 6.24e-22
C46544 a_19963_31679# EN_VIN_BSTR_N 0.004167f
C46545 a_7715_46873# VDD 0.414019f
C46546 a_n3690_38528# a_n4209_38216# 2.69e-19
C46547 a_n3420_38528# a_n3607_38528# 0.001534f
C46548 a_14097_32519# VDAC_N 2.69e-19
C46549 a_n4318_37592# a_n3420_37440# 0.001831f
C46550 a_n1630_35242# VDAC_Ni 2.54e-19
C46551 a_n784_42308# a_7754_38470# 1.35e-19
C46552 a_5932_42308# a_n3420_37984# 1.17e-19
C46553 a_20820_30879# a_22959_46660# 0.01739f
C46554 a_20202_43084# a_21542_46660# 7.08e-19
C46555 a_22591_46660# a_21076_30879# 3.06e-19
C46556 a_n2293_46634# a_n1099_45572# 0.006391f
C46557 a_n2661_46634# a_n755_45592# 4.56e-20
C46558 a_n1925_46634# a_n863_45724# 5.47e-20
C46559 a_n743_46660# a_n2293_45546# 6.76e-20
C46560 a_n1021_46688# a_n1079_45724# 4.95e-21
C46561 a_7411_46660# a_8034_45724# 6.76e-21
C46562 a_171_46873# a_n2661_45546# 7.37e-21
C46563 a_n2438_43548# a_n2956_38216# 0.020852f
C46564 a_5257_43370# a_6347_46155# 2.62e-19
C46565 a_3090_45724# a_17957_46116# 1.57e-19
C46566 a_15227_44166# a_15015_46420# 1.48e-19
C46567 a_12359_47026# a_12005_46116# 1.79e-19
C46568 a_16292_46812# a_15682_46116# 0.005299f
C46569 a_11813_46116# a_6945_45028# 1.65e-19
C46570 a_11186_47026# a_10809_44734# 3.59e-20
C46571 a_5013_44260# a_5649_42852# 1.41e-20
C46572 a_21115_43940# a_10341_43396# 1.36e-20
C46573 a_6671_43940# a_6765_43638# 2.18e-19
C46574 a_14021_43940# a_8685_43396# 0.002318f
C46575 a_10555_44260# a_10695_43548# 2.11e-20
C46576 a_n984_44318# a_n1076_43230# 6.38e-21
C46577 a_11967_42832# a_12089_42308# 0.022254f
C46578 a_n4318_40392# a_n4318_37592# 0.023213f
C46579 a_n1699_43638# a_n1821_43396# 3.16e-19
C46580 a_n447_43370# a_104_43370# 5.86e-20
C46581 a_15493_43940# a_15095_43370# 0.001144f
C46582 a_n1917_43396# VDD 0.204644f
C46583 a_4099_45572# a_n2661_43370# 0.002135f
C46584 a_15143_45578# a_14797_45144# 0.001287f
C46585 a_11688_45572# a_3232_43370# 2.05e-19
C46586 a_21363_45546# a_21188_45572# 0.233657f
C46587 a_20841_45814# a_20731_45938# 0.097745f
C46588 a_20623_45572# a_20528_45572# 0.049827f
C46589 a_n784_42308# a_768_44030# 3.1e-20
C46590 a_10835_43094# a_3090_45724# 0.008534f
C46591 a_22400_42852# a_22612_30879# 2.55e-19
C46592 a_14097_32519# a_21588_30879# 0.056136f
C46593 a_1568_43370# a_526_44458# 0.220609f
C46594 a_15493_43396# a_n443_42852# 0.025952f
C46595 a_9803_43646# a_8953_45546# 0.091141f
C46596 a_n4064_40160# w_1575_34946# 9.7e-19
C46597 a_9049_44484# a_9313_45822# 0.119007f
C46598 a_13163_45724# a_4915_47217# 1.03e-19
C46599 a_19553_46090# a_16375_45002# 2.34e-20
C46600 a_18819_46122# a_19431_46494# 3.82e-19
C46601 a_5937_45572# a_n357_42282# 1.32e-19
C46602 a_8199_44636# a_n755_45592# 5.59e-20
C46603 a_18189_46348# a_18051_46116# 0.045453f
C46604 a_18985_46122# a_19240_46482# 0.05936f
C46605 a_5066_45546# a_5527_46155# 8.1e-19
C46606 a_3483_46348# a_n443_42852# 1.96e-19
C46607 a_8791_43396# a_9127_43156# 0.007148f
C46608 a_16547_43609# a_4361_42308# 9.06e-21
C46609 a_17324_43396# a_743_42282# 8.71e-21
C46610 a_18525_43370# a_4190_30871# 0.005875f
C46611 a_3626_43646# a_14543_43071# 4.05e-22
C46612 a_n2661_42282# a_2351_42308# 8.86e-20
C46613 a_16664_43396# a_16823_43084# 0.005264f
C46614 a_15743_43084# a_19177_43646# 4.34e-19
C46615 a_11967_42832# a_18907_42674# 4.8e-21
C46616 a_22223_42860# VDD 0.250812f
C46617 en_comp VDAC_P 0.003461f
C46618 a_4099_45572# a_2998_44172# 3.68e-22
C46619 a_11787_45002# a_11827_44484# 2.02e-20
C46620 a_1307_43914# a_16922_45042# 1.8e-20
C46621 a_8696_44636# a_13857_44734# 0.004972f
C46622 a_3429_45260# a_n2661_44458# 8.32e-19
C46623 a_n1059_45260# a_8701_44490# 4.94e-19
C46624 a_n967_45348# a_n699_43396# 4.56e-20
C46625 a_327_44734# a_n1177_44458# 1.88e-21
C46626 a_n2017_45002# a_5883_43914# 8.44e-20
C46627 a_685_42968# a_n863_45724# 0.052365f
C46628 a_4743_43172# a_526_44458# 0.00549f
C46629 a_n4064_37440# w_1575_34946# 3.26e-19
C46630 a_15903_45785# a_6755_46942# 0.192397f
C46631 a_15143_45578# a_14976_45028# 0.005582f
C46632 a_14495_45572# a_15368_46634# 3.5e-20
C46633 a_6511_45714# a_765_45546# 5.27e-21
C46634 a_11682_45822# a_11735_46660# 1.59e-20
C46635 a_n2661_45010# a_n743_46660# 8.45e-21
C46636 a_6171_45002# a_12891_46348# 0.040434f
C46637 a_413_45260# a_19321_45002# 2.02e-19
C46638 a_n1059_45260# a_n2293_46634# 0.051525f
C46639 a_5691_45260# a_768_44030# 4.31e-21
C46640 a_n2956_37592# a_n2956_39768# 0.047483f
C46641 a_3232_43370# a_12549_44172# 3.99e-21
C46642 a_n2840_45002# a_n2438_43548# 0.002993f
C46643 a_n2293_45010# a_n1925_46634# 3.1e-20
C46644 a_n2017_45002# a_n2104_46634# 7.56e-20
C46645 a_2982_43646# a_13258_32519# 0.086314f
C46646 a_n2472_42826# a_n4318_38216# 0.006796f
C46647 a_n1853_43023# a_n3674_38680# 3.63e-19
C46648 a_743_42282# a_1184_42692# 0.005701f
C46649 a_10341_43396# a_10533_42308# 2.73e-21
C46650 a_3626_43646# a_19511_42282# 0.182478f
C46651 a_13678_32519# a_n784_42308# 0.009139f
C46652 a_14209_32519# COMP_P 7.77e-21
C46653 a_18985_46122# START 0.001317f
C46654 a_14275_46494# CLK 3.42e-21
C46655 a_19553_46090# RST_Z 3.65e-21
C46656 a_n4209_39590# VDD 2.06918f
C46657 a_n237_47217# a_9804_47204# 3.49e-19
C46658 a_1239_47204# a_n881_46662# 8.4e-19
C46659 a_1431_47204# a_n1613_43370# 4.26e-19
C46660 a_16241_47178# a_16327_47482# 0.185907f
C46661 a_15673_47210# a_16023_47582# 0.228897f
C46662 a_14955_47212# a_10227_46804# 0.175517f
C46663 a_15507_47210# a_16588_47582# 0.102325f
C46664 a_11599_46634# a_17591_47464# 1.03e-20
C46665 a_6575_47204# a_4883_46098# 7.51e-20
C46666 a_3160_47472# a_3315_47570# 0.005289f
C46667 a_3815_47204# a_2747_46873# 2.57e-20
C46668 a_12861_44030# a_18780_47178# 9.61e-19
C46669 a_13717_47436# a_18597_46090# 1.1e-19
C46670 a_18494_42460# a_20159_44458# 0.024732f
C46671 a_21005_45260# a_11967_42832# 3.36e-20
C46672 a_949_44458# a_n2661_43922# 0.055363f
C46673 a_2779_44458# a_n2661_42834# 0.00388f
C46674 a_10157_44484# a_9313_44734# 0.026406f
C46675 a_19778_44110# a_20640_44752# 4.84e-20
C46676 a_n2293_42834# a_n1549_44318# 7.42e-19
C46677 a_16922_45042# a_18579_44172# 1.03e-19
C46678 a_742_44458# a_n2293_43922# 1.56e-21
C46679 a_5518_44484# a_5608_44484# 0.008441f
C46680 a_5343_44458# a_5708_44484# 0.048542f
C46681 a_7499_43078# a_8229_43396# 0.001513f
C46682 a_19431_45546# a_19319_43548# 2.72e-20
C46683 a_11691_44458# a_16241_44484# 2.22e-19
C46684 a_11827_44484# a_17325_44484# 3.91e-19
C46685 a_6171_45002# a_11750_44172# 3.21e-19
C46686 a_8191_45002# a_8333_44056# 4.8e-20
C46687 a_13575_42558# a_n357_42282# 3.32e-21
C46688 a_18907_42674# a_13259_45724# 4.44e-20
C46689 a_n2216_39072# a_n2956_39304# 8.63e-19
C46690 a_n2860_39072# a_n2956_38680# 8.73e-19
C46691 a_16680_45572# VDD 0.275078f
C46692 a_20820_30879# C10_N_btm 4.87e-19
C46693 a_21076_30879# C7_N_btm 0.00198f
C46694 a_14537_43396# a_11415_45002# 0.04406f
C46695 a_13556_45296# a_12741_44636# 0.046411f
C46696 a_2382_45260# a_3699_46348# 2.18e-21
C46697 a_3065_45002# a_3147_46376# 2.49e-20
C46698 a_18587_45118# a_3090_45724# 0.039584f
C46699 a_5343_44458# a_5257_43370# 0.063407f
C46700 a_14815_43914# a_13661_43548# 0.060575f
C46701 a_13940_44484# a_768_44030# 0.003215f
C46702 a_5111_44636# a_1823_45246# 0.002758f
C46703 a_15903_45785# a_8049_45260# 0.003516f
C46704 a_3260_45572# a_3218_45724# 0.010055f
C46705 a_12016_45572# a_10586_45546# 6.73e-20
C46706 a_20273_45572# a_19900_46494# 9.45e-19
C46707 a_20107_45572# a_20708_46348# 0.007797f
C46708 a_2437_43646# a_15015_46420# 1.91e-20
C46709 a_3357_43084# a_13925_46122# 1.09e-20
C46710 a_413_45260# a_5068_46348# 2.65e-21
C46711 a_n913_45002# a_8953_45546# 0.052161f
C46712 a_n2661_42282# a_584_46384# 3.54e-21
C46713 a_n784_42308# a_6123_31319# 0.144274f
C46714 a_2713_42308# a_3318_42354# 9.16e-19
C46715 a_15597_42852# a_15803_42450# 1.45e-19
C46716 a_1067_42314# a_5932_42308# 4.34e-21
C46717 a_14097_32519# a_5742_30871# 0.004679f
C46718 a_4190_30871# C0_dummy_N_btm 1.45e-20
C46719 a_22521_40055# a_22545_38993# 0.004924f
C46720 a_22459_39145# a_22521_39511# 0.075012f
C46721 a_5807_45002# a_10623_46897# 0.005882f
C46722 a_n743_46660# a_5732_46660# 1.15e-21
C46723 a_1799_45572# a_3524_46660# 1.24e-20
C46724 a_2609_46660# a_3177_46902# 0.17072f
C46725 a_2443_46660# a_2959_46660# 0.110816f
C46726 a_n1925_46634# a_5072_46660# 0.001838f
C46727 a_2107_46812# a_3221_46660# 6.44e-19
C46728 a_9804_47204# a_8270_45546# 4.96e-19
C46729 a_n881_46662# a_11186_47026# 1.85e-19
C46730 a_11453_44696# a_19466_46812# 0.004642f
C46731 a_14311_47204# a_765_45546# 0.003681f
C46732 a_16023_47582# a_16388_46812# 0.001491f
C46733 a_16327_47482# a_16721_46634# 7.05e-19
C46734 a_13717_47436# a_19123_46287# 4.43e-21
C46735 a_12861_44030# a_18285_46348# 0.247326f
C46736 a_n746_45260# a_n1076_46494# 5.44e-19
C46737 a_n2109_47186# a_2202_46116# 6.76e-21
C46738 a_n1741_47186# a_1138_42852# 1.21e-20
C46739 a_742_44458# a_n97_42460# 0.083982f
C46740 a_n984_44318# a_175_44278# 1.1e-19
C46741 a_20193_45348# a_2982_43646# 4.86e-20
C46742 a_1307_43914# a_15743_43084# 1.61e-19
C46743 a_14539_43914# a_15037_43940# 0.054182f
C46744 a_n699_43396# a_n1917_43396# 1.68e-20
C46745 a_11823_42460# a_15785_43172# 3.45e-20
C46746 a_n2661_43922# a_11341_43940# 3.15e-19
C46747 a_13249_42308# a_13569_43230# 2.14e-19
C46748 a_n2293_45010# a_685_42968# 1.26e-20
C46749 a_n2661_45010# a_1847_42826# 1.52e-22
C46750 a_n967_45348# a_n4318_38680# 1.38e-21
C46751 a_n1059_45260# a_n1533_42852# 1.94e-19
C46752 a_n4251_37440# VDD 3.95e-19
C46753 a_17531_42308# RST_Z 1.65e-20
C46754 a_n1917_44484# VDD 0.186988f
C46755 a_7174_31319# EN_VIN_BSTR_N 0.051994f
C46756 a_20362_44736# a_12741_44636# 0.00339f
C46757 a_20835_44721# a_11415_45002# 0.002797f
C46758 a_3080_42308# a_768_44030# 1.6e-19
C46759 a_n4318_39304# a_n2442_46660# 0.023691f
C46760 a_n2661_43370# a_n452_45724# 2.54e-20
C46761 a_n2661_44458# a_8049_45260# 5.47e-19
C46762 a_45_45144# a_n443_42852# 2.99e-19
C46763 a_5883_43914# a_526_44458# 0.0033f
C46764 a_n1243_43396# a_n1613_43370# 2.95e-19
C46765 a_17364_32525# w_11334_34010# 0.016546f
C46766 a_14579_43548# a_10227_46804# 0.118896f
C46767 a_11823_42460# CLK 3.11e-20
C46768 a_n3565_39590# a_n4064_39616# 0.231239f
C46769 a_7174_31319# a_1239_39043# 7.77e-20
C46770 a_n4064_40160# a_n4251_39616# 0.001069f
C46771 a_13747_46662# VDD 3.70214f
C46772 a_18479_47436# a_n357_42282# 0.003001f
C46773 SMPL_ON_N a_20692_30879# 0.029397f
C46774 a_11453_44696# a_20205_31679# 1.75e-20
C46775 a_7411_46660# a_8016_46348# 6.73e-19
C46776 a_7715_46873# a_7920_46348# 0.080253f
C46777 a_n1925_46634# a_1431_46436# 3.57e-19
C46778 a_5807_45002# a_6347_46155# 2.63e-19
C46779 a_n2293_46634# a_n1925_42282# 0.030317f
C46780 a_16388_46812# a_16751_46987# 0.005265f
C46781 a_10554_47026# a_3483_46348# 5.06e-20
C46782 a_3090_45724# a_11415_45002# 0.16525f
C46783 a_14673_44172# a_4361_42308# 5.89e-21
C46784 a_18579_44172# a_15743_43084# 0.003564f
C46785 a_17517_44484# a_21487_43396# 9.64e-21
C46786 a_n2661_42834# a_n13_43084# 6.03e-20
C46787 a_n2293_43922# a_n901_43156# 3.99e-20
C46788 a_6109_44484# a_5755_42852# 6.71e-22
C46789 a_n356_44636# a_10835_43094# 1.71e-20
C46790 a_1307_43914# a_1606_42308# 0.003969f
C46791 a_5111_44636# a_5934_30871# 6.55e-19
C46792 a_n913_45002# a_14456_42282# 0.006851f
C46793 a_n2017_45002# a_13333_42558# 0.001525f
C46794 a_20269_44172# VDD 0.169009f
C46795 a_5263_45724# a_3537_45260# 3.44e-19
C46796 a_2711_45572# a_5147_45002# 0.003609f
C46797 a_4235_43370# a_1823_45246# 0.029154f
C46798 a_5755_42852# a_4646_46812# 5.33e-19
C46799 a_18525_43370# a_15227_44166# 2.71e-21
C46800 a_15037_43396# a_3090_45724# 1.16e-20
C46801 a_2479_44172# a_n357_42282# 0.008172f
C46802 a_9306_43218# a_n1613_43370# 0.001965f
C46803 a_20256_42852# a_16327_47482# 8.08e-21
C46804 a_1606_42308# a_n443_46116# 3.46e-19
C46805 a_1755_42282# a_4791_45118# 0.002644f
C46806 VDAC_Pi RST_Z 0.002358f
C46807 a_n3420_37984# VREF 1.33e-19
C46808 a_n4064_37984# VIN_P 0.06139f
C46809 a_n4209_37414# a_n1838_35608# 1.81e-19
C46810 a_18184_42460# RST_Z 0.001648f
C46811 a_4419_46090# VDD 0.664887f
C46812 a_2711_45572# a_n2109_47186# 0.032969f
C46813 a_n3565_39304# a_n4334_37440# 5.28e-19
C46814 a_n4209_39304# a_n3690_37440# 2.3e-19
C46815 a_n4209_38216# a_n2216_37984# 0.001433f
C46816 C8_N_btm C10_N_btm 2.07867f
C46817 a_12741_44636# a_16375_45002# 0.042457f
C46818 a_765_45546# a_n755_45592# 0.004312f
C46819 a_6165_46155# a_5066_45546# 0.041118f
C46820 a_5164_46348# a_5210_46155# 0.006879f
C46821 a_5068_46348# a_5527_46155# 6.64e-19
C46822 a_18819_46122# a_19335_46494# 0.108964f
C46823 a_18985_46122# a_19553_46090# 0.16939f
C46824 a_15682_46116# a_6945_45028# 1.56e-19
C46825 a_14840_46494# a_10809_44734# 3.79e-21
C46826 a_n1699_43638# a_n1736_43218# 1.6e-19
C46827 a_2982_43646# a_20301_43646# 9.07e-21
C46828 a_n1809_43762# a_n1991_42858# 9.16e-20
C46829 a_n97_42460# a_n901_43156# 0.011039f
C46830 a_14021_43940# a_17333_42852# 4.57e-21
C46831 a_n2293_43922# a_10533_42308# 4.97e-20
C46832 a_9313_44734# a_14113_42308# 4.32e-20
C46833 a_3080_42308# a_13678_32519# 0.002941f
C46834 a_9803_43646# a_10149_43396# 0.013377f
C46835 a_9885_43646# a_10341_43396# 0.001685f
C46836 a_9145_43396# a_14537_43646# 0.003686f
C46837 a_n356_44636# a_16269_42308# 4.62e-19
C46838 a_3422_30871# a_n1630_35242# 0.828871f
C46839 a_17730_32519# COMP_P 1.26e-20
C46840 a_8685_43396# a_13943_43396# 5.42e-19
C46841 a_n1917_43396# a_n4318_38680# 3.79e-19
C46842 VCM VSS 30.6764f
C46843 VREF_GND VSS 17.6166f
C46844 VREF VSS 8.78695f
C46845 VIN_N VSS 13.1675f
C46846 VIN_P VSS 13.143001f
C46847 CLK VSS 1.55797f
C46848 EN_OFFSET_CAL VSS 0.505642f
C46849 DATA[5] VSS 0.561058f
C46850 DATA[4] VSS 0.755679f
C46851 DATA[3] VSS 1.01838f
C46852 DATA[2] VSS 0.536983f
C46853 DATA[1] VSS 0.550109f
C46854 DATA[0] VSS 0.616231f
C46855 CLK_DATA VSS 0.488979f
C46856 SINGLE_ENDED VSS 0.60168f
C46857 START VSS 0.991673f
C46858 RST_Z VSS 11.389f
C46859 VDD VSS 0.588168p
C46860 C10_N_btm VSS 0.210692p **FLOATING
C46861 C9_N_btm VSS 79.926506f **FLOATING
C46862 C8_N_btm VSS 45.547f **FLOATING
C46863 C7_N_btm VSS 25.886099f **FLOATING
C46864 C6_N_btm VSS 15.5273f **FLOATING
C46865 C5_N_btm VSS 9.624539f **FLOATING
C46866 C4_N_btm VSS 8.794849f **FLOATING
C46867 C3_N_btm VSS 6.38289f **FLOATING
C46868 C2_N_btm VSS 5.46028f **FLOATING
C46869 C1_N_btm VSS 5.26099f **FLOATING
C46870 C0_N_btm VSS 7.20283f **FLOATING
C46871 C0_dummy_N_btm VSS 5.03035f **FLOATING
C46872 C0_dummy_P_btm VSS 5.0181f **FLOATING
C46873 C0_P_btm VSS 7.1984f **FLOATING
C46874 C1_P_btm VSS 5.27428f **FLOATING
C46875 C2_P_btm VSS 5.46972f **FLOATING
C46876 C3_P_btm VSS 6.37616f **FLOATING
C46877 C4_P_btm VSS 8.785789f **FLOATING
C46878 C5_P_btm VSS 9.614769f **FLOATING
C46879 C6_P_btm VSS 15.5172f **FLOATING
C46880 C7_P_btm VSS 25.876501f **FLOATING
C46881 C8_P_btm VSS 45.531998f **FLOATING
C46882 C9_P_btm VSS 79.8995f **FLOATING
C46883 C10_P_btm VSS 0.210676p **FLOATING
C46884 a_21589_35634# VSS 0.729455f **FLOATING
C46885 a_19864_35138# VSS 1.75392f **FLOATING
C46886 a_19120_35138# VSS 1.69667f **FLOATING
C46887 a_18194_35068# VSS 2.11801f **FLOATING
C46888 EN_VIN_BSTR_N VSS 9.04132f **FLOATING
C46889 a_11530_34132# VSS 13.9862f **FLOATING
C46890 a_n83_35174# VSS 1.72857f **FLOATING
C46891 EN_VIN_BSTR_P VSS 9.26595f **FLOATING
C46892 a_n923_35174# VSS 14.088f **FLOATING
C46893 a_n1532_35090# VSS 2.16074f **FLOATING
C46894 a_n1386_35608# VSS 1.75773f **FLOATING
C46895 a_n1838_35608# VSS 0.737725f **FLOATING
C46896 a_22717_36887# VSS 0.092029f **FLOATING
C46897 a_22717_37285# VSS 0.095943f **FLOATING
C46898 a_22705_37990# VSS 0.007968f **FLOATING
C46899 a_22609_37990# VSS 0.473213f **FLOATING
C46900 a_22705_38406# VSS 0.010928f **FLOATING
C46901 a_22609_38406# VSS 0.588255f **FLOATING
C46902 CAL_P VSS 11.418599f **FLOATING
C46903 a_22876_39857# VSS 0.00127f **FLOATING
C46904 a_22780_39857# VSS 7.39e-19 **FLOATING
C46905 a_22469_39537# VSS 2.5954f **FLOATING
C46906 a_22821_38993# VSS 0.55301f **FLOATING
C46907 a_22545_38993# VSS 0.35571f **FLOATING
C46908 a_22521_39511# VSS 1.85851f **FLOATING
C46909 a_22780_40081# VSS 0.002233f **FLOATING
C46910 a_22459_39145# VSS 2.29285f **FLOATING
C46911 a_22521_40055# VSS 1.21928f **FLOATING
C46912 a_22780_40945# VSS 0.002478f **FLOATING
C46913 a_22469_40625# VSS 1.56643f **FLOATING
C46914 a_22521_40599# VSS 1.85568f **FLOATING
C46915 CAL_N VSS 8.69238f **FLOATING
C46916 a_11206_38545# VSS 0.713084f **FLOATING
C46917 VDAC_P VSS 0.107582p **FLOATING
C46918 a_8912_37509# VSS 3.72815f **FLOATING
C46919 VDAC_N VSS 0.108181p **FLOATING
C46920 a_6886_37412# VSS 3.84457f **FLOATING
C46921 a_5700_37509# VSS 2.08109f **FLOATING
C46922 a_5088_37509# VSS 2.72043f **FLOATING
C46923 a_4338_37500# VSS 2.61369f **FLOATING
C46924 a_3726_37500# VSS 4.48332f **FLOATING
C46925 a_n3607_37440# VSS 0.002657f **FLOATING
C46926 a_n4251_37440# VSS 0.003621f **FLOATING
C46927 a_n2860_37690# VSS 0.001049f **FLOATING
C46928 a_n2302_37690# VSS 0.514508f **FLOATING
C46929 a_n4064_37440# VSS 1.7233f **FLOATING
C46930 a_n2946_37690# VSS 0.517242f **FLOATING
C46931 a_n3420_37440# VSS 5.23286f **FLOATING
C46932 a_n3690_37440# VSS 0.548488f **FLOATING
C46933 a_n3565_37414# VSS 3.16456f **FLOATING
C46934 a_n4334_37440# VSS 0.561497f **FLOATING
C46935 a_n4209_37414# VSS 3.16799f **FLOATING
C46936 a_8530_39574# VSS 2.76228f **FLOATING
C46937 a_7754_38470# VSS 3.24598f **FLOATING
C46938 a_3754_38470# VSS 4.77654f **FLOATING
C46939 VDAC_Ni VSS 2.86404f **FLOATING
C46940 a_7754_38636# VSS 0.353706f **FLOATING
C46941 a_3754_38802# VSS 0.390074f **FLOATING
C46942 a_7754_38968# VSS 0.330037f **FLOATING
C46943 a_3754_39134# VSS 0.401983f **FLOATING
C46944 a_7754_39300# VSS 0.330682f **FLOATING
C46945 a_3754_39466# VSS 0.401172f **FLOATING
C46946 a_7754_39632# VSS 0.340942f **FLOATING
C46947 VDAC_Pi VSS 3.50355f **FLOATING
C46948 a_7754_39964# VSS 2.62481f **FLOATING
C46949 a_7754_40130# VSS 2.84104f **FLOATING
C46950 a_3754_39964# VSS 0.671366f **FLOATING
C46951 a_n2860_37984# VSS 0.001049f **FLOATING
C46952 a_2113_38308# VSS 2.64372f **FLOATING
C46953 a_n3607_38304# VSS 0.002772f **FLOATING
C46954 a_n4251_38304# VSS 0.003689f **FLOATING
C46955 a_n2302_37984# VSS 0.483504f **FLOATING
C46956 a_n4064_37984# VSS 1.65074f **FLOATING
C46957 a_n2946_37984# VSS 0.485942f **FLOATING
C46958 a_n3420_37984# VSS 1.75918f **FLOATING
C46959 a_n3690_38304# VSS 0.517812f **FLOATING
C46960 a_n3565_38216# VSS 1.49258f **FLOATING
C46961 a_n4334_38304# VSS 0.529531f **FLOATING
C46962 a_n4209_38216# VSS 3.03885f **FLOATING
C46963 a_n3607_38528# VSS 0.002662f **FLOATING
C46964 a_n4251_38528# VSS 0.003622f **FLOATING
C46965 a_2684_37794# VSS 0.414596f **FLOATING
C46966 a_1177_38525# VSS 0.641945f **FLOATING
C46967 a_n2860_38778# VSS 0.001049f **FLOATING
C46968 a_n2302_38778# VSS 0.483515f **FLOATING
C46969 a_n4064_38528# VSS 1.69554f **FLOATING
C46970 a_n2946_38778# VSS 0.485895f **FLOATING
C46971 a_n3420_38528# VSS 2.03238f **FLOATING
C46972 a_n3690_38528# VSS 0.516979f **FLOATING
C46973 a_n3565_38502# VSS 1.56105f **FLOATING
C46974 a_n4334_38528# VSS 0.529888f **FLOATING
C46975 a_n4209_38502# VSS 3.0227f **FLOATING
C46976 a_2112_39137# VSS 0.414248f **FLOATING
C46977 a_n2860_39072# VSS 0.001051f **FLOATING
C46978 comp_n VSS 0.568772f **FLOATING
C46979 a_1736_39043# VSS 0.897653f **FLOATING
C46980 a_1239_39043# VSS 0.614001f **FLOATING
C46981 a_n3607_39392# VSS 0.002762f **FLOATING
C46982 a_n4251_39392# VSS 0.003686f **FLOATING
C46983 a_n2302_39072# VSS 0.483504f **FLOATING
C46984 a_n4064_39072# VSS 1.71794f **FLOATING
C46985 a_n2946_39072# VSS 0.486447f **FLOATING
C46986 a_n3420_39072# VSS 2.21624f **FLOATING
C46987 a_n3690_39392# VSS 0.517965f **FLOATING
C46988 a_n3565_39304# VSS 1.46005f **FLOATING
C46989 a_n4334_39392# VSS 0.529516f **FLOATING
C46990 a_n4209_39304# VSS 3.25385f **FLOATING
C46991 a_1343_38525# VSS 3.5734f **FLOATING
C46992 a_n3607_39616# VSS 0.002672f **FLOATING
C46993 a_n4251_39616# VSS 0.003625f **FLOATING
C46994 a_1736_39587# VSS 1.10676f **FLOATING
C46995 a_1239_39587# VSS 0.634559f **FLOATING
C46996 a_n2860_39866# VSS 0.001465f **FLOATING
C46997 a_n2302_39866# VSS 0.483537f **FLOATING
C46998 a_n4064_39616# VSS 2.1793f **FLOATING
C46999 a_n2946_39866# VSS 0.527929f **FLOATING
C47000 a_n3420_39616# VSS 2.11281f **FLOATING
C47001 a_n3690_39616# VSS 0.574329f **FLOATING
C47002 a_n3565_39590# VSS 2.12343f **FLOATING
C47003 a_n4334_39616# VSS 0.529903f **FLOATING
C47004 a_n4209_39590# VSS 4.08222f **FLOATING
C47005 a_n4251_40480# VSS 0.003684f **FLOATING
C47006 a_n2302_40160# VSS 0.522244f **FLOATING
C47007 a_n4064_40160# VSS 3.29808f **FLOATING
C47008 a_n4334_40480# VSS 0.578721f **FLOATING
C47009 a_n4315_30879# VSS 5.10683f **FLOATING
C47010 a_21973_42336# VSS 0.004685f **FLOATING
C47011 a_22465_38105# VSS 1.91115f **FLOATING
C47012 a_21421_42336# VSS 0.004685f **FLOATING
C47013 a_18997_42308# VSS 0.004143f **FLOATING
C47014 a_22775_42308# VSS 0.602961f **FLOATING
C47015 a_21613_42308# VSS 0.725408f **FLOATING
C47016 a_21887_42336# VSS 0.234022f **FLOATING
C47017 a_21335_42336# VSS 0.259392f **FLOATING
C47018 a_7174_31319# VSS 5.51208f **FLOATING
C47019 a_20712_42282# VSS 0.349662f **FLOATING
C47020 a_20107_42308# VSS 0.344464f **FLOATING
C47021 a_13258_32519# VSS 6.359931f **FLOATING
C47022 a_19647_42308# VSS 0.313304f **FLOATING
C47023 a_19511_42282# VSS 0.751141f **FLOATING
C47024 a_18548_42308# VSS 0.005248f **FLOATING
C47025 a_18310_42308# VSS 0.005141f **FLOATING
C47026 a_18220_42308# VSS 0.003723f **FLOATING
C47027 a_18214_42558# VSS 0.006283f **FLOATING
C47028 a_19332_42282# VSS 0.31505f **FLOATING
C47029 a_18907_42674# VSS 0.209311f **FLOATING
C47030 a_18727_42674# VSS 0.233526f **FLOATING
C47031 a_18057_42282# VSS 0.370712f **FLOATING
C47032 a_17531_42308# VSS 0.253358f **FLOATING
C47033 a_17303_42282# VSS 1.19698f **FLOATING
C47034 a_4958_30871# VSS 5.01459f **FLOATING
C47035 a_16269_42308# VSS 0.006939f **FLOATING
C47036 a_16197_42308# VSS 0.004992f **FLOATING
C47037 a_15761_42308# VSS 4.65e-19 **FLOATING
C47038 a_15521_42308# VSS 0.001281f **FLOATING
C47039 a_17124_42282# VSS 0.332693f **FLOATING
C47040 a_16522_42674# VSS 0.073862f **FLOATING
C47041 a_16104_42674# VSS 0.004694f **FLOATING
C47042 a_13921_42308# VSS 0.002122f **FLOATING
C47043 a_13657_42308# VSS 0.006177f **FLOATING
C47044 a_11897_42308# VSS 0.002019f **FLOATING
C47045 a_11633_42308# VSS 0.006177f **FLOATING
C47046 a_10149_42308# VSS 0.003101f **FLOATING
C47047 a_9885_42308# VSS 0.007915f **FLOATING
C47048 a_15890_42674# VSS 0.180637f **FLOATING
C47049 a_15959_42545# VSS 0.263128f **FLOATING
C47050 a_15803_42450# VSS 0.566963f **FLOATING
C47051 a_15764_42576# VSS 0.298494f **FLOATING
C47052 a_15486_42560# VSS 0.263746f **FLOATING
C47053 a_15051_42282# VSS 0.790649f **FLOATING
C47054 a_14113_42308# VSS 1.42448f **FLOATING
C47055 a_13657_42558# VSS 0.00274f **FLOATING
C47056 a_13249_42558# VSS 7.16e-20 **FLOATING
C47057 a_14456_42282# VSS 0.33927f **FLOATING
C47058 a_13575_42558# VSS 0.370369f **FLOATING
C47059 a_13070_42354# VSS 0.222095f **FLOATING
C47060 a_12563_42308# VSS 0.330976f **FLOATING
C47061 a_11633_42558# VSS 0.002749f **FLOATING
C47062 a_11551_42558# VSS 0.372919f **FLOATING
C47063 a_5742_30871# VSS 8.19455f **FLOATING
C47064 a_11323_42473# VSS 0.253445f **FLOATING
C47065 a_10723_42308# VSS 0.342975f **FLOATING
C47066 a_10533_42308# VSS 0.310658f **FLOATING
C47067 a_9885_42558# VSS 0.00274f **FLOATING
C47068 a_9377_42558# VSS 7.16e-20 **FLOATING
C47069 a_9803_42558# VSS 0.370474f **FLOATING
C47070 a_9223_42460# VSS 0.236204f **FLOATING
C47071 a_8791_42308# VSS 0.301f **FLOATING
C47072 a_8685_42308# VSS 0.163732f **FLOATING
C47073 a_8325_42308# VSS 0.316205f **FLOATING
C47074 a_4169_42308# VSS 0.00288f **FLOATING
C47075 a_3905_42308# VSS 0.007531f **FLOATING
C47076 a_8515_42308# VSS 0.250762f **FLOATING
C47077 a_5934_30871# VSS 5.17487f **FLOATING
C47078 a_7963_42308# VSS 0.256292f **FLOATING
C47079 a_6123_31319# VSS 5.02459f **FLOATING
C47080 a_7227_42308# VSS 0.359705f **FLOATING
C47081 a_6761_42308# VSS 0.447596f **FLOATING
C47082 a_5932_42308# VSS 5.11988f **FLOATING
C47083 a_6171_42473# VSS 0.257988f **FLOATING
C47084 a_5755_42308# VSS 0.314735f **FLOATING
C47085 a_5421_42558# VSS 7.16e-20 **FLOATING
C47086 a_4921_42308# VSS 0.511258f **FLOATING
C47087 a_3905_42558# VSS 0.00274f **FLOATING
C47088 a_3497_42558# VSS 7.16e-20 **FLOATING
C47089 a_5379_42460# VSS 0.564806f **FLOATING
C47090 a_5267_42460# VSS 0.204309f **FLOATING
C47091 a_3823_42558# VSS 0.381485f **FLOATING
C47092 a_3318_42354# VSS 0.238394f **FLOATING
C47093 a_2903_42308# VSS 0.340659f **FLOATING
C47094 a_2713_42308# VSS 0.31991f **FLOATING
C47095 a_n39_42308# VSS 0.006513f **FLOATING
C47096 a_n327_42308# VSS 0.002036f **FLOATING
C47097 a_2351_42308# VSS 0.210162f **FLOATING
C47098 a_2123_42473# VSS 0.21778f **FLOATING
C47099 a_1755_42282# VSS 3.17706f **FLOATING
C47100 a_1606_42308# VSS 5.2551f **FLOATING
C47101 a_1149_42558# VSS 5.47e-35 **FLOATING
C47102 a_961_42354# VSS 0.215753f **FLOATING
C47103 a_1184_42692# VSS 0.222827f **FLOATING
C47104 a_1576_42282# VSS 0.327109f **FLOATING
C47105 a_1067_42314# VSS 0.32917f **FLOATING
C47106 a_n1630_35242# VSS 10.134f **FLOATING
C47107 a_564_42282# VSS 0.36802f **FLOATING
C47108 a_n3674_37592# VSS 3.04613f **FLOATING
C47109 a_n327_42558# VSS 0.00274f **FLOATING
C47110 a_n784_42308# VSS 6.50157f **FLOATING
C47111 a_196_42282# VSS 0.343186f **FLOATING
C47112 a_n473_42460# VSS 0.366068f **FLOATING
C47113 a_n961_42308# VSS 0.328065f **FLOATING
C47114 a_n1329_42308# VSS 0.30898f **FLOATING
C47115 COMP_P VSS 11.0245f **FLOATING
C47116 a_n4318_37592# VSS 1.00428f **FLOATING
C47117 a_n1736_42282# VSS 0.320711f **FLOATING
C47118 a_n3674_38216# VSS 1.68571f **FLOATING
C47119 a_n2104_42282# VSS 0.346472f **FLOATING
C47120 a_n4318_38216# VSS 0.964502f **FLOATING
C47121 a_n2472_42282# VSS 0.335792f **FLOATING
C47122 a_n3674_38680# VSS 0.881032f **FLOATING
C47123 a_n2840_42282# VSS 0.343361f **FLOATING
C47124 a_20753_42852# VSS 0.004913f **FLOATING
C47125 a_20256_42852# VSS 1.31e-19 **FLOATING
C47126 a_14097_32519# VSS 1.90783f **FLOATING
C47127 a_22400_42852# VSS 2.02868f **FLOATING
C47128 a_20836_43172# VSS 0.003225f **FLOATING
C47129 a_20573_43172# VSS 6.53e-19 **FLOATING
C47130 a_20256_43172# VSS 0.192089f **FLOATING
C47131 a_18707_42852# VSS 0.004694f **FLOATING
C47132 a_19518_43218# VSS 0.001266f **FLOATING
C47133 a_19273_43230# VSS 4.65e-19 **FLOATING
C47134 a_18861_43218# VSS 0.00579f **FLOATING
C47135 a_17749_42852# VSS 7.16e-20 **FLOATING
C47136 a_16877_42852# VSS 0.00274f **FLOATING
C47137 a_16245_42852# VSS 0.004647f **FLOATING
C47138 a_15597_42852# VSS 0.001372f **FLOATING
C47139 a_18695_43230# VSS 0.008634f **FLOATING
C47140 a_18504_43218# VSS 0.078212f **FLOATING
C47141 a_17141_43172# VSS 0.002263f **FLOATING
C47142 a_16877_43172# VSS 0.007531f **FLOATING
C47143 a_16328_43172# VSS 0.003574f **FLOATING
C47144 a_15785_43172# VSS 0.004243f **FLOATING
C47145 a_14635_42282# VSS 0.336817f **FLOATING
C47146 a_13291_42460# VSS 0.197331f **FLOATING
C47147 a_13003_42852# VSS 0.004694f **FLOATING
C47148 a_13814_43218# VSS 0.001281f **FLOATING
C47149 a_13569_43230# VSS 4.65e-19 **FLOATING
C47150 a_11136_42852# VSS 0.004694f **FLOATING
C47151 a_13157_43218# VSS 0.004992f **FLOATING
C47152 a_12991_43230# VSS 0.006939f **FLOATING
C47153 a_12800_43218# VSS 0.073862f **FLOATING
C47154 a_11554_42852# VSS 0.073028f **FLOATING
C47155 a_11301_43218# VSS 0.006939f **FLOATING
C47156 a_11229_43218# VSS 0.004992f **FLOATING
C47157 a_10793_43218# VSS 4.65e-19 **FLOATING
C47158 a_10553_43218# VSS 0.001281f **FLOATING
C47159 a_8495_42852# VSS 0.004694f **FLOATING
C47160 a_9306_43218# VSS 0.001281f **FLOATING
C47161 a_9061_43230# VSS 4.65e-19 **FLOATING
C47162 a_8649_43218# VSS 0.004992f **FLOATING
C47163 a_7309_42852# VSS 0.003102f **FLOATING
C47164 a_5837_42852# VSS 0.00274f **FLOATING
C47165 a_5193_42852# VSS 0.00274f **FLOATING
C47166 a_4649_42852# VSS 0.006211f **FLOATING
C47167 a_3863_42891# VSS 2.7e-19 **FLOATING
C47168 a_8483_43230# VSS 0.006939f **FLOATING
C47169 a_8292_43218# VSS 0.073862f **FLOATING
C47170 a_7573_43172# VSS 0.002122f **FLOATING
C47171 a_7309_43172# VSS 0.006207f **FLOATING
C47172 a_6101_43172# VSS 0.00288f **FLOATING
C47173 a_5837_43172# VSS 0.005926f **FLOATING
C47174 a_5457_43172# VSS 0.002122f **FLOATING
C47175 a_5193_43172# VSS 0.005926f **FLOATING
C47176 a_4743_43172# VSS 0.005048f **FLOATING
C47177 a_4649_43172# VSS 0.005607f **FLOATING
C47178 a_1793_42852# VSS 1.13e-19 **FLOATING
C47179 a_1709_42852# VSS 9.12e-20 **FLOATING
C47180 a_873_42968# VSS 6.57e-20 **FLOATING
C47181 a_133_42852# VSS 0.003564f **FLOATING
C47182 a_4156_43218# VSS 0.003279f **FLOATING
C47183 a_3935_43218# VSS 0.002898f **FLOATING
C47184 a_3445_43172# VSS 0.001905f **FLOATING
C47185 a_n2293_42282# VSS 2.62914f **FLOATING
C47186 a_22959_42860# VSS 0.34332f **FLOATING
C47187 a_22223_42860# VSS 0.328988f **FLOATING
C47188 a_22165_42308# VSS 0.354098f **FLOATING
C47189 a_21671_42860# VSS 0.316857f **FLOATING
C47190 a_21195_42852# VSS 0.277519f **FLOATING
C47191 a_21356_42826# VSS 0.304166f **FLOATING
C47192 a_20922_43172# VSS 0.266814f **FLOATING
C47193 a_19987_42826# VSS 0.378798f **FLOATING
C47194 a_19164_43230# VSS 0.264863f **FLOATING
C47195 a_19339_43156# VSS 0.471496f **FLOATING
C47196 a_18599_43230# VSS 0.266382f **FLOATING
C47197 a_18817_42826# VSS 0.182139f **FLOATING
C47198 a_18249_42858# VSS 0.302863f **FLOATING
C47199 a_17333_42852# VSS 0.29982f **FLOATING
C47200 a_18083_42858# VSS 0.578693f **FLOATING
C47201 a_17701_42308# VSS 0.179963f **FLOATING
C47202 a_17595_43084# VSS 0.205109f **FLOATING
C47203 a_16795_42852# VSS 0.362281f **FLOATING
C47204 a_16414_43172# VSS 0.270304f **FLOATING
C47205 a_15567_42826# VSS 0.316627f **FLOATING
C47206 a_5342_30871# VSS 4.18155f **FLOATING
C47207 a_15279_43071# VSS 0.248252f **FLOATING
C47208 a_5534_30871# VSS 4.58471f **FLOATING
C47209 a_14543_43071# VSS 0.246071f **FLOATING
C47210 a_13460_43230# VSS 0.259861f **FLOATING
C47211 a_13635_43156# VSS 0.7696f **FLOATING
C47212 a_12895_43230# VSS 0.250159f **FLOATING
C47213 a_13113_42826# VSS 0.174096f **FLOATING
C47214 a_12545_42858# VSS 0.287468f **FLOATING
C47215 a_12089_42308# VSS 0.283874f **FLOATING
C47216 a_12379_42858# VSS 0.549229f **FLOATING
C47217 a_10341_42308# VSS 0.317389f **FLOATING
C47218 a_10922_42852# VSS 0.176112f **FLOATING
C47219 a_10991_42826# VSS 0.261283f **FLOATING
C47220 a_10796_42968# VSS 0.29877f **FLOATING
C47221 a_10835_43094# VSS 0.59174f **FLOATING
C47222 a_10518_42984# VSS 0.260322f **FLOATING
C47223 a_10083_42826# VSS 0.762957f **FLOATING
C47224 a_8952_43230# VSS 0.261046f **FLOATING
C47225 a_9127_43156# VSS 0.77314f **FLOATING
C47226 a_8387_43230# VSS 0.255573f **FLOATING
C47227 a_8605_42826# VSS 0.181157f **FLOATING
C47228 a_8037_42858# VSS 0.293593f **FLOATING
C47229 a_7765_42852# VSS 0.252651f **FLOATING
C47230 a_7871_42858# VSS 0.503534f **FLOATING
C47231 a_7227_42852# VSS 0.36607f **FLOATING
C47232 a_5755_42852# VSS 0.383967f **FLOATING
C47233 a_5111_42852# VSS 0.354197f **FLOATING
C47234 a_4520_42826# VSS 0.334784f **FLOATING
C47235 a_3935_42891# VSS 0.26911f **FLOATING
C47236 a_3681_42891# VSS 0.301094f **FLOATING
C47237 a_2905_42968# VSS 0.305424f **FLOATING
C47238 a_2075_43172# VSS 0.537699f **FLOATING
C47239 a_1847_42826# VSS 0.670072f **FLOATING
C47240 a_791_42968# VSS 0.335942f **FLOATING
C47241 a_685_42968# VSS 0.220885f **FLOATING
C47242 a_421_43172# VSS 0.006487f **FLOATING
C47243 a_133_43172# VSS 0.00288f **FLOATING
C47244 a_n1533_42852# VSS 0.004694f **FLOATING
C47245 a_n722_43218# VSS 0.001281f **FLOATING
C47246 a_n967_43230# VSS 4.65e-19 **FLOATING
C47247 a_n1379_43218# VSS 0.004992f **FLOATING
C47248 a_n1545_43230# VSS 0.006939f **FLOATING
C47249 a_n1736_43218# VSS 0.073862f **FLOATING
C47250 a_n4318_38680# VSS 1.39087f **FLOATING
C47251 a_n3674_39304# VSS 1.06639f **FLOATING
C47252 a_n13_43084# VSS 0.368998f **FLOATING
C47253 a_n1076_43230# VSS 0.263204f **FLOATING
C47254 a_n901_43156# VSS 0.76245f **FLOATING
C47255 a_n1641_43230# VSS 0.256397f **FLOATING
C47256 a_n1423_42826# VSS 0.1805f **FLOATING
C47257 a_n1991_42858# VSS 0.295941f **FLOATING
C47258 a_n1853_43023# VSS 1.30078f **FLOATING
C47259 a_n2157_42858# VSS 0.556569f **FLOATING
C47260 a_n2472_42826# VSS 0.301801f **FLOATING
C47261 a_n2840_42826# VSS 0.327636f **FLOATING
C47262 a_20749_43396# VSS 0.253248f **FLOATING
C47263 a_17364_32525# VSS 1.89398f **FLOATING
C47264 a_22959_43396# VSS 0.345439f **FLOATING
C47265 a_14209_32519# VSS 2.01016f **FLOATING
C47266 a_22591_43396# VSS 0.335697f **FLOATING
C47267 a_13887_32519# VSS 1.94312f **FLOATING
C47268 a_22223_43396# VSS 0.333609f **FLOATING
C47269 a_5649_42852# VSS 1.95364f **FLOATING
C47270 a_13678_32519# VSS 2.06126f **FLOATING
C47271 a_21855_43396# VSS 0.334538f **FLOATING
C47272 a_4361_42308# VSS 1.30251f **FLOATING
C47273 a_13467_32519# VSS 2.22551f **FLOATING
C47274 a_19095_43396# VSS 0.132304f **FLOATING
C47275 a_21487_43396# VSS 0.293844f **FLOATING
C47276 a_20556_43646# VSS 0.006736f **FLOATING
C47277 a_743_42282# VSS 1.36822f **FLOATING
C47278 a_20301_43646# VSS 0.002477f **FLOATING
C47279 a_4190_30871# VSS 7.379981f **FLOATING
C47280 a_21259_43561# VSS 0.217667f **FLOATING
C47281 a_17678_43396# VSS 0.001281f **FLOATING
C47282 a_17433_43396# VSS 4.65e-19 **FLOATING
C47283 a_16823_43084# VSS 1.23251f **FLOATING
C47284 a_17021_43396# VSS 0.004992f **FLOATING
C47285 a_16855_43396# VSS 0.006939f **FLOATING
C47286 a_15940_43402# VSS 0.003101f **FLOATING
C47287 a_15868_43402# VSS 6.07e-19 **FLOATING
C47288 a_15231_43396# VSS 0.003851f **FLOATING
C47289 a_15125_43396# VSS 0.003584f **FLOATING
C47290 a_15037_43396# VSS 0.001503f **FLOATING
C47291 a_16867_43762# VSS 0.004694f **FLOATING
C47292 a_16664_43396# VSS 0.080001f **FLOATING
C47293 a_19700_43370# VSS 0.335707f **FLOATING
C47294 a_19268_43646# VSS 0.242693f **FLOATING
C47295 a_15743_43084# VSS 1.49489f **FLOATING
C47296 a_18783_43370# VSS 0.360096f **FLOATING
C47297 a_18525_43370# VSS 0.361236f **FLOATING
C47298 a_18429_43548# VSS 0.222219f **FLOATING
C47299 a_17324_43396# VSS 0.258017f **FLOATING
C47300 a_17499_43370# VSS 0.762886f **FLOATING
C47301 a_16759_43396# VSS 0.252915f **FLOATING
C47302 a_16977_43638# VSS 0.178776f **FLOATING
C47303 a_16409_43396# VSS 0.290743f **FLOATING
C47304 a_16547_43609# VSS 0.561468f **FLOATING
C47305 a_16243_43396# VSS 0.562369f **FLOATING
C47306 a_16137_43396# VSS 0.635905f **FLOATING
C47307 a_13943_43396# VSS 0.003344f **FLOATING
C47308 a_13837_43396# VSS 0.003427f **FLOATING
C47309 a_13749_43396# VSS 0.001647f **FLOATING
C47310 a_15781_43660# VSS 0.234761f **FLOATING
C47311 a_15681_43442# VSS 0.20154f **FLOATING
C47312 a_14537_43646# VSS 7.16e-20 **FLOATING
C47313 a_10149_43396# VSS 0.003443f **FLOATING
C47314 a_9885_43396# VSS 0.006177f **FLOATING
C47315 a_8945_43396# VSS 0.002098f **FLOATING
C47316 a_8873_43396# VSS 0.001365f **FLOATING
C47317 a_12281_43396# VSS 0.691406f **FLOATING
C47318 a_10849_43646# VSS 7.16e-20 **FLOATING
C47319 a_10341_43396# VSS 0.796012f **FLOATING
C47320 a_9885_43646# VSS 0.00274f **FLOATING
C47321 a_14955_43396# VSS 0.266041f **FLOATING
C47322 a_15095_43370# VSS 0.436411f **FLOATING
C47323 a_14205_43396# VSS 0.2933f **FLOATING
C47324 a_14358_43442# VSS 0.198188f **FLOATING
C47325 a_14579_43548# VSS 0.293668f **FLOATING
C47326 a_13667_43396# VSS 0.265557f **FLOATING
C47327 a_10695_43548# VSS 0.279385f **FLOATING
C47328 a_9803_43646# VSS 0.371929f **FLOATING
C47329 a_9145_43396# VSS 0.437647f **FLOATING
C47330 a_8423_43396# VSS 0.003573f **FLOATING
C47331 a_8317_43396# VSS 0.003562f **FLOATING
C47332 a_8229_43396# VSS 0.002303f **FLOATING
C47333 a_7466_43396# VSS 0.001281f **FLOATING
C47334 a_7221_43396# VSS 4.65e-19 **FLOATING
C47335 a_8685_43396# VSS 1.0146f **FLOATING
C47336 a_6809_43396# VSS 0.004992f **FLOATING
C47337 a_6643_43396# VSS 0.006939f **FLOATING
C47338 a_5837_43396# VSS 0.001678f **FLOATING
C47339 a_5565_43396# VSS 0.00164f **FLOATING
C47340 a_4181_43396# VSS 0.001635f **FLOATING
C47341 a_3457_43396# VSS 0.379621f **FLOATING
C47342 a_2813_43396# VSS 0.412407f **FLOATING
C47343 a_2437_43396# VSS 0.001678f **FLOATING
C47344 a_6655_43762# VSS 0.004694f **FLOATING
C47345 a_6452_43396# VSS 0.073862f **FLOATING
C47346 a_9396_43370# VSS 0.338475f **FLOATING
C47347 a_8791_43396# VSS 0.235222f **FLOATING
C47348 a_8147_43396# VSS 0.256103f **FLOATING
C47349 a_7112_43396# VSS 0.256956f **FLOATING
C47350 a_7287_43370# VSS 0.754599f **FLOATING
C47351 a_6547_43396# VSS 0.253718f **FLOATING
C47352 a_6765_43638# VSS 0.174622f **FLOATING
C47353 a_6197_43396# VSS 0.290517f **FLOATING
C47354 a_6293_42852# VSS 0.473619f **FLOATING
C47355 a_6031_43396# VSS 0.541083f **FLOATING
C47356 a_1512_43396# VSS 0.003304f **FLOATING
C47357 a_648_43396# VSS 0.231254f **FLOATING
C47358 a_548_43396# VSS 0.009033f **FLOATING
C47359 a_n144_43396# VSS 0.003264f **FLOATING
C47360 a_n998_43396# VSS 0.001266f **FLOATING
C47361 a_n1243_43396# VSS 4.65e-19 **FLOATING
C47362 a_3539_42460# VSS 0.337918f **FLOATING
C47363 a_3626_43646# VSS 1.9807f **FLOATING
C47364 a_3540_43646# VSS 9.9e-19 **FLOATING
C47365 a_2982_43646# VSS 3.25953f **FLOATING
C47366 a_2896_43646# VSS 0.00155f **FLOATING
C47367 a_1987_43646# VSS 6.34e-20 **FLOATING
C47368 a_1891_43646# VSS 1.35e-19 **FLOATING
C47369 a_1427_43646# VSS 0.00568f **FLOATING
C47370 a_n1557_42282# VSS 0.870257f **FLOATING
C47371 a_766_43646# VSS 9.92e-19 **FLOATING
C47372 a_4905_42826# VSS 0.781685f **FLOATING
C47373 a_3080_42308# VSS 5.07255f **FLOATING
C47374 a_4699_43561# VSS 0.267684f **FLOATING
C47375 a_4235_43370# VSS 0.33553f **FLOATING
C47376 a_4093_43548# VSS 0.320586f **FLOATING
C47377 a_1756_43548# VSS 0.322408f **FLOATING
C47378 a_1568_43370# VSS 0.63594f **FLOATING
C47379 a_1049_43396# VSS 0.216408f **FLOATING
C47380 a_1209_43370# VSS 0.281234f **FLOATING
C47381 a_458_43396# VSS 0.252302f **FLOATING
C47382 a_n229_43646# VSS 0.004647f **FLOATING
C47383 a_n1655_43396# VSS 0.004992f **FLOATING
C47384 a_n1821_43396# VSS 0.006939f **FLOATING
C47385 a_n1809_43762# VSS 0.004697f **FLOATING
C47386 a_n2012_43396# VSS 0.073862f **FLOATING
C47387 a_104_43370# VSS 0.297328f **FLOATING
C47388 a_n97_42460# VSS 6.9914f **FLOATING
C47389 a_n447_43370# VSS 0.269574f **FLOATING
C47390 a_n1352_43396# VSS 0.260107f **FLOATING
C47391 a_n1177_43370# VSS 0.478516f **FLOATING
C47392 a_n1917_43396# VSS 0.258245f **FLOATING
C47393 a_n1699_43638# VSS 0.175452f **FLOATING
C47394 a_n2267_43396# VSS 0.297246f **FLOATING
C47395 a_n2129_43609# VSS 1.07965f **FLOATING
C47396 a_n2433_43396# VSS 0.56533f **FLOATING
C47397 a_n4318_39304# VSS 0.959585f **FLOATING
C47398 a_n2840_43370# VSS 0.316787f **FLOATING
C47399 a_17538_32519# VSS 1.88845f **FLOATING
C47400 a_20974_43370# VSS 0.458091f **FLOATING
C47401 a_14401_32519# VSS 2.32323f **FLOATING
C47402 a_21381_43940# VSS 0.358332f **FLOATING
C47403 a_19741_43940# VSS 0.007693f **FLOATING
C47404 a_21205_44306# VSS 0.004143f **FLOATING
C47405 a_18533_43940# VSS 0.00274f **FLOATING
C47406 a_19319_43548# VSS 0.229395f **FLOATING
C47407 a_19808_44306# VSS 0.005362f **FLOATING
C47408 a_18797_44260# VSS 0.002999f **FLOATING
C47409 a_18533_44260# VSS 0.007531f **FLOATING
C47410 a_15037_43940# VSS 0.00274f **FLOATING
C47411 a_13565_43940# VSS 0.00274f **FLOATING
C47412 a_9801_43940# VSS 0.006211f **FLOATING
C47413 a_9165_43940# VSS 0.001166f **FLOATING
C47414 a_7499_43940# VSS 0.004678f **FLOATING
C47415 a_6671_43940# VSS 0.004647f **FLOATING
C47416 a_5829_43940# VSS 0.001102f **FLOATING
C47417 a_5745_43940# VSS 7.11e-19 **FLOATING
C47418 a_5326_44056# VSS 9.13e-22 **FLOATING
C47419 a_3737_43940# VSS 0.001166f **FLOATING
C47420 a_3052_44056# VSS 9.13e-22 **FLOATING
C47421 a_2455_43940# VSS 7.44e-19 **FLOATING
C47422 a_2253_43940# VSS 0.001314f **FLOATING
C47423 a_1443_43940# VSS 8.96e-19 **FLOATING
C47424 a_1241_43940# VSS 0.001786f **FLOATING
C47425 a_726_44056# VSS 4.62e-19 **FLOATING
C47426 a_15301_44260# VSS 0.00288f **FLOATING
C47427 a_15037_44260# VSS 0.006076f **FLOATING
C47428 a_14761_44260# VSS 0.001738f **FLOATING
C47429 a_14485_44260# VSS 0.001738f **FLOATING
C47430 a_14021_43940# VSS 0.387813f **FLOATING
C47431 a_13829_44260# VSS 0.003443f **FLOATING
C47432 a_13565_44260# VSS 0.005972f **FLOATING
C47433 a_12710_44260# VSS 0.003489f **FLOATING
C47434 a_12603_44260# VSS 0.004224f **FLOATING
C47435 a_12495_44260# VSS 0.003836f **FLOATING
C47436 a_11816_44260# VSS 0.00475f **FLOATING
C47437 a_11173_44260# VSS 0.219946f **FLOATING
C47438 a_10555_44260# VSS 0.346315f **FLOATING
C47439 a_9895_44260# VSS 0.0063f **FLOATING
C47440 a_9801_44260# VSS 0.006656f **FLOATING
C47441 a_9248_44260# VSS 0.003866f **FLOATING
C47442 a_22959_43948# VSS 0.341565f **FLOATING
C47443 a_15493_43940# VSS 0.460801f **FLOATING
C47444 a_22223_43948# VSS 0.31992f **FLOATING
C47445 a_11341_43940# VSS 0.365183f **FLOATING
C47446 a_21115_43940# VSS 0.204633f **FLOATING
C47447 a_20935_43940# VSS 0.222887f **FLOATING
C47448 a_20623_43914# VSS 0.371294f **FLOATING
C47449 a_20365_43914# VSS 0.359455f **FLOATING
C47450 a_20269_44172# VSS 0.225063f **FLOATING
C47451 a_19862_44208# VSS 0.562087f **FLOATING
C47452 a_19478_44306# VSS 0.278384f **FLOATING
C47453 a_15493_43396# VSS 0.277875f **FLOATING
C47454 a_19328_44172# VSS 0.2031f **FLOATING
C47455 a_18451_43940# VSS 0.377396f **FLOATING
C47456 a_18326_43940# VSS 0.276559f **FLOATING
C47457 a_18079_43940# VSS 0.21121f **FLOATING
C47458 a_17973_43940# VSS 0.359917f **FLOATING
C47459 a_17737_43940# VSS 0.386318f **FLOATING
C47460 a_15682_43940# VSS 1.9643f **FLOATING
C47461 a_14955_43940# VSS 0.365393f **FLOATING
C47462 a_13483_43940# VSS 0.376442f **FLOATING
C47463 a_12429_44172# VSS 0.389129f **FLOATING
C47464 a_11750_44172# VSS 0.221782f **FLOATING
C47465 a_10807_43548# VSS 0.451031f **FLOATING
C47466 a_10949_43914# VSS 0.257331f **FLOATING
C47467 a_10729_43914# VSS 0.34307f **FLOATING
C47468 a_10405_44172# VSS 0.142993f **FLOATING
C47469 a_9672_43914# VSS 0.323006f **FLOATING
C47470 a_9028_43914# VSS 0.398016f **FLOATING
C47471 a_8333_44056# VSS 0.331632f **FLOATING
C47472 a_8018_44260# VSS 0.005204f **FLOATING
C47473 a_7911_44260# VSS 0.006364f **FLOATING
C47474 a_7584_44260# VSS 0.003279f **FLOATING
C47475 a_6756_44260# VSS 0.003243f **FLOATING
C47476 a_n2661_42282# VSS 1.51789f **FLOATING
C47477 a_6101_44260# VSS 0.001611f **FLOATING
C47478 a_5841_44260# VSS 0.001326f **FLOATING
C47479 a_3820_44260# VSS 0.004263f **FLOATING
C47480 a_3499_42826# VSS 0.380221f **FLOATING
C47481 a_2537_44260# VSS 0.001558f **FLOATING
C47482 a_2253_44260# VSS 0.002472f **FLOATING
C47483 a_1525_44260# VSS 0.001638f **FLOATING
C47484 a_1241_44260# VSS 0.001824f **FLOATING
C47485 a_261_44278# VSS 0.003386f **FLOATING
C47486 a_n1441_43940# VSS 0.004694f **FLOATING
C47487 a_n630_44306# VSS 0.002229f **FLOATING
C47488 a_n875_44318# VSS 9.68e-19 **FLOATING
C47489 a_n1287_44306# VSS 0.00579f **FLOATING
C47490 a_n1453_44318# VSS 0.008634f **FLOATING
C47491 a_n1644_44306# VSS 0.080042f **FLOATING
C47492 a_n3674_39768# VSS 0.890487f **FLOATING
C47493 a_n4318_39768# VSS 1.09976f **FLOATING
C47494 a_7845_44172# VSS 0.239173f **FLOATING
C47495 a_7542_44172# VSS 0.283767f **FLOATING
C47496 a_7281_43914# VSS 0.271121f **FLOATING
C47497 a_6453_43914# VSS 0.26639f **FLOATING
C47498 a_5663_43940# VSS 0.488325f **FLOATING
C47499 a_5495_43940# VSS 0.212229f **FLOATING
C47500 a_5013_44260# VSS 0.279924f **FLOATING
C47501 a_5244_44056# VSS 0.216368f **FLOATING
C47502 a_3905_42865# VSS 0.9893f **FLOATING
C47503 a_3600_43914# VSS 0.422049f **FLOATING
C47504 a_2998_44172# VSS 0.503048f **FLOATING
C47505 a_2889_44172# VSS 0.217034f **FLOATING
C47506 a_2675_43914# VSS 0.2974f **FLOATING
C47507 a_895_43940# VSS 0.237723f **FLOATING
C47508 a_2479_44172# VSS 0.817462f **FLOATING
C47509 a_2127_44172# VSS 0.517911f **FLOATING
C47510 a_453_43940# VSS 0.285192f **FLOATING
C47511 a_1414_42308# VSS 1.07452f **FLOATING
C47512 a_1467_44172# VSS 0.187431f **FLOATING
C47513 a_1115_44172# VSS 0.52592f **FLOATING
C47514 a_644_44056# VSS 0.227493f **FLOATING
C47515 a_175_44278# VSS 0.226801f **FLOATING
C47516 a_n984_44318# VSS 0.27358f **FLOATING
C47517 a_n809_44244# VSS 0.785904f **FLOATING
C47518 a_n1549_44318# VSS 0.264547f **FLOATING
C47519 a_n1331_43914# VSS 0.185087f **FLOATING
C47520 a_n1899_43946# VSS 0.299008f **FLOATING
C47521 a_n1761_44111# VSS 0.392075f **FLOATING
C47522 a_n2065_43946# VSS 0.658803f **FLOATING
C47523 a_n2472_43914# VSS 0.3103f **FLOATING
C47524 a_n2840_43914# VSS 0.345355f **FLOATING
C47525 a_19237_31679# VSS 1.49314f **FLOATING
C47526 a_22959_44484# VSS 0.343897f **FLOATING
C47527 a_17730_32519# VSS 2.45467f **FLOATING
C47528 a_22591_44484# VSS 0.315361f **FLOATING
C47529 a_22485_44484# VSS 0.590119f **FLOATING
C47530 a_20512_43084# VSS 0.561552f **FLOATING
C47531 a_21145_44484# VSS 0.006939f **FLOATING
C47532 a_21073_44484# VSS 0.004992f **FLOATING
C47533 a_20637_44484# VSS 4.65e-19 **FLOATING
C47534 a_20397_44484# VSS 0.001266f **FLOATING
C47535 a_22315_44484# VSS 0.238239f **FLOATING
C47536 a_3422_30871# VSS 9.021831f **FLOATING
C47537 a_21398_44850# VSS 0.073862f **FLOATING
C47538 a_20980_44850# VSS 0.004694f **FLOATING
C47539 a_19789_44512# VSS 0.003386f **FLOATING
C47540 a_18753_44484# VSS 0.006939f **FLOATING
C47541 a_18681_44484# VSS 0.004992f **FLOATING
C47542 a_18579_44172# VSS 0.812679f **FLOATING
C47543 a_18245_44484# VSS 4.65e-19 **FLOATING
C47544 a_18005_44484# VSS 0.001266f **FLOATING
C47545 a_19279_43940# VSS 1.69633f **FLOATING
C47546 a_20766_44850# VSS 0.177656f **FLOATING
C47547 a_20835_44721# VSS 0.260406f **FLOATING
C47548 a_20679_44626# VSS 0.58931f **FLOATING
C47549 a_20640_44752# VSS 0.296084f **FLOATING
C47550 a_20362_44736# VSS 0.255907f **FLOATING
C47551 a_20159_44458# VSS 0.483669f **FLOATING
C47552 a_19615_44636# VSS 0.238459f **FLOATING
C47553 a_11967_42832# VSS 6.11191f **FLOATING
C47554 a_19006_44850# VSS 0.073862f **FLOATING
C47555 a_18588_44850# VSS 0.004694f **FLOATING
C47556 a_17325_44484# VSS 0.002122f **FLOATING
C47557 a_17061_44484# VSS 0.006177f **FLOATING
C47558 a_16789_44484# VSS 0.002002f **FLOATING
C47559 a_16335_44484# VSS 0.005048f **FLOATING
C47560 a_16241_44484# VSS 0.005441f **FLOATING
C47561 a_15367_44484# VSS 0.002898f **FLOATING
C47562 a_15146_44484# VSS 0.002399f **FLOATING
C47563 a_17517_44484# VSS 0.244051f **FLOATING
C47564 a_17061_44734# VSS 0.00274f **FLOATING
C47565 a_16241_44734# VSS 0.006211f **FLOATING
C47566 a_14673_44172# VSS 0.290001f **FLOATING
C47567 a_14581_44484# VSS 0.001661f **FLOATING
C47568 a_13940_44484# VSS 0.004195f **FLOATING
C47569 a_13296_44484# VSS 0.005047f **FLOATING
C47570 a_12829_44484# VSS 0.001944f **FLOATING
C47571 a_12553_44484# VSS 0.00193f **FLOATING
C47572 a_12189_44484# VSS 0.001627f **FLOATING
C47573 a_11909_44484# VSS 0.001659f **FLOATING
C47574 a_11541_44484# VSS 0.139071f **FLOATING
C47575 a_10809_44484# VSS 0.001938f **FLOATING
C47576 a_15463_44811# VSS 2.7e-19 **FLOATING
C47577 a_15433_44458# VSS 0.301508f **FLOATING
C47578 a_14815_43914# VSS 0.445698f **FLOATING
C47579 a_13857_44734# VSS 0.001166f **FLOATING
C47580 a_13213_44734# VSS 0.001208f **FLOATING
C47581 a_n2293_43922# VSS 3.31971f **FLOATING
C47582 a_n2661_43922# VSS 1.51991f **FLOATING
C47583 a_n2661_42834# VSS 1.20196f **FLOATING
C47584 a_9159_44484# VSS 0.158168f **FLOATING
C47585 a_10617_44484# VSS 0.119149f **FLOATING
C47586 a_5708_44484# VSS 0.231649f **FLOATING
C47587 a_5608_44484# VSS 0.007818f **FLOATING
C47588 a_3363_44484# VSS 0.27629f **FLOATING
C47589 a_556_44484# VSS 0.201935f **FLOATING
C47590 a_484_44484# VSS 0.004815f **FLOATING
C47591 a_n89_44484# VSS 0.002857f **FLOATING
C47592 a_n310_44484# VSS 0.002596f **FLOATING
C47593 a_9313_44734# VSS 1.31461f **FLOATING
C47594 a_5891_43370# VSS 2.82295f **FLOATING
C47595 a_8375_44464# VSS 0.211867f **FLOATING
C47596 a_7640_43914# VSS 0.542377f **FLOATING
C47597 a_6109_44484# VSS 0.648821f **FLOATING
C47598 a_700_44734# VSS 0.001076f **FLOATING
C47599 a_n998_44484# VSS 0.002215f **FLOATING
C47600 a_n1243_44484# VSS 9.68e-19 **FLOATING
C47601 a_7_44811# VSS 2.7e-19 **FLOATING
C47602 a_n23_44458# VSS 0.278255f **FLOATING
C47603 a_n356_44636# VSS 2.91333f **FLOATING
C47604 a_n1655_44484# VSS 0.00579f **FLOATING
C47605 a_n1821_44484# VSS 0.008634f **FLOATING
C47606 a_n1809_44850# VSS 0.007269f **FLOATING
C47607 a_n2012_44484# VSS 0.080001f **FLOATING
C47608 a_18989_43940# VSS 0.423174f **FLOATING
C47609 a_18374_44850# VSS 0.179731f **FLOATING
C47610 a_18443_44721# VSS 0.253971f **FLOATING
C47611 a_18287_44626# VSS 0.507939f **FLOATING
C47612 a_18248_44752# VSS 0.294917f **FLOATING
C47613 a_17970_44736# VSS 0.26161f **FLOATING
C47614 a_17767_44458# VSS 0.474097f **FLOATING
C47615 a_16979_44734# VSS 0.363013f **FLOATING
C47616 a_14539_43914# VSS 1.18088f **FLOATING
C47617 a_16112_44458# VSS 0.326339f **FLOATING
C47618 a_15004_44636# VSS 0.254778f **FLOATING
C47619 a_13720_44458# VSS 0.403209f **FLOATING
C47620 a_13076_44458# VSS 0.38829f **FLOATING
C47621 a_12883_44458# VSS 0.287544f **FLOATING
C47622 a_12607_44458# VSS 0.499331f **FLOATING
C47623 a_8975_43940# VSS 0.652857f **FLOATING
C47624 a_10057_43914# VSS 0.654189f **FLOATING
C47625 a_10440_44484# VSS 0.210149f **FLOATING
C47626 a_10334_44484# VSS 0.210217f **FLOATING
C47627 a_10157_44484# VSS 0.208916f **FLOATING
C47628 a_9838_44484# VSS 0.276258f **FLOATING
C47629 a_5883_43914# VSS 0.792825f **FLOATING
C47630 a_8701_44490# VSS 0.358059f **FLOATING
C47631 a_8103_44636# VSS 0.340824f **FLOATING
C47632 a_6298_44484# VSS 1.93814f **FLOATING
C47633 a_5518_44484# VSS 0.242995f **FLOATING
C47634 a_5343_44458# VSS 1.28071f **FLOATING
C47635 a_4743_44484# VSS 0.327178f **FLOATING
C47636 a_n699_43396# VSS 1.82142f **FLOATING
C47637 a_4223_44672# VSS 0.659279f **FLOATING
C47638 a_2779_44458# VSS 0.532137f **FLOATING
C47639 a_949_44458# VSS 1.97734f **FLOATING
C47640 a_742_44458# VSS 1.02263f **FLOATING
C47641 a_n452_44636# VSS 0.254732f **FLOATING
C47642 a_n1352_44484# VSS 0.269853f **FLOATING
C47643 a_n1177_44458# VSS 0.493891f **FLOATING
C47644 a_n1917_44484# VSS 0.280038f **FLOATING
C47645 a_n1699_44726# VSS 0.197478f **FLOATING
C47646 a_n2267_44484# VSS 0.308908f **FLOATING
C47647 a_n2129_44697# VSS 0.307327f **FLOATING
C47648 a_n2433_44484# VSS 0.679598f **FLOATING
C47649 a_n2661_44458# VSS 0.487677f **FLOATING
C47650 a_n4318_40392# VSS 0.995833f **FLOATING
C47651 a_n2840_44458# VSS 0.316322f **FLOATING
C47652 a_19721_31679# VSS 1.6201f **FLOATING
C47653 a_18114_32519# VSS 3.11255f **FLOATING
C47654 a_17801_45144# VSS 8.35e-20 **FLOATING
C47655 a_16237_45028# VSS 0.017944f **FLOATING
C47656 a_20193_45348# VSS 1.70015f **FLOATING
C47657 a_11691_44458# VSS 1.78467f **FLOATING
C47658 a_19113_45348# VSS 0.367248f **FLOATING
C47659 a_22959_45036# VSS 0.345334f **FLOATING
C47660 a_22223_45036# VSS 0.354178f **FLOATING
C47661 a_11827_44484# VSS 1.28091f **FLOATING
C47662 a_21359_45002# VSS 0.397791f **FLOATING
C47663 a_21101_45002# VSS 0.35202f **FLOATING
C47664 a_21005_45260# VSS 0.212992f **FLOATING
C47665 a_20567_45036# VSS 0.31908f **FLOATING
C47666 a_18494_42460# VSS 1.15626f **FLOATING
C47667 a_18184_42460# VSS 0.838573f **FLOATING
C47668 a_19778_44110# VSS 0.599421f **FLOATING
C47669 a_18911_45144# VSS 0.307008f **FLOATING
C47670 a_18587_45118# VSS 0.214925f **FLOATING
C47671 a_18315_45260# VSS 0.334834f **FLOATING
C47672 a_17719_45144# VSS 0.331229f **FLOATING
C47673 a_17613_45144# VSS 0.244364f **FLOATING
C47674 a_17023_45118# VSS 0.20885f **FLOATING
C47675 a_16922_45042# VSS 0.818675f **FLOATING
C47676 a_16501_45348# VSS 0.005461f **FLOATING
C47677 a_16405_45348# VSS 0.003038f **FLOATING
C47678 a_16321_45348# VSS 0.002956f **FLOATING
C47679 a_14309_45028# VSS 0.006587f **FLOATING
C47680 a_13807_45067# VSS 2.7e-19 **FLOATING
C47681 a_15685_45394# VSS 0.003883f **FLOATING
C47682 a_15060_45348# VSS 0.006388f **FLOATING
C47683 a_14976_45348# VSS 0.005191f **FLOATING
C47684 a_14403_45348# VSS 0.006612f **FLOATING
C47685 a_14309_45348# VSS 0.006958f **FLOATING
C47686 a_13711_45394# VSS 0.002898f **FLOATING
C47687 a_13490_45394# VSS 0.002596f **FLOATING
C47688 a_13105_45348# VSS 0.001738f **FLOATING
C47689 a_11915_45394# VSS 0.004143f **FLOATING
C47690 a_n2661_43370# VSS 0.820606f **FLOATING
C47691 a_11361_45348# VSS 0.001666f **FLOATING
C47692 a_7735_45067# VSS 2.7e-19 **FLOATING
C47693 a_10903_45394# VSS 0.004143f **FLOATING
C47694 a_8560_45348# VSS 0.185033f **FLOATING
C47695 a_8488_45348# VSS 0.003218f **FLOATING
C47696 a_8137_45348# VSS 0.001684f **FLOATING
C47697 a_n2293_42834# VSS 1.1151f **FLOATING
C47698 a_7639_45394# VSS 0.002898f **FLOATING
C47699 a_7418_45394# VSS 0.002596f **FLOATING
C47700 a_6945_45348# VSS 0.001738f **FLOATING
C47701 a_5837_45028# VSS 0.00274f **FLOATING
C47702 a_5093_45028# VSS 0.001102f **FLOATING
C47703 a_5009_45028# VSS 7.39e-19 **FLOATING
C47704 a_2809_45028# VSS 0.00638f **FLOATING
C47705 a_2448_45028# VSS 1.19e-20 **FLOATING
C47706 a_6517_45366# VSS 0.003386f **FLOATING
C47707 a_6125_45348# VSS 0.007531f **FLOATING
C47708 a_5837_45348# VSS 0.002999f **FLOATING
C47709 a_5365_45348# VSS 0.002387f **FLOATING
C47710 a_5105_45348# VSS 0.001558f **FLOATING
C47711 a_4640_45348# VSS 0.006141f **FLOATING
C47712 a_4185_45348# VSS 0.001865f **FLOATING
C47713 a_3602_45348# VSS 0.005184f **FLOATING
C47714 a_3495_45348# VSS 0.006372f **FLOATING
C47715 a_2903_45348# VSS 0.005166f **FLOATING
C47716 a_2809_45348# VSS 0.006958f **FLOATING
C47717 a_2304_45348# VSS 0.182367f **FLOATING
C47718 a_2232_45348# VSS 0.004649f **FLOATING
C47719 a_1423_45028# VSS 0.980773f **FLOATING
C47720 a_1145_45348# VSS 0.001816f **FLOATING
C47721 a_626_44172# VSS 0.67926f **FLOATING
C47722 a_501_45348# VSS 0.001778f **FLOATING
C47723 a_375_42282# VSS 0.447027f **FLOATING
C47724 a_16751_45260# VSS 0.316547f **FLOATING
C47725 a_1307_43914# VSS 2.30311f **FLOATING
C47726 a_16019_45002# VSS 0.25377f **FLOATING
C47727 a_15595_45028# VSS 0.214111f **FLOATING
C47728 a_15415_45028# VSS 0.221991f **FLOATING
C47729 a_14797_45144# VSS 0.249222f **FLOATING
C47730 a_14537_43396# VSS 1.73146f **FLOATING
C47731 a_14180_45002# VSS 0.327485f **FLOATING
C47732 a_13777_45326# VSS 0.272936f **FLOATING
C47733 a_13556_45296# VSS 1.01916f **FLOATING
C47734 a_9482_43914# VSS 3.42654f **FLOATING
C47735 a_13348_45260# VSS 0.243533f **FLOATING
C47736 a_13159_45002# VSS 0.265737f **FLOATING
C47737 a_13017_45260# VSS 0.362048f **FLOATING
C47738 a_11963_45334# VSS 0.226884f **FLOATING
C47739 a_11787_45002# VSS 0.212512f **FLOATING
C47740 a_10951_45334# VSS 0.228638f **FLOATING
C47741 a_10775_45002# VSS 0.204487f **FLOATING
C47742 a_8953_45002# VSS 1.94941f **FLOATING
C47743 a_8191_45002# VSS 0.325964f **FLOATING
C47744 a_7705_45326# VSS 0.273009f **FLOATING
C47745 a_6709_45028# VSS 0.354418f **FLOATING
C47746 a_7229_43940# VSS 0.786182f **FLOATING
C47747 a_7276_45260# VSS 0.251523f **FLOATING
C47748 a_5205_44484# VSS 0.546179f **FLOATING
C47749 a_6431_45366# VSS 0.233718f **FLOATING
C47750 a_6171_45002# VSS 0.700605f **FLOATING
C47751 a_3232_43370# VSS 2.99721f **FLOATING
C47752 a_5691_45260# VSS 0.370273f **FLOATING
C47753 a_4927_45028# VSS 0.520892f **FLOATING
C47754 a_5111_44636# VSS 3.44603f **FLOATING
C47755 a_5147_45002# VSS 0.803306f **FLOATING
C47756 a_4558_45348# VSS 0.446148f **FLOATING
C47757 a_4574_45260# VSS 0.208274f **FLOATING
C47758 a_3537_45260# VSS 2.45782f **FLOATING
C47759 a_3429_45260# VSS 0.274034f **FLOATING
C47760 a_3065_45002# VSS 0.864786f **FLOATING
C47761 a_2680_45002# VSS 0.321351f **FLOATING
C47762 a_2382_45260# VSS 1.03422f **FLOATING
C47763 a_2274_45254# VSS 0.187307f **FLOATING
C47764 a_1667_45002# VSS 0.345429f **FLOATING
C47765 a_327_44734# VSS 0.419171f **FLOATING
C47766 a_413_45260# VSS 4.87522f **FLOATING
C47767 a_n37_45144# VSS 0.321746f **FLOATING
C47768 a_n143_45144# VSS 0.209896f **FLOATING
C47769 a_n467_45028# VSS 0.311181f **FLOATING
C47770 a_n659_45366# VSS 0.004685f **FLOATING
C47771 a_n967_45348# VSS 0.453992f **FLOATING
C47772 en_comp VSS 7.869411f **FLOATING
C47773 a_n2956_37592# VSS 2.90302f **FLOATING
C47774 a_n2810_45028# VSS 1.52635f **FLOATING
C47775 a_n745_45366# VSS 0.257282f **FLOATING
C47776 a_n913_45002# VSS 5.04726f **FLOATING
C47777 a_n1059_45260# VSS 2.30619f **FLOATING
C47778 a_n2017_45002# VSS 1.09013f **FLOATING
C47779 a_n2109_45247# VSS 0.252392f **FLOATING
C47780 a_n2293_45010# VSS 0.614925f **FLOATING
C47781 a_n2472_45002# VSS 0.298945f **FLOATING
C47782 a_n2661_45010# VSS 0.839496f **FLOATING
C47783 a_n2840_45002# VSS 0.340687f **FLOATING
C47784 a_21542_45572# VSS 0.002215f **FLOATING
C47785 a_21297_45572# VSS 9.68e-19 **FLOATING
C47786 a_20447_31679# VSS 1.49316f **FLOATING
C47787 a_22959_45572# VSS 0.34535f **FLOATING
C47788 a_19963_31679# VSS 1.43962f **FLOATING
C47789 a_22591_45572# VSS 0.363695f **FLOATING
C47790 a_3357_43084# VSS 2.42707f **FLOATING
C47791 a_19479_31679# VSS 1.67418f **FLOATING
C47792 a_22223_45572# VSS 0.334964f **FLOATING
C47793 a_2437_43646# VSS 6.25635f **FLOATING
C47794 a_21513_45002# VSS 0.669089f **FLOATING
C47795 a_20885_45572# VSS 0.004992f **FLOATING
C47796 a_20719_45572# VSS 0.006939f **FLOATING
C47797 a_19610_45572# VSS 0.002215f **FLOATING
C47798 a_19365_45572# VSS 4.65e-19 **FLOATING
C47799 a_20731_45938# VSS 0.004694f **FLOATING
C47800 a_20528_45572# VSS 0.073082f **FLOATING
C47801 a_21188_45572# VSS 0.284872f **FLOATING
C47802 a_21363_45546# VSS 0.515994f **FLOATING
C47803 a_20623_45572# VSS 0.256236f **FLOATING
C47804 a_20841_45814# VSS 0.180037f **FLOATING
C47805 a_20273_45572# VSS 0.288513f **FLOATING
C47806 a_20107_45572# VSS 0.541125f **FLOATING
C47807 a_18953_45572# VSS 0.004992f **FLOATING
C47808 a_18787_45572# VSS 0.006939f **FLOATING
C47809 a_17668_45572# VSS 0.217142f **FLOATING
C47810 a_17568_45572# VSS 0.005817f **FLOATING
C47811 a_17034_45572# VSS 0.001266f **FLOATING
C47812 a_16789_45572# VSS 4.65e-19 **FLOATING
C47813 a_18799_45938# VSS 0.004694f **FLOATING
C47814 a_18596_45572# VSS 0.073862f **FLOATING
C47815 a_19256_45572# VSS 0.257674f **FLOATING
C47816 a_19431_45546# VSS 0.487121f **FLOATING
C47817 a_18691_45572# VSS 0.255356f **FLOATING
C47818 a_18909_45814# VSS 0.178658f **FLOATING
C47819 a_18341_45572# VSS 0.291608f **FLOATING
C47820 a_18479_45785# VSS 1.15946f **FLOATING
C47821 a_18175_45572# VSS 0.516981f **FLOATING
C47822 a_16147_45260# VSS 0.506229f **FLOATING
C47823 a_16377_45572# VSS 0.004992f **FLOATING
C47824 a_16211_45572# VSS 0.006939f **FLOATING
C47825 a_14127_45572# VSS 0.006612f **FLOATING
C47826 a_14033_45572# VSS 0.006958f **FLOATING
C47827 a_13485_45572# VSS 0.001696f **FLOATING
C47828 a_13385_45572# VSS 0.004208f **FLOATING
C47829 a_13297_45572# VSS 0.004404f **FLOATING
C47830 a_12749_45572# VSS 0.00153f **FLOATING
C47831 a_12649_45572# VSS 0.005051f **FLOATING
C47832 a_12561_45572# VSS 0.005505f **FLOATING
C47833 a_16223_45938# VSS 0.004694f **FLOATING
C47834 a_16020_45572# VSS 0.073862f **FLOATING
C47835 a_17478_45572# VSS 0.232341f **FLOATING
C47836 a_15861_45028# VSS 0.449058f **FLOATING
C47837 a_8696_44636# VSS 0.917254f **FLOATING
C47838 a_16680_45572# VSS 0.258674f **FLOATING
C47839 a_16855_45546# VSS 0.471485f **FLOATING
C47840 a_16115_45572# VSS 0.253972f **FLOATING
C47841 a_16333_45814# VSS 0.178165f **FLOATING
C47842 a_15765_45572# VSS 0.291326f **FLOATING
C47843 a_15903_45785# VSS 0.4164f **FLOATING
C47844 a_15599_45572# VSS 0.50233f **FLOATING
C47845 a_15037_45618# VSS 0.209713f **FLOATING
C47846 a_14033_45822# VSS 0.006541f **FLOATING
C47847 a_12016_45572# VSS 0.005248f **FLOATING
C47848 a_11778_45572# VSS 0.003039f **FLOATING
C47849 a_11688_45572# VSS 0.002091f **FLOATING
C47850 a_11136_45572# VSS 0.17156f **FLOATING
C47851 a_11064_45572# VSS 0.003188f **FLOATING
C47852 a_10544_45572# VSS 0.006484f **FLOATING
C47853 a_10306_45572# VSS 0.004928f **FLOATING
C47854 a_10216_45572# VSS 0.003935f **FLOATING
C47855 a_9159_45572# VSS 0.151638f **FLOATING
C47856 a_8791_45572# VSS 0.00583f **FLOATING
C47857 a_8697_45572# VSS 0.005152f **FLOATING
C47858 a_8192_45572# VSS 0.17002f **FLOATING
C47859 a_8120_45572# VSS 0.004768f **FLOATING
C47860 a_11682_45822# VSS 0.010374f **FLOATING
C47861 a_10907_45822# VSS 0.547001f **FLOATING
C47862 a_10210_45822# VSS 0.012573f **FLOATING
C47863 a_8697_45822# VSS 0.006221f **FLOATING
C47864 a_6977_45572# VSS 0.008634f **FLOATING
C47865 a_6905_45572# VSS 0.00579f **FLOATING
C47866 a_6469_45572# VSS 9.68e-19 **FLOATING
C47867 a_6229_45572# VSS 0.002215f **FLOATING
C47868 a_15143_45578# VSS 0.315994f **FLOATING
C47869 a_14495_45572# VSS 0.325874f **FLOATING
C47870 a_13249_42308# VSS 1.08648f **FLOATING
C47871 a_13904_45546# VSS 0.327907f **FLOATING
C47872 a_13527_45546# VSS 0.245514f **FLOATING
C47873 a_13163_45724# VSS 0.180841f **FLOATING
C47874 a_12791_45546# VSS 0.237787f **FLOATING
C47875 a_11823_42460# VSS 2.45644f **FLOATING
C47876 a_12427_45724# VSS 0.190531f **FLOATING
C47877 a_11962_45724# VSS 0.218739f **FLOATING
C47878 a_11652_45724# VSS 0.258015f **FLOATING
C47879 a_11525_45546# VSS 0.346102f **FLOATING
C47880 a_11322_45546# VSS 0.62914f **FLOATING
C47881 a_10490_45724# VSS 0.972668f **FLOATING
C47882 a_8746_45002# VSS 0.547616f **FLOATING
C47883 a_10193_42453# VSS 3.59848f **FLOATING
C47884 a_10180_45724# VSS 0.281135f **FLOATING
C47885 a_10053_45546# VSS 0.373668f **FLOATING
C47886 a_9049_44484# VSS 0.249658f **FLOATING
C47887 a_7499_43078# VSS 3.22587f **FLOATING
C47888 a_8568_45546# VSS 0.317032f **FLOATING
C47889 a_8162_45546# VSS 0.376225f **FLOATING
C47890 a_7230_45938# VSS 0.078992f **FLOATING
C47891 a_6812_45938# VSS 0.004694f **FLOATING
C47892 a_5437_45600# VSS 0.004685f **FLOATING
C47893 a_4880_45572# VSS 0.182839f **FLOATING
C47894 a_4808_45572# VSS 0.004805f **FLOATING
C47895 a_5024_45822# VSS 2.99e-19 **FLOATING
C47896 a_3260_45572# VSS 0.003272f **FLOATING
C47897 a_2211_45572# VSS 0.002983f **FLOATING
C47898 a_1990_45572# VSS 0.00263f **FLOATING
C47899 a_3775_45552# VSS 0.209244f **FLOATING
C47900 a_7227_45028# VSS 0.439395f **FLOATING
C47901 a_6598_45938# VSS 0.185967f **FLOATING
C47902 a_6667_45809# VSS 0.264656f **FLOATING
C47903 a_6511_45714# VSS 0.647716f **FLOATING
C47904 a_6472_45840# VSS 0.310105f **FLOATING
C47905 a_6194_45824# VSS 0.2717f **FLOATING
C47906 a_5907_45546# VSS 0.592148f **FLOATING
C47907 a_5263_45724# VSS 0.250928f **FLOATING
C47908 a_4099_45572# VSS 0.33915f **FLOATING
C47909 a_3175_45822# VSS 0.004647f **FLOATING
C47910 a_2711_45572# VSS 1.77517f **FLOATING
C47911 a_1609_45572# VSS 0.001977f **FLOATING
C47912 a_1260_45572# VSS 0.006784f **FLOATING
C47913 a_1176_45572# VSS 0.005484f **FLOATING
C47914 a_603_45572# VSS 0.008207f **FLOATING
C47915 a_509_45572# VSS 0.005519f **FLOATING
C47916 a_n89_45572# VSS 0.003313f **FLOATING
C47917 a_n310_45572# VSS 0.002596f **FLOATING
C47918 a_2307_45899# VSS 3.38e-19 **FLOATING
C47919 a_1990_45899# VSS 1.9e-19 **FLOATING
C47920 a_2277_45546# VSS 0.303704f **FLOATING
C47921 a_1609_45822# VSS 0.5528f **FLOATING
C47922 a_n443_42852# VSS 4.64762f **FLOATING
C47923 a_509_45822# VSS 0.010571f **FLOATING
C47924 a_n906_45572# VSS 0.006201f **FLOATING
C47925 a_n1013_45572# VSS 0.008252f **FLOATING
C47926 a_7_45899# VSS 2.7e-19 **FLOATING
C47927 a_n23_45546# VSS 0.281189f **FLOATING
C47928 a_n356_45724# VSS 0.32306f **FLOATING
C47929 a_3503_45724# VSS 0.322319f **FLOATING
C47930 a_3316_45546# VSS 0.336134f **FLOATING
C47931 a_3218_45724# VSS 0.379893f **FLOATING
C47932 a_2957_45546# VSS 0.276358f **FLOATING
C47933 a_1848_45724# VSS 0.245258f **FLOATING
C47934 a_997_45618# VSS 0.248122f **FLOATING
C47935 a_n755_45592# VSS 5.8889f **FLOATING
C47936 a_n357_42282# VSS 2.46134f **FLOATING
C47937 a_310_45028# VSS 0.207165f **FLOATING
C47938 a_n1099_45572# VSS 0.339525f **FLOATING
C47939 a_380_45546# VSS 0.337145f **FLOATING
C47940 a_n452_45724# VSS 0.253614f **FLOATING
C47941 a_n863_45724# VSS 3.49288f **FLOATING
C47942 a_n1079_45724# VSS 0.289271f **FLOATING
C47943 a_n2293_45546# VSS 0.879703f **FLOATING
C47944 a_n2956_38216# VSS 1.49846f **FLOATING
C47945 a_n2472_45546# VSS 0.340801f **FLOATING
C47946 a_n2661_45546# VSS 1.58481f **FLOATING
C47947 a_n2810_45572# VSS 1.43198f **FLOATING
C47948 a_n2840_45546# VSS 0.344757f **FLOATING
C47949 a_21167_46155# VSS 2.7e-19 **FLOATING
C47950 a_20692_30879# VSS 1.61586f **FLOATING
C47951 a_20205_31679# VSS 1.45878f **FLOATING
C47952 a_21071_46482# VSS 0.003313f **FLOATING
C47953 a_20850_46482# VSS 0.003279f **FLOATING
C47954 a_19443_46116# VSS 0.004694f **FLOATING
C47955 a_20254_46482# VSS 0.001266f **FLOATING
C47956 a_20009_46494# VSS 4.65e-19 **FLOATING
C47957 a_19597_46482# VSS 0.004992f **FLOATING
C47958 a_18051_46116# VSS 0.006211f **FLOATING
C47959 a_19431_46494# VSS 0.006939f **FLOATING
C47960 a_19240_46482# VSS 0.073862f **FLOATING
C47961 a_16375_45002# VSS 1.44161f **FLOATING
C47962 a_18243_46436# VSS 0.005441f **FLOATING
C47963 a_18147_46436# VSS 0.005048f **FLOATING
C47964 a_13259_45724# VSS 4.49011f **FLOATING
C47965 a_14383_46116# VSS 0.00471f **FLOATING
C47966 a_15194_46482# VSS 0.001266f **FLOATING
C47967 a_14949_46494# VSS 9.68e-19 **FLOATING
C47968 a_14537_46482# VSS 0.004992f **FLOATING
C47969 a_12839_46116# VSS 0.001465f **FLOATING
C47970 a_11315_46155# VSS 2.7e-19 **FLOATING
C47971 a_14371_46494# VSS 0.006939f **FLOATING
C47972 a_14180_46482# VSS 0.073862f **FLOATING
C47973 a_12638_46436# VSS 0.162178f **FLOATING
C47974 a_12379_46436# VSS 0.275423f **FLOATING
C47975 a_12005_46436# VSS 0.001661f **FLOATING
C47976 a_9751_46155# VSS 2.7e-19 **FLOATING
C47977 a_11608_46482# VSS 0.003279f **FLOATING
C47978 a_11387_46482# VSS 0.002827f **FLOATING
C47979 a_10586_45546# VSS 0.542658f **FLOATING
C47980 a_8379_46155# VSS 2.7e-19 **FLOATING
C47981 a_10044_46482# VSS 0.003279f **FLOATING
C47982 a_9823_46482# VSS 0.002827f **FLOATING
C47983 a_9241_46436# VSS 0.001883f **FLOATING
C47984 a_8049_45260# VSS 0.741927f **FLOATING
C47985 a_8781_46436# VSS 0.00189f **FLOATING
C47986 a_6347_46155# VSS 2.7e-19 **FLOATING
C47987 a_8034_45724# VSS 0.299594f **FLOATING
C47988 a_8283_46482# VSS 0.002857f **FLOATING
C47989 a_8062_46482# VSS 0.003279f **FLOATING
C47990 a_5527_46155# VSS 2.7e-19 **FLOATING
C47991 a_6640_46482# VSS 0.003279f **FLOATING
C47992 a_6419_46482# VSS 0.003313f **FLOATING
C47993 a_5066_45546# VSS 0.436834f **FLOATING
C47994 a_5431_46482# VSS 0.003543f **FLOATING
C47995 a_5210_46482# VSS 0.003279f **FLOATING
C47996 a_4365_46436# VSS 0.001655f **FLOATING
C47997 a_1337_46116# VSS 0.007537f **FLOATING
C47998 a_835_46155# VSS 0.001095f **FLOATING
C47999 a_518_46155# VSS 4.91e-19 **FLOATING
C48000 a_3873_46454# VSS 0.00338f **FLOATING
C48001 a_n1925_42282# VSS 1.34109f **FLOATING
C48002 a_526_44458# VSS 6.44493f **FLOATING
C48003 a_2981_46116# VSS 0.091491f **FLOATING
C48004 a_1431_46436# VSS 0.005311f **FLOATING
C48005 a_1337_46436# VSS 0.005657f **FLOATING
C48006 a_739_46482# VSS 0.004344f **FLOATING
C48007 a_518_46482# VSS 0.003651f **FLOATING
C48008 a_n1533_46116# VSS 0.006086f **FLOATING
C48009 a_n722_46482# VSS 0.001281f **FLOATING
C48010 a_n967_46494# VSS 4.65e-19 **FLOATING
C48011 a_n1379_46482# VSS 0.004992f **FLOATING
C48012 a_n1545_46494# VSS 0.006939f **FLOATING
C48013 a_n1736_46482# VSS 0.07565f **FLOATING
C48014 a_n2956_38680# VSS 1.34225f **FLOATING
C48015 a_n2956_39304# VSS 1.60721f **FLOATING
C48016 a_22959_46124# VSS 0.345245f **FLOATING
C48017 a_10809_44734# VSS 1.05002f **FLOATING
C48018 a_22223_46124# VSS 0.354467f **FLOATING
C48019 a_6945_45028# VSS 0.978274f **FLOATING
C48020 a_21137_46414# VSS 0.340736f **FLOATING
C48021 a_20708_46348# VSS 0.268156f **FLOATING
C48022 a_19900_46494# VSS 0.26164f **FLOATING
C48023 a_20075_46420# VSS 0.475201f **FLOATING
C48024 a_19335_46494# VSS 0.260378f **FLOATING
C48025 a_19553_46090# VSS 0.179968f **FLOATING
C48026 a_18985_46122# VSS 0.297132f **FLOATING
C48027 a_18819_46122# VSS 0.545109f **FLOATING
C48028 a_17957_46116# VSS 0.309446f **FLOATING
C48029 a_18189_46348# VSS 0.296366f **FLOATING
C48030 a_17715_44484# VSS 0.55862f **FLOATING
C48031 a_17583_46090# VSS 0.307562f **FLOATING
C48032 a_15682_46116# VSS 1.96743f **FLOATING
C48033 a_2324_44458# VSS 6.12227f **FLOATING
C48034 a_14840_46494# VSS 0.263367f **FLOATING
C48035 a_15015_46420# VSS 0.472948f **FLOATING
C48036 a_14275_46494# VSS 0.258968f **FLOATING
C48037 a_14493_46090# VSS 0.176122f **FLOATING
C48038 a_13925_46122# VSS 0.294602f **FLOATING
C48039 a_13759_46122# VSS 0.518292f **FLOATING
C48040 a_13351_46090# VSS 0.304427f **FLOATING
C48041 a_12594_46348# VSS 0.284494f **FLOATING
C48042 a_12005_46116# VSS 0.381711f **FLOATING
C48043 a_10903_43370# VSS 2.66576f **FLOATING
C48044 a_11387_46155# VSS 0.260117f **FLOATING
C48045 a_11133_46155# VSS 0.299642f **FLOATING
C48046 a_11189_46129# VSS 0.32558f **FLOATING
C48047 a_9290_44172# VSS 4.78398f **FLOATING
C48048 a_10355_46116# VSS 0.290668f **FLOATING
C48049 a_9823_46155# VSS 0.261206f **FLOATING
C48050 a_9569_46155# VSS 0.304755f **FLOATING
C48051 a_9625_46129# VSS 0.369694f **FLOATING
C48052 a_8953_45546# VSS 1.00397f **FLOATING
C48053 a_5937_45572# VSS 1.8333f **FLOATING
C48054 a_8199_44636# VSS 2.29742f **FLOATING
C48055 a_8349_46414# VSS 0.273442f **FLOATING
C48056 a_8016_46348# VSS 0.539696f **FLOATING
C48057 a_7920_46348# VSS 0.269852f **FLOATING
C48058 a_6419_46155# VSS 0.273686f **FLOATING
C48059 a_6165_46155# VSS 0.303989f **FLOATING
C48060 a_5497_46414# VSS 0.304684f **FLOATING
C48061 a_5204_45822# VSS 0.338817f **FLOATING
C48062 a_5164_46348# VSS 0.419282f **FLOATING
C48063 a_5068_46348# VSS 0.25855f **FLOATING
C48064 a_4704_46090# VSS 0.296767f **FLOATING
C48065 a_4419_46090# VSS 0.357571f **FLOATING
C48066 a_4185_45028# VSS 2.50501f **FLOATING
C48067 a_3699_46348# VSS 0.226584f **FLOATING
C48068 a_3483_46348# VSS 4.80498f **FLOATING
C48069 a_3147_46376# VSS 0.52775f **FLOATING
C48070 a_2804_46116# VSS 0.222855f **FLOATING
C48071 a_2698_46116# VSS 0.215567f **FLOATING
C48072 a_2521_46116# VSS 0.220999f **FLOATING
C48073 a_167_45260# VSS 1.32487f **FLOATING
C48074 a_2202_46116# VSS 0.273578f **FLOATING
C48075 a_1823_45246# VSS 2.36307f **FLOATING
C48076 a_1138_42852# VSS 0.456566f **FLOATING
C48077 a_1176_45822# VSS 0.278365f **FLOATING
C48078 a_1208_46090# VSS 0.348206f **FLOATING
C48079 a_805_46414# VSS 0.27506f **FLOATING
C48080 a_472_46348# VSS 0.32751f **FLOATING
C48081 a_376_46348# VSS 0.285607f **FLOATING
C48082 a_n1076_46494# VSS 0.262147f **FLOATING
C48083 a_n901_46420# VSS 0.762523f **FLOATING
C48084 a_n1641_46494# VSS 0.256945f **FLOATING
C48085 a_n1423_46090# VSS 0.176189f **FLOATING
C48086 a_n1991_46122# VSS 0.305274f **FLOATING
C48087 a_n1853_46287# VSS 0.341802f **FLOATING
C48088 a_n2157_46122# VSS 0.525314f **FLOATING
C48089 a_n2293_46098# VSS 0.690447f **FLOATING
C48090 a_n2472_46090# VSS 0.290925f **FLOATING
C48091 a_n2840_46090# VSS 0.340313f **FLOATING
C48092 a_21542_46660# VSS 0.002215f **FLOATING
C48093 a_21297_46660# VSS 9.68e-19 **FLOATING
C48094 a_21076_30879# VSS 2.07961f **FLOATING
C48095 a_22959_46660# VSS 0.338967f **FLOATING
C48096 a_12741_44636# VSS 0.979225f **FLOATING
C48097 a_20820_30879# VSS 1.68292f **FLOATING
C48098 a_22591_46660# VSS 0.292786f **FLOATING
C48099 a_11415_45002# VSS 1.63684f **FLOATING
C48100 a_20202_43084# VSS 1.05073f **FLOATING
C48101 a_22365_46825# VSS 0.208388f **FLOATING
C48102 a_20885_46660# VSS 0.004992f **FLOATING
C48103 a_20719_46660# VSS 0.006939f **FLOATING
C48104 a_19636_46660# VSS 0.003657f **FLOATING
C48105 a_18900_46660# VSS 0.006141f **FLOATING
C48106 a_18280_46660# VSS 0.29316f **FLOATING
C48107 a_17639_46660# VSS 0.308795f **FLOATING
C48108 a_16655_46660# VSS 0.003226f **FLOATING
C48109 a_16434_46660# VSS 0.003279f **FLOATING
C48110 a_20731_47026# VSS 0.004694f **FLOATING
C48111 a_20528_46660# VSS 0.07565f **FLOATING
C48112 a_22000_46634# VSS 0.295895f **FLOATING
C48113 a_21188_46660# VSS 0.261124f **FLOATING
C48114 a_21363_46634# VSS 0.488515f **FLOATING
C48115 a_20623_46660# VSS 0.258464f **FLOATING
C48116 a_20841_46902# VSS 0.180869f **FLOATING
C48117 a_20273_46660# VSS 0.309206f **FLOATING
C48118 a_20411_46873# VSS 0.393328f **FLOATING
C48119 a_20107_46660# VSS 0.575208f **FLOATING
C48120 a_19551_46910# VSS 0.005326f **FLOATING
C48121 a_19123_46287# VSS 0.477642f **FLOATING
C48122 a_18285_46348# VSS 0.577053f **FLOATING
C48123 a_17829_46910# VSS 3.25e-20 **FLOATING
C48124 a_765_45546# VSS 0.902406f **FLOATING
C48125 a_17339_46660# VSS 0.927636f **FLOATING
C48126 a_15312_46660# VSS 0.003243f **FLOATING
C48127 a_14447_46660# VSS 0.002898f **FLOATING
C48128 a_14226_46660# VSS 0.002596f **FLOATING
C48129 a_16751_46987# VSS 2.7e-19 **FLOATING
C48130 a_16721_46634# VSS 0.305539f **FLOATING
C48131 a_16388_46812# VSS 1.42609f **FLOATING
C48132 a_13059_46348# VSS 2.36107f **FLOATING
C48133 a_15227_46910# VSS 0.004775f **FLOATING
C48134 a_13693_46688# VSS 0.003947f **FLOATING
C48135 a_14543_46987# VSS 2.7e-19 **FLOATING
C48136 a_14513_46634# VSS 0.29862f **FLOATING
C48137 a_14180_46812# VSS 0.368158f **FLOATING
C48138 a_14035_46660# VSS 0.322858f **FLOATING
C48139 a_13885_46660# VSS 0.297377f **FLOATING
C48140 a_13170_46660# VSS 0.001266f **FLOATING
C48141 a_12925_46660# VSS 4.65e-19 **FLOATING
C48142 a_12513_46660# VSS 0.004992f **FLOATING
C48143 a_12347_46660# VSS 0.006939f **FLOATING
C48144 a_10933_46660# VSS 0.008634f **FLOATING
C48145 a_10861_46660# VSS 0.00579f **FLOATING
C48146 a_12359_47026# VSS 0.007095f **FLOATING
C48147 a_12156_46660# VSS 0.074642f **FLOATING
C48148 a_10425_46660# VSS 9.68e-19 **FLOATING
C48149 a_10185_46660# VSS 0.002215f **FLOATING
C48150 a_19692_46634# VSS 1.97188f **FLOATING
C48151 a_19466_46812# VSS 0.675335f **FLOATING
C48152 a_19333_46634# VSS 0.289568f **FLOATING
C48153 a_15227_44166# VSS 2.80559f **FLOATING
C48154 a_18834_46812# VSS 0.198054f **FLOATING
C48155 a_17609_46634# VSS 0.205547f **FLOATING
C48156 a_16292_46812# VSS 0.271203f **FLOATING
C48157 a_15559_46634# VSS 0.394779f **FLOATING
C48158 a_15368_46634# VSS 0.278142f **FLOATING
C48159 a_14976_45028# VSS 0.479565f **FLOATING
C48160 a_3090_45724# VSS 2.6372f **FLOATING
C48161 a_15009_46634# VSS 0.270859f **FLOATING
C48162 a_14084_46812# VSS 0.251005f **FLOATING
C48163 a_13607_46688# VSS 0.218935f **FLOATING
C48164 a_12816_46660# VSS 0.260317f **FLOATING
C48165 a_12991_46634# VSS 0.475827f **FLOATING
C48166 a_12251_46660# VSS 0.270927f **FLOATING
C48167 a_12469_46902# VSS 0.193369f **FLOATING
C48168 a_11901_46660# VSS 0.303844f **FLOATING
C48169 a_11813_46116# VSS 0.563718f **FLOATING
C48170 a_11735_46660# VSS 0.520568f **FLOATING
C48171 a_11186_47026# VSS 0.078586f **FLOATING
C48172 a_10768_47026# VSS 0.006047f **FLOATING
C48173 a_8846_46660# VSS 0.002215f **FLOATING
C48174 a_8601_46660# VSS 9.68e-19 **FLOATING
C48175 a_8270_45546# VSS 0.779033f **FLOATING
C48176 a_8189_46660# VSS 0.004992f **FLOATING
C48177 a_8023_46660# VSS 0.006939f **FLOATING
C48178 a_6903_46660# VSS 0.002857f **FLOATING
C48179 a_6682_46660# VSS 0.002596f **FLOATING
C48180 a_8035_47026# VSS 0.004694f **FLOATING
C48181 a_7832_46660# VSS 0.073862f **FLOATING
C48182 a_6086_46660# VSS 0.001266f **FLOATING
C48183 a_5841_46660# VSS 4.65e-19 **FLOATING
C48184 a_6999_46987# VSS 2.7e-19 **FLOATING
C48185 a_6969_46634# VSS 0.289597f **FLOATING
C48186 a_6755_46942# VSS 3.33348f **FLOATING
C48187 a_10249_46116# VSS 0.414443f **FLOATING
C48188 a_10554_47026# VSS 0.191251f **FLOATING
C48189 a_10623_46897# VSS 0.283572f **FLOATING
C48190 a_10467_46802# VSS 0.523954f **FLOATING
C48191 a_10428_46928# VSS 0.314538f **FLOATING
C48192 a_10150_46912# VSS 0.276624f **FLOATING
C48193 a_9863_46634# VSS 0.607398f **FLOATING
C48194 a_8492_46660# VSS 0.283316f **FLOATING
C48195 a_8667_46634# VSS 0.596387f **FLOATING
C48196 a_7927_46660# VSS 0.269867f **FLOATING
C48197 a_8145_46902# VSS 0.179735f **FLOATING
C48198 a_7577_46660# VSS 0.314978f **FLOATING
C48199 a_7715_46873# VSS 0.546182f **FLOATING
C48200 a_7411_46660# VSS 0.532412f **FLOATING
C48201 a_5257_43370# VSS 1.42323f **FLOATING
C48202 a_5429_46660# VSS 0.004992f **FLOATING
C48203 a_5263_46660# VSS 0.006939f **FLOATING
C48204 a_3878_46660# VSS 0.002215f **FLOATING
C48205 a_3633_46660# VSS 9.68e-19 **FLOATING
C48206 a_5275_47026# VSS 0.005488f **FLOATING
C48207 a_5072_46660# VSS 0.073862f **FLOATING
C48208 a_6540_46812# VSS 0.248814f **FLOATING
C48209 a_5732_46660# VSS 0.260482f **FLOATING
C48210 a_5907_46634# VSS 0.473347f **FLOATING
C48211 a_5167_46660# VSS 0.263586f **FLOATING
C48212 a_5385_46902# VSS 0.17737f **FLOATING
C48213 a_4817_46660# VSS 0.296797f **FLOATING
C48214 a_4955_46873# VSS 0.365781f **FLOATING
C48215 a_4651_46660# VSS 0.548065f **FLOATING
C48216 a_4646_46812# VSS 2.12519f **FLOATING
C48217 a_3877_44458# VSS 2.8543f **FLOATING
C48218 a_3221_46660# VSS 0.00579f **FLOATING
C48219 a_3055_46660# VSS 0.008634f **FLOATING
C48220 a_2162_46660# VSS 0.006278f **FLOATING
C48221 a_1302_46660# VSS 0.001378f **FLOATING
C48222 a_1057_46660# VSS 5.58e-19 **FLOATING
C48223 a_3067_47026# VSS 0.004694f **FLOATING
C48224 a_2864_46660# VSS 0.080001f **FLOATING
C48225 a_3524_46660# VSS 0.267612f **FLOATING
C48226 a_3699_46634# VSS 0.499647f **FLOATING
C48227 a_2959_46660# VSS 0.261026f **FLOATING
C48228 a_3177_46902# VSS 0.184239f **FLOATING
C48229 a_2609_46660# VSS 0.302878f **FLOATING
C48230 a_2443_46660# VSS 0.657702f **FLOATING
C48231 a_n2661_46098# VSS 2.05975f **FLOATING
C48232 a_1799_45572# VSS 0.30194f **FLOATING
C48233 a_645_46660# VSS 0.006691f **FLOATING
C48234 a_479_46660# VSS 0.008994f **FLOATING
C48235 a_1110_47026# VSS 8.17e-20 **FLOATING
C48236 a_n935_46688# VSS 0.004685f **FLOATING
C48237 a_491_47026# VSS 0.010533f **FLOATING
C48238 a_288_46660# VSS 0.075217f **FLOATING
C48239 a_1983_46706# VSS 0.205951f **FLOATING
C48240 a_2107_46812# VSS 1.13475f **FLOATING
C48241 a_948_46660# VSS 0.263413f **FLOATING
C48242 a_1123_46634# VSS 0.776627f **FLOATING
C48243 a_383_46660# VSS 0.269735f **FLOATING
C48244 a_601_46902# VSS 0.192316f **FLOATING
C48245 a_33_46660# VSS 0.309712f **FLOATING
C48246 a_171_46873# VSS 0.579977f **FLOATING
C48247 a_n133_46660# VSS 0.576523f **FLOATING
C48248 a_n2438_43548# VSS 2.99787f **FLOATING
C48249 a_n743_46660# VSS 3.29885f **FLOATING
C48250 a_n1021_46688# VSS 0.271211f **FLOATING
C48251 a_n1925_46634# VSS 1.33202f **FLOATING
C48252 a_n2312_38680# VSS 2.0221f **FLOATING
C48253 a_n2104_46634# VSS 0.340006f **FLOATING
C48254 a_n2293_46634# VSS 1.52366f **FLOATING
C48255 a_n2442_46660# VSS 1.32617f **FLOATING
C48256 a_n2472_46634# VSS 0.323981f **FLOATING
C48257 a_n2661_46634# VSS 0.742038f **FLOATING
C48258 a_n2956_39768# VSS 1.30197f **FLOATING
C48259 a_n2840_46634# VSS 0.328049f **FLOATING
C48260 a_22612_30879# VSS 3.44324f **FLOATING
C48261 a_21588_30879# VSS 2.81091f **FLOATING
C48262 a_20916_46384# VSS 0.827544f **FLOATING
C48263 a_20843_47204# VSS 0.121976f **FLOATING
C48264 a_19594_46812# VSS 0.277274f **FLOATING
C48265 a_19321_45002# VSS 1.15234f **FLOATING
C48266 a_19452_47524# VSS 0.006141f **FLOATING
C48267 a_13747_46662# VSS 2.11905f **FLOATING
C48268 a_13661_43548# VSS 2.82749f **FLOATING
C48269 a_5807_45002# VSS 2.5828f **FLOATING
C48270 a_16131_47204# VSS 0.004694f **FLOATING
C48271 a_16942_47570# VSS 0.001266f **FLOATING
C48272 a_16697_47582# VSS 4.65e-19 **FLOATING
C48273 a_16285_47570# VSS 0.004992f **FLOATING
C48274 a_16119_47582# VSS 0.006939f **FLOATING
C48275 a_15928_47570# VSS 0.075455f **FLOATING
C48276 a_768_44030# VSS 3.03052f **FLOATING
C48277 a_12549_44172# VSS 2.68201f **FLOATING
C48278 a_12891_46348# VSS 1.22195f **FLOATING
C48279 a_11309_47204# VSS 0.423399f **FLOATING
C48280 a_11117_47542# VSS 0.003386f **FLOATING
C48281 a_10037_47542# VSS 0.004685f **FLOATING
C48282 a_9804_47204# VSS 0.528639f **FLOATING
C48283 a_8128_46384# VSS 0.573494f **FLOATING
C48284 a_5159_47243# VSS 2.7e-19 **FLOATING
C48285 a_7989_47542# VSS 0.004685f **FLOATING
C48286 a_n881_46662# VSS 4.56296f **FLOATING
C48287 a_n1613_43370# VSS 4.90074f **FLOATING
C48288 a_3411_47243# VSS 4.87e-19 **FLOATING
C48289 a_3094_47243# VSS 3.78e-19 **FLOATING
C48290 a_5063_47570# VSS 0.003543f **FLOATING
C48291 a_4842_47570# VSS 0.003279f **FLOATING
C48292 a_2583_47243# VSS 2.7e-19 **FLOATING
C48293 a_2266_47243# VSS 6.13e-20 **FLOATING
C48294 a_3315_47570# VSS 0.003543f **FLOATING
C48295 a_3094_47570# VSS 0.003279f **FLOATING
C48296 a_7_47243# VSS 2.7e-19 **FLOATING
C48297 a_2747_46873# VSS 0.287894f **FLOATING
C48298 a_2487_47570# VSS 0.003543f **FLOATING
C48299 a_2266_47570# VSS 0.003328f **FLOATING
C48300 a_n89_47570# VSS 0.002898f **FLOATING
C48301 a_n310_47570# VSS 0.003279f **FLOATING
C48302 a_n2312_39304# VSS 1.49307f **FLOATING
C48303 a_n2312_40392# VSS 2.25565f **FLOATING
C48304 a_22959_47212# VSS 0.322938f **FLOATING
C48305 a_11453_44696# VSS 0.689179f **FLOATING
C48306 SMPL_ON_N VSS 2.60102f **FLOATING
C48307 a_22731_47423# VSS 0.227778f **FLOATING
C48308 a_22223_47212# VSS 0.332189f **FLOATING
C48309 a_12465_44636# VSS 5.61685f **FLOATING
C48310 a_21811_47423# VSS 0.23358f **FLOATING
C48311 a_4883_46098# VSS 1.54736f **FLOATING
C48312 a_21496_47436# VSS 0.249536f **FLOATING
C48313 a_13507_46334# VSS 4.83849f **FLOATING
C48314 a_21177_47436# VSS 0.223524f **FLOATING
C48315 a_20990_47178# VSS 0.224581f **FLOATING
C48316 a_20894_47436# VSS 0.233111f **FLOATING
C48317 a_19787_47423# VSS 0.258015f **FLOATING
C48318 a_19386_47436# VSS 0.209882f **FLOATING
C48319 a_18597_46090# VSS 2.82344f **FLOATING
C48320 a_18780_47178# VSS 0.319719f **FLOATING
C48321 a_18479_47436# VSS 1.19826f **FLOATING
C48322 a_18143_47464# VSS 0.579061f **FLOATING
C48323 a_10227_46804# VSS 8.12328f **FLOATING
C48324 a_17591_47464# VSS 0.576556f **FLOATING
C48325 a_16588_47582# VSS 0.263715f **FLOATING
C48326 a_16763_47508# VSS 0.587861f **FLOATING
C48327 a_16023_47582# VSS 0.264352f **FLOATING
C48328 a_16327_47482# VSS 5.17799f **FLOATING
C48329 a_16241_47178# VSS 0.18232f **FLOATING
C48330 a_15673_47210# VSS 0.315684f **FLOATING
C48331 a_15811_47375# VSS 0.349499f **FLOATING
C48332 a_15507_47210# VSS 0.556554f **FLOATING
C48333 a_11599_46634# VSS 2.84967f **FLOATING
C48334 a_14955_47212# VSS 0.358339f **FLOATING
C48335 a_14311_47204# VSS 0.248858f **FLOATING
C48336 a_13487_47204# VSS 0.643275f **FLOATING
C48337 a_12861_44030# VSS 3.64545f **FLOATING
C48338 a_13717_47436# VSS 1.02478f **FLOATING
C48339 a_n1435_47204# VSS 9.72476f **FLOATING
C48340 a_13381_47204# VSS 0.225132f **FLOATING
C48341 a_11459_47204# VSS 0.553679f **FLOATING
C48342 a_9313_45822# VSS 1.04727f **FLOATING
C48343 a_11031_47542# VSS 0.247302f **FLOATING
C48344 a_9863_47436# VSS 0.265619f **FLOATING
C48345 a_9067_47204# VSS 0.606182f **FLOATING
C48346 a_6575_47204# VSS 0.798434f **FLOATING
C48347 a_7903_47542# VSS 0.258657f **FLOATING
C48348 a_7227_47204# VSS 0.610401f **FLOATING
C48349 a_6851_47204# VSS 0.346433f **FLOATING
C48350 a_6491_46660# VSS 0.343406f **FLOATING
C48351 a_6545_47178# VSS 0.597936f **FLOATING
C48352 a_6151_47436# VSS 2.12954f **FLOATING
C48353 a_5815_47464# VSS 0.594449f **FLOATING
C48354 a_5129_47502# VSS 0.361487f **FLOATING
C48355 a_4915_47217# VSS 2.79467f **FLOATING
C48356 a_n443_46116# VSS 4.167f **FLOATING
C48357 a_4791_45118# VSS 2.65418f **FLOATING
C48358 a_4700_47436# VSS 0.271201f **FLOATING
C48359 a_4007_47204# VSS 0.628996f **FLOATING
C48360 a_3815_47204# VSS 0.440491f **FLOATING
C48361 a_3785_47178# VSS 0.541893f **FLOATING
C48362 a_3381_47502# VSS 0.320926f **FLOATING
C48363 a_n1151_42308# VSS 3.78206f **FLOATING
C48364 a_3160_47472# VSS 0.607125f **FLOATING
C48365 a_2905_45572# VSS 0.47073f **FLOATING
C48366 a_2952_47436# VSS 0.275026f **FLOATING
C48367 a_2553_47502# VSS 0.294118f **FLOATING
C48368 a_2063_45854# VSS 1.92678f **FLOATING
C48369 a_584_46384# VSS 2.10508f **FLOATING
C48370 a_2124_47436# VSS 0.276508f **FLOATING
C48371 a_1431_47204# VSS 0.595895f **FLOATING
C48372 a_1239_47204# VSS 0.33333f **FLOATING
C48373 a_1209_47178# VSS 0.474725f **FLOATING
C48374 a_327_47204# VSS 0.581187f **FLOATING
C48375 a_n785_47204# VSS 0.361759f **FLOATING
C48376 a_n23_47502# VSS 0.278861f **FLOATING
C48377 a_n237_47217# VSS 3.05697f **FLOATING
C48378 a_n746_45260# VSS 0.993718f **FLOATING
C48379 a_n971_45724# VSS 4.81311f **FLOATING
C48380 a_n452_47436# VSS 0.28781f **FLOATING
C48381 a_n815_47178# VSS 0.513835f **FLOATING
C48382 a_n1605_47204# VSS 0.250546f **FLOATING
C48383 SMPL_ON_P VSS 4.94844f **FLOATING
C48384 a_n1741_47186# VSS 1.81488f **FLOATING
C48385 a_n1920_47178# VSS 0.310881f **FLOATING
C48386 a_n2109_47186# VSS 0.936844f **FLOATING
C48387 a_n2288_47178# VSS 0.346995f **FLOATING
C48388 a_n2497_47436# VSS 2.31207f **FLOATING
C48389 a_n2833_47464# VSS 0.602779f **FLOATING
C48390 w_11334_34010# VSS 51.3801f **FLOATING
C48391 w_1575_34946# VSS 51.6622f **FLOATING
.ends
