magic
tech sky130A
magscale 1 2
timestamp 1711312488
<< metal3 >>
rect -1436 812 1436 840
rect -1436 -812 1352 812
rect 1416 -812 1436 812
rect -1436 -840 1436 -812
<< via3 >>
rect 1352 -812 1416 812
<< mimcap >>
rect -1396 760 1104 800
rect -1396 -760 -1356 760
rect 1064 -760 1104 760
rect -1396 -800 1104 -760
<< mimcapcontact >>
rect -1356 -760 1064 760
<< metal4 >>
rect 1336 812 1432 828
rect -1357 760 1065 761
rect -1357 -760 -1356 760
rect 1064 -760 1065 760
rect -1357 -761 1065 -760
rect 1336 -812 1352 812
rect 1416 -812 1432 812
rect 1336 -828 1432 -812
<< properties >>
string FIXED_BBOX -1436 -840 1144 840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12.5 l 8 val 207.79 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
