* SPICE3 file created from CDAC_mim_12bit_flat.ext - technology: sky130A
* Changed subckt name to match symbol

.subckt CDAC_12bit C0_dummy C0 C1 C2 C3 C4 C5 C6 C7 C8 C9 C10 Ctop VSS
C0 C9 C8 27.029099f
C1 C10 C9 37.3538f
C2 C0_dummy Ctop 0.86078f
C3 C0 Ctop 0.86078f
C4 C0 C0_dummy 0.843585f
C5 C2 Ctop 3.44648f
C6 C2 C0_dummy 1.21947f
C7 C1 Ctop 1.72211f
C8 C2 C0 0.375889f
C9 C3 Ctop 6.89425f
C10 C4 Ctop 13.79f
C11 C1 C0 0.843585f
C12 C1 C2 0.410234f
C13 C5 Ctop 27.5919f
C14 C3 C2 1.13411f
C15 C6 Ctop 55.199303f
C16 C4 C2 1.25611f
C17 C3 C1 1.632f
C18 C7 Ctop 0.110397p
C19 C8 Ctop 0.220888p
C20 C4 C3 4.70302f
C21 C9 Ctop 0.441826p
C22 C10 Ctop 0.883365p
C23 C5 C4 7.15914f
C24 C6 C5 10.395f
C25 C7 C6 14.374f
C26 C8 C7 19.122501f
C27 Ctop VSS 85.3252f
C28 C0_dummy VSS 1.24206f
C29 C0 VSS 1.24206f
C30 C2 VSS 1.59764f
C31 C1 VSS 1.35955f
C32 C3 VSS 2.08631f
C33 C4 VSS 5.19193f
C34 C5 VSS 6.00823f
C35 C6 VSS 12.0184f
C36 C7 VSS 21.763699f
C37 C8 VSS 41.6382f
C38 C9 VSS 74.623505f
C39 C10 VSS 0.199576p
.ends
