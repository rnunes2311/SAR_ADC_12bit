magic
tech sky130A
magscale 1 2
timestamp 1711974700
<< pwell >>
rect 12750 3370 12830 3450
rect 10150 3230 10370 3270
rect 10380 3230 10540 3290
rect 12510 3240 12590 3320
rect 10150 3140 10540 3230
rect 10200 3130 10280 3140
rect 10370 3120 10540 3140
rect 10370 3100 10650 3120
rect 10380 3040 10650 3100
rect 12430 3060 12510 3140
rect 12670 3060 12750 3140
rect 10520 3030 10650 3040
rect 10570 2960 10650 3030
rect 10700 2880 10860 3040
rect 10910 2800 11070 2960
rect 12600 2900 12680 2980
<< locali >>
rect -130 3950 5570 3960
rect -130 3900 -80 3950
rect 5520 3900 5570 3950
rect -130 3890 5570 3900
rect 5630 3950 13470 3960
rect 5630 3910 5710 3950
rect 13370 3910 13470 3950
rect 5630 3890 13470 3910
rect -130 3860 -50 3890
rect -130 2100 -110 3860
rect -70 2100 -50 3860
rect -130 2060 -50 2100
rect 5630 3860 5700 3890
rect 5630 2100 5650 3860
rect 5690 2100 5700 3860
rect 5630 2060 5700 2100
rect 13410 3850 13470 3890
rect 13410 2090 13420 3850
rect 13460 2090 13470 3850
rect 13410 2060 13470 2090
rect -130 2050 5530 2060
rect -130 2010 10 2050
rect 5490 2010 5530 2050
rect -130 1990 5530 2010
rect 5630 2050 13470 2060
rect 5630 2010 5730 2050
rect 13390 2010 13470 2050
rect 5630 1990 13470 2010
<< viali >>
rect -80 3900 5520 3950
rect 5710 3910 13370 3950
rect -110 2100 -70 3860
rect 5650 2100 5690 3860
rect 13420 2090 13460 3850
rect 10 2010 5490 2050
rect 5730 2010 13390 2050
<< metal1 >>
rect -130 3950 5570 3960
rect -130 3900 -80 3950
rect 5520 3900 5570 3950
rect -130 3890 5570 3900
rect 5630 3950 13470 3960
rect 5630 3910 5710 3950
rect 13370 3910 13470 3950
rect 5630 3890 13470 3910
rect -130 3860 -50 3890
rect -130 3550 -110 3860
rect -70 3550 -50 3860
rect 5630 3860 5700 3890
rect 60 3780 70 3840
rect 130 3831 140 3840
rect 130 3781 2060 3831
rect 2110 3830 2120 3840
rect 130 3780 140 3781
rect 2100 3780 2120 3830
rect 2180 3830 2190 3840
rect 2180 3780 3090 3830
rect 3130 3780 3140 3840
rect 3200 3830 3210 3840
rect 3650 3830 3660 3840
rect 3200 3780 3600 3830
rect 3640 3780 3660 3830
rect 3720 3830 3730 3840
rect 3720 3780 3850 3830
rect 3900 3780 3910 3840
rect 3970 3780 3980 3840
rect 4140 3780 4150 3840
rect 4210 3780 4220 3840
rect 4390 3780 4400 3840
rect 4460 3780 4470 3840
rect 4630 3780 4640 3840
rect 4700 3780 4710 3840
rect 4870 3780 4880 3840
rect 4940 3780 4950 3840
rect 5120 3780 5130 3840
rect 5190 3780 5200 3840
rect 5350 3780 5360 3840
rect 5420 3780 5430 3840
rect -130 3490 -120 3550
rect -60 3490 -50 3550
rect -130 3400 -110 3490
rect -70 3400 -50 3490
rect -130 3340 -120 3400
rect -60 3340 -50 3400
rect -130 3250 -110 3340
rect -70 3250 -50 3340
rect -130 3190 -120 3250
rect -60 3190 -50 3250
rect 4000 3200 4010 3680
rect -130 2100 -110 3190
rect -70 2100 -50 3190
rect -10 3030 0 3090
rect 60 3030 70 3090
rect 250 3030 260 3090
rect 320 3030 330 3090
rect 510 3030 520 3090
rect 580 3030 590 3090
rect 760 3030 770 3090
rect 830 3030 840 3090
rect 1020 3030 1030 3090
rect 1090 3030 1100 3090
rect 1270 3030 1280 3090
rect 1340 3030 1350 3090
rect 1530 3030 1540 3090
rect 1600 3030 1610 3090
rect 1790 3030 1800 3090
rect 1860 3030 1870 3090
rect 2040 3030 2050 3090
rect 2110 3030 2120 3090
rect 2300 3030 2310 3090
rect 2370 3030 2380 3090
rect 2550 3030 2560 3090
rect 2620 3030 2630 3090
rect 2810 3030 2820 3090
rect 2880 3030 2890 3090
rect 3070 3030 3080 3090
rect 3140 3030 3150 3090
rect 3320 3030 3330 3090
rect 3390 3030 3400 3090
rect 3580 3030 3590 3090
rect 3650 3030 3660 3090
rect 3840 3030 3850 3090
rect 3910 3030 3920 3090
rect 4080 3030 4090 3090
rect 4150 3030 4160 3090
rect 4320 3030 4330 3090
rect 4390 3030 4400 3090
rect 4560 3030 4570 3090
rect 4630 3030 4640 3090
rect 4810 3030 4820 3090
rect 4880 3030 4890 3090
rect 5050 3030 5060 3090
rect 5120 3030 5130 3090
rect 5290 3030 5300 3090
rect 5360 3030 5370 3090
rect 120 2160 130 2220
rect 190 2160 200 2220
rect 380 2160 390 2220
rect 450 2160 460 2220
rect 640 2160 650 2220
rect 710 2160 720 2220
rect 890 2160 900 2220
rect 960 2160 970 2220
rect 1150 2160 1160 2220
rect 1220 2160 1230 2220
rect 1400 2160 1410 2220
rect 1470 2160 1480 2220
rect 1660 2160 1670 2220
rect 1730 2160 1740 2220
rect 1920 2160 1930 2220
rect 1990 2160 2000 2220
rect 2170 2160 2180 2220
rect 2240 2160 2250 2220
rect 2430 2160 2440 2220
rect 2500 2160 2510 2220
rect 2680 2160 2690 2220
rect 2750 2160 2760 2220
rect 2940 2160 2950 2220
rect 3010 2160 3020 2220
rect 3190 2160 3200 2220
rect 3260 2160 3270 2220
rect 3450 2160 3460 2220
rect 3520 2160 3530 2220
rect 3710 2160 3720 2220
rect 3780 2160 3790 2220
rect 3960 2160 3970 2220
rect 4030 2160 4040 2220
rect 4230 2190 4270 3020
rect 4470 2190 4510 3020
rect 4710 2190 4750 3020
rect 4960 2190 5000 3030
rect 5200 2190 5240 3030
rect 5440 2190 5480 3030
rect 5630 2970 5650 3860
rect 5690 2970 5700 3860
rect 13410 3850 13470 3890
rect 5900 3760 5910 3820
rect 5970 3810 5980 3820
rect 5970 3760 6560 3810
rect 6670 3760 6680 3820
rect 6740 3810 6750 3820
rect 6740 3760 6940 3810
rect 7060 3760 7070 3820
rect 7130 3760 7140 3820
rect 7230 3760 7240 3820
rect 7300 3760 7310 3820
rect 7450 3760 7460 3820
rect 7520 3760 7710 3820
rect 7870 3760 7880 3820
rect 7940 3760 8530 3820
rect 8640 3760 8650 3820
rect 8710 3760 9290 3820
rect 9410 3760 9420 3820
rect 9480 3760 9670 3820
rect 9790 3760 9800 3820
rect 9860 3760 9870 3820
rect 9980 3760 9990 3820
rect 10050 3760 10060 3820
rect 10190 3760 10200 3820
rect 10260 3760 10270 3820
rect 10380 3760 10390 3820
rect 10450 3760 10460 3820
rect 10500 3760 10510 3820
rect 10570 3760 10580 3820
rect 10710 3760 10720 3820
rect 10780 3760 10790 3820
rect 10920 3760 10930 3820
rect 10990 3760 11000 3820
rect 11130 3760 11140 3820
rect 11200 3760 11210 3820
rect 11340 3760 11350 3820
rect 11410 3760 11420 3820
rect 12860 3800 13070 3840
rect 7730 3640 7740 3700
rect 7800 3640 7810 3700
rect 7920 3640 7930 3700
rect 7990 3640 8000 3700
rect 8110 3640 8120 3700
rect 8180 3640 8190 3700
rect 8300 3640 8310 3700
rect 8370 3640 8380 3700
rect 8500 3640 8510 3700
rect 8570 3640 8580 3700
rect 8690 3640 8700 3700
rect 8760 3640 8770 3700
rect 8880 3640 8890 3700
rect 8950 3640 8960 3700
rect 9070 3640 9080 3700
rect 9140 3640 9150 3700
rect 9270 3640 9280 3700
rect 9340 3640 9350 3700
rect 9460 3640 9470 3700
rect 9530 3640 9540 3700
rect 9650 3640 9660 3700
rect 9720 3640 9730 3700
rect 9840 3640 9850 3700
rect 9910 3640 9920 3700
rect 10050 3540 10060 3600
rect 10120 3540 10130 3600
rect 10240 3540 10250 3600
rect 10310 3540 10320 3600
rect 10450 3540 10460 3600
rect 10520 3540 10530 3600
rect 10660 3540 10670 3600
rect 10730 3540 10740 3600
rect 10870 3540 10880 3600
rect 10940 3540 10950 3600
rect 11080 3540 11090 3600
rect 11150 3540 11160 3600
rect 11290 3540 11300 3600
rect 11360 3540 11370 3600
rect 7830 3440 7840 3500
rect 7900 3440 7910 3500
rect 8020 3440 8030 3500
rect 8090 3440 8100 3500
rect 8210 3440 8220 3500
rect 8280 3440 8290 3500
rect 8400 3440 8410 3500
rect 8470 3440 8480 3500
rect 10150 3370 10160 3430
rect 10220 3370 10230 3430
rect 10340 3370 10350 3430
rect 10410 3370 10420 3430
rect 10550 3370 10560 3430
rect 10620 3370 10630 3430
rect 10760 3370 10770 3430
rect 10830 3370 10840 3430
rect 10970 3370 10980 3430
rect 11040 3370 11050 3430
rect 11180 3380 11190 3440
rect 11250 3380 11260 3440
rect 11390 3380 11400 3440
rect 11460 3380 11470 3440
rect 12860 3430 12910 3800
rect 12940 3630 12950 3690
rect 13010 3630 13020 3690
rect 13300 3630 13310 3650
rect 13090 3600 13310 3630
rect 13300 3590 13310 3600
rect 13370 3590 13380 3650
rect 12860 3390 13070 3430
rect 11240 3230 11250 3290
rect 11310 3280 11320 3290
rect 12860 3280 12910 3390
rect 11310 3240 12910 3280
rect 11310 3230 11320 3240
rect 12030 3200 12040 3210
rect 10200 3140 10210 3200
rect 10270 3160 12040 3200
rect 10270 3140 10280 3160
rect 12030 3150 12040 3160
rect 12100 3150 12110 3210
rect 10390 3070 10400 3130
rect 10460 3120 10470 3130
rect 11870 3120 11880 3130
rect 10460 3080 11880 3120
rect 10460 3070 10470 3080
rect 11870 3070 11880 3080
rect 11940 3070 11950 3130
rect 10500 2990 10510 3050
rect 10570 3040 10580 3050
rect 11710 3040 11720 3050
rect 10570 3000 11720 3040
rect 10570 2990 10580 3000
rect 11710 2990 11720 3000
rect 11780 2990 11790 3050
rect 12860 3000 12910 3240
rect 12940 3220 12950 3280
rect 13010 3220 13020 3280
rect 13220 3230 13230 3250
rect 13090 3200 13230 3230
rect 13220 3190 13230 3200
rect 13290 3190 13300 3250
rect 5630 2910 5640 2970
rect 5700 2910 5710 2970
rect 10710 2910 10720 2970
rect 10780 2960 10790 2970
rect 11950 2960 11960 2970
rect 10780 2920 11960 2960
rect 10780 2910 10790 2920
rect 11950 2910 11960 2920
rect 12020 2910 12030 2970
rect 12860 2960 13070 3000
rect 5630 2810 5650 2910
rect 5690 2810 5700 2910
rect 10920 2830 10930 2890
rect 10990 2880 11000 2890
rect 11790 2880 11800 2890
rect 10990 2840 11800 2880
rect 10990 2830 11000 2840
rect 11790 2830 11800 2840
rect 11860 2830 11870 2890
rect 5630 2750 5640 2810
rect 5700 2750 5710 2810
rect 11130 2750 11140 2810
rect 11200 2800 11210 2810
rect 11630 2800 11640 2810
rect 11200 2760 11640 2800
rect 11200 2750 11210 2760
rect 11630 2750 11640 2760
rect 11700 2750 11710 2810
rect 5630 2680 5650 2750
rect 5690 2680 5700 2750
rect 5630 2620 5640 2680
rect 5700 2620 5710 2680
rect 5760 2620 5770 2680
rect 5830 2620 5840 2680
rect 5950 2620 5960 2680
rect 6020 2620 6030 2680
rect 6140 2620 6150 2680
rect 6210 2620 6220 2680
rect 6340 2620 6350 2680
rect 6410 2620 6420 2680
rect 6530 2620 6540 2680
rect 6600 2620 6610 2680
rect 6720 2620 6730 2680
rect 6790 2620 6800 2680
rect 6910 2620 6920 2680
rect 6980 2620 6990 2680
rect 7100 2620 7110 2680
rect 7170 2620 7180 2680
rect 11340 2670 11350 2730
rect 11410 2720 11420 2730
rect 11470 2720 11480 2730
rect 11410 2680 11480 2720
rect 11410 2670 11420 2680
rect 11470 2670 11480 2680
rect 11540 2670 11550 2730
rect 12860 2620 12910 2960
rect 12940 2790 12950 2850
rect 13010 2790 13020 2850
rect 13140 2780 13150 2800
rect 13090 2750 13150 2780
rect 13140 2740 13150 2750
rect 13210 2740 13220 2800
rect 4210 2130 4220 2190
rect 4280 2130 4290 2190
rect 4450 2130 4460 2190
rect 4520 2130 4530 2190
rect 4690 2130 4700 2190
rect 4760 2130 4770 2190
rect 4940 2130 4950 2190
rect 5010 2130 5020 2190
rect 5180 2130 5190 2190
rect 5250 2130 5260 2190
rect 5420 2130 5430 2190
rect 5490 2130 5500 2190
rect -130 2060 -50 2100
rect 5630 2100 5650 2620
rect 5690 2100 5700 2620
rect 10200 2560 10210 2620
rect 10270 2560 10280 2620
rect 10390 2560 10400 2620
rect 10460 2560 10470 2620
rect 10500 2560 10510 2620
rect 10570 2560 10580 2620
rect 10710 2560 10720 2620
rect 10780 2560 10790 2620
rect 10920 2560 10930 2620
rect 10990 2560 11000 2620
rect 11130 2560 11140 2620
rect 11200 2560 11210 2620
rect 11340 2560 11350 2620
rect 11410 2560 11420 2620
rect 11550 2560 11560 2620
rect 11620 2560 11630 2620
rect 11860 2570 13070 2620
rect 7310 2490 7320 2550
rect 7380 2490 7390 2550
rect 7500 2490 7510 2550
rect 7570 2490 7580 2550
rect 10050 2450 10060 2510
rect 10120 2450 10130 2510
rect 10240 2450 10250 2510
rect 10310 2450 10320 2510
rect 10450 2450 10460 2510
rect 10520 2450 10530 2510
rect 10660 2450 10670 2510
rect 10730 2450 10740 2510
rect 10870 2450 10880 2510
rect 10940 2450 10950 2510
rect 11080 2450 11090 2510
rect 11150 2450 11160 2510
rect 11290 2450 11300 2510
rect 11360 2450 11370 2510
rect 11500 2450 11510 2510
rect 11570 2450 11580 2510
rect 11710 2450 11720 2510
rect 11780 2450 11790 2510
rect 11900 2450 11910 2510
rect 11970 2450 11980 2510
rect 12210 2450 12220 2510
rect 12280 2450 12290 2510
rect 12420 2450 12430 2510
rect 12490 2450 12500 2510
rect 12630 2450 12640 2510
rect 12700 2450 12710 2510
rect 12840 2450 12850 2510
rect 12910 2450 12920 2510
rect 13050 2450 13060 2510
rect 13120 2450 13130 2510
rect 12110 2340 12120 2400
rect 12180 2340 12190 2400
rect 12320 2340 12330 2400
rect 12390 2340 12400 2400
rect 12530 2340 12540 2400
rect 12600 2340 12610 2400
rect 12740 2340 12750 2400
rect 12810 2340 12820 2400
rect 12950 2340 12960 2400
rect 13020 2340 13030 2400
rect 5860 2180 5870 2240
rect 5930 2180 5940 2240
rect 6050 2180 6060 2240
rect 6120 2180 6130 2240
rect 6240 2180 6250 2240
rect 6310 2180 6320 2240
rect 6430 2180 6440 2240
rect 6500 2180 6510 2240
rect 6620 2180 6630 2240
rect 6690 2180 6700 2240
rect 6820 2180 6830 2240
rect 6890 2180 6900 2240
rect 7010 2180 7020 2240
rect 7080 2180 7090 2240
rect 7200 2180 7210 2240
rect 7270 2180 7280 2240
rect 7410 2180 7420 2240
rect 7480 2180 7490 2240
rect 7600 2180 7610 2240
rect 7670 2180 7680 2240
rect 8590 2150 8600 2210
rect 8660 2150 8670 2210
rect 8790 2150 8800 2210
rect 8860 2150 8870 2210
rect 8980 2150 8990 2210
rect 9050 2150 9060 2210
rect 9170 2150 9180 2210
rect 9240 2150 9250 2210
rect 9360 2150 9370 2210
rect 9430 2150 9440 2210
rect 9550 2150 9560 2210
rect 9620 2150 9630 2210
rect 9750 2150 9760 2210
rect 9820 2150 9830 2210
rect 9940 2150 9950 2210
rect 10010 2150 10020 2210
rect 10150 2190 10160 2250
rect 10220 2190 10230 2250
rect 10340 2190 10350 2250
rect 10410 2190 10420 2250
rect 10550 2190 10560 2250
rect 10620 2190 10630 2250
rect 10760 2190 10770 2250
rect 10830 2190 10840 2250
rect 10970 2190 10980 2250
rect 11040 2190 11050 2250
rect 11180 2190 11190 2250
rect 11250 2190 11260 2250
rect 11390 2190 11400 2250
rect 11460 2190 11470 2250
rect 11600 2190 11610 2250
rect 11670 2190 11680 2250
rect 11810 2160 11820 2220
rect 11880 2160 11890 2220
rect 12000 2160 12010 2220
rect 12070 2160 12080 2220
rect 5630 2060 5700 2100
rect 13410 2090 13420 3850
rect 13460 2090 13470 3850
rect 13410 2060 13470 2090
rect -130 2050 5530 2060
rect -130 2010 10 2050
rect 5490 2010 5530 2050
rect -130 1990 5530 2010
rect 5630 2050 13470 2060
rect 5630 2010 5730 2050
rect 13390 2010 13470 2050
rect 5630 1990 13470 2010
rect 120 1855 130 1915
rect 190 1900 200 1915
rect 5860 1900 5870 1915
rect 190 1870 5870 1900
rect 190 1855 200 1870
rect 5860 1855 5870 1870
rect 5930 1900 5940 1915
rect 7410 1900 7420 1915
rect 5930 1870 7420 1900
rect 5930 1855 5940 1870
rect 7410 1855 7420 1870
rect 7480 1900 7490 1915
rect 8590 1900 8600 1915
rect 7480 1870 8600 1900
rect 7480 1855 7490 1870
rect 8590 1855 8600 1870
rect 8660 1900 8670 1915
rect 8660 1870 13440 1900
rect 8660 1855 8670 1870
rect 2170 1765 2180 1825
rect 2240 1810 2250 1825
rect 6620 1810 6630 1825
rect 2240 1780 6630 1810
rect 2240 1765 2250 1780
rect 6620 1765 6630 1780
rect 6690 1810 6700 1825
rect 7600 1810 7610 1825
rect 6690 1780 7610 1810
rect 6690 1765 6700 1780
rect 7600 1765 7610 1780
rect 7670 1810 7680 1825
rect 9360 1810 9370 1825
rect 7670 1780 9370 1810
rect 7670 1765 7680 1780
rect 9360 1765 9370 1780
rect 9430 1810 9440 1825
rect 9430 1780 13440 1810
rect 9430 1765 9440 1780
rect 3190 1675 3200 1735
rect 3260 1720 3270 1735
rect 7010 1720 7020 1735
rect 3260 1690 7020 1720
rect 3260 1675 3270 1690
rect 7010 1675 7020 1690
rect 7080 1720 7090 1735
rect 9740 1720 9750 1735
rect 7080 1690 9750 1720
rect 7080 1675 7090 1690
rect 9740 1675 9750 1690
rect 9810 1720 9820 1735
rect 11810 1720 11820 1735
rect 9810 1690 11820 1720
rect 9810 1675 9820 1690
rect 11810 1675 11820 1690
rect 11880 1720 11890 1735
rect 11880 1690 13440 1720
rect 11880 1675 11890 1690
rect 3710 1585 3720 1645
rect 3780 1630 3790 1645
rect 7200 1630 7210 1645
rect 3780 1600 7210 1630
rect 3780 1585 3790 1600
rect 7200 1585 7210 1600
rect 7270 1630 7280 1645
rect 9940 1630 9950 1645
rect 7270 1600 9950 1630
rect 7270 1585 7280 1600
rect 9940 1585 9950 1600
rect 10010 1630 10020 1645
rect 12000 1630 12010 1645
rect 10010 1600 12010 1630
rect 10010 1585 10020 1600
rect 12000 1585 12010 1600
rect 12070 1630 12080 1645
rect 12070 1600 13440 1630
rect 12070 1585 12080 1600
rect 3960 1495 3970 1555
rect 4030 1540 4040 1555
rect 10150 1540 10160 1555
rect 4030 1510 10160 1540
rect 4030 1495 4040 1510
rect 10150 1495 10160 1510
rect 10220 1540 10230 1555
rect 12110 1540 12120 1555
rect 10220 1510 12120 1540
rect 10220 1495 10230 1510
rect 12110 1495 12120 1510
rect 12180 1540 12190 1555
rect 12180 1510 13440 1540
rect 12180 1495 12190 1510
rect 4210 1405 4220 1465
rect 4280 1450 4290 1465
rect 10340 1450 10350 1465
rect 4280 1420 10350 1450
rect 4280 1405 4290 1420
rect 10340 1405 10350 1420
rect 10410 1450 10420 1465
rect 12320 1450 12330 1465
rect 10410 1420 12330 1450
rect 10410 1405 10420 1420
rect 12320 1405 12330 1420
rect 12390 1450 12400 1465
rect 12390 1420 13440 1450
rect 12390 1405 12400 1420
rect 4450 1315 4460 1375
rect 4520 1360 4530 1375
rect 10550 1360 10560 1375
rect 4520 1330 10560 1360
rect 4520 1315 4530 1330
rect 10550 1315 10560 1330
rect 10620 1360 10630 1375
rect 12530 1360 12540 1375
rect 10620 1330 12540 1360
rect 10620 1315 10630 1330
rect 12530 1315 12540 1330
rect 12600 1360 12610 1375
rect 12600 1330 13440 1360
rect 12600 1315 12610 1330
rect 4690 1225 4700 1285
rect 4760 1270 4770 1285
rect 10760 1270 10770 1285
rect 4760 1240 10770 1270
rect 4760 1225 4770 1240
rect 10760 1225 10770 1240
rect 10830 1270 10840 1285
rect 13140 1270 13150 1285
rect 10830 1240 13150 1270
rect 10830 1225 10840 1240
rect 13140 1225 13150 1240
rect 13210 1270 13220 1285
rect 13210 1240 13440 1270
rect 13210 1225 13220 1240
rect 4940 1135 4950 1195
rect 5010 1180 5020 1195
rect 10970 1180 10980 1195
rect 5010 1150 10980 1180
rect 5010 1135 5020 1150
rect 10970 1135 10980 1150
rect 11040 1180 11050 1195
rect 12740 1180 12750 1195
rect 11040 1150 12750 1180
rect 11040 1135 11050 1150
rect 12740 1135 12750 1150
rect 12810 1180 12820 1195
rect 12810 1150 13440 1180
rect 12810 1135 12820 1150
rect 5180 1045 5190 1105
rect 5250 1090 5260 1105
rect 11180 1090 11190 1105
rect 5250 1060 11190 1090
rect 5250 1045 5260 1060
rect 11180 1045 11190 1060
rect 11250 1090 11260 1105
rect 13220 1090 13230 1105
rect 11250 1060 13230 1090
rect 11250 1045 11260 1060
rect 13220 1045 13230 1060
rect 13290 1090 13300 1105
rect 13290 1060 13440 1090
rect 13290 1045 13300 1060
rect 5420 955 5430 1015
rect 5490 1000 5500 1015
rect 11390 1000 11400 1015
rect 5490 970 11400 1000
rect 5490 955 5500 970
rect 11390 955 11400 970
rect 11460 1000 11470 1015
rect 12950 1000 12960 1015
rect 11460 970 12960 1000
rect 11460 955 11470 970
rect 12950 955 12960 970
rect 13020 1000 13030 1015
rect 13020 970 13440 1000
rect 13020 955 13030 970
rect 11600 865 11610 925
rect 11670 910 11680 925
rect 13300 910 13310 925
rect 11670 880 13310 910
rect 11670 865 11680 880
rect 13300 865 13310 880
rect 13370 910 13380 925
rect 13370 880 13440 910
rect 13370 865 13380 880
<< via1 >>
rect 70 3780 130 3840
rect 2120 3780 2180 3840
rect 3140 3780 3200 3840
rect 3660 3780 3720 3840
rect 3910 3780 3970 3840
rect 4150 3780 4210 3840
rect 4400 3780 4460 3840
rect 4640 3780 4700 3840
rect 4880 3780 4940 3840
rect 5130 3780 5190 3840
rect 5360 3780 5420 3840
rect -120 3490 -110 3550
rect -110 3490 -70 3550
rect -70 3490 -60 3550
rect -120 3340 -110 3400
rect -110 3340 -70 3400
rect -70 3340 -60 3400
rect -120 3190 -110 3250
rect -110 3190 -70 3250
rect -70 3190 -60 3250
rect 0 3030 60 3090
rect 260 3030 320 3090
rect 520 3030 580 3090
rect 770 3030 830 3090
rect 1030 3030 1090 3090
rect 1280 3030 1340 3090
rect 1540 3030 1600 3090
rect 1800 3030 1860 3090
rect 2050 3030 2110 3090
rect 2310 3030 2370 3090
rect 2560 3030 2620 3090
rect 2820 3030 2880 3090
rect 3080 3030 3140 3090
rect 3330 3030 3390 3090
rect 3590 3030 3650 3090
rect 3850 3030 3910 3090
rect 4090 3030 4150 3090
rect 4330 3030 4390 3090
rect 4570 3030 4630 3090
rect 4820 3030 4880 3090
rect 5060 3030 5120 3090
rect 5300 3030 5360 3090
rect 130 2160 190 2220
rect 390 2160 450 2220
rect 650 2160 710 2220
rect 900 2160 960 2220
rect 1160 2160 1220 2220
rect 1410 2160 1470 2220
rect 1670 2160 1730 2220
rect 1930 2160 1990 2220
rect 2180 2160 2240 2220
rect 2440 2160 2500 2220
rect 2690 2160 2750 2220
rect 2950 2160 3010 2220
rect 3200 2160 3260 2220
rect 3460 2160 3520 2220
rect 3720 2160 3780 2220
rect 3970 2160 4030 2220
rect 5910 3760 5970 3820
rect 6680 3760 6740 3820
rect 7070 3760 7130 3820
rect 7240 3760 7300 3820
rect 7460 3760 7520 3820
rect 7880 3760 7940 3820
rect 8650 3760 8710 3820
rect 9420 3760 9480 3820
rect 9800 3760 9860 3820
rect 9990 3760 10050 3820
rect 10200 3760 10260 3820
rect 10390 3760 10450 3820
rect 10510 3760 10570 3820
rect 10720 3760 10780 3820
rect 10930 3760 10990 3820
rect 11140 3760 11200 3820
rect 11350 3760 11410 3820
rect 7740 3640 7800 3700
rect 7930 3640 7990 3700
rect 8120 3640 8180 3700
rect 8310 3640 8370 3700
rect 8510 3640 8570 3700
rect 8700 3640 8760 3700
rect 8890 3640 8950 3700
rect 9080 3640 9140 3700
rect 9280 3640 9340 3700
rect 9470 3640 9530 3700
rect 9660 3640 9720 3700
rect 9850 3640 9910 3700
rect 10060 3540 10120 3600
rect 10250 3540 10310 3600
rect 10460 3540 10520 3600
rect 10670 3540 10730 3600
rect 10880 3540 10940 3600
rect 11090 3540 11150 3600
rect 11300 3540 11360 3600
rect 7840 3440 7900 3500
rect 8030 3440 8090 3500
rect 8220 3440 8280 3500
rect 8410 3440 8470 3500
rect 10160 3370 10220 3430
rect 10350 3370 10410 3430
rect 10560 3370 10620 3430
rect 10770 3370 10830 3430
rect 10980 3370 11040 3430
rect 11190 3380 11250 3440
rect 11400 3380 11460 3440
rect 12950 3630 13010 3690
rect 13310 3590 13370 3650
rect 11250 3230 11310 3290
rect 10210 3140 10270 3200
rect 12040 3150 12100 3210
rect 10400 3070 10460 3130
rect 11880 3070 11940 3130
rect 10510 2990 10570 3050
rect 11720 2990 11780 3050
rect 12950 3220 13010 3280
rect 13230 3190 13290 3250
rect 5640 2910 5650 2970
rect 5650 2910 5690 2970
rect 5690 2910 5700 2970
rect 10720 2910 10780 2970
rect 11960 2910 12020 2970
rect 10930 2830 10990 2890
rect 11800 2830 11860 2890
rect 5640 2750 5650 2810
rect 5650 2750 5690 2810
rect 5690 2750 5700 2810
rect 11140 2750 11200 2810
rect 11640 2750 11700 2810
rect 5640 2620 5650 2680
rect 5650 2620 5690 2680
rect 5690 2620 5700 2680
rect 5770 2620 5830 2680
rect 5960 2620 6020 2680
rect 6150 2620 6210 2680
rect 6350 2620 6410 2680
rect 6540 2620 6600 2680
rect 6730 2620 6790 2680
rect 6920 2620 6980 2680
rect 7110 2620 7170 2680
rect 11350 2670 11410 2730
rect 11480 2670 11540 2730
rect 12950 2790 13010 2850
rect 13150 2740 13210 2800
rect 4220 2130 4280 2190
rect 4460 2130 4520 2190
rect 4700 2130 4760 2190
rect 4950 2130 5010 2190
rect 5190 2130 5250 2190
rect 5430 2130 5490 2190
rect 10210 2560 10270 2620
rect 10400 2560 10460 2620
rect 10510 2560 10570 2620
rect 10720 2560 10780 2620
rect 10930 2560 10990 2620
rect 11140 2560 11200 2620
rect 11350 2560 11410 2620
rect 11560 2560 11620 2620
rect 7320 2490 7380 2550
rect 7510 2490 7570 2550
rect 10060 2450 10120 2510
rect 10250 2450 10310 2510
rect 10460 2450 10520 2510
rect 10670 2450 10730 2510
rect 10880 2450 10940 2510
rect 11090 2450 11150 2510
rect 11300 2450 11360 2510
rect 11510 2450 11570 2510
rect 11720 2450 11780 2510
rect 11910 2450 11970 2510
rect 12220 2450 12280 2510
rect 12430 2450 12490 2510
rect 12640 2450 12700 2510
rect 12850 2450 12910 2510
rect 13060 2450 13120 2510
rect 12120 2340 12180 2400
rect 12330 2340 12390 2400
rect 12540 2340 12600 2400
rect 12750 2340 12810 2400
rect 12960 2340 13020 2400
rect 5870 2180 5930 2240
rect 6060 2180 6120 2240
rect 6250 2180 6310 2240
rect 6440 2180 6500 2240
rect 6630 2180 6690 2240
rect 6830 2180 6890 2240
rect 7020 2180 7080 2240
rect 7210 2180 7270 2240
rect 7420 2180 7480 2240
rect 7610 2180 7670 2240
rect 8600 2150 8660 2210
rect 8800 2150 8860 2210
rect 8990 2150 9050 2210
rect 9180 2150 9240 2210
rect 9370 2150 9430 2210
rect 9560 2150 9620 2210
rect 9760 2150 9820 2210
rect 9950 2150 10010 2210
rect 10160 2190 10220 2250
rect 10350 2190 10410 2250
rect 10560 2190 10620 2250
rect 10770 2190 10830 2250
rect 10980 2190 11040 2250
rect 11190 2190 11250 2250
rect 11400 2190 11460 2250
rect 11610 2190 11670 2250
rect 11820 2160 11880 2220
rect 12010 2160 12070 2220
rect 130 1855 190 1915
rect 5870 1855 5930 1915
rect 7420 1855 7480 1915
rect 8600 1855 8660 1915
rect 2180 1765 2240 1825
rect 6630 1765 6690 1825
rect 7610 1765 7670 1825
rect 9370 1765 9430 1825
rect 3200 1675 3260 1735
rect 7020 1675 7080 1735
rect 9750 1675 9810 1735
rect 11820 1675 11880 1735
rect 3720 1585 3780 1645
rect 7210 1585 7270 1645
rect 9950 1585 10010 1645
rect 12010 1585 12070 1645
rect 3970 1495 4030 1555
rect 10160 1495 10220 1555
rect 12120 1495 12180 1555
rect 4220 1405 4280 1465
rect 10350 1405 10410 1465
rect 12330 1405 12390 1465
rect 4460 1315 4520 1375
rect 10560 1315 10620 1375
rect 12540 1315 12600 1375
rect 4700 1225 4760 1285
rect 10770 1225 10830 1285
rect 13150 1225 13210 1285
rect 4950 1135 5010 1195
rect 10980 1135 11040 1195
rect 12750 1135 12810 1195
rect 5190 1045 5250 1105
rect 11190 1045 11250 1105
rect 13230 1045 13290 1105
rect 5430 955 5490 1015
rect 11400 955 11460 1015
rect 12960 955 13020 1015
rect 11610 865 11670 925
rect 13310 865 13370 925
<< metal2 >>
rect 80 3850 120 4020
rect 2135 3850 2175 4090
rect 3150 3850 3190 4090
rect 3670 3850 3710 4090
rect 3920 3850 3960 4090
rect 4160 3850 4200 4090
rect 4410 3850 4450 4090
rect 4650 3850 4690 4090
rect 4890 3850 4930 4090
rect 5140 3850 5180 4090
rect 5370 3850 5410 4090
rect 60 3840 140 3850
rect 60 3780 70 3840
rect 130 3780 140 3840
rect 60 3770 140 3780
rect 2120 3840 2180 3850
rect 2120 3770 2180 3780
rect 3140 3840 3200 3850
rect 3140 3770 3200 3780
rect 3660 3840 3720 3850
rect 3660 3770 3720 3780
rect 3910 3840 3970 3850
rect 3910 3770 3970 3780
rect 4150 3840 4210 3850
rect 4150 3770 4210 3780
rect 4400 3840 4460 3850
rect 4400 3770 4460 3780
rect 4640 3840 4700 3850
rect 4640 3770 4700 3780
rect 4880 3840 4940 3850
rect 4880 3770 4940 3780
rect 5130 3840 5190 3850
rect 5130 3770 5190 3780
rect 5360 3840 5420 3850
rect 5920 3830 5960 4090
rect 6690 3830 6730 4090
rect 7080 3830 7120 4090
rect 7250 3830 7290 4090
rect 7470 3830 7510 4090
rect 7890 3830 7930 4090
rect 8660 3830 8700 4090
rect 9430 3830 9470 4090
rect 9810 3830 9850 4090
rect 10000 3830 10040 4090
rect 10210 3830 10250 4090
rect 10400 3830 10440 4090
rect 10520 3830 10560 4090
rect 10730 3830 10770 4090
rect 10940 3830 10980 4090
rect 11150 3830 11190 4090
rect 11360 3830 11400 4090
rect 5360 3770 5420 3780
rect 5910 3820 5970 3830
rect 5910 3750 5970 3760
rect 6680 3820 6740 3830
rect 6680 3750 6740 3760
rect 7070 3820 7130 3830
rect 7070 3750 7130 3760
rect 7240 3820 7300 3830
rect 7240 3750 7300 3760
rect 7460 3820 7520 3830
rect 7460 3750 7520 3760
rect 7880 3820 7940 3830
rect 7880 3750 7940 3760
rect 8650 3820 8710 3830
rect 8650 3750 8710 3760
rect 9420 3820 9480 3830
rect 9420 3750 9480 3760
rect 9800 3820 9860 3830
rect 9800 3750 9860 3760
rect 9990 3820 10050 3830
rect 9990 3750 10050 3760
rect 10200 3820 10260 3830
rect 10200 3750 10260 3760
rect 10390 3820 10450 3830
rect 10390 3750 10450 3760
rect 10510 3820 10570 3830
rect 10510 3750 10570 3760
rect 10720 3820 10780 3830
rect 10720 3750 10780 3760
rect 10930 3820 10990 3830
rect 10930 3750 10990 3760
rect 11140 3820 11200 3830
rect 11140 3750 11200 3760
rect 11350 3820 11410 3830
rect 11350 3750 11410 3760
rect 7740 3700 7800 3710
rect -200 3650 7740 3690
rect 7930 3700 7990 3710
rect 7800 3650 7930 3690
rect 7740 3630 7800 3640
rect 8120 3700 8180 3710
rect 7990 3650 8120 3690
rect 7930 3630 7990 3640
rect 8310 3700 8370 3710
rect 8180 3650 8310 3690
rect 8120 3630 8180 3640
rect 8510 3700 8570 3710
rect 8370 3650 8510 3690
rect 8310 3630 8370 3640
rect 8700 3700 8760 3710
rect 8570 3650 8700 3690
rect 8510 3630 8570 3640
rect 8890 3700 8950 3710
rect 8760 3650 8890 3690
rect 8700 3630 8760 3640
rect 9080 3700 9140 3710
rect 8950 3650 9080 3690
rect 8890 3630 8950 3640
rect 9280 3700 9340 3710
rect 9140 3650 9280 3690
rect 9080 3630 9140 3640
rect 9470 3700 9530 3710
rect 9340 3650 9470 3690
rect 9280 3630 9340 3640
rect 9660 3700 9720 3710
rect 9530 3650 9660 3690
rect 9470 3630 9530 3640
rect 9850 3700 9910 3710
rect 9720 3650 9850 3690
rect 9850 3630 9910 3640
rect 9660 3620 9720 3630
rect 10060 3600 10120 3610
rect 9850 3580 10060 3590
rect -120 3550 -60 3560
rect 9910 3540 10060 3580
rect 10250 3600 10310 3610
rect 10120 3550 10250 3590
rect 10070 3530 10120 3540
rect 10460 3600 10520 3610
rect 10310 3550 10460 3590
rect 10250 3530 10310 3540
rect 10670 3600 10730 3610
rect 10520 3550 10670 3590
rect 10460 3530 10520 3540
rect 10880 3600 10940 3610
rect 10730 3550 10880 3590
rect 10670 3530 10730 3540
rect 11090 3600 11150 3610
rect 10940 3550 11090 3590
rect 10880 3530 10940 3540
rect 11300 3600 11360 3610
rect 11150 3550 11300 3590
rect 11090 3530 11150 3540
rect 11300 3530 11360 3540
rect 9850 3510 9910 3520
rect -120 3400 -60 3490
rect 7840 3500 7900 3510
rect 8030 3500 8090 3510
rect 7900 3450 8030 3490
rect 7840 3430 7900 3440
rect 8130 3500 8190 3510
rect 8090 3450 8130 3490
rect 8030 3430 8090 3440
rect 8220 3500 8280 3510
rect 8190 3450 8220 3490
rect 8130 3430 8190 3440
rect 8410 3500 8470 3510
rect 8280 3450 8410 3490
rect 8220 3430 8280 3440
rect 11190 3440 11250 3450
rect 8410 3430 8470 3440
rect 10160 3430 10220 3440
rect -180 3350 -120 3390
rect 10160 3360 10220 3370
rect 10350 3430 10410 3440
rect 10350 3360 10410 3370
rect 10560 3430 10620 3440
rect 10560 3360 10620 3370
rect 10770 3430 10830 3440
rect 10770 3360 10830 3370
rect 10980 3430 11040 3440
rect 11190 3370 11250 3380
rect 11400 3440 11460 3450
rect 11400 3370 11460 3380
rect 10980 3360 11040 3370
rect -120 3250 -60 3340
rect 7460 3290 7520 3300
rect 11250 3290 11310 3300
rect 7520 3240 11250 3280
rect 7460 3220 7520 3230
rect 11250 3220 11310 3230
rect -120 3180 -60 3190
rect 10210 3200 10270 3210
rect 10210 3130 10270 3140
rect 10400 3130 10460 3140
rect 0 3090 60 3100
rect -180 3040 0 3080
rect 260 3090 320 3100
rect 60 3040 260 3080
rect 0 3020 60 3030
rect 520 3090 580 3100
rect 320 3040 520 3080
rect 260 3020 320 3030
rect 770 3090 830 3100
rect 580 3040 770 3080
rect 520 3020 580 3030
rect 1030 3090 1090 3100
rect 830 3040 1030 3080
rect 770 3020 830 3030
rect 1280 3090 1340 3100
rect 1090 3040 1280 3080
rect 1030 3020 1090 3030
rect 1540 3090 1600 3100
rect 1340 3040 1540 3080
rect 1280 3020 1340 3030
rect 1800 3090 1860 3100
rect 1600 3040 1800 3080
rect 1540 3020 1600 3030
rect 2050 3090 2110 3100
rect 1860 3040 2050 3080
rect 1800 3020 1860 3030
rect 2310 3090 2370 3100
rect 2110 3040 2310 3080
rect 2050 3020 2110 3030
rect 2560 3090 2620 3100
rect 2370 3040 2560 3080
rect 2310 3020 2370 3030
rect 2820 3090 2880 3100
rect 2620 3040 2820 3080
rect 2560 3020 2620 3030
rect 3080 3090 3140 3100
rect 2880 3040 3080 3080
rect 2820 3020 2880 3030
rect 3330 3090 3390 3100
rect 3140 3040 3330 3080
rect 3080 3020 3140 3030
rect 3590 3090 3650 3100
rect 3390 3040 3590 3080
rect 3330 3020 3390 3030
rect 3850 3090 3910 3100
rect 3650 3040 3850 3080
rect 3590 3020 3650 3030
rect 4090 3090 4150 3100
rect 3910 3040 4090 3080
rect 3850 3020 3910 3030
rect 4330 3090 4390 3100
rect 4150 3040 4330 3080
rect 4090 3020 4150 3030
rect 4570 3090 4630 3100
rect 4390 3040 4570 3080
rect 4330 3020 4390 3030
rect 4820 3090 4880 3100
rect 4630 3040 4820 3080
rect 4570 3020 4630 3030
rect 5060 3090 5120 3100
rect 4880 3040 5060 3080
rect 4820 3020 4880 3030
rect 5300 3090 5360 3100
rect 5120 3040 5300 3080
rect 5060 3020 5120 3030
rect 5300 3020 5360 3030
rect 7110 3060 7170 3070
rect 9850 3060 9910 3070
rect 7170 3010 9850 3050
rect 7110 2990 7170 3000
rect 9850 2990 9910 3000
rect 5640 2970 5700 2980
rect 5640 2810 5700 2910
rect 5640 2680 5700 2750
rect -200 2630 5640 2670
rect 5770 2680 5830 2690
rect 5700 2630 5770 2670
rect 5640 2610 5700 2620
rect 5960 2680 6020 2690
rect 5830 2630 5960 2670
rect 5770 2610 5830 2620
rect 6150 2680 6210 2690
rect 6020 2630 6150 2670
rect 5960 2610 6020 2620
rect 6350 2680 6410 2690
rect 6210 2630 6350 2670
rect 6150 2610 6210 2620
rect 6540 2680 6600 2690
rect 6410 2630 6540 2670
rect 6350 2610 6410 2620
rect 6730 2680 6790 2690
rect 6600 2630 6730 2670
rect 6540 2610 6600 2620
rect 6920 2680 6980 2690
rect 6790 2630 6920 2670
rect 6730 2610 6790 2620
rect 7110 2680 7170 2690
rect 6980 2630 7110 2670
rect 6920 2610 6980 2620
rect 10220 2630 10260 3130
rect 10400 3060 10460 3070
rect 10410 2630 10450 3060
rect 10510 3050 10570 3060
rect 10510 2980 10570 2990
rect 10520 2630 10560 2980
rect 10720 2970 10780 2980
rect 10720 2900 10780 2910
rect 10730 2630 10770 2900
rect 10930 2890 10990 2900
rect 10930 2820 10990 2830
rect 10940 2630 10980 2820
rect 11140 2810 11200 2820
rect 11140 2740 11200 2750
rect 11490 2740 11530 4090
rect 11150 2630 11190 2740
rect 11350 2730 11410 2740
rect 11350 2660 11410 2670
rect 11480 2730 11540 2740
rect 11480 2660 11540 2670
rect 11360 2630 11400 2660
rect 11570 2630 11610 4090
rect 11650 2820 11690 4090
rect 11730 3060 11770 4090
rect 11720 3050 11780 3060
rect 11720 2980 11780 2990
rect 11810 2900 11850 4090
rect 11890 3140 11930 4090
rect 11880 3130 11940 3140
rect 11880 3060 11940 3070
rect 11970 2980 12010 4090
rect 12050 3220 12090 4090
rect 12950 3690 13010 3700
rect 12950 3620 13010 3630
rect 13310 3650 13370 3660
rect 12960 3290 12990 3620
rect 13310 3580 13370 3590
rect 12950 3280 13010 3290
rect 12040 3210 12100 3220
rect 12950 3210 13010 3220
rect 13230 3250 13290 3260
rect 12040 3140 12100 3150
rect 11960 2970 12020 2980
rect 11960 2900 12020 2910
rect 11800 2890 11860 2900
rect 12960 2860 12990 3210
rect 13230 3180 13290 3190
rect 11800 2820 11860 2830
rect 12950 2850 13010 2860
rect 11640 2810 11700 2820
rect 12950 2780 13010 2790
rect 13150 2800 13210 2810
rect 11640 2740 11700 2750
rect 7110 2610 7170 2620
rect 10210 2620 10270 2630
rect 7320 2550 7380 2560
rect -200 2500 7320 2540
rect 7510 2550 7570 2560
rect 10210 2550 10270 2560
rect 10400 2620 10460 2630
rect 10400 2550 10460 2560
rect 10510 2620 10570 2630
rect 10510 2550 10570 2560
rect 10720 2620 10780 2630
rect 10720 2550 10780 2560
rect 10930 2620 10990 2630
rect 10930 2550 10990 2560
rect 11140 2620 11200 2630
rect 11140 2550 11200 2560
rect 11350 2620 11410 2630
rect 11350 2550 11410 2560
rect 11560 2620 11620 2630
rect 11560 2550 11620 2560
rect 7380 2500 7510 2540
rect 7320 2480 7380 2490
rect 7505 2490 7510 2500
rect 7505 2480 7570 2490
rect 9660 2510 9720 2520
rect 10060 2510 10120 2520
rect 10250 2510 10310 2520
rect 10460 2510 10520 2520
rect 10670 2510 10730 2520
rect 10880 2510 10940 2520
rect 11090 2510 11150 2520
rect 11300 2510 11360 2520
rect 11510 2510 11570 2520
rect 7505 2370 7555 2480
rect 9720 2450 10060 2510
rect 10120 2450 10250 2510
rect 10310 2450 10460 2510
rect 10520 2450 10670 2510
rect 10730 2450 10880 2510
rect 10940 2450 11090 2510
rect 11150 2450 11300 2510
rect 11360 2450 11510 2510
rect 9660 2440 9720 2450
rect 10060 2440 10120 2450
rect 10250 2440 10310 2450
rect 10460 2440 10520 2450
rect 10670 2440 10730 2450
rect 10880 2440 10940 2450
rect 11090 2440 11150 2450
rect 11300 2440 11360 2450
rect 11510 2440 11570 2450
rect 11720 2510 11780 2520
rect 11910 2510 11970 2520
rect 11780 2460 11910 2500
rect 11720 2440 11780 2450
rect 12220 2510 12280 2520
rect 11970 2460 12220 2500
rect 11910 2440 11970 2450
rect 12430 2510 12490 2520
rect 12280 2460 12430 2500
rect 12220 2440 12280 2450
rect 12640 2510 12700 2520
rect 12490 2460 12640 2500
rect 12430 2440 12490 2450
rect 12850 2510 12910 2520
rect 12700 2460 12850 2500
rect 12640 2440 12700 2450
rect 12960 2500 12990 2780
rect 13150 2730 13210 2740
rect 13060 2510 13120 2520
rect 12910 2460 13060 2500
rect 12850 2440 12910 2450
rect 13060 2440 13120 2450
rect 11740 2370 11770 2440
rect 7505 2320 11770 2370
rect 12120 2400 12180 2410
rect 12120 2330 12180 2340
rect 12330 2400 12390 2410
rect 12330 2330 12390 2340
rect 12540 2400 12600 2410
rect 12540 2330 12600 2340
rect 12750 2400 12810 2410
rect 12750 2330 12810 2340
rect 12960 2400 13020 2410
rect 12960 2330 13020 2340
rect 10160 2250 10220 2260
rect 5870 2240 5930 2250
rect 130 2220 190 2230
rect 390 2220 450 2230
rect 190 2170 390 2210
rect 130 2150 190 2160
rect 650 2220 710 2230
rect 450 2170 650 2210
rect 390 2150 450 2160
rect 900 2220 960 2230
rect 710 2170 900 2210
rect 650 2150 710 2160
rect 1160 2220 1220 2230
rect 960 2170 1160 2210
rect 900 2150 960 2160
rect 1410 2220 1470 2230
rect 1220 2170 1410 2210
rect 1160 2150 1220 2160
rect 1670 2220 1730 2230
rect 1470 2170 1670 2210
rect 1410 2150 1470 2160
rect 1930 2220 1990 2230
rect 1730 2170 1930 2210
rect 1670 2150 1730 2160
rect 1930 2150 1990 2160
rect 2180 2220 2240 2230
rect 2440 2220 2500 2230
rect 2240 2170 2440 2210
rect 2180 2150 2240 2160
rect 2690 2220 2750 2230
rect 2500 2170 2690 2210
rect 2440 2150 2500 2160
rect 2950 2220 3010 2230
rect 2750 2170 2950 2210
rect 2690 2150 2750 2160
rect 2950 2150 3010 2160
rect 3200 2220 3260 2230
rect 3460 2220 3520 2230
rect 3260 2170 3460 2210
rect 3200 2150 3260 2160
rect 3460 2150 3520 2160
rect 3720 2220 3780 2230
rect 3720 2150 3780 2160
rect 3970 2220 4030 2230
rect 3970 2150 4030 2160
rect 4220 2190 4280 2200
rect 140 1925 180 2150
rect 130 1915 190 1925
rect 130 1845 190 1855
rect 2190 1835 2230 2150
rect 2180 1825 2240 1835
rect 2180 1755 2240 1765
rect 3210 1745 3250 2150
rect 3200 1735 3260 1745
rect 3200 1665 3260 1675
rect 3730 1655 3770 2150
rect 3720 1645 3780 1655
rect 3720 1575 3780 1585
rect 3980 1565 4020 2150
rect 4220 2120 4280 2130
rect 4460 2190 4520 2200
rect 4460 2120 4520 2130
rect 4700 2190 4760 2200
rect 4700 2120 4760 2130
rect 4950 2190 5010 2200
rect 4950 2120 5010 2130
rect 5190 2190 5250 2200
rect 5190 2120 5250 2130
rect 5430 2190 5490 2200
rect 6060 2240 6120 2250
rect 5930 2190 6060 2230
rect 5870 2170 5930 2180
rect 6250 2240 6310 2250
rect 6120 2190 6250 2230
rect 6060 2170 6120 2180
rect 6440 2240 6500 2250
rect 6310 2190 6440 2230
rect 6250 2170 6310 2180
rect 6440 2170 6500 2180
rect 6630 2240 6690 2250
rect 6830 2240 6890 2250
rect 6690 2190 6830 2230
rect 6630 2170 6690 2180
rect 6830 2170 6890 2180
rect 7020 2240 7080 2250
rect 7020 2170 7080 2180
rect 7210 2240 7270 2250
rect 7210 2170 7270 2180
rect 7420 2240 7480 2250
rect 7420 2170 7480 2180
rect 7610 2240 7670 2250
rect 7610 2170 7670 2180
rect 8600 2210 8660 2220
rect 5430 2120 5490 2130
rect 3970 1555 4030 1565
rect 3970 1485 4030 1495
rect 4230 1475 4270 2120
rect 4220 1465 4280 1475
rect 4220 1395 4280 1405
rect 4470 1385 4510 2120
rect 4460 1375 4520 1385
rect 4460 1305 4520 1315
rect 4710 1295 4750 2120
rect 4700 1285 4760 1295
rect 4700 1215 4760 1225
rect 4960 1205 5000 2120
rect 4950 1195 5010 1205
rect 4950 1125 5010 1135
rect 5200 1115 5240 2120
rect 5190 1105 5250 1115
rect 5190 1035 5250 1045
rect 5440 1025 5480 2120
rect 5880 1925 5920 2170
rect 5870 1915 5930 1925
rect 5870 1845 5930 1855
rect 6640 1835 6680 2170
rect 6630 1825 6690 1835
rect 6630 1755 6690 1765
rect 7030 1745 7070 2170
rect 7020 1735 7080 1745
rect 7020 1665 7080 1675
rect 7220 1655 7260 2170
rect 7430 1925 7470 2170
rect 7420 1915 7480 1925
rect 7420 1845 7480 1855
rect 7620 1835 7660 2170
rect 8800 2210 8860 2220
rect 8660 2160 8800 2200
rect 8600 2140 8660 2150
rect 8990 2210 9050 2220
rect 8860 2160 8990 2200
rect 8800 2140 8860 2150
rect 9180 2210 9240 2220
rect 9050 2160 9180 2200
rect 8990 2140 9050 2150
rect 9180 2140 9240 2150
rect 9370 2210 9430 2220
rect 9560 2210 9620 2220
rect 9430 2160 9560 2200
rect 9370 2140 9430 2150
rect 9560 2140 9620 2150
rect 9760 2210 9820 2220
rect 9760 2140 9820 2150
rect 9950 2210 10010 2220
rect 10160 2180 10220 2190
rect 10350 2250 10410 2260
rect 10350 2180 10410 2190
rect 10560 2250 10620 2260
rect 10560 2180 10620 2190
rect 10770 2250 10830 2260
rect 10770 2180 10830 2190
rect 10980 2250 11040 2260
rect 10980 2180 11040 2190
rect 11190 2250 11250 2260
rect 11190 2180 11250 2190
rect 11400 2250 11460 2260
rect 11400 2180 11460 2190
rect 11610 2250 11670 2260
rect 11610 2180 11670 2190
rect 11820 2220 11880 2230
rect 9950 2140 10010 2150
rect 8610 1925 8650 2140
rect 8600 1915 8660 1925
rect 8600 1845 8660 1855
rect 9380 1835 9420 2140
rect 7610 1825 7670 1835
rect 7610 1755 7670 1765
rect 9370 1825 9430 1835
rect 9370 1755 9430 1765
rect 9760 1745 9800 2140
rect 9750 1735 9810 1745
rect 9750 1665 9810 1675
rect 9960 1655 10000 2140
rect 7210 1645 7270 1655
rect 7210 1575 7270 1585
rect 9950 1645 10010 1655
rect 9950 1575 10010 1585
rect 10170 1565 10210 2180
rect 10160 1555 10220 1565
rect 10160 1485 10220 1495
rect 10360 1475 10400 2180
rect 10350 1465 10410 1475
rect 10350 1395 10410 1405
rect 10570 1385 10610 2180
rect 10560 1375 10620 1385
rect 10560 1305 10620 1315
rect 10780 1295 10820 2180
rect 10770 1285 10830 1295
rect 10770 1215 10830 1225
rect 10990 1205 11030 2180
rect 10980 1195 11040 1205
rect 10980 1125 11040 1135
rect 11200 1115 11240 2180
rect 11190 1105 11250 1115
rect 11190 1035 11250 1045
rect 11410 1025 11450 2180
rect 5430 1015 5490 1025
rect 5430 945 5490 955
rect 11400 1015 11460 1025
rect 11400 945 11460 955
rect 11620 935 11660 2180
rect 11820 2150 11880 2160
rect 12010 2220 12070 2230
rect 12010 2150 12070 2160
rect 11830 1745 11870 2150
rect 11820 1735 11880 1745
rect 11820 1665 11880 1675
rect 12020 1655 12060 2150
rect 12010 1645 12070 1655
rect 12010 1575 12070 1585
rect 12130 1565 12170 2330
rect 12120 1555 12180 1565
rect 12120 1485 12180 1495
rect 12340 1475 12380 2330
rect 12330 1465 12390 1475
rect 12330 1395 12390 1405
rect 12550 1385 12590 2330
rect 12540 1375 12600 1385
rect 12540 1305 12600 1315
rect 12760 1205 12800 2330
rect 12750 1195 12810 1205
rect 12750 1125 12810 1135
rect 12970 1025 13010 2330
rect 13160 1295 13200 2730
rect 13150 1285 13210 1295
rect 13150 1215 13210 1225
rect 13240 1115 13280 3180
rect 13230 1105 13290 1115
rect 13230 1035 13290 1045
rect 12960 1015 13020 1025
rect 12960 945 13020 955
rect 13320 935 13360 3580
rect 11610 925 11670 935
rect 11610 855 11670 865
rect 13310 925 13370 935
rect 13310 855 13370 865
<< via2 >>
rect 7460 3760 7520 3820
rect 9660 3640 9720 3700
rect 9660 3630 9720 3640
rect 9850 3520 9910 3580
rect 8130 3440 8190 3500
rect 10160 3370 10220 3430
rect 10350 3370 10410 3430
rect 10560 3370 10620 3430
rect 10770 3370 10830 3430
rect 10980 3370 11040 3430
rect 11190 3380 11250 3440
rect 11400 3380 11460 3440
rect 7460 3230 7520 3290
rect 7110 3000 7170 3060
rect 9850 3000 9910 3060
rect 7110 2620 7170 2680
rect 9660 2450 9720 2510
rect 10160 2190 10220 2250
rect 10350 2190 10410 2250
rect 10560 2190 10620 2250
rect 10770 2190 10830 2250
rect 10980 2190 11040 2250
rect 11190 2190 11250 2250
rect 11400 2190 11460 2250
<< metal3 >>
rect 7450 3820 7530 3825
rect 7450 3760 7460 3820
rect 7520 3760 7530 3820
rect 7450 3290 7530 3760
rect 9650 3700 9730 3705
rect 9650 3630 9660 3700
rect 9720 3630 9730 3700
rect 8110 3510 8210 3520
rect 8110 3430 8120 3510
rect 8200 3430 8210 3510
rect 8110 3420 8210 3430
rect 7450 3230 7460 3290
rect 7520 3230 7530 3290
rect 7450 3220 7530 3230
rect 7100 3060 7180 3070
rect 7100 3000 7110 3060
rect 7170 3000 7180 3060
rect 7100 2680 7180 3000
rect 7100 2620 7110 2680
rect 7170 2620 7180 2680
rect 7100 2610 7180 2620
rect 9650 2510 9730 3630
rect 9840 3580 9920 3585
rect 9840 3520 9850 3580
rect 9910 3520 9920 3580
rect 9840 3060 9920 3520
rect 11180 3440 11260 3445
rect 9840 3000 9850 3060
rect 9910 3000 9920 3060
rect 9840 2990 9920 3000
rect 10150 3430 10230 3440
rect 10150 3370 10160 3430
rect 10220 3370 10230 3430
rect 9650 2450 9660 2510
rect 9720 2450 9730 2510
rect 9650 2440 9730 2450
rect 10150 2250 10230 3370
rect 10150 2190 10160 2250
rect 10220 2190 10230 2250
rect 10150 2180 10230 2190
rect 10340 3430 10420 3440
rect 10340 3370 10350 3430
rect 10410 3370 10420 3430
rect 10340 2250 10420 3370
rect 10340 2190 10350 2250
rect 10410 2190 10420 2250
rect 10340 2180 10420 2190
rect 10550 3430 10630 3440
rect 10550 3370 10560 3430
rect 10620 3370 10630 3430
rect 10550 2250 10630 3370
rect 10550 2190 10560 2250
rect 10620 2190 10630 2250
rect 10550 2180 10630 2190
rect 10760 3430 10840 3440
rect 10760 3370 10770 3430
rect 10830 3370 10840 3430
rect 10760 2250 10840 3370
rect 10760 2190 10770 2250
rect 10830 2190 10840 2250
rect 10760 2180 10840 2190
rect 10970 3430 11050 3440
rect 10970 3370 10980 3430
rect 11040 3370 11050 3430
rect 10970 2250 11050 3370
rect 10970 2190 10980 2250
rect 11040 2190 11050 2250
rect 10970 2180 11050 2190
rect 11180 3380 11190 3440
rect 11250 3380 11260 3440
rect 11180 2250 11260 3380
rect 11180 2190 11190 2250
rect 11250 2190 11260 2250
rect 11180 2180 11260 2190
rect 11390 3440 11470 3445
rect 11390 3380 11400 3440
rect 11460 3380 11470 3440
rect 11390 2250 11470 3380
rect 11390 2190 11400 2250
rect 11460 2190 11470 2250
rect 11390 2180 11470 2190
<< via3 >>
rect 8120 3500 8200 3510
rect 8120 3440 8130 3500
rect 8130 3440 8190 3500
rect 8190 3440 8200 3500
rect 8120 3430 8200 3440
<< metal4 >>
rect 8110 3510 8210 3520
rect 8110 3430 8120 3510
rect 8200 3430 8210 3510
rect 8110 3420 8210 3430
use sky130_fd_pr__nfet_01v8_4AP47J  sky130_fd_pr__nfet_01v8_4AP47J_0
timestamp 1711821647
transform 1 0 12932 0 1 2289
box -812 18 182 1558
use sky130_fd_pr__nfet_01v8_BG2JC8  sky130_fd_pr__nfet_01v8_BG2JC8_0
timestamp 1711813427
transform 1 0 11893 0 1 2333
box -173 -226 245 299
use sky130_fd_pr__nfet_01v8_BG2JC8  sky130_fd_pr__nfet_01v8_BG2JC8_1
timestamp 1711813427
transform 1 0 10233 0 1 3532
box -173 -226 245 299
use sky130_fd_pr__nfet_01v8_CA2JC5  sky130_fd_pr__nfet_01v8_CA2JC5_0
timestamp 1711802150
transform 1 0 7497 0 1 2932
box -173 -826 215 901
use sky130_fd_pr__nfet_01v8_D6PFL8  sky130_fd_pr__nfet_01v8_D6PFL8_0
timestamp 1711827946
transform 1 0 6520 0 1 2932
box -887 -940 6957 1030
use sky130_fd_pr__nfet_01v8_KJP4PL  sky130_fd_pr__nfet_01v8_KJP4PL_0
timestamp 1711814111
transform 1 0 11062 0 1 3532
box -602 -226 392 288
use sky130_fd_pr__nfet_01v8_lvt_HYT5PW  sky130_fd_pr__nfet_01v8_lvt_HYT5PW_0
timestamp 1711813510
transform 1 0 10233 0 1 2332
box -173 -226 234 294
use sky130_fd_pr__nfet_01v8_lvt_KJGFCE  sky130_fd_pr__nfet_01v8_lvt_KJGFCE_0
timestamp 1711814111
transform 1 0 11062 0 1 2332
box -602 -226 602 292
use sky130_fd_pr__nfet_01v8_lvt_PPAFQT  sky130_fd_pr__nfet_01v8_lvt_PPAFQT_0
timestamp 1711802774
transform 1 0 8873 0 1 2932
box -1133 -826 1209 905
use sky130_fd_pr__pfet_01v8_lvt_BA634A  sky130_fd_pr__pfet_01v8_lvt_BA634A_0
timestamp 1711799238
transform 1 0 4790 0 1 3376
box -734 -498 734 464
use sky130_fd_pr__pfet_01v8_lvt_D3D366  sky130_fd_pr__pfet_01v8_lvt_D3D366_0
timestamp 1711827888
transform 1 0 2020 0 1 2976
box -2151 -986 3611 984
<< labels >>
rlabel metal2 3150 4050 3190 4090 1 EN_VREF_Z[8]
port 3 n
rlabel metal2 3670 4050 3710 4090 1 EN_VREF_Z[7]
port 4 n
rlabel metal2 3920 4050 3960 4090 1 EN_VREF_Z[6]
port 5 n
rlabel metal2 4160 4050 4200 4090 1 EN_VREF_Z[5]
port 6 n
rlabel metal2 4410 4050 4450 4090 1 EN_VREF_Z[4]
port 7 n
rlabel metal2 4650 4050 4690 4090 1 EN_VREF_Z[3]
port 8 n
rlabel metal2 4890 4050 4930 4090 1 EN_VREF_Z[2]
port 9 n
rlabel metal2 5140 4050 5180 4090 1 EN_VREF_Z[1]
port 10 n
rlabel metal2 5370 4050 5410 4090 1 EN_VREF_Z[0]
port 11 n
rlabel metal1 13400 880 13430 910 1 Cbtm_0_dummy
port 12 n
rlabel metal1 13400 970 13430 1000 1 Cbtm_0
port 13 n
rlabel metal1 13400 1060 13430 1090 1 Cbtm_1
port 14 n
rlabel metal1 13400 1150 13430 1180 1 Cbtm_2
port 15 n
rlabel metal1 13400 1240 13430 1270 1 Cbtm_3
port 16 n
rlabel metal1 13400 1330 13430 1360 1 Cbtm_4
port 17 n
rlabel metal1 13400 1420 13430 1450 1 Cbtm_5
port 18 n
rlabel metal1 13400 1510 13430 1540 1 Cbtm_6
port 19 n
rlabel metal1 13400 1600 13430 1630 1 Cbtm_7
port 20 n
rlabel metal1 13400 1690 13430 1720 1 Cbtm_8
port 21 n
rlabel metal1 13400 1780 13430 1810 1 Cbtm_9
port 22 n
rlabel metal1 13400 1870 13430 1900 1 Cbtm_10
port 23 n
rlabel metal2 5920 4050 5960 4090 1 EN_VSS[10]
port 28 n
rlabel metal2 6690 4050 6730 4090 1 EN_VSS[9]
port 29 n
rlabel metal2 7080 4050 7120 4090 1 EN_VSS[8]
port 30 n
rlabel metal2 7250 4050 7290 4090 1 EN_VSS[7]
port 31 n
rlabel metal2 7470 4050 7510 4090 1 EN_VIN
port 32 n
rlabel metal2 7890 4050 7930 4090 1 EN_VCM_SW
port 33 n
rlabel metal2 8660 4050 8700 4090 1 EN_VCM[10]
port 34 n
rlabel metal2 9430 4050 9470 4090 1 EN_VCM[9]
port 35 n
rlabel metal2 9810 4050 9850 4090 1 EN_VCM[8]
port 36 n
rlabel metal2 10000 4050 10040 4090 1 EN_VCM[7]
port 37 n
rlabel metal2 10210 4050 10250 4090 1 EN_VSS[6]
port 38 n
rlabel metal2 10400 4050 10440 4090 1 EN_VSS[5]
port 39 n
rlabel metal2 10520 4050 10560 4090 1 EN_VSS[4]
port 40 n
rlabel metal2 10730 4050 10770 4090 1 EN_VSS[3]
port 41 n
rlabel metal2 10940 4050 10980 4090 1 EN_VSS[2]
port 42 n
rlabel metal2 11150 4050 11190 4090 1 EN_VSS[1]
port 43 n
rlabel metal2 11360 4050 11400 4090 1 EN_VSS[0]
port 44 n
rlabel metal2 11490 4050 11530 4090 1 EN_VCM[0]
port 45 n
rlabel metal2 11570 4050 11610 4090 1 EN_VCM_DUMMY
port 46 n
rlabel metal2 11650 4050 11690 4090 1 EN_VCM[1]
port 47 n
rlabel metal2 11730 4050 11770 4090 1 EN_VCM[4]
port 48 n
rlabel metal2 11810 4050 11850 4090 1 EN_VCM[2]
port 49 n
rlabel metal2 11890 4050 11930 4090 1 EN_VCM[5]
port 50 n
rlabel metal2 11970 4050 12010 4090 1 EN_VCM[3]
port 51 n
rlabel metal2 12050 4050 12090 4090 1 EN_VCM[6]
port 52 n
rlabel metal4 8120 3430 8200 3510 1 VDAC
port 54 n
rlabel metal2 2135 4050 2175 4090 1 EN_VREF_Z[9]
port 2 n
rlabel metal2 -180 3350 -140 3390 1 VDD
port 53 n
rlabel metal2 -200 3650 -160 3690 1 VCM
port 27 n
rlabel metal2 -180 3040 -140 3080 1 VREF
port 26 n
rlabel metal2 -200 2630 -160 2670 1 VSS
port 25 n
rlabel metal2 -200 2500 -160 2540 1 VIN
port 24 n
rlabel metal2 80 3980 120 4020 1 EN_VREF_Z[10]
port 1 n
<< end >>
