magic
tech sky130A
magscale 1 2
timestamp 1711883479
<< error_p >>
rect 19 872 77 878
rect 19 838 31 872
rect 19 832 77 838
rect -77 -838 -19 -832
rect -77 -872 -65 -838
rect -77 -878 -19 -872
<< pwell >>
rect -263 -1010 263 1010
<< nmos >>
rect -63 -800 -33 800
rect 33 -800 63 800
<< ndiff >>
rect -125 788 -63 800
rect -125 -788 -113 788
rect -79 -788 -63 788
rect -125 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 125 800
rect 63 -788 79 788
rect 113 -788 125 788
rect 63 -800 125 -788
<< ndiffc >>
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
<< psubdiff >>
rect -227 940 -131 974
rect 131 940 227 974
rect -227 878 -193 940
rect 193 878 227 940
rect -227 -940 -193 -878
rect 193 -940 227 -878
rect -227 -974 -131 -940
rect 131 -974 227 -940
<< psubdiffcont >>
rect -131 940 131 974
rect -227 -878 -193 878
rect 193 -878 227 878
rect -131 -974 131 -940
<< poly >>
rect 15 872 81 888
rect 15 838 31 872
rect 65 838 81 872
rect -63 800 -33 826
rect 15 822 81 838
rect 33 800 63 822
rect -63 -822 -33 -800
rect -81 -838 -15 -822
rect 33 -826 63 -800
rect -81 -872 -65 -838
rect -31 -872 -15 -838
rect -81 -888 -15 -872
<< polycont >>
rect 31 838 65 872
rect -65 -872 -31 -838
<< locali >>
rect -227 940 -131 974
rect 131 940 227 974
rect -227 878 -193 940
rect 193 878 227 940
rect 15 838 31 872
rect 65 838 81 872
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect -81 -872 -65 -838
rect -31 -872 -15 -838
rect -227 -940 -193 -878
rect 193 -940 227 -878
rect -227 -974 -131 -940
rect 131 -974 227 -940
<< viali >>
rect 31 838 65 872
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect -65 -872 -31 -838
<< metal1 >>
rect 19 872 77 878
rect 19 838 31 872
rect 65 838 77 872
rect 19 832 77 838
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect -77 -838 -19 -832
rect -77 -872 -65 -838
rect -31 -872 -19 -838
rect -77 -878 -19 -872
<< properties >>
string FIXED_BBOX -210 -957 210 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8.0 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
