magic
tech sky130A
magscale 1 2
timestamp 1711883049
<< error_p >>
rect -77 272 -19 278
rect 115 272 173 278
rect -77 238 -65 272
rect 115 238 127 272
rect -77 232 -19 238
rect 115 232 173 238
rect -173 -238 -115 -232
rect 19 -238 77 -232
rect -173 -272 -161 -238
rect 19 -272 31 -238
rect -173 -278 -115 -272
rect 19 -278 77 -272
<< pwell >>
rect -359 -410 359 410
<< nmos >>
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
<< ndiff >>
rect -221 188 -159 200
rect -221 -188 -209 188
rect -175 -188 -159 188
rect -221 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 221 200
rect 159 -188 175 188
rect 209 -188 221 188
rect 159 -200 221 -188
<< ndiffc >>
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
<< psubdiff >>
rect -323 340 -227 374
rect 227 340 323 374
rect -323 278 -289 340
rect 289 278 323 340
rect -323 -340 -289 -278
rect 289 -340 323 -278
rect -323 -374 -227 -340
rect 227 -374 323 -340
<< psubdiffcont >>
rect -227 340 227 374
rect -323 -278 -289 278
rect 289 -278 323 278
rect -227 -374 227 -340
<< poly >>
rect -81 272 -15 288
rect -81 238 -65 272
rect -31 238 -15 272
rect -159 200 -129 226
rect -81 222 -15 238
rect 111 272 177 288
rect 111 238 127 272
rect 161 238 177 272
rect -63 200 -33 222
rect 33 200 63 226
rect 111 222 177 238
rect 129 200 159 222
rect -159 -222 -129 -200
rect -177 -238 -111 -222
rect -63 -226 -33 -200
rect 33 -222 63 -200
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect -177 -288 -111 -272
rect 15 -238 81 -222
rect 129 -226 159 -200
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 15 -288 81 -272
<< polycont >>
rect -65 238 -31 272
rect 127 238 161 272
rect -161 -272 -127 -238
rect 31 -272 65 -238
<< locali >>
rect -323 340 -227 374
rect 227 340 323 374
rect -323 278 -289 340
rect 289 278 323 340
rect -81 238 -65 272
rect -31 238 -15 272
rect 111 238 127 272
rect 161 238 177 272
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect 15 -272 31 -238
rect 65 -272 81 -238
rect -323 -340 -289 -278
rect 289 -340 323 -278
rect -323 -374 -227 -340
rect 227 -374 323 -340
<< viali >>
rect -65 238 -31 272
rect 127 238 161 272
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect -161 -272 -127 -238
rect 31 -272 65 -238
<< metal1 >>
rect -77 272 -19 278
rect -77 238 -65 272
rect -31 238 -19 272
rect -77 232 -19 238
rect 115 272 173 278
rect 115 238 127 272
rect 161 238 173 272
rect 115 232 173 238
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect -173 -238 -115 -232
rect -173 -272 -161 -238
rect -127 -272 -115 -238
rect -173 -278 -115 -272
rect 19 -238 77 -232
rect 19 -272 31 -238
rect 65 -272 77 -238
rect 19 -278 77 -272
<< properties >>
string FIXED_BBOX -306 -357 306 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
