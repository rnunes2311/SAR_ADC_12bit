magic
tech sky130A
magscale 1 2
timestamp 1711798895
<< error_p >>
rect -351 445 -289 451
rect -223 445 -161 451
rect -95 445 -33 451
rect 33 445 95 451
rect 161 445 223 451
rect 289 445 351 451
rect -351 411 -339 445
rect -223 411 -211 445
rect -95 411 -83 445
rect 33 411 45 445
rect 161 411 173 445
rect 289 411 301 445
rect -351 405 -289 411
rect -223 405 -161 411
rect -95 405 -33 411
rect 33 405 95 411
rect 161 405 223 411
rect 289 405 351 411
<< nwell >>
rect -449 -498 449 464
<< pmoslvt >>
rect -355 -436 -285 364
rect -227 -436 -157 364
rect -99 -436 -29 364
rect 29 -436 99 364
rect 157 -436 227 364
rect 285 -436 355 364
<< pdiff >>
rect -413 352 -355 364
rect -413 -424 -401 352
rect -367 -424 -355 352
rect -413 -436 -355 -424
rect -285 352 -227 364
rect -285 -424 -273 352
rect -239 -424 -227 352
rect -285 -436 -227 -424
rect -157 352 -99 364
rect -157 -424 -145 352
rect -111 -424 -99 352
rect -157 -436 -99 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 99 352 157 364
rect 99 -424 111 352
rect 145 -424 157 352
rect 99 -436 157 -424
rect 227 352 285 364
rect 227 -424 239 352
rect 273 -424 285 352
rect 227 -436 285 -424
rect 355 352 413 364
rect 355 -424 367 352
rect 401 -424 413 352
rect 355 -436 413 -424
<< pdiffc >>
rect -401 -424 -367 352
rect -273 -424 -239 352
rect -145 -424 -111 352
rect -17 -424 17 352
rect 111 -424 145 352
rect 239 -424 273 352
rect 367 -424 401 352
<< poly >>
rect -355 445 -285 461
rect -355 411 -339 445
rect -301 411 -285 445
rect -355 364 -285 411
rect -227 445 -157 461
rect -227 411 -211 445
rect -173 411 -157 445
rect -227 364 -157 411
rect -99 445 -29 461
rect -99 411 -83 445
rect -45 411 -29 445
rect -99 364 -29 411
rect 29 445 99 461
rect 29 411 45 445
rect 83 411 99 445
rect 29 364 99 411
rect 157 445 227 461
rect 157 411 173 445
rect 211 411 227 445
rect 157 364 227 411
rect 285 445 355 461
rect 285 411 301 445
rect 339 411 355 445
rect 285 364 355 411
rect -355 -462 -285 -436
rect -227 -462 -157 -436
rect -99 -462 -29 -436
rect 29 -462 99 -436
rect 157 -462 227 -436
rect 285 -462 355 -436
<< polycont >>
rect -339 411 -301 445
rect -211 411 -173 445
rect -83 411 -45 445
rect 45 411 83 445
rect 173 411 211 445
rect 301 411 339 445
<< locali >>
rect -355 411 -339 445
rect -301 411 -285 445
rect -227 411 -211 445
rect -173 411 -157 445
rect -99 411 -83 445
rect -45 411 -29 445
rect 29 411 45 445
rect 83 411 99 445
rect 157 411 173 445
rect 211 411 227 445
rect 285 411 301 445
rect 339 411 355 445
rect -401 352 -367 368
rect -401 -440 -367 -424
rect -273 352 -239 368
rect -273 -440 -239 -424
rect -145 352 -111 368
rect -145 -440 -111 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 111 352 145 368
rect 111 -440 145 -424
rect 239 352 273 368
rect 239 -440 273 -424
rect 367 352 401 368
rect 367 -440 401 -424
<< viali >>
rect -339 411 -301 445
rect -211 411 -173 445
rect -83 411 -45 445
rect 45 411 83 445
rect 173 411 211 445
rect 301 411 339 445
rect -401 -424 -367 352
rect -273 -424 -239 352
rect -145 -424 -111 352
rect -17 -424 17 352
rect 111 -424 145 352
rect 239 -424 273 352
rect 367 -424 401 352
<< metal1 >>
rect -351 445 -289 451
rect -351 411 -339 445
rect -301 411 -289 445
rect -351 405 -289 411
rect -223 445 -161 451
rect -223 411 -211 445
rect -173 411 -161 445
rect -223 405 -161 411
rect -95 445 -33 451
rect -95 411 -83 445
rect -45 411 -33 445
rect -95 405 -33 411
rect 33 445 95 451
rect 33 411 45 445
rect 83 411 95 445
rect 33 405 95 411
rect 161 445 223 451
rect 161 411 173 445
rect 211 411 223 445
rect 161 405 223 411
rect 289 445 351 451
rect 289 411 301 445
rect 339 411 351 445
rect 289 405 351 411
rect -407 352 -361 364
rect -407 -424 -401 352
rect -367 -424 -361 352
rect -407 -436 -361 -424
rect -279 352 -233 364
rect -279 -424 -273 352
rect -239 -424 -233 352
rect -279 -436 -233 -424
rect -151 352 -105 364
rect -151 -424 -145 352
rect -111 -424 -105 352
rect -151 -436 -105 -424
rect -23 352 23 364
rect -23 -424 -17 352
rect 17 -424 23 352
rect -23 -436 23 -424
rect 105 352 151 364
rect 105 -424 111 352
rect 145 -424 151 352
rect 105 -436 151 -424
rect 233 352 279 364
rect 233 -424 239 352
rect 273 -424 279 352
rect 233 -436 279 -424
rect 361 352 407 364
rect 361 -424 367 352
rect 401 -424 407 352
rect 361 -436 407 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 0.35 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
