magic
tech sky130A
magscale 1 2
timestamp 1711802774
<< error_p >>
rect -989 872 -931 878
rect -797 872 -739 878
rect -605 872 -547 878
rect -413 872 -355 878
rect -221 872 -163 878
rect -29 872 29 878
rect 163 872 221 878
rect 355 872 413 878
rect 547 872 605 878
rect 739 872 797 878
rect 931 872 989 878
rect 1123 872 1181 878
rect -989 838 -977 872
rect -797 838 -785 872
rect -605 838 -593 872
rect -413 838 -401 872
rect -221 838 -209 872
rect -29 838 -17 872
rect 163 838 175 872
rect 355 838 367 872
rect 547 838 559 872
rect 739 838 751 872
rect 931 838 943 872
rect 1123 838 1135 872
rect -989 832 -931 838
rect -797 832 -739 838
rect -605 832 -547 838
rect -413 832 -355 838
rect -221 832 -163 838
rect -29 832 29 838
rect 163 832 221 838
rect 355 832 413 838
rect 547 832 605 838
rect 739 832 797 838
rect 931 832 989 838
rect 1123 832 1181 838
<< pwell >>
rect 1022 819 1209 905
rect 1135 811 1178 819
<< nmoslvt >>
rect -1071 -800 -1041 800
rect -975 -800 -945 800
rect -879 -800 -849 800
rect -783 -800 -753 800
rect -687 -800 -657 800
rect -591 -800 -561 800
rect -495 -800 -465 800
rect -399 -800 -369 800
rect -303 -800 -273 800
rect -207 -800 -177 800
rect -111 -800 -81 800
rect -15 -800 15 800
rect 81 -800 111 800
rect 177 -800 207 800
rect 273 -800 303 800
rect 369 -800 399 800
rect 465 -800 495 800
rect 561 -800 591 800
rect 657 -800 687 800
rect 753 -800 783 800
rect 849 -800 879 800
rect 945 -800 975 800
rect 1041 -800 1071 800
<< ndiff >>
rect -1133 788 -1071 800
rect -1133 -788 -1121 788
rect -1087 -788 -1071 788
rect -1133 -800 -1071 -788
rect -1041 788 -975 800
rect -1041 -788 -1025 788
rect -991 -788 -975 788
rect -1041 -800 -975 -788
rect -945 788 -879 800
rect -945 -788 -929 788
rect -895 -788 -879 788
rect -945 -800 -879 -788
rect -849 788 -783 800
rect -849 -788 -833 788
rect -799 -788 -783 788
rect -849 -800 -783 -788
rect -753 788 -687 800
rect -753 -788 -737 788
rect -703 -788 -687 788
rect -753 -800 -687 -788
rect -657 788 -591 800
rect -657 -788 -641 788
rect -607 -788 -591 788
rect -657 -800 -591 -788
rect -561 788 -495 800
rect -561 -788 -545 788
rect -511 -788 -495 788
rect -561 -800 -495 -788
rect -465 788 -399 800
rect -465 -788 -449 788
rect -415 -788 -399 788
rect -465 -800 -399 -788
rect -369 788 -303 800
rect -369 -788 -353 788
rect -319 -788 -303 788
rect -369 -800 -303 -788
rect -273 788 -207 800
rect -273 -788 -257 788
rect -223 -788 -207 788
rect -273 -800 -207 -788
rect -177 788 -111 800
rect -177 -788 -161 788
rect -127 -788 -111 788
rect -177 -800 -111 -788
rect -81 788 -15 800
rect -81 -788 -65 788
rect -31 -788 -15 788
rect -81 -800 -15 -788
rect 15 788 81 800
rect 15 -788 31 788
rect 65 -788 81 788
rect 15 -800 81 -788
rect 111 788 177 800
rect 111 -788 127 788
rect 161 -788 177 788
rect 111 -800 177 -788
rect 207 788 273 800
rect 207 -788 223 788
rect 257 -788 273 788
rect 207 -800 273 -788
rect 303 788 369 800
rect 303 -788 319 788
rect 353 -788 369 788
rect 303 -800 369 -788
rect 399 788 465 800
rect 399 -788 415 788
rect 449 -788 465 788
rect 399 -800 465 -788
rect 495 788 561 800
rect 495 -788 511 788
rect 545 -788 561 788
rect 495 -800 561 -788
rect 591 788 657 800
rect 591 -788 607 788
rect 641 -788 657 788
rect 591 -800 657 -788
rect 687 788 753 800
rect 687 -788 703 788
rect 737 -788 753 788
rect 687 -800 753 -788
rect 783 788 849 800
rect 783 -788 799 788
rect 833 -788 849 788
rect 783 -800 849 -788
rect 879 788 945 800
rect 879 -788 895 788
rect 929 -788 945 788
rect 879 -800 945 -788
rect 975 788 1041 800
rect 975 -788 991 788
rect 1025 -788 1041 788
rect 975 -800 1041 -788
rect 1071 788 1133 800
rect 1071 -788 1087 788
rect 1121 -788 1133 788
rect 1071 -800 1133 -788
<< ndiffc >>
rect -1121 -788 -1087 788
rect -1025 -788 -991 788
rect -929 -788 -895 788
rect -833 -788 -799 788
rect -737 -788 -703 788
rect -641 -788 -607 788
rect -545 -788 -511 788
rect -449 -788 -415 788
rect -353 -788 -319 788
rect -257 -788 -223 788
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
rect 223 -788 257 788
rect 319 -788 353 788
rect 415 -788 449 788
rect 511 -788 545 788
rect 607 -788 641 788
rect 703 -788 737 788
rect 799 -788 833 788
rect 895 -788 929 788
rect 991 -788 1025 788
rect 1087 -788 1121 788
<< poly >>
rect -993 872 -927 888
rect -993 869 -977 872
rect -1071 838 -977 869
rect -943 869 -927 872
rect -801 872 -735 888
rect -801 869 -785 872
rect -943 838 -785 869
rect -751 869 -735 872
rect -609 872 -543 888
rect -609 869 -593 872
rect -751 838 -593 869
rect -559 869 -543 872
rect -417 872 -351 888
rect -417 869 -401 872
rect -559 838 -401 869
rect -367 838 -351 872
rect -225 872 -159 888
rect -225 869 -209 872
rect -1071 826 -351 838
rect -1071 800 -1041 826
rect -993 822 -927 826
rect -975 800 -945 822
rect -879 800 -849 826
rect -801 822 -735 826
rect -783 800 -753 822
rect -687 800 -657 826
rect -609 822 -543 826
rect -591 800 -561 822
rect -495 800 -465 826
rect -417 822 -351 826
rect -303 838 -209 869
rect -175 869 -159 872
rect -33 872 33 888
rect -33 869 -17 872
rect -175 838 -17 869
rect 17 869 33 872
rect 159 872 225 888
rect 159 869 175 872
rect 17 838 175 869
rect 209 869 225 872
rect 351 872 417 888
rect 351 869 367 872
rect 209 838 367 869
rect 401 838 417 872
rect 543 872 609 888
rect 543 869 559 872
rect -303 826 417 838
rect -399 800 -369 822
rect -303 800 -273 826
rect -225 822 -159 826
rect -207 800 -177 822
rect -111 800 -81 826
rect -33 822 33 826
rect -15 800 15 822
rect 81 800 111 826
rect 159 822 225 826
rect 177 800 207 822
rect 273 800 303 826
rect 351 822 417 826
rect 465 838 559 869
rect 593 869 609 872
rect 735 872 801 888
rect 735 869 751 872
rect 593 838 751 869
rect 785 838 801 872
rect 927 872 993 888
rect 927 869 943 872
rect 465 826 801 838
rect 369 800 399 822
rect 465 800 495 826
rect 543 822 609 826
rect 561 800 591 822
rect 657 800 687 826
rect 735 822 801 826
rect 849 838 943 869
rect 977 838 993 872
rect 1119 872 1185 888
rect 1119 869 1135 872
rect 849 826 993 838
rect 753 800 783 822
rect 849 800 879 826
rect 927 822 993 826
rect 1041 838 1135 869
rect 1169 838 1185 872
rect 1041 826 1185 838
rect 945 800 975 822
rect 1041 800 1071 826
rect 1119 822 1185 826
rect -1071 -826 -1041 -800
rect -975 -826 -945 -800
rect -879 -826 -849 -800
rect -783 -826 -753 -800
rect -687 -826 -657 -800
rect -591 -826 -561 -800
rect -495 -826 -465 -800
rect -399 -826 -369 -800
rect -303 -826 -273 -800
rect -207 -826 -177 -800
rect -111 -826 -81 -800
rect -15 -826 15 -800
rect 81 -826 111 -800
rect 177 -826 207 -800
rect 273 -826 303 -800
rect 369 -826 399 -800
rect 465 -826 495 -800
rect 561 -826 591 -800
rect 657 -826 687 -800
rect 753 -826 783 -800
rect 849 -826 879 -800
rect 945 -826 975 -800
rect 1041 -826 1071 -800
<< polycont >>
rect -977 838 -943 872
rect -785 838 -751 872
rect -593 838 -559 872
rect -401 838 -367 872
rect -209 838 -175 872
rect -17 838 17 872
rect 175 838 209 872
rect 367 838 401 872
rect 559 838 593 872
rect 751 838 785 872
rect 943 838 977 872
rect 1135 838 1169 872
<< locali >>
rect -993 838 -977 872
rect -943 838 -927 872
rect -801 838 -785 872
rect -751 838 -735 872
rect -609 838 -593 872
rect -559 838 -543 872
rect -417 838 -401 872
rect -367 838 -351 872
rect -225 838 -209 872
rect -175 838 -159 872
rect -33 838 -17 872
rect 17 838 33 872
rect 159 838 175 872
rect 209 838 225 872
rect 351 838 367 872
rect 401 838 417 872
rect 543 838 559 872
rect 593 838 609 872
rect 735 838 751 872
rect 785 838 801 872
rect 927 838 943 872
rect 977 838 993 872
rect 1119 838 1135 872
rect 1169 838 1185 872
rect -1121 788 -1087 804
rect -1121 -804 -1087 -788
rect -1025 788 -991 804
rect -1025 -804 -991 -788
rect -929 788 -895 804
rect -929 -804 -895 -788
rect -833 788 -799 804
rect -833 -804 -799 -788
rect -737 788 -703 804
rect -737 -804 -703 -788
rect -641 788 -607 804
rect -641 -804 -607 -788
rect -545 788 -511 804
rect -545 -804 -511 -788
rect -449 788 -415 804
rect -449 -804 -415 -788
rect -353 788 -319 804
rect -353 -804 -319 -788
rect -257 788 -223 804
rect -257 -804 -223 -788
rect -161 788 -127 804
rect -161 -804 -127 -788
rect -65 788 -31 804
rect -65 -804 -31 -788
rect 31 788 65 804
rect 31 -804 65 -788
rect 127 788 161 804
rect 127 -804 161 -788
rect 223 788 257 804
rect 223 -804 257 -788
rect 319 788 353 804
rect 319 -804 353 -788
rect 415 788 449 804
rect 415 -804 449 -788
rect 511 788 545 804
rect 511 -804 545 -788
rect 607 788 641 804
rect 607 -804 641 -788
rect 703 788 737 804
rect 703 -804 737 -788
rect 799 788 833 804
rect 799 -804 833 -788
rect 895 788 929 804
rect 895 -804 929 -788
rect 991 788 1025 804
rect 991 -804 1025 -788
rect 1087 788 1121 804
rect 1087 -804 1121 -788
<< viali >>
rect -977 838 -943 872
rect -785 838 -751 872
rect -593 838 -559 872
rect -401 838 -367 872
rect -209 838 -175 872
rect -17 838 17 872
rect 175 838 209 872
rect 367 838 401 872
rect 559 838 593 872
rect 751 838 785 872
rect 943 838 977 872
rect 1135 838 1169 872
rect -1121 -788 -1087 788
rect -1025 -788 -991 788
rect -929 -788 -895 788
rect -833 -788 -799 788
rect -737 -788 -703 788
rect -641 -788 -607 788
rect -545 -788 -511 788
rect -449 -788 -415 788
rect -353 -788 -319 788
rect -257 -788 -223 788
rect -161 -788 -127 788
rect -65 -788 -31 788
rect 31 -788 65 788
rect 127 -788 161 788
rect 223 -788 257 788
rect 319 -788 353 788
rect 415 -788 449 788
rect 511 -788 545 788
rect 607 -788 641 788
rect 703 -788 737 788
rect 799 -788 833 788
rect 895 -788 929 788
rect 991 -788 1025 788
rect 1087 -788 1121 788
<< metal1 >>
rect -989 872 -931 878
rect -989 838 -977 872
rect -943 838 -931 872
rect -989 832 -931 838
rect -797 872 -739 878
rect -797 838 -785 872
rect -751 838 -739 872
rect -797 832 -739 838
rect -605 872 -547 878
rect -605 838 -593 872
rect -559 838 -547 872
rect -605 832 -547 838
rect -413 872 -355 878
rect -413 838 -401 872
rect -367 838 -355 872
rect -413 832 -355 838
rect -221 872 -163 878
rect -221 838 -209 872
rect -175 838 -163 872
rect -221 832 -163 838
rect -29 872 29 878
rect -29 838 -17 872
rect 17 838 29 872
rect -29 832 29 838
rect 163 872 221 878
rect 163 838 175 872
rect 209 838 221 872
rect 163 832 221 838
rect 355 872 413 878
rect 355 838 367 872
rect 401 838 413 872
rect 355 832 413 838
rect 547 872 605 878
rect 547 838 559 872
rect 593 838 605 872
rect 547 832 605 838
rect 739 872 797 878
rect 739 838 751 872
rect 785 838 797 872
rect 739 832 797 838
rect 931 872 989 878
rect 931 838 943 872
rect 977 838 989 872
rect 931 832 989 838
rect 1123 872 1181 878
rect 1123 838 1135 872
rect 1169 838 1181 872
rect 1123 832 1181 838
rect -1127 788 -1081 800
rect -1127 -788 -1121 788
rect -1087 -788 -1081 788
rect -1127 -800 -1081 -788
rect -1031 788 -985 800
rect -1031 -788 -1025 788
rect -991 -788 -985 788
rect -1031 -800 -985 -788
rect -935 788 -889 800
rect -935 -788 -929 788
rect -895 -788 -889 788
rect -935 -800 -889 -788
rect -839 788 -793 800
rect -839 -788 -833 788
rect -799 -788 -793 788
rect -839 -800 -793 -788
rect -743 788 -697 800
rect -743 -788 -737 788
rect -703 -788 -697 788
rect -743 -800 -697 -788
rect -647 788 -601 800
rect -647 -788 -641 788
rect -607 -788 -601 788
rect -647 -800 -601 -788
rect -551 788 -505 800
rect -551 -788 -545 788
rect -511 -788 -505 788
rect -551 -800 -505 -788
rect -455 788 -409 800
rect -455 -788 -449 788
rect -415 -788 -409 788
rect -455 -800 -409 -788
rect -359 788 -313 800
rect -359 -788 -353 788
rect -319 -788 -313 788
rect -359 -800 -313 -788
rect -263 788 -217 800
rect -263 -788 -257 788
rect -223 -788 -217 788
rect -263 -800 -217 -788
rect -167 788 -121 800
rect -167 -788 -161 788
rect -127 -788 -121 788
rect -167 -800 -121 -788
rect -71 788 -25 800
rect -71 -788 -65 788
rect -31 -788 -25 788
rect -71 -800 -25 -788
rect 25 788 71 800
rect 25 -788 31 788
rect 65 -788 71 788
rect 25 -800 71 -788
rect 121 788 167 800
rect 121 -788 127 788
rect 161 -788 167 788
rect 121 -800 167 -788
rect 217 788 263 800
rect 217 -788 223 788
rect 257 -788 263 788
rect 217 -800 263 -788
rect 313 788 359 800
rect 313 -788 319 788
rect 353 -788 359 788
rect 313 -800 359 -788
rect 409 788 455 800
rect 409 -788 415 788
rect 449 -788 455 788
rect 409 -800 455 -788
rect 505 788 551 800
rect 505 -788 511 788
rect 545 -788 551 788
rect 505 -800 551 -788
rect 601 788 647 800
rect 601 -788 607 788
rect 641 -788 647 788
rect 601 -800 647 -788
rect 697 788 743 800
rect 697 -788 703 788
rect 737 -788 743 788
rect 697 -800 743 -788
rect 793 788 839 800
rect 793 -788 799 788
rect 833 -788 839 788
rect 793 -800 839 -788
rect 889 788 935 800
rect 889 -788 895 788
rect 929 -788 935 788
rect 889 -800 935 -788
rect 985 788 1031 800
rect 985 -788 991 788
rect 1025 -788 1031 788
rect 985 -800 1031 -788
rect 1081 788 1127 800
rect 1081 -788 1087 788
rect 1121 -788 1127 788
rect 1081 -800 1127 -788
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8 l 0.150 m 1 nf 23 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
