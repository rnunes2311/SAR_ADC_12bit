magic
tech sky130A
magscale 1 2
timestamp 1711994201
<< nwell >>
rect -1196 -4573 1196 4573
<< pmoslvt >>
rect -1000 2354 1000 4354
rect -1000 118 1000 2118
rect -1000 -2118 1000 -118
rect -1000 -4354 1000 -2354
<< pdiff >>
rect -1058 4342 -1000 4354
rect -1058 2366 -1046 4342
rect -1012 2366 -1000 4342
rect -1058 2354 -1000 2366
rect 1000 4342 1058 4354
rect 1000 2366 1012 4342
rect 1046 2366 1058 4342
rect 1000 2354 1058 2366
rect -1058 2106 -1000 2118
rect -1058 130 -1046 2106
rect -1012 130 -1000 2106
rect -1058 118 -1000 130
rect 1000 2106 1058 2118
rect 1000 130 1012 2106
rect 1046 130 1058 2106
rect 1000 118 1058 130
rect -1058 -130 -1000 -118
rect -1058 -2106 -1046 -130
rect -1012 -2106 -1000 -130
rect -1058 -2118 -1000 -2106
rect 1000 -130 1058 -118
rect 1000 -2106 1012 -130
rect 1046 -2106 1058 -130
rect 1000 -2118 1058 -2106
rect -1058 -2366 -1000 -2354
rect -1058 -4342 -1046 -2366
rect -1012 -4342 -1000 -2366
rect -1058 -4354 -1000 -4342
rect 1000 -2366 1058 -2354
rect 1000 -4342 1012 -2366
rect 1046 -4342 1058 -2366
rect 1000 -4354 1058 -4342
<< pdiffc >>
rect -1046 2366 -1012 4342
rect 1012 2366 1046 4342
rect -1046 130 -1012 2106
rect 1012 130 1046 2106
rect -1046 -2106 -1012 -130
rect 1012 -2106 1046 -130
rect -1046 -4342 -1012 -2366
rect 1012 -4342 1046 -2366
<< nsubdiff >>
rect -1160 4503 -1064 4537
rect 1064 4503 1160 4537
rect -1160 4441 -1126 4503
rect 1126 4441 1160 4503
rect -1160 -4503 -1126 -4441
rect 1126 -4503 1160 -4441
rect -1160 -4537 -1064 -4503
rect 1064 -4537 1160 -4503
<< nsubdiffcont >>
rect -1064 4503 1064 4537
rect -1160 -4441 -1126 4441
rect 1126 -4441 1160 4441
rect -1064 -4537 1064 -4503
<< poly >>
rect -1000 4435 1000 4451
rect -1000 4401 -984 4435
rect 984 4401 1000 4435
rect -1000 4354 1000 4401
rect -1000 2307 1000 2354
rect -1000 2273 -984 2307
rect 984 2273 1000 2307
rect -1000 2257 1000 2273
rect -1000 2199 1000 2215
rect -1000 2165 -984 2199
rect 984 2165 1000 2199
rect -1000 2118 1000 2165
rect -1000 71 1000 118
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 21 1000 37
rect -1000 -37 1000 -21
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1000 -118 1000 -71
rect -1000 -2165 1000 -2118
rect -1000 -2199 -984 -2165
rect 984 -2199 1000 -2165
rect -1000 -2215 1000 -2199
rect -1000 -2273 1000 -2257
rect -1000 -2307 -984 -2273
rect 984 -2307 1000 -2273
rect -1000 -2354 1000 -2307
rect -1000 -4401 1000 -4354
rect -1000 -4435 -984 -4401
rect 984 -4435 1000 -4401
rect -1000 -4451 1000 -4435
<< polycont >>
rect -984 4401 984 4435
rect -984 2273 984 2307
rect -984 2165 984 2199
rect -984 37 984 71
rect -984 -71 984 -37
rect -984 -2199 984 -2165
rect -984 -2307 984 -2273
rect -984 -4435 984 -4401
<< locali >>
rect -1160 4503 -1064 4537
rect 1064 4503 1160 4537
rect -1160 4441 -1126 4503
rect 1126 4441 1160 4503
rect -1000 4401 -984 4435
rect 984 4401 1000 4435
rect -1046 4342 -1012 4358
rect -1046 2350 -1012 2366
rect 1012 4342 1046 4358
rect 1012 2350 1046 2366
rect -1000 2273 -984 2307
rect 984 2273 1000 2307
rect -1000 2165 -984 2199
rect 984 2165 1000 2199
rect -1046 2106 -1012 2122
rect -1046 114 -1012 130
rect 1012 2106 1046 2122
rect 1012 114 1046 130
rect -1000 37 -984 71
rect 984 37 1000 71
rect -1000 -71 -984 -37
rect 984 -71 1000 -37
rect -1046 -130 -1012 -114
rect -1046 -2122 -1012 -2106
rect 1012 -130 1046 -114
rect 1012 -2122 1046 -2106
rect -1000 -2199 -984 -2165
rect 984 -2199 1000 -2165
rect -1000 -2307 -984 -2273
rect 984 -2307 1000 -2273
rect -1046 -2366 -1012 -2350
rect -1046 -4358 -1012 -4342
rect 1012 -2366 1046 -2350
rect 1012 -4358 1046 -4342
rect -1000 -4435 -984 -4401
rect 984 -4435 1000 -4401
rect -1160 -4503 -1126 -4441
rect 1126 -4503 1160 -4441
rect -1160 -4537 -1064 -4503
rect 1064 -4537 1160 -4503
<< viali >>
rect -984 4401 984 4435
rect -1046 2366 -1012 4342
rect 1012 2366 1046 4342
rect -984 2273 984 2307
rect -984 2165 984 2199
rect -1046 130 -1012 2106
rect 1012 130 1046 2106
rect -984 37 984 71
rect -984 -71 984 -37
rect -1046 -2106 -1012 -130
rect 1012 -2106 1046 -130
rect -984 -2199 984 -2165
rect -984 -2307 984 -2273
rect -1046 -4342 -1012 -2366
rect 1012 -4342 1046 -2366
rect -984 -4435 984 -4401
<< metal1 >>
rect -996 4435 996 4441
rect -996 4401 -984 4435
rect 984 4401 996 4435
rect -996 4395 996 4401
rect -1052 4342 -1006 4354
rect -1052 2366 -1046 4342
rect -1012 2366 -1006 4342
rect -1052 2354 -1006 2366
rect 1006 4342 1052 4354
rect 1006 2366 1012 4342
rect 1046 2366 1052 4342
rect 1006 2354 1052 2366
rect -996 2307 996 2313
rect -996 2273 -984 2307
rect 984 2273 996 2307
rect -996 2267 996 2273
rect -996 2199 996 2205
rect -996 2165 -984 2199
rect 984 2165 996 2199
rect -996 2159 996 2165
rect -1052 2106 -1006 2118
rect -1052 130 -1046 2106
rect -1012 130 -1006 2106
rect -1052 118 -1006 130
rect 1006 2106 1052 2118
rect 1006 130 1012 2106
rect 1046 130 1052 2106
rect 1006 118 1052 130
rect -996 71 996 77
rect -996 37 -984 71
rect 984 37 996 71
rect -996 31 996 37
rect -996 -37 996 -31
rect -996 -71 -984 -37
rect 984 -71 996 -37
rect -996 -77 996 -71
rect -1052 -130 -1006 -118
rect -1052 -2106 -1046 -130
rect -1012 -2106 -1006 -130
rect -1052 -2118 -1006 -2106
rect 1006 -130 1052 -118
rect 1006 -2106 1012 -130
rect 1046 -2106 1052 -130
rect 1006 -2118 1052 -2106
rect -996 -2165 996 -2159
rect -996 -2199 -984 -2165
rect 984 -2199 996 -2165
rect -996 -2205 996 -2199
rect -996 -2273 996 -2267
rect -996 -2307 -984 -2273
rect 984 -2307 996 -2273
rect -996 -2313 996 -2307
rect -1052 -2366 -1006 -2354
rect -1052 -4342 -1046 -2366
rect -1012 -4342 -1006 -2366
rect -1052 -4354 -1006 -4342
rect 1006 -2366 1052 -2354
rect 1006 -4342 1012 -2366
rect 1046 -4342 1052 -2366
rect 1006 -4354 1052 -4342
rect -996 -4401 996 -4395
rect -996 -4435 -984 -4401
rect 984 -4435 996 -4401
rect -996 -4441 996 -4435
<< properties >>
string FIXED_BBOX -1143 -4520 1143 4520
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 10.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
