* NGSPICE file created from SAR_ADC_12bit_flat.ext - technology: sky130A

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START EN_OFFSET_CAL CLK VREF_GND
+ SINGLE_ENDED
X0 a_13076_44458# a_13259_45724.t13 a_13296_44484# VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_8912_37509.t15 VDAC_P.t23 a_5088_37509.t10 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2 VSS.t42 a_12427_45724# a_10490_45724# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VDD.t3173 a_2324_44458.t62 a_949_44458# VDD.t3172 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VDD.t227 VSS.t3732 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5 a_5088_37509.t13 VDAC_P.t21 a_8912_37509.t2 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6 VDD.t3430 CAL_N.t3 VDD.t3430 VDD.t1753 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X7 VDD.t46 a_2903_42308# a_3080_42308.t1 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8 VDD.t3189 a_12861_44030.t25 a_17829_46910# VDD.t3188 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VSS.t7 a_1209_43370# a_n1557_42282# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_16237_45028# a_16147_45260# a_16019_45002# VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_2075_43172# a_526_44458.t25 VSS.t3402 VSS.t3401 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VDD.t3436 a_n755_45592.t8 a_1176_45822# VDD.t3435 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X13 a_6756_44260# a_5937_45572.t18 a_6453_43914# VSS.t3500 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X14 a_15868_43402# a_15681_43442# a_15781_43660# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X15 a_n1533_42852# a_n1613_43370.t8 VDD.t3364 VDD.t3363 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X16 a_8103_44636# a_8375_44464# a_8333_44734# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 VSS.t3366 a_16327_47482.t23 a_16377_45572# VSS.t3365 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 a_2437_43646.t0 a_n443_46116.t19 a_2437_43396# VSS.t3051 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_5088_37509.t17 VSS.t3738 VDAC_Ni.t1 VDD.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X20 a_n2810_45028.t3 a_n2840_45002# VSS.t85 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X21 a_2113_38308# VDAC_Ni.t9 a_2112_39137# VSS.t3347 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X22 VDD.t3559 a_3626_43646.t6 a_19647_42308# VDD.t3558 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 VSS.t93 a_10334_44484# a_10440_44484# VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_1576_42282# a_1755_42282# VSS.t97 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X25 a_10933_46660# a_10554_47026# a_10861_46660# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 a_14021_43940.t0 a_13483_43940# VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X27 a_16867_43762# a_16327_47482.t43 VDD.t3358 VDD.t3357 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VREF.t1 a_21076_30879.t4 C8_N_btm.t1 VDD.t3554 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X29 VSS.t111 a_n2946_37690# a_n3565_37414.t7 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_n913_45002.t11 a_1307_43914.t8 a_2075_43172# VSS.t3483 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_n2840_43370# a_n2661_43370.t3 VSS.t2821 VSS.t1732 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X32 a_3457_43396# a_584_46384.t8 VSS.t2773 VSS.t2772 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X33 a_14180_46482# a_14035_46660# VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X34 VSS.t119 a_18989_43940# a_19006_44850# VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X35 VSS.t121 a_9672_43914# a_2107_46812.t1 VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X36 a_n1059_45260.t7 a_17499_43370# VSS.t129 VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_n1696_34930.t7 a_n1794_35082.t4 VSS.t2837 VSS.t2836 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VSS.t133 a_10695_43548# a_10057_43914# VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X39 a_n2104_42282# a_n1925_42282.t3 VSS.t2835 VSS.t2834 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X40 a_20749_43396# a_12549_44172.t30 a_743_42282.t1 VSS.t2722 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X41 VDD.t318 a_3877_44458# a_2382_45260# VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_n1699_44726# a_n1917_44484# VSS.t157 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X43 VSS.t162 a_n4334_39616# a_n4064_39616.t7 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X44 a_9241_45822# a_5066_45546# VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X45 VDD.t346 a_12883_44458# a_n2293_43922.t0 VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X46 a_11909_44484# a_3232_43370.t17 a_11827_44484# VSS.t2828 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X47 a_835_46155# a_584_46384.t21 a_376_46348# VDD.t3008 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X48 VSS.t2714 a_1666_39043.t3 a_1169_39043# VSS.t1799 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X49 a_5210_46155# a_5164_46348# VDD.t360 VDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X50 VDD.t364 a_n3690_39392# a_n3420_39072.t2 VDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X51 VDD.t374 a_167_45260# a_1609_45822# VDD.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X52 VSS.t3413 a_526_44458.t33 a_3363_44484# VSS.t3412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 a_19268_43646# a_19319_43548# a_19095_43396# VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X54 VSS.t219 a_22959_44484# a_19237_31679.t3 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 a_n2216_39072# a_n2312_39304.t4 a_n2302_39072# VDD.t2877 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X56 a_19987_42826# a_10193_42453.t13 VDD.t3022 VDD.t3021 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X57 a_6151_47436.t0 a_14311_47204# VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X58 a_8145_46902# a_7927_46660# VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X59 VCM.t2 a_4190_30871.t15 C10_N_btm.t0 VSS.t2813 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X60 a_14275_46494# a_13925_46122# a_14180_46482# VDD.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X61 a_20512_43084# a_11967_42832.t48 VSS.t2943 VSS.t2942 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X62 a_14539_43914# a_17701_42308# VSS.t814 VSS.t813 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 a_6298_44484# a_2324_44458.t46 VSS.t3007 VSS.t3006 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X64 a_644_44056# a_626_44172# VSS.t855 VSS.t854 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X65 a_10949_43914# a_12429_44172# VDD.t1041 VDD.t1040 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X66 VSS.t861 a_n2302_39866# a_n4209_39590.t7 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X67 VSS.t865 a_21811_47423# a_20916_46384# VSS.t864 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X68 VDD.t1056 a_3699_46634# a_3686_47026# VDD.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 VSS.t872 a_15682_46116# a_11599_46634.t28 VSS.t871 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X70 a_8035_47026# a_7411_46660# a_7927_46660# VDD.t1094 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X71 a_5691_45260# a_5111_44636# a_5837_45348# VSS.t749 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X72 VDD.t3542 a_1307_43914.t33 a_1241_43940# VDD.t3541 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X73 a_5088_37509.t14 VDAC_P.t17 a_8912_37509.t3 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X74 a_18249_42858# a_18083_42858# VSS.t923 VSS.t922 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 VDD.t1126 a_104_43370# a_n971_45724.t0 VDD.t1125 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X76 VDD.t418 a_n2833_47464# CLK_DATA.t0 VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X77 a_3363_44484# a_1823_45246# a_3232_43370.t4 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X78 a_n1331_43914# a_n1549_44318# VDD.t446 VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X79 VCM.t34 a_4958_30871.t7 C9_P_btm.t7 VSS.t2695 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X80 VSS.t3529 a_n3565_39590.t8 a_n3607_39616# VSS.t3521 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X81 VSS.t265 a_12281_43396# a_12563_42308# VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X82 VSS.t271 a_18780_47178# a_13661_43548.t3 VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X83 a_n4318_39768.t3 a_n2840_43914# VSS.t277 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X84 DATA[5].t3 a_11459_47204# VDD.t466 VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X85 a_7230_45938# a_6472_45840# a_6667_45809# VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X86 VDD.t3100 a_8049_45260.t3 a_22959_45572# VDD.t3099 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X87 a_2324_44458.t22 a_8953_45002# VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X88 a_8746_45002# a_7499_43078# VSS.t326 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 a_15004_44636# a_11691_44458.t4 a_15146_44484# VSS.t2885 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 a_16223_45938# a_15599_45572# a_16115_45572# VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X91 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS.t354 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X92 a_n809_44244# a_n1613_43370.t45 VDD.t3400 VDD.t3399 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X93 a_n4064_39616.t6 a_n4334_39616# VSS.t164 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X94 a_17124_42282# a_17303_42282# VSS.t367 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X95 VDD.t1076 a_15682_46116# a_11599_46634.t2 VDD.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X96 VSS.t373 a_3065_45002# a_2680_45002# VSS.t372 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X97 a_5193_42852# a_5111_44636# VDD.t1106 VDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X98 VDD.t568 a_6969_46634# a_6999_46987# VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X99 VDD.t570 a_10623_46897# a_10554_47026# VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X100 a_16137_43396# a_15781_43660# VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X101 VDD.t576 a_n2472_46634# a_n2442_46660.t1 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X102 VDD.t1892 a_4185_45028.t3 a_22959_45036# VDD.t1891 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X103 a_15225_45822# a_15037_45618# a_15143_45578# VDD.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X104 VSS.t2672 a_3537_45260.t21 a_4640_45348# VSS.t2671 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 a_n2012_43396# a_n2129_43609# VDD.t583 VDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X106 VDD.t585 a_n13_43084# a_n1853_43023# VDD.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X107 a_5068_46348# a_n1151_42308.t4 a_5210_46155# VDD.t1880 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X108 a_873_42968# a_685_42968# a_791_42968# VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X109 a_17730_32519.t1 a_22591_44484# VDD.t594 VDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X110 a_11967_42832.t25 a_15682_43940# VSS.t440 VSS.t439 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 VDD.t630 a_22485_44484# a_20974_43370# VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X112 a_n1021_46688# a_n1151_42308.t17 VDD.t1887 VDD.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X113 VSS.t2961 a_11599_46634.t46 a_11735_46660# VSS.t2960 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X114 a_13163_45724# a_13259_45724.t21 VDD.t248 VDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X115 C9_P_btm.t5 a_4958_30871.t8 VCM.t35 VSS.t2696 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X116 a_11599_46634.t29 a_15682_46116# VSS.t896 VSS.t895 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X117 a_n2012_44484# a_n2129_44697# VSS.t462 VSS.t461 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X118 VIN_N.t3 EN_VIN_BSTR_N.t22 a_10890_34112.t1 VSS.t2927 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X119 a_13940_44484# a_13556_45296# VSS.t465 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X120 VSS.t475 a_1414_42308# a_1525_44260# VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X121 a_8487_44056# a_4223_44672.t4 a_8415_44056# VDD.t2895 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X122 VDAC_P.t3 a_3422_30871.t15 VCM.t53 VSS.t3516 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X123 a_16434_46660# a_16388_46812# VSS.t477 VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X124 a_22613_38993# a_22527_39145# VDD.t661 VDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X125 a_3315_47570# a_n1151_42308.t13 a_2952_47436# VSS.t1660 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X126 a_2680_45002# a_1823_45246# a_2903_45348# VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X127 a_1307_43914.t1 a_2779_44458# VDD.t667 VDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X128 a_22731_47423# SMPL_ON_N.t8 VDD.t3573 VDD.t3572 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X129 VDD.t3538 a_1307_43914.t31 a_3681_42891# VDD.t3537 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X130 a_n863_45724# a_1667_45002# VSS.t499 VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 VDD.t464 a_11459_47204# DATA[5].t2 VDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X132 VSS.t307 a_8953_45002# a_2324_44458.t21 VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X133 a_4646_46812.t1 a_6298_44484# VDD.t1011 VDD.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X134 VSS.t3157 VDD.t3826 VSS.t3156 VSS.t3155 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X135 VREF_GND.t10 a_18114_32519.t5 C10_N_btm.t25 VSS.t2648 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X136 a_n4209_38216.t3 a_n2302_37984# VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X137 a_10467_46802# a_11599_46634.t45 VDD.t3163 VDD.t3162 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X138 VDD.t3083 a_13747_46662.t3 a_19862_44208# VDD.t3082 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X139 a_n2946_39866# a_n2956_39768.t4 VSS.t2871 VSS.t1734 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X140 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X141 VSS.t546 a_15279_43071# a_14579_43548# VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X142 DATA[3].t3 a_7227_47204# VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X143 VSS.t2877 a_8049_45260.t4 a_22959_45572# VSS.t1665 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X144 a_7584_44260# a_7542_44172# a_7281_43914# VSS.t557 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X145 a_n97_42460.t3 a_19700_43370# VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X146 VDD.t262 a_19647_42308# a_13258_32519.t1 VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X147 a_3754_39466# a_7754_39300# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X148 VSS.t485 a_2952_47436# a_2747_46873# VSS.t484 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X149 VDD.t751 a_16751_45260# a_6171_45002.t0 VDD.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X150 a_18326_43940# a_18079_43940# VDD.t753 VDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X151 a_9248_44260# a_8270_45546# VSS.t574 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X152 a_3503_45724# a_3775_45552# a_3733_45822# VDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X153 a_n2017_45002.t1 a_19987_42826# VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X154 a_288_46660# a_171_46873# VSS.t584 VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X155 a_10037_46155# a_9804_47204# a_9823_46155# VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X156 a_20075_46420# a_16327_47482.t29 VDD.t3425 VDD.t3424 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X157 VDD.t774 a_196_42282# a_n3674_37592.t1 VDD.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X158 VSS.t597 a_14513_46634# a_14447_46660# VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 a_n4064_39072.t3 a_n4334_39392# VDD.t782 VDD.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X160 a_1149_42558# a_961_42354# a_1067_42314# VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 a_13569_47204# a_13381_47204# a_13487_47204# VDD.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X162 VDD.t798 a_14840_46494# a_15015_46420# VDD.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 C6_P_btm.t2 a_n3565_39304.t8 VREF.t65 VDD.t3604 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X164 VDD.t223 VSS.t3764 VDD.t222 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X165 a_2324_44458.t20 a_8953_45002# VSS.t297 VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X166 a_14537_43396# a_14358_43442# VSS.t620 VSS.t619 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X167 VDD.t809 a_14955_47212# a_10227_46804.t0 VDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X168 VDD.t3589 a_7754_40130.t9 a_11206_38545.t3 VDD.t3588 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X169 a_n3565_39590.t1 a_n2946_39866# VDD.t722 VDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_n901_43156# a_n1613_43370.t23 VDD.t3374 VDD.t3373 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X171 a_17668_45572# a_3090_45724.t6 VSS.t1583 VSS.t1582 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X172 a_n2438_43548.t29 a_949_44458# VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X173 a_15493_43396.t1 a_14955_43396# VSS.t641 VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X174 a_7309_43172# a_5891_43370.t8 VSS.t1649 VSS.t1648 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X175 VDD.t825 a_1138_42852# a_1337_46116# VDD.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X176 a_1427_43646# a_1568_43370# VDD.t827 VDD.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X177 a_18184_42460.t0 a_15743_43084# VSS.t650 VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X178 VDD.t837 a_13351_46090# a_10903_43370.t1 VDD.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X179 a_8379_46155# a_8128_46384# a_7920_46348# VDD.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X180 VSS.t3081 a_3483_46348.t13 a_17325_44484# VSS.t3080 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X181 VDD.t3279 a_9290_44172.t28 a_10949_43914# VDD.t3278 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X182 VSS.t3543 a_11823_42460.t21 a_14358_43442# VSS.t3542 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X183 a_18310_42308# a_10193_42453.t21 a_18220_42308# VSS.t2797 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X184 VDD.t846 a_n2288_47178# a_n2312_40392.t1 VDD.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X185 a_17719_45144# a_16375_45002# VSS.t666 VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X186 VDD.t1816 a_5891_43370.t23 a_5147_45002# VDD.t1815 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X187 a_7287_43370# a_n1613_43370.t43 VDD.t3398 VDD.t3397 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X188 a_11173_44260# a_2063_45854.t11 VSS.t1642 VSS.t1641 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X189 a_11897_42308# a_11823_42460.t27 a_11551_42558# VSS.t3548 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X190 VDD.t3199 a_12861_44030.t33 a_13759_47204# VDD.t3198 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X191 a_19466_46812# a_19778_44110# VSS.t688 VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X192 a_9049_44484# a_8701_44490# VSS.t695 VSS.t694 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X193 a_n3565_38502.t7 a_n2946_38778# VSS.t700 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X194 VDD.t887 a_16588_47582# a_16763_47508# VDD.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X195 a_9396_43370# a_4883_46098.t3 VSS.t1631 VSS.t1630 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X196 C0_P_btm.t1 a_n784_42308.t4 VCM.t60 VSS.t3530 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X197 a_n1736_42282# a_n1557_42282# VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X198 VDD.t903 a_14113_42308# a_16522_42674# VDD.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X199 a_10651_43940# a_3090_45724.t19 a_10555_43940# VDD.t1823 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X200 VDD.t907 a_8667_46634# a_n237_47217.t0 VDD.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 a_6123_31319.t3 a_7227_42308# VSS.t729 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X202 a_7499_43078# a_10083_42826# VSS.t732 VSS.t731 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X203 VSS.t3388 a_n755_45592.t25 a_1145_45348# VSS.t3387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X204 C7_P_btm.t1 a_5534_30871.t4 VCM.t40 VSS.t3025 sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X205 VREF.t27 a_22612_30879.t19 C10_N_btm.t23 VDD.t1954 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X206 VSS.t3024 a_n4064_37984.t8 a_n2302_37984# VSS.t1787 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VSS.t17 a_949_44458# a_n2438_43548.t24 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X208 a_3581_42558# a_3539_42460# a_3497_42558# VDD.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X209 a_n3674_38680.t1 a_n2840_42282# VDD.t926 VDD.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X210 VSS.t752 a_5907_45546# a_5937_45572.t2 VSS.t751 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X211 VDD.t937 a_22589_40055# a_22527_39145# VDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X212 a_18783_43370# a_15743_43084# VSS.t648 VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X213 VSS.t758 a_1799_45572# a_1983_46706# VSS.t757 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X214 VDD.t947 a_22959_46660# a_21076_30879.t1 VDD.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X215 a_13467_32519.t1 a_21487_43396# VDD.t949 VDD.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X216 C10_P_btm.t14 a_n4064_40160.t11 VREF_GND.t37 VSS.t2684 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X217 a_2864_46660# a_2747_46873# VSS.t566 VSS.t565 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X218 VDD.t179 VSS.t3752 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X219 a_8199_44636# a_10355_46116# VSS.t769 VSS.t768 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X220 a_14403_45348# a_13259_45724.t15 a_14309_45348# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X221 a_556_44484# a_742_44458# VSS.t789 VSS.t788 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X222 VSS.t795 a_15433_44458# a_15367_44484# VSS.t794 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X223 a_n1794_35082.t0 a_564_42282# VDD.t982 VDD.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X224 a_n2840_43370# a_n2661_43370.t4 VDD.t3035 VDD.t1762 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X225 w_1575_34786.t7 a_n1696_34930.t10 EN_VIN_BSTR_P.t6 w_1575_34786.t6 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X226 VSS.t2864 a_13747_46662.t7 a_13693_46688# VSS.t2863 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_18245_44484# a_17767_44458# VSS.t803 VSS.t802 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X228 a_19741_43940# a_19862_44208# VDD.t715 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X229 a_16855_43396# a_16409_43396# a_16759_43396# VSS.t804 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X230 a_13113_42826# a_12895_43230# VSS.t1316 VSS.t1315 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X231 VSS.t1319 a_22365_46825# a_20202_43084# VSS.t1318 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X232 a_n1079_45724# a_n755_45592.t19 VSS.t3381 VSS.t3380 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X233 a_19386_47436# a_19321_45002# VDD.t1538 VDD.t1537 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X234 a_4646_46812.t23 a_6298_44484# VSS.t835 VSS.t834 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 VSS.t3415 a_526_44458.t35 a_2075_43172# VSS.t3414 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X236 a_n89_47570# a_n237_47217.t10 a_n452_47436# VSS.t3034 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X237 VDD.t115 VSS.t3759 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X238 a_1176_45822# a_167_45260# VDD.t372 VDD.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X239 a_10341_43396.t1 a_9803_43646# VSS.t1339 VSS.t1338 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X240 VDD.t2920 a_n4209_38502.t8 a_n4334_38528# VDD.t1970 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X241 a_5111_42852# a_4905_42826# a_5193_43172# VSS.t1352 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X242 a_13887_32519.t3 a_22223_43396# VSS.t1355 VSS.t1235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X243 a_5437_45600# a_n881_46662.t4 VSS.t1556 VSS.t1555 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X244 a_18953_45572# a_18909_45814# a_18787_45572# VSS.t1356 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X245 VDD.t2003 a_4791_45118.t4 a_6165_46155# VDD.t2002 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X246 VDD.t1568 a_3429_45260# a_3316_45546# VDD.t1567 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X247 VCM.t57 a_3422_30871.t19 VDAC_P.t6 VSS.t3520 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X248 a_n3607_39616# a_n3674_39768.t4 a_n3690_39616# VSS.t2640 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X249 a_4842_47570# a_4791_45118.t21 VSS.t1767 VSS.t1766 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X250 a_1337_46116# a_n881_46662.t21 VDD.t1798 VDD.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X251 a_11136_45572# a_11322_45546# VSS.t1367 VSS.t1366 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X252 a_n2661_42834.t1 a_10809_44734.t3 a_12189_44484# VSS.t3570 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X253 VSS.t1371 a_10249_46116# a_11186_47026# VSS.t1370 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X254 a_16655_46660# a_n743_46660.t2 a_16292_46812# VSS.t3552 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X255 a_n1991_46122# a_n2157_46122# VSS.t1376 VSS.t1375 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 VREF_GND.t5 a_n3420_39072.t9 C6_P_btm.t1 VSS.t1843 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X257 a_n3565_37414.t6 a_n2946_37690# VSS.t107 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 VDD.t272 a_1576_42282# a_1606_42308.t1 VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X259 a_5159_47243# a_n443_46116.t23 a_4700_47436# VDD.t3257 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X260 VSS.t1581 a_5891_43370.t25 a_8375_44464# VSS.t1580 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 a_2075_43172# a_526_44458.t31 VSS.t3411 VSS.t3410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X262 VDD.t237 a_13076_44458# a_12883_44458# VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X263 VSS.t819 a_14539_43914# a_14485_44260# VSS.t818 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 C0_N_btm.t1 EN_VIN_BSTR_N.t23 VIN_N.t8 VSS.t2925 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X265 a_15297_45822# a_11823_42460.t17 a_15225_45822# VDD.t3629 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X266 VSS.t3698 a_18194_34908.t8 a_10890_34112.t2 VSS.t3697 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X267 VDD.t354 a_1169_39043# comp_n VDD.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X268 a_18479_47436# a_20075_46420# VDD.t770 VDD.t769 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X269 a_1423_45028.t1 a_167_45260# VDD.t380 VDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X270 a_2382_45260# a_3877_44458# VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X271 a_8103_44636# a_8199_44636# VSS.t775 VSS.t774 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X272 a_n1899_43946# a_n2065_43946# VSS.t1389 VSS.t1388 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X273 a_6765_43638# a_6547_43396# VDD.t1605 VDD.t1604 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X274 VSS.t1396 a_22400_42852# a_22848_40945# VSS.t1395 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X275 a_n2293_43922.t1 a_12741_44636.t3 VDD.t1976 VDD.t1975 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X276 a_n3565_38216.t7 a_n2946_37984# VSS.t1404 VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X277 VDD.t368 a_n3690_39392# a_n3420_39072.t3 VDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X278 a_945_42968# a_n1059_45260.t21 a_873_42968# VDD.t2994 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X279 VDD.t1618 a_3785_47178# a_3815_47204# VDD.t1617 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X280 VDD.t1623 a_14084_46812# a_14035_46660# VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X281 a_765_45546.t1 a_12549_44172.t20 a_17829_46910# VDD.t2943 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X282 VDD.t634 a_20974_43370# a_20556_43646# VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X283 a_14275_46494# a_13759_46122# a_14180_46482# VSS.t1415 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X284 VSS.t1418 a_15051_42282# a_11823_42460.t6 VSS.t1417 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X285 a_1609_45822# a_n443_46116.t25 VDD.t3260 VDD.t3259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X286 a_17517_44484.t0 a_16979_44734# VDD.t1639 VDD.t1638 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X287 VDD.t3755 a_4915_47217.t5 a_12891_46348# VDD.t3754 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 a_20679_44626# a_11967_42832.t46 VSS.t2941 VSS.t2940 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X289 VSS.t1722 a_1423_45028.t5 a_9838_44484# VSS.t1721 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X290 a_13921_42308# a_13259_45724.t19 a_13575_42558# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X291 VCM.t61 a_n784_42308.t6 C0_N_btm.t3 VSS.t1673 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X292 VSS.t2953 a_11599_46634.t39 a_13759_46122# VSS.t2952 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X293 a_14127_45572# a_11823_42460.t19 a_14033_45572# VSS.t3539 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X294 VSS.t1449 a_19998_34978# a_21753_35474# VSS.t1448 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X295 a_13569_43230# a_12379_42858# a_13460_43230# VSS.t1461 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X296 a_5072_46660# a_4955_46873# VSS.t1464 VSS.t1463 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X297 VCM.t58 a_3422_30871.t21 VDAC_P.t7 VSS.t3523 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X298 a_8037_42858# a_7871_42858# VSS.t1466 VSS.t1465 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X299 VSS.t1474 a_22591_46660# a_20820_30879.t3 VSS.t1473 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 VDD.t422 a_n2833_47464# CLK_DATA.t3 VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X301 a_3686_47026# a_2609_46660# a_3524_46660# VDD.t1685 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X302 a_9672_43914# a_10057_43914# a_9801_43940# VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X303 VDD.t1689 a_18429_43548# a_16823_43084# VDD.t1688 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X304 a_17339_46660# a_12861_44030.t35 VDD.t3203 VDD.t3202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 VSS.t1730 a_1606_42308.t6 a_2351_42308# VSS.t1729 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X306 a_16409_43396# a_16243_43396# VSS.t1488 VSS.t1487 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 VSS.t1492 a_9625_46129# a_10044_46482# VSS.t1491 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X308 VDD.t3760 a_n4209_37414.t8 a_n4334_37440# VDD.t3094 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X309 a_13468_44734# a_768_44030.t8 a_13213_44734# VDD.t3679 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X310 VSS.t225 a_n2302_39072# a_n4209_39304.t5 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_2124_47436# a_584_46384.t17 a_2266_47570# VSS.t2781 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X312 VDD.t1930 a_n971_45724.t27 a_2809_45028# VDD.t1929 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X313 a_10809_44734.t2 a_2063_45854.t12 a_10809_44484# VSS.t1643 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X314 a_7577_46660# a_7411_46660# VSS.t904 VSS.t903 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4921_42308# a_4791_45118.t15 VSS.t1761 VSS.t1760 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_16023_47582# a_15507_47210# a_15928_47570# VSS.t1512 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X317 a_12791_45546# a_12861_44030.t31 VDD.t3195 VDD.t3194 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X318 a_10193_42453.t2 a_20712_42282# VSS.t1517 VSS.t1516 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X319 VSS.t1569 a_n881_46662.t15 a_n659_45366# VSS.t1568 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 a_6481_42558# a_n913_45002.t31 a_1755_42282# VDD.t2969 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X321 a_n2956_38680.t3 a_n2472_46090# VSS.t1521 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X322 a_14955_43940# a_14537_43396# a_15037_44260# VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X323 VREF_GND.t32 a_14097_32519.t4 C4_N_btm.t2 VSS.t2678 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X324 VDD.t1736 a_21188_45572# a_21363_45546# VDD.t1735 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 VDD.t486 a_8953_45002# a_2324_44458.t1 VDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X326 a_15682_43940# a_2324_44458.t56 VSS.t3019 VSS.t3018 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 a_18907_42674# a_18727_42674# VDD.t1742 VDD.t1741 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X328 a_12545_42858# a_12379_42858# VSS.t1459 VSS.t1458 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_11967_42832.t29 a_15682_43940# VSS.t430 VSS.t429 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X330 C9_P_btm.t0 a_n4064_39616.t11 VREF_GND.t0 VSS.t2848 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X331 VDAC_P.t4 a_3422_30871.t17 VCM.t55 VSS.t3518 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X332 a_13720_44458# a_9482_43914# VSS.t1096 VSS.t1095 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X333 a_15125_43396# a_15095_43370# a_15037_43396# VSS.t1103 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X334 VREF.t32 a_20692_30879.t4 C6_N_btm.t1 VDD.t2001 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X335 a_2998_44172# a_584_46384.t19 VDD.t3005 VDD.t3004 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X336 a_20974_43370# a_22485_44484# VDD.t632 VDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X337 a_18548_42308# a_18494_42460# a_18057_42282# VSS.t1110 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X338 a_n875_44318# a_n2065_43946# a_n984_44318# VSS.t1391 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X339 a_n2293_42834.t0 a_8049_45260.t5 VDD.t3102 VDD.t3101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X340 VSS.t1116 a_4743_44484# a_4791_45118.t2 VSS.t1115 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X341 a_3626_43646.t5 a_3232_43370.t23 VDD.t3050 VDD.t2914 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X342 VSS.t3678 a_n2438_43548.t41 a_n2433_44484# VSS.t3677 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X343 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD.t1321 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X344 VDD.t1329 a_17973_43940# a_18079_43940# VDD.t1328 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X345 C9_N_btm.t12 a_21588_30879.t5 VREF.t5 VDD.t1774 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X346 VREF_GND.t30 a_17538_32519.t4 C8_N_btm.t6 VSS.t2645 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X347 VDD.t1333 a_22223_46124# a_20205_31679.t1 VDD.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X348 a_4646_46812.t8 a_6298_44484# VDD.t1023 VDD.t1022 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X349 a_4704_46090# a_4883_46098.t4 VDD.t1858 VDD.t1857 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X350 a_5815_47464# a_6151_47436.t8 VDD.t2977 VDD.t2976 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X351 a_17478_45572# a_n881_46662.t19 VDD.t1794 VDD.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X352 DATA[3].t1 a_7227_47204# VDD.t739 VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X353 VDD.t3065 a_n1794_35082.t13 a_18194_34908.t3 VDD.t3064 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 VDD.t202 VSS.t3716 VDD.t201 VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X355 a_17034_45572# a_16327_47482.t41 VSS.t3306 VSS.t3305 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X356 VSS.t2642 a_n3420_39616.t8 a_n2946_39866# VSS.t2641 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X357 a_133_42852# a_n97_42460.t21 a_n13_43084# VDD.t1904 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X358 VDD.t195 VSS.t3762 VDD.t194 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X359 a_n1925_46634.t1 a_8162_45546# VDD.t1349 VDD.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X360 a_21350_47026# a_20273_46660# a_21188_46660# VDD.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X361 VDD.t1355 a_2713_42308# a_2903_42308# VDD.t1354 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X362 a_n3674_39304.t1 a_n2840_42826# VDD.t1357 VDD.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X363 a_13565_43940# a_13059_46348# VDD.t1363 VDD.t1362 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X364 a_n4315_30879.t5 a_n2302_40160# VSS.t1172 VSS.t1171 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 VDD.t430 a_1823_45246# a_2202_46116# VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X366 VSS.t1180 a_n3690_38304# a_n3420_37984.t7 VSS.t1179 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X367 VSS.t3210 VDD.t3784 VSS.t3209 VSS.t3208 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X368 a_2211_45572# a_2063_45854.t13 a_1848_45724# VSS.t1644 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X369 VSS.t1190 a_16112_44458# a_14673_44172# VSS.t1189 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X370 VSS.t1361 a_3316_45546# a_3260_45572# VSS.t1360 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X371 VDD.t3256 a_n443_46116.t21 a_2896_43646# VDD.t3255 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X372 a_n310_47570# a_n971_45724.t29 VSS.t1702 VSS.t1701 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X373 a_21177_47436# a_13507_46334.t7 VSS.t1741 VSS.t1740 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X374 VSS.t3067 a_9290_44172.t20 a_13943_43396# VSS.t3066 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X375 a_n3674_37592.t0 a_196_42282# VDD.t772 VDD.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X376 a_18780_47178# a_18597_46090# VDD.t1396 VDD.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X377 VDD.t176 VSS.t3714 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X378 VSS.t1205 a_8791_42308# a_5934_30871.t3 VSS.t1204 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X379 a_421_43172# a_n97_42460.t15 a_n13_43084# VSS.t1678 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X380 VDD.t1694 a_17339_46660# a_18051_46116# VDD.t1693 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X381 VDD.t1015 a_6298_44484# a_4646_46812.t9 VDD.t1014 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X382 VSS.t1206 a_n2840_46090# a_n2956_39304.t3 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X383 a_n2661_43370.t0 a_10907_45822# VDD.t1410 VDD.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X384 a_9396_43370# a_4883_46098.t5 VDD.t1860 VDD.t1859 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X385 VDD.t1412 a_19333_46634# a_19123_46287# VDD.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X386 a_n2438_43548.t21 a_949_44458# VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X387 a_5755_42852# a_n97_42460.t19 a_5837_43172# VSS.t1680 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X388 a_n4251_39392# a_n4318_39304.t4 a_n4334_39392# VSS.t1664 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X389 a_805_46414# a_472_46348# VSS.t1219 VSS.t1218 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X390 VDD.t1327 a_n1076_43230# a_n901_43156# VDD.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X391 a_21845_43940# a_12549_44172.t28 a_19692_46634.t2 VDD.t2950 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X392 VDD.t1424 a_4520_42826# a_4093_43548# VDD.t1423 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X393 a_12469_46902# a_12251_46660# VSS.t1226 VSS.t1225 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X394 a_15415_45028# a_15227_44166.t17 VSS.t3595 VSS.t3594 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X395 a_19479_31679.t1 a_22223_45572# VDD.t1433 VDD.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X396 a_7542_44172# a_7499_43078# VDD.t522 VDD.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X397 a_3080_42308.t2 a_2903_42308# VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X398 VSS.t1232 a_22165_42308# a_22223_42860# VSS.t1231 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X399 VDD.t1583 a_10249_46116# a_11186_47026# VDD.t1582 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X400 a_3905_42558# a_2382_45260# a_3823_42558# VDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X401 a_12347_46660# a_11901_46660# a_12251_46660# VSS.t1239 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X402 VSS.t386 a_16137_43396# a_16414_43172# VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X403 a_5066_45546# a_4791_45118.t23 VSS.t1771 VSS.t1770 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X404 a_14581_44484# a_13249_42308# VSS.t1246 VSS.t1245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X405 VREF.t57 a_n4209_39590.t12 C9_P_btm.t13 VDD.t3075 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X406 a_2113_38308# a_1273_38525.t9 VSS.t1806 VSS.t1805 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X407 a_n473_42460# a_n755_45592.t23 a_n327_42558# VDD.t3450 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X408 VDD.t1454 a_n1699_43638# a_n1809_43762# VDD.t1453 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X409 a_13759_47204# a_13717_47436.t2 a_13675_47204# VDD.t2886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X410 a_n3420_39616.t4 a_n3690_39616# VSS.t1362 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X411 C4_N_btm.t0 EN_VIN_BSTR_N.t20 VIN_N.t15 VSS.t2926 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X412 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS.t1377 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X413 a_2779_44458# a_1423_45028.t6 VSS.t1724 VSS.t1723 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X414 VDD.t390 a_19319_43548# a_19268_43646# VDD.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X415 C10_P_btm.t3 a_4190_30871.t19 VCM.t13 VSS.t2816 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X416 VDD.t1460 a_9127_43156# a_5891_43370.t1 VDD.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X417 a_1123_46634# a_948_46660# a_1302_46660# VSS.t1262 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X418 a_n755_45592.t6 a_n809_44244# VSS.t359 VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X419 a_2952_47436# a_3160_47472# a_3094_47570# VSS.t1273 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X420 a_5807_45002# a_16763_47508# VDD.t889 VDD.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X421 a_3726_37500# a_3754_38470.t3 VDAC_Ni.t5 VSS.t2632 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X422 a_6293_42852# a_5755_42852# VSS.t1215 VSS.t1214 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X423 a_8120_45572# a_8034_45724# a_n1925_46634.t3 VSS.t1285 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X424 a_11541_44484# a_11691_44458.t6 VSS.t2889 VSS.t2888 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X425 C10_P_btm.t29 a_n4315_30879.t23 VREF.t47 VDD.t2083 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X426 VSS.t736 a_10083_42826# a_7499_43078# VSS.t735 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X427 a_5257_43370# a_5907_46634# VDD.t1497 VDD.t1496 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X428 a_4880_45572# a_5066_45546# VSS.t170 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X429 VIN_P.t2 EN_VIN_BSTR_P.t23 C0_P_btm.t3 VSS.t3574 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X430 C9_P_btm.t15 a_n4209_39590.t13 VREF.t58 VDD.t3076 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X431 a_3497_42558# a_1823_45246# VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X432 VSS.t1266 a_1123_46634# a_584_46384.t6 VSS.t1265 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 a_16223_45938# a_16327_47482.t19 VDD.t3413 VDD.t3412 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X434 a_4883_46098.t0 a_21363_46634# VDD.t1510 VDD.t1509 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X435 a_2711_45572.t1 a_768_44030.t23 VDD.t3692 VDD.t3691 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X436 VSS.t1304 a_2553_47502# a_2487_47570# VSS.t1303 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X437 VDD.t1430 a_12469_46902# a_12359_47026# VDD.t1429 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X438 a_6453_43914# a_6109_44484# VSS.t1306 VSS.t1305 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X439 a_7765_42852# a_7227_42852# VDD.t1517 VDD.t1516 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X440 VDD.t182 VSS.t3735 VDD.t181 VDD.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X441 a_17786_45822# a_15861_45028# a_17478_45572# VDD.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X442 a_18450_45144# a_15227_44166.t23 VDD.t3676 VDD.t3675 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X443 a_6765_43638# a_6547_43396# VSS.t1393 VSS.t1392 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X444 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD.t1591 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X445 VSS.t2062 a_n4334_40480# a_n4064_40160.t5 VSS.t2061 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X446 a_12089_42308# a_11551_42558# VDD.t866 VDD.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X447 a_16547_43609# a_16414_43172# VDD.t1446 VDD.t1445 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X448 a_3221_46660# a_3177_46902# a_3055_46660# VSS.t2073 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X449 a_6667_45809# a_6472_45840# a_6977_45572# VSS.t286 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X450 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD.t2328 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X451 a_6643_43396# a_6197_43396# a_6547_43396# VSS.t2078 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X452 a_5837_45348# a_5807_45002# VSS.t1279 VSS.t1278 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X453 a_5565_43396# a_4905_42826# VSS.t1351 VSS.t1350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X454 a_7418_45067# a_7229_43940# VDD.t2336 VDD.t2335 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X455 a_1307_43914.t5 a_2779_44458# VSS.t487 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X456 a_1793_42852# a_742_44458# a_1709_42852# VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 VDD.t1854 a_10227_46804.t31 a_10083_42826# VDD.t1853 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 a_11301_43218# a_10922_42852# a_11229_43218# VSS.t2083 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X459 VSS.t2085 a_13291_42460# a_13249_42308# VSS.t2084 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X460 a_18341_45572# a_18175_45572# VDD.t2342 VDD.t2341 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X461 w_1575_34786.t12 a_n1057_35014.t4 w_1575_34786.t11 w_1575_34786.t10 sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X462 a_19113_45348# a_19321_45002# VSS.t1330 VSS.t1329 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X463 VDD.t214 VSS.t3730 VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X464 a_8696_44636.t1 a_16855_45546# VSS.t2094 VSS.t2093 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X465 a_12189_44484# a_8975_43940# VSS.t2096 VSS.t2095 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X466 a_n1736_46482# a_n1853_46287# VDD.t2353 VDD.t2352 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X467 a_1239_47204# a_1209_47178# VDD.t2357 VDD.t2356 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X468 VSS.t3476 a_n1696_34930.t11 a_n217_35014# VSS.t3475 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X469 VDD.t3403 VDAC_Ni.t10 a_6886_37412# VSS.t3348 sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X470 a_n4064_37984.t6 a_n4334_38304# VSS.t2111 VSS.t1346 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X471 a_1606_42308.t0 a_1576_42282# VDD.t274 VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X472 VDD.t3717 a_n443_42852.t19 a_6481_42558# VDD.t3716 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X473 VDD.t2367 a_12005_46116# a_n1741_47186.t3 VDD.t2366 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X474 a_18315_45260# a_18587_45118# VSS.t2116 VSS.t2115 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 VSS.t3623 a_768_44030.t25 a_3600_43914# VSS.t3622 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X476 VDD.t2925 a_4958_30871.t9 a_17531_42308# VDD.t2924 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X477 a_16795_42852# a_n97_42460.t23 a_16877_42852# VDD.t1906 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X478 a_18900_46660# a_18834_46812# a_18285_46348# VSS.t2125 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X479 VDD.t90 VSS.t3705 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X480 a_17973_43940# a_17737_43940# VSS.t2129 VSS.t2128 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X481 a_6419_46155# a_5257_43370# a_6347_46155# VDD.t1504 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X482 a_18597_46090# a_19431_45546# VSS.t2133 VSS.t2132 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X483 a_3737_43940# a_3537_45260.t27 VDD.t2915 VDD.t2914 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X484 comp_n a_1169_39043# VDD.t356 VDD.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 VDD.t424 a_1823_45246# a_4419_46090# VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X486 a_22848_40945# COMP_P.t8 a_22589_40599# VSS.t1705 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X487 VDD.t2396 a_4007_47204# DATA[2].t3 VDD.t2395 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X488 VSS.t2151 a_21496_47436# a_13507_46334.t1 VSS.t2150 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X489 VDD.t2404 a_n2002_35448# SMPL_ON_P.t3 VDD.t2403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X490 VSS.t2163 a_10723_42308# a_5742_30871.t3 VSS.t2162 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X491 a_22737_36887# a_22527_39145# a_22629_37990# VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X492 a_11823_42460.t4 a_15051_42282# VSS.t1424 VSS.t1423 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 VSS.t2874 a_n4209_38216.t9 a_n4251_38304# VSS.t2679 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X494 a_12891_46348# a_4915_47217.t6 VDD.t3757 VDD.t3756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 VSS.t1440 a_20679_44626# a_20640_44752# VSS.t1439 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X496 a_21115_43940# a_20935_43940# VDD.t2418 VDD.t2417 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X497 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS.t2074 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X498 VSS.t3107 VDD.t3808 VSS.t3106 VSS.t3105 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X499 VDD.t2424 a_10951_45334# a_10775_45002# VDD.t2423 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X500 a_20850_46155# a_19692_46634.t7 VDD.t2064 VDD.t2063 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X501 VDD.t3123 a_13661_43548.t23 a_18587_45118# VDD.t3122 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X502 a_11649_44734# a_3232_43370.t19 a_n2661_44458.t0 VDD.t3047 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X503 a_20820_30879.t2 a_22591_46660# VSS.t1472 VSS.t1471 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X504 VSS.t2175 a_21359_45002# a_21101_45002# VSS.t2174 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X505 EN_VIN_BSTR_N.t3 a_18194_34908.t11 w_10694_33990.t17 w_10694_33990.t16 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X506 a_17364_32525.t3 a_22959_43396# VSS.t2179 VSS.t2178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X507 a_18989_43940# a_18451_43940# VSS.t2183 VSS.t2182 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X508 a_6197_43396# a_6031_43396# VSS.t2185 VSS.t2184 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 VDD.t1642 a_12891_46348# a_13213_44734# VDD.t1641 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X510 a_8912_37509.t16 VDAC_N.t8 a_5700_37509.t9 VDD.t69 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X511 VREF_GND.t44 a_13467_32519.t4 C1_N_btm.t1 VSS.t1731 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X512 VDD.t3001 a_584_46384.t13 a_3540_43646# VDD.t3000 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X513 a_8873_43396# a_5891_43370.t17 a_8791_43396# VSS.t1575 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X514 C10_N_btm.t21 a_22612_30879.t17 VREF.t25 VDD.t1952 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X515 VSS.t600 a_n4334_39392# a_n4064_39072.t7 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X516 C9_P_btm.t4 a_4958_30871.t11 VCM.t37 VSS.t2698 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X517 a_10809_44484# a_10057_43914# VSS.t135 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X518 C6_N_btm.t4 a_5742_30871.t5 VCM.t25 VSS.t1553 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X519 a_6545_47178# a_6419_46155# VDD.t2383 VDD.t2382 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X520 a_11599_46634.t13 a_15682_46116# VDD.t1062 VDD.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X521 a_6109_44484# a_5518_44484# VDD.t2446 VDD.t2445 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X522 a_n4318_38216.t3 a_n2472_42282# VSS.t2197 VSS.t2196 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X523 VDD.t2452 a_n901_46420# a_n443_46116.t0 VDD.t2451 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X524 a_13258_32519.t3 a_19647_42308# VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X525 VDD.t3154 a_11599_46634.t35 a_18819_46122# VDD.t3153 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X526 a_18194_34908.t5 a_n1794_35082.t15 VSS.t2855 VSS.t2854 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X527 a_n1435_47204.t0 a_n1605_47204# VDD.t2466 VDD.t2465 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X528 VDD.t482 a_8953_45002# a_2324_44458.t5 VDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X529 a_15682_43940# a_2324_44458.t54 VSS.t3017 VSS.t3016 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X530 C10_P_btm.t15 a_n4064_40160.t13 VREF_GND.t38 VSS.t2685 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X531 a_14113_42308# a_13575_42558# VDD.t1653 VDD.t1652 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X532 VSS.t2876 a_4646_46812.t33 a_4651_46660# VSS.t2875 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X533 a_13381_47204# a_12549_44172.t31 VDD.t2954 VDD.t2953 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X534 VSS.t1520 a_n2472_46090# a_n2956_38680.t2 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X535 a_4958_30871.t0 a_17124_42282# VDD.t560 VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X536 VSS.t1234 a_22223_42860# a_22400_42852# VSS.t1233 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X537 C0_P_btm.t0 a_n3565_37414.t8 VREF.t53 VDD.t2955 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X538 VDD.t2472 a_1208_46090# a_472_46348# VDD.t2471 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X539 VSS.t1387 a_18479_47436# a_19452_47524# VSS.t1386 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 VSS.t221 a_n2302_39072# a_n4209_39304.t6 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X541 a_5088_37509.t15 VDAC_P.t10 a_8912_37509.t4 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X542 a_n443_46116.t1 a_n901_46420# VDD.t2456 VDD.t2455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X543 a_20623_45572# a_20107_45572# a_20528_45572# VSS.t2225 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X544 a_12281_43396# a_9290_44172.t26 VSS.t3071 VSS.t3070 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X545 VSS.t2843 a_n1794_35082.t11 a_18194_34908.t6 VSS.t2842 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X546 C1_P_btm.t2 a_n4209_37414.t9 VREF.t72 VDD.t3761 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X547 VSS.t3522 a_n3565_39304.t9 a_n3607_39392# VSS.t3521 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X548 a_15486_42560# a_15764_42576# a_15720_42674# VDD.t2480 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X549 VSS.t3332 a_n1613_43370.t29 a_8649_43218# VSS.t3331 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X550 a_15765_45572# a_15599_45572# VDD.t537 VDD.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X551 VSS.t535 a_n2946_39866# a_n3565_39590.t4 VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X552 a_n1613_43370.t2 a_5815_47464# VDD.t1345 VDD.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X553 VSS.t2236 a_14495_45572# a_n881_46662.t3 VSS.t2235 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X554 a_4646_46812.t10 a_6298_44484# VDD.t1009 VDD.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X555 a_10617_44484# a_10440_44484# VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X556 VDD.t1104 a_5111_44636# a_8487_44056# VDD.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X557 VREF.t59 a_n4209_39590.t15 C9_P_btm.t10 VDD.t3078 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X558 VCM.t20 a_5932_42308.t4 C3_N_btm.t3 VSS.t1802 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X559 a_20708_46348# a_15227_44166.t13 a_20850_46155# VDD.t3666 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X560 a_n2267_44484# a_n2433_44484# VSS.t1120 VSS.t1119 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X561 a_4646_46812.t14 a_6298_44484# VDD.t1027 VDD.t1026 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X562 a_1115_44172# a_453_43940# VSS.t2242 VSS.t2241 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X563 VSS.t1707 COMP_P.t9 a_n1329_42308# VSS.t1706 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X564 VSS.t2252 a_1847_42826# a_2905_42968# VSS.t2251 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X565 VSS.t1312 a_15861_45028# a_17023_45118# VSS.t1311 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X566 a_16292_46812# a_5807_45002# a_16434_46660# VSS.t1282 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X567 a_17325_44484# a_15227_44166.t21 a_16979_44734# VSS.t3599 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X568 a_n4064_39072.t6 a_n4334_39392# VSS.t599 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X569 a_15803_42450# a_11967_42832.t45 VDD.t3148 VDD.t3147 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X570 a_5534_30871.t1 a_12563_42308# VDD.t454 VDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X571 VSS.t2262 a_3381_47502# a_3315_47570# VSS.t2261 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X572 VDD.t2512 a_9863_46634# a_2063_45854.t0 VDD.t2511 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X573 VDD.t290 a_n2840_43370# a_n4318_39304.t1 VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X574 VSS.t2775 a_584_46384.t11 a_3457_43396# VSS.t2774 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X575 VIN_N.t10 EN_VIN_BSTR_N.t19 C3_N_btm.t0 VSS.t2925 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X576 a_3863_42891# a_3681_42891# VDD.t677 VDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X577 VDD.t877 a_9049_44484# a_9313_45822# VDD.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X578 VDD.t350 a_376_46348# a_171_46873# VDD.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X579 a_11541_44484# a_11453_44696.t2 a_n2661_44458.t1 VSS.t3632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X580 VDD.t2113 a_1431_47204# DATA[1].t0 VDD.t2112 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X581 a_19553_46090# a_19335_46494# VSS.t1860 VSS.t1859 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X582 a_n1613_43370.t5 a_5815_47464# VSS.t1140 VSS.t1139 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X583 a_18727_42674# a_n1059_45260.t17 VSS.t2768 VSS.t2767 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X584 a_n1925_42282.t0 a_4185_45028.t4 VDD.t1894 VDD.t1893 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X585 VDD.t705 a_n2302_37984# a_n4209_38216.t1 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X586 VSS.t1863 a_17591_47464# a_16327_47482.t5 VSS.t1862 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X587 VSS.t1184 a_n3690_38304# a_n3420_37984.t6 VSS.t1183 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X588 VDD.t2133 a_19164_43230# a_19339_43156# VDD.t2132 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X589 a_2479_44172# a_2905_42968# VSS.t2254 VSS.t2253 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X590 VSS.t1794 a_4361_42308.t2 a_21855_43396# VSS.t1793 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X591 a_n1741_47186.t0 a_12891_46348# a_12839_46116# VDD.t1644 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X592 VDD.t1 a_8103_44636# a_7640_43914# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X593 a_8192_45572# a_8162_45546# a_8120_45572# VSS.t1149 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X594 a_5009_45028# a_3090_45724.t15 a_4927_45028# VDD.t1819 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X595 a_12549_44172.t2 a_20567_45036# VSS.t1889 VSS.t1888 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X596 VSS.t746 a_n2840_42282# a_n3674_38680.t3 VSS.t745 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X597 a_5129_47502# a_4791_45118.t17 VSS.t1763 VSS.t1762 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X598 a_14840_46494# a_13759_46122# a_14493_46090# VDD.t1627 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X599 VSS.t3005 a_2324_44458.t44 a_949_44458# VSS.t3004 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X600 VDD.t3133 EN_VIN_BSTR_N.t13 w_10694_33990.t1 w_10694_33990.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X601 VSS.t2739 a_n913_45002.t25 a_2713_42308# VSS.t2738 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X602 VDD.t689 a_n863_45724# a_1221_42558# VDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X603 a_8601_46660# a_7411_46660# a_8492_46660# VSS.t906 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X604 a_2307_45899# a_n237_47217.t11 a_1848_45724# VDD.t3241 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X605 VDD.t3591 a_7754_40130.t10 a_8912_37509.t35 VDD.t3590 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X606 VDD.t1971 a_n4209_39304.t10 a_n4334_39392# VDD.t1970 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X607 VSS.t3254 VDD.t3801 VSS.t3253 VSS.t3144 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X608 a_n2946_39072# a_n2956_39304.t4 VSS.t1735 VSS.t1734 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X609 a_15861_45028# a_15595_45028# VSS.t1901 VSS.t1900 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X610 VSS.t3140 VDD.t3819 VSS.t3139 VSS.t3138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X611 VSS.t3342 a_n1613_43370.t39 a_3221_46660# VSS.t3341 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X612 a_1756_43548# a_768_44030.t21 a_1987_43646# VDD.t3690 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X613 a_3754_39134# a_7754_39300# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X614 VSS.t3134 VDD.t3817 VSS.t3133 VSS.t3132 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X615 a_n4318_40392.t3 a_n2840_44458# VSS.t1903 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X616 a_5700_37509.t17 VDAC_N.t21 a_8912_37509.t29 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X617 VSS.t1906 a_18143_47464# a_12861_44030.t4 VSS.t1905 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X618 a_19332_42282# a_19511_42282# VSS.t1914 VSS.t1913 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X619 VSS.t1922 a_17583_46090# a_13259_45724.t3 VSS.t1921 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 VSS.t3249 VDD.t3799 VSS.t3248 VSS.t3247 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X621 a_20623_43914# a_19321_45002# VDD.t1540 VDD.t1539 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X622 VSS.t131 a_17499_43370# a_n1059_45260.t6 VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X623 VSS.t1931 a_7754_38470# a_6886_37412# VSS.t1930 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X624 a_n3420_39616.t5 a_n3690_39616# VSS.t1364 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X625 a_4185_45348# a_3065_45002# VSS.t375 VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X626 a_n2661_46634.t0 a_13017_45260# VDD.t2190 VDD.t2189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X627 VDD.t1542 a_19321_45002# a_20567_45036# VDD.t1541 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X628 VDD.t2444 a_6545_47178# a_6575_47204# VDD.t2443 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X629 VDD.t2379 a_18285_46348# a_18051_46116# VDD.t2378 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X630 a_2864_46660# a_2747_46873# VDD.t749 VDD.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X631 VSS.t365 a_n809_44244# a_n755_45592.t4 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X632 VSS.t3243 VDD.t3797 VSS.t3242 VSS.t3228 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X633 VDD.t3536 a_1307_43914.t29 a_2253_43940# VDD.t3535 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X634 a_n2002_35448# a_n1550_35448# VDD.t2194 VDD.t2193 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X635 a_13351_46090# a_13507_46334.t9 VSS.t1743 VSS.t1742 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X636 a_18374_44850# a_18248_44752# a_17970_44736# VSS.t1945 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X637 a_n913_45002.t10 a_1307_43914.t19 a_2075_43172# VSS.t3462 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X638 VDD.t628 a_15682_43940# a_11967_42832.t2 VDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X639 a_13657_42308# a_11823_42460.t29 VSS.t3551 VSS.t3550 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X640 a_375_42282# a_413_45260.t2 VDD.t2104 VDD.t2103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 a_3090_45724.t0 a_19321_45002# VDD.t1536 VDD.t1535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X642 a_n1696_34930.t6 a_n1794_35082.t9 VSS.t2841 VSS.t2840 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X643 a_10334_44484# a_10157_44484# VDD.t2206 VDD.t2205 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X644 VSS.t3097 a_10903_43370.t12 a_10057_43914# VSS.t3096 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X645 a_5700_37509.t2 VSS.t3743 VDAC_Pi.t2 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X646 a_2113_38308# a_2113_38308# a_2113_38308# VSS.t86 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X647 VSS.t3674 a_n2438_43548.t37 a_n133_46660# VSS.t3673 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X648 a_584_46384.t5 a_1123_46634# VSS.t1272 VSS.t1271 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 VSS.t1957 a_22959_46124# a_20692_30879.t3 VSS.t760 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 a_n3674_39768.t1 a_n2472_43914# VDD.t2214 VDD.t2213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X651 VREF.t31 a_n4209_39304.t11 C7_P_btm.t3 VDD.t1972 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X652 VSS.t1963 a_20107_42308# a_7174_31319.t3 VSS.t1962 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X653 a_n4209_39590.t4 a_n2302_39866# VSS.t862 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 a_526_44458.t4 a_3147_46376# VSS.t1971 VSS.t1970 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X655 VREF_GND.t39 a_n4064_40160.t15 C10_P_btm.t12 VSS.t2688 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X656 a_20301_43646# a_19692_46634.t8 a_20556_43646# VDD.t2065 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X657 VDD.t2454 a_n901_46420# a_n914_46116# VDD.t2453 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X658 a_n971_45724.t1 a_104_43370# VDD.t1124 VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X659 a_20447_31679.t1 a_22959_45572# VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X660 VSS.t1975 a_13348_45260# a_13159_45002# VSS.t1974 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X661 a_n4334_38304# a_n4318_38216.t4 VDD.t2044 VDD.t2043 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X662 VSS.t1571 a_n881_46662.t17 a_6517_45366# VSS.t1570 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X663 a_8685_42308# a_8515_42308# VDD.t2234 VDD.t2233 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X664 VSS.t1983 a_6491_46660# a_6851_47204# VSS.t1982 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X665 a_768_44030.t2 a_13487_47204# VDD.t796 VDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X666 VDD.t2156 a_14493_46090# a_14383_46116# VDD.t2155 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X667 a_n327_42308# a_n357_42282.t16 VSS.t1837 VSS.t1836 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X668 a_22485_44484# a_22315_44484# VDD.t2243 VDD.t2242 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X669 a_15673_47210# a_15507_47210# VSS.t1510 VSS.t1509 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X670 a_8605_42826# a_8387_43230# VSS.t1993 VSS.t1992 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X671 a_1709_42852# a_n863_45724# VDD.t697 VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 a_5700_37509.t4 VDAC_N.t17 a_8912_37509.t25 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X673 VDD.t901 a_n1736_42282# a_n4318_37592.t1 VDD.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X674 VREF.t71 a_19721_31679.t4 C2_N_btm.t3 VDD.t3702 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X675 VSS.t1996 a_895_43940# a_2537_44260# VSS.t1995 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X676 VSS.t3180 VDD.t3773 VSS.t3179 VSS.t3178 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X677 a_17609_46634# a_12861_44030.t29 VDD.t3193 VDD.t3192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X678 VDD.t3156 a_11599_46634.t36 a_18175_45572# VDD.t3155 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X679 a_8945_43396# a_3537_45260.t17 a_8873_43396# VSS.t2669 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X680 a_13249_42308# a_10903_43370.t20 VSS.t3101 VSS.t3100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X681 a_601_46902# a_383_46660# VSS.t2000 VSS.t1999 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X682 a_4640_45348# a_4574_45260# a_4558_45348# VSS.t2002 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X683 a_n467_45028# a_n745_45366# VDD.t2263 VDD.t2262 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X684 a_1208_46090# a_765_45546.t8 a_1337_46116# VDD.t3763 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X685 a_3820_44260# a_2382_45260# VSS.t151 VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X686 VSS.t514 a_n863_45724# a_2905_42968# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X687 VSS.t2009 a_16721_46634# a_16655_46660# VSS.t2008 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X688 C5_P_btm.t3 a_n4064_38528.t8 VREF_GND.t26 VSS.t1786 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X689 a_21588_30879.t1 a_22223_47212# VDD.t2270 VDD.t2269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X690 a_16877_42852# a_16823_43084# a_16795_42852# VDD.t1690 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X691 a_11967_42832.t22 a_15682_43940# VSS.t436 VSS.t435 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X692 VSS.t2017 a_17715_44484# a_17737_43940# VSS.t2016 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X693 a_16241_47178# a_16023_47582# VDD.t1723 VDD.t1722 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X694 a_12359_47026# a_11735_46660# a_12251_46660# VDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X695 VDD.t109 VSS.t3719 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X696 a_5883_43914# a_8333_44056# VDD.t2278 VDD.t2277 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X697 a_16759_43396# a_16409_43396# a_16664_43396# VDD.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X698 VDD.t3612 a_n3565_39590.t11 a_n3690_39616# VDD.t3611 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X699 a_17665_42852# a_17595_43084# a_14539_43914# VDD.t2281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X700 VSS.t3670 a_n2438_43548.t35 a_n2157_42858# VSS.t3669 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X701 VDD.t2394 a_4007_47204# DATA[2].t0 VDD.t2393 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X702 a_1990_45572# a_167_45260# VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X703 a_2324_44458.t9 a_8953_45002# VDD.t496 VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X704 a_5072_46660# a_4955_46873# VDD.t1673 VDD.t1672 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X705 a_22889_38993# a_22400_42852# VSS.t1398 VSS.t1397 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X706 VDD.t2046 a_3357_43084.t3 a_22591_45572# VDD.t2045 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X707 VSS.t1410 a_3815_47204# a_4007_47204# VSS.t1409 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X708 a_1666_39587.t1 a_1666_39043.t4 a_2112_39137# VSS.t2715 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X709 a_15803_42450# a_11967_42832.t35 VSS.t2931 VSS.t2930 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X710 a_20528_46660# a_20411_46873# VDD.t2289 VDD.t2288 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 a_n3607_39392# a_n3674_39304.t4 a_n3690_39392# VSS.t2640 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X712 VDD.t3063 a_n4064_39616.t12 a_n2216_39866# VDD.t2922 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X713 a_21421_42336# a_16327_47482.t27 a_21335_42336# VSS.t3367 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X714 a_6655_43762# a_n1613_43370.t27 VDD.t3378 VDD.t3377 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X715 a_14371_46494# a_13925_46122# a_14275_46494# VSS.t809 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X716 VSS.t3186 VDD.t3775 VSS.t3185 VSS.t3184 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X717 VDD.t761 a_3503_45724# a_3218_45724# VDD.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X718 VDD.t460 a_n2840_43914# a_n4318_39768.t1 VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X719 a_15037_43940# a_13556_45296# a_14955_43940# VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X720 VSS.t639 a_n901_43156# a_n443_42852.t7 VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VDD.t712 a_10467_46802# a_10428_46928# VDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X722 a_15060_45348# a_13661_43548.t13 a_14976_45348# VSS.t2895 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X723 a_9895_44260# a_9290_44172.t16 a_9801_44260# VSS.t3063 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X724 VDD.t2297 a_6171_42473# a_5379_42460# VDD.t2296 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X725 a_5009_45028# a_5147_45002# a_5093_45028# VDD.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X726 a_13904_45546# a_10903_43370.t14 a_14127_45572# VSS.t3098 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X727 a_3537_45260.t7 a_7287_43370# VSS.t676 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X728 SMPL_ON_N.t3 a_21753_35474# VDD.t1661 VDD.t1660 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X729 a_19900_46494# a_18985_46122# a_19553_46090# VSS.t2044 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X730 VDD.t1956 a_8696_44636.t4 a_17478_45572# VDD.t1955 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X731 C10_P_btm.t6 a_4190_30871.t21 VCM.t16 VSS.t2818 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X732 a_3935_42891# a_3905_42865# a_3863_42891# VDD.t2305 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X733 DATA[0].t3 a_327_47204# VDD.t2316 VDD.t2315 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X734 VSS.t1565 a_n881_46662.t11 a_11117_47542# VSS.t1564 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X735 C3_P_btm.t2 EN_VIN_BSTR_P.t20 VIN_P.t7 VSS.t3574 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X736 VSS.t160 a_n4334_39616# a_n4064_39616.t4 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X737 DATA[2].t5 a_4007_47204# VSS.t2147 VSS.t2146 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X738 a_15682_46116# a_2324_44458.t41 VDD.t3213 VDD.t3212 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X739 a_1057_46660# a_n133_46660# a_948_46660# VSS.t1955 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X740 VREF.t49 a_n4315_30879.t25 C10_P_btm.t31 VDD.t2085 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X741 a_11599_46634.t0 a_15682_46116# VDD.t1066 VDD.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X742 VSS.t1783 a_2982_43646.t6 a_21487_43396# VSS.t1782 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X743 a_21363_45546# a_21188_45572# a_21542_45572# VSS.t1524 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X744 VSS.t3536 a_11823_42460.t15 a_11322_45546# VSS.t3535 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_18204_44850# a_17767_44458# VDD.t988 VDD.t987 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X746 a_n447_43370# a_n2497_47436# VSS.t2394 VSS.t2393 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X747 a_17324_43396# a_16409_43396# a_16977_43638# VSS.t805 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X748 VSS.t1788 a_n4064_38528.t9 a_n2302_38778# VSS.t1787 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 a_n443_42852.t6 a_n901_43156# VSS.t637 VSS.t636 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X750 a_15095_43370# a_15567_42826# VSS.t2404 VSS.t2403 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X751 a_10150_46912# a_10428_46928# a_10384_47026# VDD.t2295 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X752 VSS.t2199 a_n2472_42282# a_n4318_38216.t2 VSS.t2198 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X753 VDD.t1659 a_21753_35474# SMPL_ON_N.t0 VDD.t1658 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X754 a_8492_46660# a_7577_46660# a_8145_46902# VSS.t1505 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X755 a_5649_42852.t1 a_5111_42852# VSS.t1353 VSS.t1292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X756 VDD.t2657 a_18287_44626# a_18248_44752# VDD.t2656 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X757 a_20894_47436# a_20990_47178# VDD.t2660 VDD.t2659 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X758 a_19636_46660# a_19594_46812# a_19333_46634# VSS.t2414 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X759 a_10249_46116# a_9823_46155# VSS.t587 VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X760 VDD.t168 VSS.t3755 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X761 a_10227_46804.t1 a_14955_47212# VDD.t811 VDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X762 a_739_46482# a_n743_46660.t6 a_376_46348# VSS.t3556 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X763 VSS.t2173 a_10775_45002# a_10180_45724# VSS.t2172 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X764 a_2896_43646# a_2479_44172# a_2982_43646.t5 VDD.t2139 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X765 VSS.t890 a_15682_46116# a_11599_46634.t17 VSS.t889 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X766 a_12791_45546# a_12861_44030.t19 VSS.t2980 VSS.t2979 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X767 VSS.t1275 a_5807_45002# a_11691_44458.t3 VSS.t1274 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X768 VSS.t1797 a_3357_43084.t4 a_22591_45572# VSS.t1796 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X769 VSS.t153 a_2382_45260# a_2304_45348# VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X770 a_n4315_30879.t0 a_n2302_40160# VDD.t1374 VDD.t1048 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X771 VDD.t2458 a_n901_46420# a_n443_46116.t2 VDD.t2457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X772 a_6298_44484# a_2324_44458.t39 VDD.t3209 VDD.t3208 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 a_949_44458# a_2324_44458.t37 VSS.t2999 VSS.t2998 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X774 VDD.t1128 a_2277_45546# a_2307_45899# VDD.t1127 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X775 a_10053_45546# a_8746_45002# a_10306_45572# VSS.t344 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X776 a_18194_34908.t4 a_n1794_35082.t7 VSS.t2839 VSS.t2838 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X777 a_n2956_39768.t1 a_n2840_46634# VDD.t1134 VDD.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X778 VDD.t2042 a_4361_42308.t3 a_21855_43396# VDD.t2041 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X779 VDD.t2129 a_17591_47464# a_16327_47482.t2 VDD.t2128 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X780 VSS.t1824 a_6945_45028.t3 a_22223_46124# VSS.t1823 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X781 VDD.t1499 a_5257_43370# a_5263_45724# VDD.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X782 a_n3565_39590.t3 a_n2946_39866# VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X783 VDD.t121 VSS.t3750 VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X784 VDAC_Ni.t3 VSS.t3748 a_5088_37509.t19 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X785 a_18494_42460# a_18907_42674# VSS.t1531 VSS.t1530 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X786 VDD.t136 VSS.t3746 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X787 a_n1151_42308.t0 a_n1329_42308# VDD.t2497 VDD.t2496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X788 a_16763_47508# a_16327_47482.t21 VDD.t3415 VDD.t3414 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X789 a_21259_43561# a_4190_30871.t17 VDD.t3032 VDD.t2419 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X790 a_8349_46414# a_8016_46348# VDD.t1140 VDD.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X791 VDD.t2119 a_1431_47204# DATA[1].t3 VDD.t2118 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X792 a_17970_44736# a_18287_44626# a_18245_44484# VSS.t2409 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X793 a_1123_46634# a_n1613_43370.t37 VDD.t3388 VDD.t3387 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X794 a_n237_47217.t1 a_8667_46634# VDD.t909 VDD.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X795 a_5837_42852# a_3537_45260.t19 a_5755_42852# VDD.t1717 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X796 VSS.t1816 a_19692_46634.t10 a_19636_46660# VSS.t1815 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X797 a_8697_45572# a_3483_46348.t21 VSS.t3088 VSS.t3087 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X798 a_1145_45348# a_n863_45724# a_626_44172# VSS.t508 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X799 VSS.t3611 a_5934_30871.t5 a_8515_42308# VSS.t3610 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X800 VSS.t2104 a_1239_47204# a_1431_47204# VSS.t2103 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X801 VSS.t1869 a_17591_47464# a_16327_47482.t4 VSS.t1868 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X802 a_11173_44260# a_10729_43914# VSS.t950 VSS.t949 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X803 VDD.t2361 a_n4334_38304# a_n4064_37984.t1 VDD.t1709 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X804 a_22165_42308# a_21887_42336# VSS.t954 VSS.t953 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X805 a_5244_44056# a_5147_45002# VSS.t671 VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X806 VSS.t1779 a_n4064_37440.t8 a_n2302_37690# VSS.t1778 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X807 VDD.t1156 a_8952_43230# a_9127_43156# VDD.t1155 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X808 a_n2956_37592.t1 a_n2472_45002# VDD.t1158 VDD.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X809 VSS.t971 a_2127_44172# a_n2661_45010# VSS.t970 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X810 VSS.t975 a_15493_43940# a_22959_43948# VSS.t974 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X811 a_n3565_38502.t6 a_n2946_38778# VSS.t698 VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X812 VSS.t3230 VDD.t3792 VSS.t3229 VSS.t3228 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X813 VSS.t35 a_949_44458# a_n2438_43548.t19 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X814 a_19339_43156# a_16327_47482.t25 VDD.t3421 VDD.t3420 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X815 VDD.t1172 a_n1920_47178# a_n2312_39304.t1 VDD.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X816 VDD.t1178 a_n1177_44458# a_n1190_44850# VDD.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X817 VDD.t1585 a_16292_46812# a_15811_47375# VDD.t1584 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X818 a_5164_46348# a_4927_45028# VDD.t2148 VDD.t2147 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X819 a_9482_43914# a_9838_44484# VDD.t1651 VDD.t1650 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X820 a_20835_44721# a_20679_44626# a_20980_44850# VDD.t1646 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X821 VSS.t3499 a_5937_45572.t16 a_8781_46436# VSS.t3498 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 a_5837_42852# a_5891_43370.t15 VDD.t1804 VDD.t1803 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X823 a_10037_47542# a_n881_46662.t9 VSS.t1561 VSS.t1560 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X824 a_7221_43396# a_6031_43396# a_7112_43396# VSS.t2187 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X825 VSS.t3496 a_5937_45572.t12 a_8560_45348# VSS.t3495 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X826 C7_N_btm.t3 a_20820_30879.t4 VREF.t28 VDD.t1963 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X827 VSS.t992 a_15559_46634# a_13059_46348# VSS.t991 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X828 a_5385_46902# a_5167_46660# VSS.t996 VSS.t995 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X829 VDD.t266 a_10334_44484# a_10440_44484# VDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X830 a_19597_46482# a_19553_46090# a_19431_46494# VSS.t1861 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X831 VDD.t707 a_n2302_37984# a_n4209_38216.t2 VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 a_18051_46116# a_18189_46348# VDD.t1194 VDD.t1193 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X833 a_15493_43940# a_14955_43940# VSS.t1523 VSS.t1522 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X834 a_19250_34978# VDD.t3786 EN_VIN_BSTR_N.t0 VSS.t3212 sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X835 a_16414_43172# a_n1059_45260.t15 a_16328_43172# VSS.t2766 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X836 a_21297_46660# a_20107_46660# a_21188_46660# VSS.t1000 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X837 a_11813_46116# a_11387_46155# VDD.t1200 VDD.t1199 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X838 VSS.t1800 a_1666_39587.t3 a_1169_39587# VSS.t1799 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X839 VSS.t1704 SMPL_ON_P.t9 a_n1605_47204# VSS.t1703 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X840 DATA[4].t3 a_9067_47204# VDD.t1216 VDD.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X841 a_5894_47026# a_4817_46660# a_5732_46660# VDD.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X842 VDD.t1224 a_4699_43561# a_3539_42460# VDD.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X843 VSS.t2800 a_n3420_39072.t11 a_n2946_39072# VSS.t2641 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X844 VDD.t1900 a_n97_42460.t17 a_16245_42852# VDD.t1899 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X845 VDD.t644 a_13163_45724# a_11962_45724# VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X846 a_15433_44458# a_9482_43914# VSS.t1098 VSS.t1097 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X847 VDD.t3350 a_16327_47482.t33 a_20980_44850# VDD.t3349 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X848 a_18114_32519.t3 a_22223_45036# VSS.t1028 VSS.t1027 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X849 a_n452_44636# a_n1151_42308.t11 a_n310_44484# VSS.t1659 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X850 VDD.t2432 a_22959_43396# a_17364_32525.t1 VDD.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X851 a_n4064_37984.t3 a_n4334_38304# VDD.t2363 VDD.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X852 VDD.t3534 a_1307_43914.t27 a_4149_42891# VDD.t3533 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X853 VSS.t1835 a_n357_42282.t12 a_7573_43172# VSS.t1834 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X854 VDD.t1233 a_9863_47436# a_9804_47204# VDD.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X855 a_3754_39134# a_7754_38968# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X856 a_4649_43172# a_526_44458.t29 VSS.t3408 VSS.t3407 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X857 a_526_44458.t2 a_3147_46376# VDD.t2226 VDD.t2225 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X858 VSS.t1188 a_1848_45724# a_1799_45572# VSS.t1187 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X859 a_22485_38105# a_22775_42308# VSS.t1034 VSS.t1033 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X860 a_20885_45572# a_20841_45814# a_20719_45572# VSS.t1042 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X861 a_10554_47026# a_10428_46928# a_10150_46912# VSS.t2037 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X862 a_n746_45260# a_n1177_44458# VDD.t1176 VDD.t1175 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X863 a_7_44811# a_n1151_42308.t9 a_n452_44636# VDD.t1883 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X864 VDD.t3207 a_2324_44458.t35 a_15682_43940# VDD.t3206 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X865 VDD.t955 a_10355_46116# a_8199_44636# VDD.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X866 a_4181_43396# a_4093_43548# a_n2661_45546.t1 VSS.t1224 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X867 VDD.t3245 a_2437_43646.t3 a_22223_45572# VDD.t2086 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X868 a_21005_45260# a_21101_45002# VDD.t2430 VDD.t2429 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X869 VCM.t10 a_4190_30871.t13 C10_P_btm.t0 VSS.t2811 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X870 a_n3565_37414.t5 a_n2946_37690# VSS.t109 VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X871 a_3754_38802# a_7754_38968# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X872 a_2075_43172# a_1307_43914.t21 a_n913_45002.t9 VSS.t3463 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X873 VSS.t127 a_17499_43370# a_n1059_45260.t4 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X874 VSS.t2988 a_12861_44030.t27 a_17339_46660# VSS.t2987 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X875 VDD.t258 a_n2840_45002# a_n2810_45028.t1 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X876 a_10057_43914# a_10807_43548# VSS.t1054 VSS.t1053 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X877 a_5343_44458# a_7963_42308# VSS.t1056 VSS.t1055 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X878 a_n1423_42826# a_n1641_43230# VSS.t1062 VSS.t1061 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X879 a_526_44458.t5 a_3147_46376# VSS.t1967 VSS.t1966 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X880 VDD.t348 a_11827_44484# a_22223_45036# VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X881 VDD.t2216 a_n2472_43914# a_n3674_39768.t0 VDD.t2215 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X882 VDD.t602 a_15682_43940# a_11967_42832.t11 VDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X883 a_6945_45028.t1 a_5937_45572.t15 a_6945_45348# VSS.t3497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X884 VSS.t426 a_15682_43940# a_11967_42832.t30 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X885 a_20301_43646# a_13661_43548.t21 a_743_42282.t6 VDD.t3121 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X886 VDD.t1578 a_n3690_39616# a_n3420_39616.t2 VDD.t1577 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X887 a_n2216_39866# a_n2442_46660.t4 a_n2302_39866# VDD.t1876 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X888 VDD.t1266 a_22000_46634# a_15227_44166.t0 VDD.t1265 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X889 VSS.t1068 a_2889_44172# a_413_45260.t1 VSS.t1067 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X890 VSS.t1672 a_n97_42460.t11 a_n144_43396# VSS.t1671 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X891 a_n3674_38216.t1 a_n2104_42282# VDD.t312 VDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X892 a_16321_45348# a_1307_43914.t17 a_16019_45002# VSS.t3459 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X893 VSS.t843 a_6298_44484# a_4646_46812.t18 VSS.t842 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X894 VDD.t3275 a_9290_44172.t24 a_13070_42354# VDD.t3274 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X895 a_133_42852# a_n357_42282.t14 VDD.t2097 VDD.t2096 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X896 VSS.t3215 VDD.t3787 VSS.t3214 VSS.t3213 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X897 a_n3420_39072.t4 a_n3690_39392# VSS.t192 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X898 a_n2860_38778# a_n2956_38680.t4 a_n2946_38778# VDD.t1962 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X899 a_22485_38105# a_22775_42308# VDD.t1237 VDD.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X900 a_6517_45366# a_5937_45572.t9 a_6431_45366# VSS.t3494 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X901 a_10555_44260# a_10729_43914# VSS.t952 VSS.t951 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X902 VDD.t1096 a_5111_44636# a_5837_45028# VDD.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X903 a_14401_32519.t3 a_22223_43948# VSS.t1076 VSS.t1075 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X904 VSS.t3065 a_9290_44172.t18 a_13070_42354# VSS.t3064 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X905 VSS.t404 a_5068_46348# a_4955_46873# VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X906 VDD.t3273 a_9290_44172.t22 a_10586_45546# VDD.t3272 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X907 a_16751_45260# a_8696_44636.t5 VSS.t1712 VSS.t1711 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X908 a_1666_39587.t0 a_1666_39043.t5 VDD.t2945 VDD.t2944 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X909 a_n913_45002.t2 a_526_44458.t21 VDD.t3471 VDD.t3470 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X910 VSS.t2951 a_11599_46634.t38 a_15507_47210# VSS.t2950 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X911 VSS.t3609 a_768_44030.t15 a_644_44056# VSS.t3608 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X912 a_12465_44636# a_5807_45002# VDD.t1483 VDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X913 VDD.t2099 a_n357_42282.t15 a_16877_42852# VDD.t2098 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X914 a_5193_43172# a_3905_42865# VSS.t2050 VSS.t2049 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X915 VSS.t756 a_18783_43370# a_18525_43370# VSS.t755 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X916 a_3540_43646# a_1414_42308# a_3626_43646.t1 VDD.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X917 a_21363_45546# a_16327_47482.t45 VDD.t3362 VDD.t3361 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X918 VSS.t2276 a_n3690_38528# a_n3420_38528.t7 VSS.t1179 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X919 a_5421_42558# a_5379_42460# a_5337_42558# VDD.t2298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X920 VDD.t3185 a_12861_44030.t21 a_17609_46634# VDD.t3184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X921 a_n2956_38216.t3 a_n2472_45546# VSS.t2278 VSS.t968 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X922 a_13885_46660# a_13607_46688# VSS.t2280 VSS.t2279 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X923 VCM.t39 a_4958_30871.t13 C9_N_btm.t3 VSS.t2700 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X924 a_2232_45348# a_1609_45822# a_n2293_45546.t2 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X925 a_5691_45260# a_6171_45002.t2 a_5837_45028# VDD.t3606 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X926 a_9801_44260# a_3483_46348.t15 VSS.t3084 VSS.t3083 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X927 VCM.t0 a_3080_42308.t6 C2_N_btm.t0 VSS.t1539 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X928 a_327_44734# a_526_44458.t17 VDD.t3465 VDD.t3464 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X929 VSS.t331 a_7499_43078# a_8746_45002# VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X930 a_11967_42832.t23 a_15682_43940# VSS.t420 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X931 a_15743_43084# a_19339_43156# VDD.t2135 VDD.t2134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X932 VSS.t2287 a_22591_43396# a_14209_32519.t3 VSS.t2286 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X933 VSS.t3040 a_2437_43646.t4 a_22223_45572# VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X934 a_6547_43396# a_6197_43396# a_6452_43396# VDD.t2332 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X935 a_20556_43646# a_12549_44172.t18 VDD.t2940 VDD.t2939 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X936 a_1987_43646# a_742_44458# a_1891_43646# VDD.t978 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X937 a_4646_46812.t21 a_6298_44484# VSS.t845 VSS.t844 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X938 a_648_43396# a_584_46384.t18 VSS.t2783 VSS.t2782 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X939 VDD.t2537 a_n23_47502# a_7_47243# VDD.t2536 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X940 a_17609_46634# a_12549_44172.t24 VDD.t2949 VDD.t2948 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X941 a_3602_45348# a_3537_45260.t23 a_3495_45348# VSS.t2673 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X942 VDD.t3695 CLK.t1 a_8953_45002# VDD.t3694 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X943 VDD.t2032 a_2982_43646.t7 a_21487_43396# VDD.t2031 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X944 a_13661_43548.t0 a_18780_47178# VDD.t458 VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X945 VDD.t81 VSS.t3709 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X946 a_9313_44734.t1 a_3232_43370.t15 a_9159_44484# VSS.t2826 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X947 C6_P_btm.t4 a_5742_30871.t6 VCM.t26 VSS.t1844 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X948 a_11323_42473# a_5742_30871.t7 VSS.t1846 VSS.t1845 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X949 a_14383_46116# a_13759_46122# a_14275_46494# VDD.t1626 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X950 a_2813_43396# a_2479_44172# VSS.t1879 VSS.t1878 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X951 a_16721_46634# a_16388_46812# VSS.t479 VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X952 VSS.t312 a_8953_45002# a_2324_44458.t17 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X953 VDD.t3461 a_526_44458.t15 a_9885_43646# VDD.t3460 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X954 VSS.t2292 a_22537_40625# a_22737_36887# VSS.t2138 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X955 VREF.t29 a_20820_30879.t5 C7_N_btm.t2 VDD.t1964 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X956 VDD.t50 a_15681_43442# a_15781_43660# VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X957 a_6125_45348# a_3232_43370.t13 a_5691_45260# VSS.t2825 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X958 VSS.t3171 VDD.t3770 VSS.t3170 VSS.t3169 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X959 a_10907_45822# a_3483_46348.t19 VDD.t3297 VDD.t3296 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X960 a_14955_43396# a_9145_43396.t2 VDD.t1765 VDD.t1764 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X961 a_8128_46384# a_7903_47542# VDD.t2542 VDD.t2541 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X962 a_3429_45260# a_n971_45724.t17 VSS.t1691 VSS.t1690 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X963 VDD.t3674 a_15227_44166.t19 a_17969_45144# VDD.t3673 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X964 DATA[0].t1 a_327_47204# VDD.t2310 VDD.t2309 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X965 a_n2860_37690# a_n2956_37592.t4 a_n2946_37690# VDD.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X966 a_15682_46116# a_2324_44458.t61 VDD.t3171 VDD.t3170 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X967 VSS.t682 a_7287_43370# a_3537_45260.t5 VSS.t681 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X968 C4_P_btm.t3 a_n3420_38528.t8 VREF_GND.t24 VSS.t1775 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X969 a_18599_43230# a_18083_42858# a_18504_43218# VSS.t924 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X970 DATA[2].t4 a_4007_47204# VSS.t2143 VSS.t2142 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X971 a_18057_42282# a_18494_42460# a_18214_42558# VDD.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X972 a_11117_47542# a_4915_47217.t7 a_11031_47542# VSS.t3683 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X973 w_10694_33990.t15 a_18194_34908.t15 EN_VIN_BSTR_N.t6 w_10694_33990.t14 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X974 a_7112_43396# a_6197_43396# a_6765_43638# VSS.t2077 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X975 a_584_46384.t0 a_1123_46634# VDD.t1472 VDD.t1471 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X976 VSS.t2306 a_n3690_37440# a_n3420_37440.t7 VSS.t2305 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X977 VSS.t633 a_n901_43156# a_n443_42852.t4 VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X978 a_19240_46482# a_19123_46287# VDD.t1414 VDD.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X979 VCM.t27 a_5742_30871.t8 C6_N_btm.t5 VSS.t1554 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X980 VSS.t2796 a_10193_42453.t19 a_10149_42308# VSS.t2795 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X981 VDD.t3030 a_10193_42453.t23 a_10210_45822# VDD.t3029 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X982 VSS.t3015 a_2324_44458.t53 a_15682_46116# VSS.t3014 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X983 EN_VIN_BSTR_N.t1 VDD.t3825 a_19250_34978# VSS.t3154 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X984 VSS.t2308 a_n967_45348# a_n961_42308# VSS.t2307 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X985 a_564_42282# a_743_42282.t9 VDD.t3546 VDD.t3545 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X986 a_21195_42852# a_20922_43172# VDD.t2558 VDD.t2557 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X987 VDD.t2192 a_6575_47204# a_9067_47204# VDD.t2191 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X988 a_22612_30879.t0 a_22959_47212# VDD.t2562 VDD.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X989 a_21188_46660# a_20273_46660# a_20841_46902# VSS.t1151 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X990 a_13749_43396# a_13661_43548.t19 a_13667_43396# VSS.t2901 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X991 VSS.t2325 a_n2840_45546# a_n2810_45572.t3 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 a_13490_45394# a_9482_43914# VSS.t1088 VSS.t1087 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X993 a_n2840_43914# a_n2661_43922.t3 VDD.t1763 VDD.t1762 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X994 a_n822_43940# a_n1899_43946# a_n984_44318# VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X995 a_21613_42308# a_21335_42336# VSS.t2035 VSS.t2034 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X996 a_7112_43396# a_6031_43396# a_6765_43638# VDD.t2438 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X997 a_14537_43396# a_13059_46348# VSS.t1161 VSS.t1160 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X998 VDAC_Pi.t7 a_3754_38470.t5 a_4338_37500.t5 VSS.t2634 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X999 a_n4064_39616.t3 a_n4334_39616# VDD.t336 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1000 a_n23_47502# a_n971_45724.t23 VSS.t1698 VSS.t1697 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1001 a_n2438_43548.t18 a_949_44458# VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1002 a_14543_43071# a_5534_30871.t6 VDD.t3232 VDD.t2766 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1003 VSS.t886 a_15682_46116# a_11599_46634.t21 VSS.t885 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1004 VDD.t2304 a_19900_46494# a_20075_46420# VDD.t2303 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1005 VDD.t2574 a_7227_45028# a_7230_45938# VDD.t2573 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1006 VSS.t3371 a_16327_47482.t31 a_19597_46482# VSS.t3370 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1007 a_9823_46155# a_n743_46660.t7 a_9751_46155# VDD.t3641 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1008 VDD.t1168 a_22959_43948# a_17538_32519.t1 VDD.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1009 a_18214_42558# a_16137_43396# a_18057_42282# VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1010 a_n3690_38304# a_n3674_38216.t4 VDD.t2026 VDD.t2025 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1011 a_15009_46634# a_3090_45724.t13 VSS.t1595 VSS.t1594 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1012 a_17591_47464# a_10227_46804.t29 VDD.t1852 VDD.t1851 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1013 VSS.t1627 a_10227_46804.t33 a_15521_42308# VSS.t1626 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1014 VDD.t100 VSS.t3728 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1015 a_22485_44484# a_22315_44484# VSS.t1989 VSS.t1988 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1016 a_n1644_44306# a_n1761_44111# VDD.t2578 VDD.t2577 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1017 VDD.t1767 RST_Z.t0 a_8530_39574# VDD.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1018 VDD.t2499 a_n1329_42308# a_n1151_42308.t1 VDD.t2498 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1019 VSS.t1747 a_13507_46334.t11 a_18184_42460.t2 VSS.t1746 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1020 a_n630_44306# a_n1613_43370.t21 VSS.t3324 VSS.t3323 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1021 a_18783_43370# a_15743_43084# VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1022 a_n4064_38528.t7 a_n4334_38528# VSS.t1347 VSS.t1346 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1023 a_8325_42308# a_n913_45002.t21 a_8337_42558# VDD.t2963 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1024 VDD.t1754 CAL_P.t3 VDD.t1754 VDD.t1753 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X1025 a_21973_42336# a_20202_43084# a_21887_42336# VSS.t1324 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1026 VSS.t3340 a_n1613_43370.t35 a_645_46660# VSS.t3339 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1027 a_10341_42308# a_9803_42558# VDD.t2582 VDD.t2581 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1028 a_n1920_47178# a_n1741_47186.t8 VSS.t1848 VSS.t1847 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1029 VSS.t3360 a_16327_47482.t17 a_20885_45572# VSS.t3359 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1030 VSS.t1052 a_10807_43548# a_11173_44260# VSS.t1051 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1031 VSS.t1291 a_5257_43370# a_3905_42865# VSS.t1290 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1032 a_9127_43156# a_n1613_43370.t25 VDD.t3376 VDD.t3375 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1033 VDD.t1160 a_n2472_45002# a_n2956_37592.t0 VDD.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1034 VSS.t1896 a_n2946_39072# a_n3565_39304.t5 VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1035 a_13259_45724.t1 a_17583_46090# VDD.t2186 VDD.t2185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1036 VSS.t1078 a_10586_45546# a_10544_45572# VSS.t1077 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X1037 a_16751_45260# a_17023_45118# VSS.t2256 VSS.t2255 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1038 a_n2438_43548.t0 a_949_44458# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1039 VSS.t2680 a_n4209_38502.t10 a_n4251_38528# VSS.t2679 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1040 VSS.t730 a_7227_42308# a_6123_31319.t2 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1041 VSS.t740 a_10083_42826# a_7499_43078# VSS.t739 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 a_n2840_42826# a_n2661_42834.t3 VDD.t1982 VDD.t1981 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1043 a_1302_46660# a_n1613_43370.t33 VSS.t3336 VSS.t3335 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1044 a_5907_45546# a_6194_45824# VDD.t2586 VDD.t2585 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1045 a_13059_46348# a_15559_46634# VSS.t994 VSS.t993 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1046 a_n2302_37984# a_n2810_45572.t4 VSS.t1541 VSS.t1540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1047 VREF_GND.t23 a_14209_32519.t4 C5_N_btm.t3 VSS.t1774 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1048 a_3065_45002# a_3318_42354# a_3581_42558# VDD.t2587 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1049 a_16023_47582# a_15673_47210# a_15928_47570# VDD.t2244 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1050 VSS.t1563 a_n881_46662.t10 a_n935_46688# VSS.t1562 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1051 VDD.t149 VSS.t3713 VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1052 C6_N_btm.t0 EN_VIN_BSTR_N.t14 VIN_N.t14 VSS.t2920 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1053 VDD.t951 a_21487_43396# a_13467_32519.t0 VDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1054 a_2553_47502# a_n971_45724.t13 VSS.t1687 VSS.t1686 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1055 VDD.t3713 a_n443_42852.t17 a_997_45618# VDD.t3712 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1056 a_8568_45546# a_8199_44636# a_8791_45572# VSS.t778 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1057 a_4338_37500.t4 a_3754_38470.t6 VDAC_Pi.t6 VSS.t2635 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1058 a_13635_43156# a_10227_46804.t27 VDD.t1848 VDD.t1847 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1059 a_11967_42832.t10 a_15682_43940# VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1060 VDD.t984 a_564_42282# a_n1794_35082.t1 VDD.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1061 a_n473_42460# a_n971_45724.t21 a_n327_42308# VSS.t1696 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1062 a_16335_44484# a_13661_43548.t25 a_16241_44484# VSS.t2905 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1063 VDD.t1521 a_15861_45028# a_17023_45118# VDD.t1520 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1064 a_5205_44734# a_5111_44636# VDD.t1112 VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1065 a_7499_43078# a_10083_42826# VDD.t919 VDD.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1066 VSS.t1268 a_1123_46634# a_1057_46660# VSS.t1267 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1067 a_5700_37509.t3 VSS.t3711 VDAC_Pi.t3 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1068 a_n4064_37440.t4 a_n4334_37440# VSS.t1500 VSS.t1499 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1069 VSS.t67 a_13259_45724.t11 a_18315_45260# VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 a_22737_37285# a_22527_39145# a_22629_38406# VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1071 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS.t353 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1072 VSS.t1400 a_22400_42852# a_22848_40081# VSS.t1399 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1073 VSS.t1354 a_22223_43396# a_13887_32519.t2 VSS.t1233 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1074 a_11682_45822# a_11322_45546# a_11525_45546# VDD.t1579 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1075 VDD.t2287 a_22591_45572# a_19963_31679.t1 VDD.t2286 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1076 a_5934_30871.t2 a_8791_42308# VSS.t1203 VSS.t1202 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1077 a_18429_43548# a_18525_43370# VSS.t2272 VSS.t2271 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1078 a_509_45822# a_n1099_45572# VDD.t728 VDD.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1079 a_20980_44850# a_20766_44850# VDD.t2605 VDD.t2604 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1080 a_4190_30871.t0 a_19332_42282# VDD.t2180 VDD.t2179 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1081 a_3381_47502# a_2905_45572# VDD.t2607 VDD.t2606 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1082 VDD.t2908 a_3537_45260.t15 a_4649_42852# VDD.t2907 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1083 a_6682_46660# a_n971_45724.t15 VSS.t1689 VSS.t1688 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1084 a_20273_45572# a_20107_45572# VDD.t2474 VDD.t2473 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1085 VDD.t2613 a_11963_45334# a_11787_45002# VDD.t2612 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1086 VDD.t1974 a_1423_45028.t7 a_9838_44484# VDD.t1973 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1087 a_19256_45572# a_18175_45572# a_18909_45814# VDD.t2340 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1088 a_n755_45592.t0 a_n809_44244# VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1089 VSS.t870 a_3699_46634# a_3633_46660# VSS.t869 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1090 VSS.t3493 a_5937_45572.t7 a_9159_44484# VSS.t3492 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 a_14226_46987# a_14180_46812# VDD.t2621 VDD.t2620 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1092 VSS.t3672 a_n2438_43548.t36 a_n2157_46122# VSS.t3671 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1093 VSS.t2379 a_8953_45546# a_9241_46436# VSS.t2378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1094 a_n2840_45002# a_n2661_45010# VSS.t973 VSS.t972 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1095 a_n722_43218# a_n1613_43370.t47 VSS.t3346 VSS.t3345 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1096 a_12005_46436# a_2063_45854.t9 VSS.t1640 VSS.t1639 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1097 a_9885_43396# a_8270_45546# VSS.t578 VSS.t577 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1098 VSS.t3688 a_n4209_37414.t10 a_n4251_37440# VSS.t3687 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1099 VDD.t1576 a_n3690_39616# a_n3420_39616.t0 VDD.t1575 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1100 a_18817_42826# a_18599_43230# VDD.t2544 VDD.t2543 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1101 VDD.t384 a_167_45260# a_1423_45028.t0 VDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1102 VDAC_Pi.t0 VSS.t3717 a_5700_37509.t0 VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1103 VSS.t1138 a_4704_46090# a_1823_45246# VSS.t1137 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1104 a_16886_45144# a_8696_44636.t6 VDD.t1958 VDD.t1957 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X1105 a_11688_45572# a_11652_45724# VSS.t2382 VSS.t2381 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X1106 a_8953_45002# CLK.t2 VDD.t3697 VDD.t3696 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1107 VSS.t849 a_6298_44484# a_4646_46812.t29 VSS.t848 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1108 a_4520_42826# a_1823_45246# a_4743_43172# VSS.t246 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1109 a_949_44458# a_2324_44458.t57 VDD.t3227 VDD.t3226 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1110 a_n3420_39072.t7 a_n3690_39392# VSS.t196 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1111 VSS.t2027 a_22889_38993# a_22944_39857# VSS.t2026 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 VIN_P.t9 EN_VIN_BSTR_P.t16 a_n1057_35014.t2 VSS.t3568 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1113 VDD.t314 a_n2104_42282# a_n3674_38216.t0 VDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1114 VDD.t1769 RST_Z.t1 a_14311_47204# VDD.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1115 a_19721_31679.t3 a_22959_45036# VSS.t391 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1116 a_458_43396# a_526_44458.t13 VDD.t3459 VDD.t3458 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X1117 a_19339_43156# a_19164_43230# a_19518_43218# VSS.t1870 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1118 a_11453_44696.t0 a_17719_45144# VDD.t851 VDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1119 VDD.t2888 a_n3420_37984.t10 a_n2860_37984# VDD.t2887 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1120 a_13711_45394# a_12891_46348# a_13348_45260# VSS.t1431 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1121 a_16664_43396# a_16547_43609# VSS.t2072 VSS.t2071 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1122 a_1138_42852# a_791_42968# VSS.t408 VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1123 a_21259_43561# a_4190_30871.t9 VSS.t2807 VSS.t2806 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1124 a_10586_45546# a_9290_44172.t25 VDD.t3277 VDD.t3276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1125 VSS.t2949 a_11599_46634.t33 a_15599_45572# VSS.t2948 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1126 VSS.t2274 a_n3690_38528# a_n3420_38528.t6 VSS.t1183 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1127 a_11599_46634.t14 a_15682_46116# VDD.t1070 VDD.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1128 a_8912_37509.t5 VDAC_P.t18 a_5088_37509.t0 VDD.t69 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1129 a_196_42282# a_375_42282# VDD.t2204 VDD.t2203 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1130 VSS.t1567 a_n881_46662.t12 a_7989_47542# VSS.t1566 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1131 a_7832_46660# a_7715_46873# VSS.t2386 VSS.t2385 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1132 VDD.t2635 a_n2109_45247# en_comp VDD.t2634 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1133 VREF.t7 a_21588_30879.t7 C9_N_btm.t14 VDD.t1776 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1134 a_15928_47570# a_15811_47375# VSS.t987 VSS.t986 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1135 a_3633_46660# a_2443_46660# a_3524_46660# VSS.t2540 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1136 VSS.t2277 a_n2472_45546# a_n2956_38216.t2 VSS.t966 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1137 a_2127_44172# a_2675_43914# VSS.t2545 VSS.t2544 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1138 a_9885_43646# a_5111_44636# VDD.t1110 VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1139 a_n2472_43914# a_n2293_43922.t3 VDD.t3052 VDD.t3051 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1140 VDD.t2803 a_12991_46634# a_12978_47026# VDD.t2802 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1141 VDD.t681 a_1667_45002# a_n863_45724# VDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1142 a_n4209_39304.t4 a_n2302_39072# VSS.t227 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1143 a_14084_46812# a_n1151_42308.t6 a_14226_46987# VDD.t1881 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1144 a_5837_45028# a_3232_43370.t11 a_5691_45260# VDD.t3044 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X1145 a_21753_35474# a_19998_34978# VDD.t1657 VDD.t1656 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1146 VDD.t2560 a_21195_42852# a_21671_42860# VDD.t2559 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1147 C10_N_btm.t19 a_22612_30879.t15 VREF.t23 VDD.t1950 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1148 a_12427_45724# a_12791_45546# a_12749_45572# VSS.t1515 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1149 VSS.t2733 a_n913_45002.t19 a_4921_42308# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1150 a_14209_32519.t2 a_22591_43396# VSS.t2285 VSS.t2284 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1151 a_4646_46812.t30 a_6298_44484# VSS.t837 VSS.t836 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1152 a_12553_44484# a_12465_44636# a_n2661_43922.t1 VSS.t1082 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1153 C9_N_btm.t13 a_21588_30879.t9 VREF.t9 VDD.t1778 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1154 a_5829_43940# a_1307_43914.t15 VDD.t3525 VDD.t3524 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1155 a_16237_45028# a_n743_46660.t9 VDD.t3644 VDD.t3643 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1156 VDD.t578 a_22959_45036# a_19721_31679.t1 VDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1157 a_14761_44260# a_14673_44172# a_n2293_46634.t1 VSS.t1191 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 VSS.t3316 a_n1613_43370.t17 a_5429_46660# VSS.t3315 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1159 CAL_P.t0 a_22485_38105# VDD.t1243 VDD.t1242 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1160 VSS.t1300 a_21363_46634# a_21297_46660# VSS.t1299 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1161 VDD.t2811 a_n452_45724# a_n1853_46287# VDD.t2810 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1162 VDD.t3010 a_584_46384.t22 a_2998_44172# VDD.t3009 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 VSS.t1023 a_4699_43561# a_3539_42460# VSS.t1022 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1164 VDD.t2813 a_15959_42545# a_15890_42674# VDD.t2812 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1165 VSS.t1615 a_10227_46804.t19 a_13157_43218# VSS.t1614 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1166 a_n4209_38502.t1 a_n2302_38778# VDD.t2650 VDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1167 VSS.t539 a_n2946_39866# a_n3565_39590.t5 VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1168 a_11599_46634.t25 a_15682_46116# VSS.t884 VSS.t883 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1169 a_17538_32519.t3 a_22959_43948# VSS.t976 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1170 a_n144_43396# a_n971_45724.t11 a_n447_43370# VSS.t1685 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1171 a_16680_45572# a_15599_45572# a_16333_45814# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1172 VSS.t3491 a_5937_45572.t5 a_6101_44260# VSS.t3490 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1173 a_9672_43914# a_8199_44636# a_9895_44260# VSS.t785 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1174 a_15231_43396# a_9145_43396.t3 a_15125_43396# VSS.t1550 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1175 a_8387_43230# a_7871_42858# a_8292_43218# VSS.t1468 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1176 VDD.t675 a_22731_47423# a_13717_47436.t0 VDD.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1177 VDD.t3281 a_9290_44172.t29 a_13667_43396# VDD.t3280 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1178 a_n3420_37984.t0 a_n3690_38304# VDD.t1380 VDD.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1179 VDD.t3319 a_10903_43370.t18 a_13163_45724# VDD.t3318 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X1180 VDD.t986 a_17767_44458# a_17715_44484# VDD.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1181 VDD.t2821 a_7845_44172# a_7542_44172# VDD.t2820 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X1182 a_n2840_44458# a_n2661_44458.t3 VDD.t3709 VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1183 a_22400_42852# a_22223_42860# VDD.t1440 VDD.t1439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1184 VDD.t693 a_n863_45724# a_945_42968# VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1185 VSS.t1090 a_9482_43914# a_10157_44484# VSS.t1089 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1186 VDD.t2936 a_12549_44172.t14 a_10949_43914# VDD.t2935 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X1187 a_4933_42558# a_4791_45118.t11 VDD.t2012 VDD.t2011 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1188 a_19333_46634# a_19466_46812# VSS.t691 VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1189 a_13565_44260# a_12891_46348# VSS.t1433 VSS.t1432 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 VSS.t2304 a_n3690_37440# a_n3420_37440.t6 VSS.t2303 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1191 a_2324_44458.t12 a_8953_45002# VDD.t504 VDD.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1192 a_n2293_46098.t1 a_5663_43940# VSS.t2563 VSS.t2562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1193 EN_VIN_BSTR_P.t2 VDD.t3824 a_n217_35014# VSS.t3153 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1194 VSS.t3634 a_11453_44696.t3 a_22959_47212# VSS.t3633 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1195 VSS.t269 a_12563_42308# a_5534_30871.t3 VSS.t268 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1196 a_n2472_42826# a_n2293_42834.t3 VDD.t1986 VDD.t1985 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1197 a_7920_46348# a_8128_46384# a_8062_46482# VSS.t658 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1198 a_5088_37509.t1 VDAC_P.t14 a_8912_37509.t6 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1199 a_n13_43084# a_n443_42852.t15 a_133_42852# VDD.t3711 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1200 a_2698_46116# a_2521_46116# VDD.t2827 VDD.t2826 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1201 a_15785_43172# a_15743_43084# a_15095_43370# VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1202 a_8654_47026# a_7577_46660# a_8492_46660# VDD.t1716 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 VDD.t1512 a_21363_46634# a_21350_47026# VDD.t1511 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1204 a_n2438_43548.t17 a_949_44458# VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1205 VDD.t548 a_n809_44244# a_n822_43940# VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1206 a_766_43646# a_626_44172# a_458_43396# VDD.t1036 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X1207 a_n784_42308.t1 a_n961_42308# VDD.t2556 VDD.t2555 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1208 a_12895_43230# a_12379_42858# a_12800_43218# VSS.t1460 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1209 VSS.t1221 a_805_46414# a_739_46482# VSS.t1220 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1210 VSS.t2573 a_8191_45002# a_8137_45348# VSS.t2572 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1211 a_15959_42545# a_15803_42450# a_16104_42674# VDD.t2508 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1212 a_5210_46482# a_5164_46348# VSS.t188 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1213 a_11341_43940.t1 a_3232_43370.t9 a_11173_44260# VSS.t2822 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1214 VDD.t2833 a_7705_45326# a_7735_45067# VDD.t2832 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1215 a_13720_44458# a_13661_43548.t11 a_13940_44484# VSS.t2894 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1216 a_2162_46660# a_2107_46812.t2 VSS.t2820 VSS.t2819 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1217 VSS.t598 a_n4334_39392# a_n4064_39072.t5 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1218 a_n1423_42826# a_n1641_43230# VDD.t1264 VDD.t1263 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1219 a_n2956_39304.t2 a_n2840_46090# VSS.t1207 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1220 VDD.t2835 a_11415_45002# a_n2661_43370.t1 VDD.t2834 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1221 a_15037_43940# a_15227_44166.t25 VDD.t3678 VDD.t3677 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1222 VDD.t1980 a_1606_42308.t4 a_2351_42308# VDD.t1979 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1223 a_2277_45546# a_167_45260# VDD.t376 VDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1224 VCM.t52 a_3422_30871.t13 VDAC_N.t1 VSS.t3515 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1225 a_6903_46660# a_6755_46942# a_6540_46812# VSS.t2585 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1226 VDD.t2850 a_14180_45002# a_13017_45260# VDD.t2849 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1227 a_3232_43370.t3 a_1823_45246# VDD.t436 VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1228 VDD.t1375 a_n2302_40160# a_n4315_30879.t2 VDD.t1046 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1229 VDD.t957 a_8199_44636# a_8191_45002# VDD.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1230 a_n4209_37414.t0 a_n2302_37690# VDD.t1152 VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1231 a_1576_42282# a_1755_42282# VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1232 a_7573_43172# a_7499_43078# a_7227_42852# VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1233 VSS.t1883 a_21855_43396# a_13678_32519.t3 VSS.t1882 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1234 VDD.t294 a_18989_43940# a_19006_44850# VDD.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1235 VSS.t2587 a_6540_46812# a_6491_46660# VSS.t2586 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 VSS.t3110 VDD.t3809 VSS.t3109 VSS.t3108 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1237 VDD.t1434 a_22223_45572# a_19479_31679.t0 VDD.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1238 VIN_N.t6 EN_VIN_BSTR_N.t17 C0_dummy_N_btm.t0 VSS.t2923 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1239 VSS.t50 a_2903_42308# a_3080_42308.t3 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1240 VSS.t510 a_n863_45724# a_n906_45572# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1241 a_n2840_44458# a_n2661_44458.t4 VSS.t3640 VSS.t1542 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1242 a_22629_37990# a_22581_37893# CAL_P.t2 VDD.t3480 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1243 a_3823_42558# a_3065_45002# a_3905_42558# VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1244 VSS.t489 a_2779_44458# a_1307_43914.t7 VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1245 VSS.t940 a_5263_45724# a_5204_45822# VSS.t939 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1246 VDD.t1714 a_2124_47436# a_1209_47178# VDD.t1713 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1247 a_12925_46660# a_11735_46660# a_12816_46660# VSS.t455 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1248 VSS.t3420 a_2957_45546# a_2905_45572# VSS.t3419 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1249 a_376_46348# a_n743_46660.t4 a_518_46155# VDD.t3640 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1250 a_11415_45002# a_4915_47217.t9 a_14581_44484# VSS.t3686 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1251 VDD.t3594 a_7754_40130.t11 VDD.t3593 VDD.t3592 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X1252 a_n2104_42282# a_n1925_42282.t4 VDD.t3054 VDD.t3053 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1253 a_n2472_45002# a_n2293_45010# VSS.t3421 VSS.t1772 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1254 a_21398_44850# a_20679_44626# a_20835_44721# VSS.t1441 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1255 VDD.t2817 a_16333_45814# a_16223_45938# VDD.t2816 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1256 a_16241_44484# a_2711_45572.t6 VSS.t3656 VSS.t3655 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1257 a_3905_42865# a_5257_43370# VSS.t1296 VSS.t1295 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1258 VSS.t2607 a_8685_43396.t2 a_15231_43396# VSS.t2606 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1259 VSS.t382 a_10623_46897# a_10554_47026# VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1260 a_13485_45572# a_12549_44172.t22 a_13385_45572# VSS.t2716 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1261 C3_P_btm.t0 a_n4209_38216.t10 VREF.t62 VDD.t3096 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1262 VSS.t291 a_22959_45572# a_20447_31679.t3 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1263 a_22848_39857# a_22485_38105# a_22581_37893# VSS.t1041 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1264 VDD.t406 a_19987_42826# a_n2017_45002.t0 VDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X1265 a_9028_43914# a_9482_43914# a_9420_43940# VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1266 VSS.t1130 a_17973_43940# a_18079_43940# VSS.t1129 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1267 a_n2860_39072# a_n2956_39304.t5 a_n2946_39072# VDD.t1962 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1268 a_9290_44172.t4 a_13635_43156# VSS.t2358 VSS.t2357 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1269 a_3059_42968# a_742_44458# a_2987_42968# VDD.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1270 a_n452_44636# a_n467_45028# a_n310_44811# VDD.t2264 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1271 VREF.t10 a_21588_30879.t10 C9_N_btm.t15 VDD.t1779 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1272 VDD.t3685 a_768_44030.t13 a_2711_45572.t0 VDD.t3684 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1273 a_11967_42832.t9 a_15682_43940# VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1274 VDD.t450 a_12281_43396# a_12563_42308# VDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1275 VDD.t1978 a_12741_44636.t4 a_22959_46660# VDD.t1977 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1276 a_8333_44734# a_3537_45260.t26 a_8238_44734# VDD.t2913 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1277 VDD.t36 a_949_44458# a_n2438_43548.t11 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1278 a_17124_42282# a_17303_42282# VDD.t556 VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1279 a_12156_46660# a_11813_46116# VSS.t1006 VSS.t1005 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1280 VDD.t3646 a_10809_44734.t4 a_22959_46124# VDD.t3099 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1281 VSS.t2244 a_1115_44172# a_n2293_45010# VSS.t2243 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1282 a_5013_44260# a_1307_43914.t11 VSS.t3486 VSS.t3485 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1283 VDD.t2643 a_n447_43370# a_n2129_43609# VDD.t2642 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1284 a_3357_43084.t1 a_5257_43370# a_5565_43396# VSS.t1292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1285 a_1568_43370# a_1847_42826# a_1793_42852# VDD.t2500 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1286 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS.t1125 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1287 a_11682_45822# a_10586_45546# VDD.t1280 VDD.t1279 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1288 a_18315_45260# a_15227_44166.t11 VSS.t3593 VSS.t3592 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1289 a_n2012_44484# a_n2129_44697# VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1290 a_14543_43071# a_5534_30871.t7 VSS.t3028 VSS.t3027 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1291 a_16147_45260# a_17478_45572# VDD.t1347 VDD.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1292 a_22848_40081# en_comp a_22589_40055# VSS.t1041 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 a_19963_31679.t0 a_22591_45572# VDD.t2285 VDD.t2284 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1294 a_n967_45348# a_n1059_45260.t11 VSS.t2762 VSS.t2761 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1295 VDD.t1064 a_15682_46116# a_11599_46634.t5 VDD.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1296 VDD.t3165 a_11599_46634.t47 a_20107_45572# VDD.t3164 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1297 VSS.t3427 a_7276_45260# a_7227_45028# VSS.t3426 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1298 a_1241_44260# a_584_46384.t12 VSS.t2777 VSS.t2776 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1299 VDD.t554 a_n809_44244# a_n755_45592.t2 VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1300 VSS.t3431 a_n815_47178# a_n785_47204# VSS.t3430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1301 a_n4334_40480# a_n4318_40392.t4 VDD.t2106 VDD.t1889 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1302 a_3175_45822# a_3090_45724.t11 a_2957_45546# VDD.t1817 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1303 a_14621_43646# a_14579_43548# a_14537_43646# VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1304 VDD.t1616 a_n2946_37984# a_n3565_38216.t2 VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1305 VREF.t51 a_20205_31679.t4 C4_N_btm.t3 VDD.t2893 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1306 VSS.t3601 a_15227_44166.t22 a_18900_46660# VSS.t3600 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1307 a_n310_44811# a_n356_44636.t2 VDD.t3653 VDD.t3652 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1308 VDD.t2645 a_16977_43638# a_16867_43762# VDD.t2644 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1309 VDD.t3660 a_15227_44166.t7 a_17749_42852# VDD.t3659 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1310 a_3147_46376# a_3483_46348.t23 VSS.t3090 VSS.t3089 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1311 a_12638_46436# a_12594_46348# a_12379_46436# VSS.t3435 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1312 a_n2438_43548.t8 a_949_44458# VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1313 VSS.t3013 a_2324_44458.t52 a_6298_44484# VSS.t3012 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1314 a_2324_44458.t13 a_8953_45002# VDD.t484 VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1315 VSS.t831 a_6298_44484# a_4646_46812.t16 VSS.t830 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1316 a_21071_46482# a_15227_44166.t6 a_20708_46348# VSS.t3587 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1317 a_n1059_45260.t5 a_17499_43370# VSS.t125 VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1318 VDD.t2057 a_1273_38525.t10 a_2684_37794# VDD.t2056 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1319 a_961_42354# a_n1059_45260.t18 VDD.t2991 VDD.t2990 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1320 a_9127_43156# a_8952_43230# a_9306_43218# VSS.t965 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1321 VSS.t1726 a_12741_44636.t5 a_22959_46660# VSS.t1725 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1322 VSS.t948 a_8349_46414# a_8283_46482# VSS.t947 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1323 VSS.t2370 a_11787_45002# a_11652_45724# VSS.t2369 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1324 a_4223_44672.t2 a_3537_45260.t11 VSS.t2666 VSS.t2665 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1325 a_509_45822# a_n357_42282.t9 VDD.t2091 VDD.t2090 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1326 a_16119_47582# a_15673_47210# a_16023_47582# VSS.t1991 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1327 a_6452_43396# a_6293_42852# VSS.t1284 VSS.t1283 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1328 VSS.t3627 CLK.t3 a_8953_45002# VSS.t3626 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 a_6194_45824# a_6472_45840# a_6428_45938# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1330 a_3754_38802# a_7754_38636# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X1331 a_11599_46634.t15 a_15682_46116# VDD.t1074 VDD.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1332 C9_P_btm.t9 a_n4209_39590.t17 VREF.t61 VDD.t3080 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1333 VDD.t1790 a_n881_46662.t16 a_11031_47542# VDD.t1789 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1334 VSS.t2102 a_1209_47178# a_1239_47204# VSS.t2101 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1335 a_15559_46634# a_13507_46334.t5 VDD.t1996 VDD.t1995 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1336 a_12429_44172# a_12861_44030.t17 VDD.t3183 VDD.t3182 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1337 VDAC_N.t3 a_3422_30871.t11 VCM.t50 VSS.t3513 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1338 a_11229_43218# a_10227_46804.t25 VSS.t1623 VSS.t1622 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1339 a_16020_45572# a_15903_45785# VSS.t3437 VSS.t3436 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1340 C3_P_btm.t3 a_5932_42308.t6 VCM.t21 VSS.t1803 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1341 a_10149_42308# a_9290_44172.t9 a_9803_42558# VSS.t3057 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1342 VSS.t2238 a_20708_46348# a_20411_46873# VSS.t2237 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1343 VDD.t229 VSS.t3727 VDD.t228 VDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1344 C9_N_btm.t2 a_4958_30871.t4 VCM.t32 VSS.t2691 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1345 a_10793_43218# a_10083_42826# VSS.t734 VSS.t733 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1346 a_n863_45724# a_1667_45002# VDD.t679 VDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1347 a_13635_43156# a_13460_43230# a_13814_43218# VSS.t1462 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1348 a_12379_46436# a_12594_46348# a_12638_46436# VSS.t3434 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1349 VREF.t41 a_n4315_30879.t15 C10_P_btm.t23 VDD.t2075 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1350 VDD.t494 a_8953_45002# a_2324_44458.t8 VDD.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1351 a_1209_43370# a_1049_43396# VSS.t3439 VSS.t3438 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1352 a_2982_43646.t3 a_3232_43370.t18 a_2813_43396# VSS.t2829 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1353 a_n443_46116.t3 a_n901_46420# VDD.t2460 VDD.t2459 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1354 a_21542_45572# a_16327_47482.t15 VSS.t3358 VSS.t3357 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1355 VSS.t89 a_19647_42308# a_13258_32519.t2 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1356 a_18985_46122# a_18819_46122# VDD.t2462 VDD.t2461 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1357 VSS.t2853 a_n1794_35082.t14 a_18194_34908.t7 VSS.t2852 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1358 a_12839_46116# a_13059_46348# VDD.t1367 VDD.t1366 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1359 VDD.t3740 a_n2438_43548.t34 a_2443_46660# VDD.t3739 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1360 VDD.t3491 a_9028_43914# a_8975_43940# VDD.t3490 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1361 VDD.t558 a_17124_42282# a_4958_30871.t1 VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1362 VSS.t934 a_10053_45546# a_9625_46129# VSS.t933 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X1363 a_17639_46660# a_17609_46634# a_765_45546.t5 VSS.t1998 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1364 VSS.t3441 a_380_45546# a_n356_45724# VSS.t3440 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1365 VSS.t3447 a_20193_45348# a_21973_42336# VSS.t3446 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1366 VSS.t593 a_196_42282# a_n3674_37592.t3 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1367 VDD.t1506 a_5257_43370# a_5826_44734# VDD.t1505 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X1368 a_9803_42558# a_n97_42460.t9 a_9885_42308# VSS.t1670 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1369 a_11599_46634.t16 a_15682_46116# VSS.t876 VSS.t875 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1370 VSS.t1611 a_10227_46804.t15 a_10553_43218# VSS.t1610 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1371 VSS.t1199 a_18597_46090# a_16375_45002# VSS.t1198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1372 VSS.t2735 a_n913_45002.t20 a_12281_43396# VSS.t2734 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1373 a_12816_46660# a_11901_46660# a_12469_46902# VSS.t1240 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1374 a_n3565_39590.t7 a_n2946_39866# VSS.t537 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1375 a_20205_45028# a_18184_42460.t6 VDD.t3734 VDD.t3733 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1376 a_n3420_37984.t3 a_n3690_38304# VDD.t1384 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1377 VDD.t254 a_13259_45724.t9 a_13667_43396# VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1378 a_n1736_42282# a_n1557_42282# VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1379 a_13747_46662.t0 a_19386_47436# VDD.t1546 VDD.t1545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1380 VSS.t1755 a_4791_45118.t9 a_6165_46155# VSS.t1754 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X1381 a_261_44278# a_n863_45724# a_175_44278# VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1382 a_2324_44458.t3 a_8953_45002# VDD.t492 VDD.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1383 a_8325_42308# a_5891_43370.t13 VSS.t1655 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1384 a_10623_46897# a_10467_46802# a_10768_47026# VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1385 a_17957_46116# a_765_45546.t10 VSS.t3693 VSS.t3692 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1386 a_2675_43914# a_2998_44172# VSS.t1105 VSS.t1104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 a_18695_43230# a_18249_42858# a_18599_43230# VSS.t925 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1388 a_17613_45144# a_8696_44636.t2 VSS.t1709 VSS.t1708 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1389 a_n4318_39304.t0 a_n2840_43370# VDD.t288 VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1390 a_18799_45938# a_16327_47482.t16 VDD.t3411 VDD.t3410 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1391 VSS.t531 a_19862_44208# a_20922_43172# VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1392 a_6151_47436.t1 a_14311_47204# VSS.t233 VSS.t232 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1393 a_5700_37509.t14 VDAC_N.t13 a_8912_37509.t21 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1394 VSS.t1893 a_5129_47502# a_5063_47570# VSS.t1892 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1395 VSS.t211 a_167_45260# a_2521_46116# VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1396 a_3733_45822# a_n755_45592.t14 a_3638_45822# VDD.t3443 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1397 a_16333_45814# a_16115_45572# VSS.t352 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1398 VDD.t187 VSS.t3721 VDD.t186 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1399 a_1337_46116# a_1176_45822# VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1400 a_13163_45724# a_13527_45546# a_13485_45572# VSS.t1532 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1401 a_8605_42826# a_8387_43230# VDD.t2247 VDD.t2246 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1402 VDD.t2389 a_4419_46090# a_n1925_42282.t2 VDD.t2388 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1403 a_n4209_38216.t0 a_n2302_37984# VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1404 a_20712_42282# a_n357_42282.t7 VSS.t1831 VSS.t1830 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1405 VSS.t3125 VDD.t3814 VSS.t3124 VSS.t3123 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1406 a_1241_43940# a_1467_44172# a_1443_43940# VDD.t3523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1407 a_9145_43396.t0 a_8791_43396# VDD.t2440 VDD.t2439 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1408 VDD.t2554 a_n961_42308# a_n784_42308.t0 VDD.t2553 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1409 a_7227_42852# a_n97_42460.t10 a_7309_42852# VDD.t1898 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1410 a_14976_45348# a_13059_46348# VSS.t1159 VSS.t1158 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1411 a_9863_47436# a_n881_46662.t22 VDD.t1800 VDD.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1412 a_743_42282.t2 a_19692_46634.t5 VSS.t1812 VSS.t1811 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1413 a_4915_47217.t0 a_12991_46634# VDD.t2805 VDD.t2804 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1414 VSS.t1430 a_12891_46348# a_12638_46436# VSS.t1429 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1415 a_n3674_38680.t2 a_n2840_42282# VSS.t744 VSS.t743 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1416 VCM.t38 a_4958_30871.t12 C9_N_btm.t0 VSS.t2699 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1417 VSS.t742 a_3539_42460# a_3065_45002# VSS.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 a_17801_45144# a_17613_45144# a_17719_45144# VDD.t3522 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1419 VDD.t3077 a_n4209_39590.t14 a_n4334_39616# VDD.t2078 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1420 a_18787_45572# a_18341_45572# a_18691_45572# VSS.t2090 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1421 a_10922_42852# a_10796_42968# a_10518_42984# VSS.t3270 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1422 VSS.t3206 VDD.t3782 VSS.t3205 VSS.t3135 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1423 a_3754_39964# a_7754_40130.t3 VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X1424 VDD.t2318 a_n4334_40480# a_n4064_40160.t2 VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1425 VDD.t3457 a_526_44458.t11 a_3232_43370.t0 VDD.t3456 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1426 a_n1794_35082.t3 a_564_42282# VSS.t797 VSS.t796 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1427 a_167_45260# a_2202_46116# VSS.t1178 VSS.t1177 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1428 VDD.t3137 a_11967_42832.t33 a_20512_43084# VDD.t3136 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1429 VDD.t56 a_16019_45002# a_15903_45785# VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1430 a_2896_43646# a_n443_46116.t18 VDD.t3254 VDD.t3253 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1431 VSS.t1018 a_9067_47204# DATA[4].t6 VSS.t1017 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1432 a_n2312_38680.t1 a_n2104_46634# VDD.t3331 VDD.t3330 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1433 a_12005_46116# a_10903_43370.t23 a_12005_46436# VSS.t3104 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1434 a_n2288_47178# a_n2109_47186.t2 VSS.t3579 VSS.t3578 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1435 VREF.t19 a_22612_30879.t11 C10_N_btm.t15 VDD.t1946 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1436 a_14097_32519.t1 a_22959_42860# VDD.t3333 VDD.t3332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1437 a_6999_46987# a_3877_44458# a_6540_46812# VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1438 a_8199_44636# a_10355_46116# VDD.t953 VDD.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1439 a_3429_45260# a_n971_45724.t9 VDD.t1912 VDD.t1911 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1440 C8_N_btm.t8 EN_VIN_BSTR_N.t7 VIN_N.t1 VSS.t2914 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1441 a_4338_37500.t1 VSS.t58 VSS.t60 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X1442 a_9293_42558# a_9223_42460# a_8953_45546# VDD.t3336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1443 VDD.t1548 a_n452_47436# a_n815_47178# VDD.t1547 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1444 VDD.t1373 a_n2302_40160# a_n4315_30879.t3 VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 a_14309_45348# a_2711_45572.t9 VSS.t3658 VSS.t3657 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1446 a_13807_45067# a_13556_45296# a_13348_45260# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1447 a_2981_46116# a_2804_46116# VDD.t3338 VDD.t3337 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1448 a_1176_45822# a_997_45618# a_1260_45572# VSS.t2346 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X1449 a_4185_45028.t1 a_3877_44458# a_4185_45348# VSS.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 VDD.t2232 a_13159_45002# a_n2661_46634.t2 VDD.t2231 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1451 VSS.t3284 a_20269_44172# a_19319_43548# VSS.t3283 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1452 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS.t1250 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1453 a_16104_42674# a_15890_42674# VDD.t2815 VDD.t2814 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1454 a_5700_37509.t13 VDAC_N.t11 a_8912_37509.t19 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1455 a_22731_47423# SMPL_ON_N.t9 VSS.t3504 VSS.t3503 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1456 a_n722_46482# a_n1613_43370.t20 VSS.t3322 VSS.t3321 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1457 VSS.t3643 a_n443_42852.t13 a_997_45618# VSS.t3642 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1458 a_6945_45348# a_5205_44484# VSS.t3286 VSS.t3285 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1459 a_21513_45002# a_21363_45546# VSS.t1528 VSS.t1527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1460 a_4791_45118.t1 a_4743_44484# VDD.t1313 VDD.t1312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1461 VSS.t99 a_1576_42282# a_1606_42308.t3 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1462 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD.t1588 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1463 a_15227_44166.t1 a_22000_46634# VDD.t1268 VDD.t1267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1464 a_n743_46660.t0 a_n1021_46688# VDD.t638 VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1465 a_n4064_40160.t3 a_n4334_40480# VDD.t2317 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1466 a_2075_43172# a_1307_43914.t10 a_n913_45002.t8 VSS.t3484 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1467 VSS.t3288 a_5205_44484# a_6756_44260# VSS.t3287 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1468 VDD.t2531 a_327_44734# a_375_42282# VDD.t2530 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1469 VDD.t1544 a_19321_45002# a_3090_45724.t1 VDD.t1543 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1470 VSS.t3086 a_3483_46348.t17 a_13829_44260# VSS.t3085 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1471 VDD.t3585 a_7754_40130.t7 a_11206_38545.t2 VDD.t3584 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1472 VDD.t26 a_949_44458# a_n2438_43548.t2 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1473 VDD.t3567 a_5937_45572.t11 a_6671_43940# VDD.t3566 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1474 VDD.t685 a_n863_45724# a_458_43396# VDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1475 VDD.t2362 a_n4334_38304# a_n4064_37984.t0 VDD.t1711 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1476 VDD.t3455 a_526_44458.t10 a_n913_45002.t3 VDD.t3454 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1477 VDD.t2166 a_1756_43548# a_1467_44172# VDD.t2165 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X1478 VDD.t2014 a_4791_45118.t12 a_5066_45546# VDD.t2013 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1479 VDD.t38 a_949_44458# a_n2438_43548.t15 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1480 a_20269_44172# a_20365_43914# VDD.t2668 VDD.t2667 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1481 VDD.t2670 a_14976_45028# a_15227_46910# VDD.t2669 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1482 VSS.t2042 a_13904_45546# a_12594_46348# VSS.t2041 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1483 VREF_GND.t13 a_18114_32519.t7 C10_N_btm.t27 VSS.t2650 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1484 VSS.t2376 a_8953_45546# a_8568_45546# VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1485 VDAC_Pi.t5 a_3754_38470.t7 a_4338_37500.t3 VSS.t2636 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1486 a_16112_44458# a_15227_44166.t4 a_16335_44484# VSS.t3586 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1487 VSS.t3350 a_16327_47482.t8 a_17021_43396# VSS.t3349 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1488 a_n913_45002.t4 a_1307_43914.t20 VDD.t3527 VDD.t3526 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1489 VSS.t450 a_20974_43370# a_20749_43396# VSS.t449 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1490 a_16388_46812# a_17957_46116# VDD.t3521 VDD.t3520 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1491 VSS.t2421 a_20159_44458# a_19321_45002# VSS.t2420 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1492 VDD.t296 a_9672_43914# a_2107_46812.t0 VDD.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1493 VSS.t2139 a_22589_40599# a_22737_37285# VSS.t2138 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1494 a_n4318_37592.t0 a_n1736_42282# VDD.t899 VDD.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1495 VSS.t2756 a_6151_47436.t11 a_8189_46660# VSS.t2755 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1496 VDD.t2938 a_12549_44172.t15 a_17609_46634# VDD.t2937 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1497 a_6229_45572# a_6194_45824# a_5907_45546# VSS.t2343 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1498 VDD.t745 a_19700_43370# a_n97_42460.t1 VDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1499 a_6851_47204# a_6491_46660# VDD.t2239 VDD.t2238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1500 VDD.t2676 a_19615_44636# a_18579_44172# VDD.t2675 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1501 a_8423_43396# a_n443_42852.t11 a_8317_43396# VSS.t3641 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1502 VDD.t517 a_7499_43078# a_8697_45822# VDD.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1503 a_18799_45938# a_18175_45572# a_18691_45572# VDD.t2343 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1504 a_1755_42282# a_n913_45002.t18 VSS.t2732 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 a_n1741_47186.t5 a_12005_46116# a_12379_46436# VSS.t2114 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X1506 VSS.t3001 a_2324_44458.t38 a_6298_44484# VSS.t3000 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1507 VDD.t1607 a_6765_43638# a_6655_43762# VDD.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1508 a_5700_37509.t12 VDAC_N.t10 a_8912_37509.t18 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1509 a_n4209_39304.t3 a_n2302_39072# VDD.t400 VDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1510 VDD.t2268 a_22223_47212# a_21588_30879.t0 VDD.t2267 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1511 a_n2438_43548.t4 a_949_44458# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1512 a_685_42968# a_n443_42852.t18 VDD.t3715 VDD.t3714 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1513 a_10467_46802# a_11599_46634.t44 VSS.t2959 VSS.t2958 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1514 VDD.t3719 a_n443_42852.t20 a_15781_43660# VDD.t3718 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1515 a_17749_42852# a_17701_42308# a_17665_42852# VDD.t999 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1516 a_18599_43230# a_18249_42858# a_18504_43218# VDD.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1517 CLK_DATA.t2 a_n2833_47464# VDD.t420 VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1518 VDD.t842 a_7920_46348# a_7715_46873# VDD.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1519 a_3537_45260.t4 a_7287_43370# VSS.t684 VSS.t683 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1520 a_2809_45028# a_526_44458.t20 VDD.t3469 VDD.t3468 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1521 a_7832_46660# a_7715_46873# VDD.t2633 VDD.t2632 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1522 a_3873_46454# a_n881_46662.t8 VSS.t1559 VSS.t1558 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1523 VDD.t232 VSS.t3744 VDD.t231 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1524 VSS.t1349 a_4905_42826# a_4520_42826# VSS.t1348 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1525 a_6709_45028# a_6431_45366# VDD.t1273 VDD.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1526 VSS.t1323 a_20202_43084# a_21421_42336# VSS.t1322 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1527 VSS.t322 a_8953_45002# a_2324_44458.t24 VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 a_20623_43914# a_19321_45002# VSS.t1326 VSS.t1325 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1529 a_20193_45348# a_18494_42460# a_20205_45028# VDD.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1530 VSS.t2270 a_9313_45822# a_11459_47204# VSS.t2269 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1531 a_n4318_39768.t0 a_n2840_43914# VDD.t459 VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1532 a_n443_42852.t5 a_n901_43156# VSS.t635 VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 a_6428_45938# a_5907_45546# VDD.t930 VDD.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1534 C10_N_btm.t5 a_4190_30871.t7 VCM.t7 VSS.t2804 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1535 a_1273_38525.t0 a_1107_38525# VDD.t2687 VDD.t2686 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1536 a_n2104_46634# a_n1925_46634.t4 VDD.t1988 VDD.t1987 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1537 VDD.t162 VSS.t3761 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1538 VSS.t680 a_7287_43370# a_3537_45260.t6 VSS.t679 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 a_2987_42968# a_1847_42826# a_2905_42968# VDD.t2501 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1540 a_11031_47542# a_4915_47217.t2 VDD.t3752 VDD.t3751 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1541 VSS.t2547 a_12991_46634# a_12925_46660# VSS.t2546 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1542 VSS.t434 a_15682_43940# a_11967_42832.t24 VSS.t433 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1543 VDAC_Ni.t4 a_7754_38636# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X1544 VSS.t2413 a_20894_47436# a_20843_47204# VSS.t2412 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 a_13076_44458# a_9482_43914# a_13468_44734# VDD.t1289 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1546 a_10752_42852# a_10083_42826# VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1547 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD.t2691 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1548 a_17970_44736# a_18248_44752# a_18204_44850# VDD.t2198 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1549 a_5663_43940# a_5883_43914# a_5841_44260# VSS.t2021 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1550 a_n2302_38778# a_n2312_38680.t4 VSS.t2616 VSS.t1540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 a_16588_47582# a_15507_47210# a_16241_47178# VDD.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1552 VSS.t2442 a_4099_45572# a_3483_46348.t2 VSS.t2441 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1553 VSS.t817 a_14539_43914# a_16112_44458# VSS.t816 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1554 a_16867_43762# a_16243_43396# a_16759_43396# VDD.t1699 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1555 VDD.t2683 a_1107_38525# a_1273_38525.t3 VDD.t2682 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1556 a_n745_45366# a_n746_45260# VDD.t1250 VDD.t1249 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1557 a_10518_42984# a_10835_43094# a_10793_43218# VSS.t2446 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1558 C2_P_btm.t2 a_n3420_37984.t9 VREF_GND.t27 VSS.t2631 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1559 VIN_P.t8 EN_VIN_BSTR_P.t13 C5_P_btm.t0 VSS.t3565 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1560 a_n37_45144# a_n443_42852.t14 VSS.t3645 VSS.t3644 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1561 a_18287_44626# a_11967_42832.t41 VDD.t3143 VDD.t3142 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1562 a_20159_44458# a_20362_44736# VDD.t2703 VDD.t2702 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1563 VSS.t3585 a_11341_43940.t3 a_22223_43948# VSS.t3584 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1564 VSS.t2336 a_8530_39574# a_3754_38470.t1 VSS.t1546 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1565 DATA[5].t0 a_11459_47204# VDD.t468 VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1566 a_6969_46634# a_n971_45724.t7 VDD.t1908 VDD.t1907 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 VDD.t1025 a_6298_44484# a_4646_46812.t3 VDD.t1024 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1568 a_2324_44458.t25 a_8953_45002# VSS.t299 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1569 a_18861_43218# a_18817_42826# a_18695_43230# VSS.t2380 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1570 a_11322_45546# a_11823_42460.t26 VDD.t3637 VDD.t3636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1571 a_n3674_37592.t2 a_196_42282# VSS.t595 VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1572 a_n1809_43762# a_n1613_43370.t13 VDD.t3370 VDD.t3369 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1573 a_4419_46090# a_526_44458.t32 VDD.t3477 VDD.t3476 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1574 VDD.t2705 a_11189_46129# a_11133_46155# VDD.t2704 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1575 VDD.t733 a_7227_47204# DATA[3].t2 VDD.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1576 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS.t1379 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1577 VSS.t1885 a_7640_43914# a_7584_44260# VSS.t1884 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1578 VSS.t1455 a_21753_35474# SMPL_ON_N.t7 VSS.t1454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 a_15959_42545# a_15764_42576# a_16269_42308# VSS.t2228 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1580 a_16375_45002# a_18597_46090# VSS.t1201 VSS.t1200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1581 VDD.t332 a_n1699_44726# a_n1809_44850# VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1582 a_4235_43370# a_3935_42891# VSS.t2052 VSS.t2051 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1583 a_21177_47436# a_13507_46334.t4 VDD.t1994 VDD.t1993 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1584 a_7418_45394# a_7229_43940# VSS.t2082 VSS.t2081 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1585 a_22000_46634# a_13507_46334.t2 VDD.t1990 VDD.t1989 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1586 VDD.t741 a_7542_44172# a_7499_43940# VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1587 VCM.t48 a_3422_30871.t9 VDAC_P.t1 VSS.t3511 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1588 a_11309_47204# a_11031_47542# VDD.t2546 VDD.t2545 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1589 VDD.t3540 a_1307_43914.t32 a_3353_43940# VDD.t3539 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1590 a_3905_42308# a_2382_45260# VSS.t155 VSS.t154 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1591 a_8483_43230# a_8037_42858# a_8387_43230# VSS.t1470 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1592 a_n2104_46634# a_n1925_46634.t5 VSS.t1739 VSS.t1738 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1593 a_453_43940# a_175_44278# VSS.t3451 VSS.t3450 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1594 a_7281_43914# a_3090_45724.t8 VSS.t1587 VSS.t1586 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1595 a_9028_43914# a_9290_44172.t15 a_9248_44260# VSS.t3062 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1596 EN_VIN_BSTR_P.t0 VDD.t3783 a_n1550_35448# VSS.t3207 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X1597 VDD.t2649 a_n2302_38778# a_n4209_38502.t3 VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1598 VDD.t1593 a_4700_47436# a_3785_47178# VDD.t1592 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1599 a_18909_45814# a_18691_45572# VDD.t3323 VDD.t3322 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1600 a_15521_42308# a_15486_42560# a_15051_42282# VSS.t2230 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1601 a_11551_42558# a_n97_42460.t16 a_11633_42308# VSS.t1679 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1602 VSS.t283 a_11459_47204# DATA[5].t4 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1603 VDD.t3662 a_15227_44166.t9 a_15415_45028# VDD.t3661 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1604 VSS.t3354 a_16327_47482.t10 a_20397_44484# VSS.t3353 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1605 a_n809_44244# a_n984_44318# a_n630_44306# VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1606 VDD.t757 a_8270_45546# a_9165_43940# VDD.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1607 VDD.t1468 a_948_46660# a_1123_46634# VDD.t1467 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1608 VDD.t2576 a_15009_46634# a_14180_46812# VDD.t2575 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1609 a_20766_44850# a_20679_44626# a_20362_44736# VDD.t1649 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1610 C10_N_btm.t28 a_18114_32519.t8 VREF_GND.t11 VSS.t2651 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1611 a_13385_45572# a_10903_43370.t21 a_13297_45572# VSS.t3102 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1612 VDD.t2716 a_13777_45326# a_13807_45067# VDD.t2715 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1613 VSS.t3378 a_n755_45592.t16 a_n39_42308# VSS.t3377 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1614 a_14976_45028# a_14797_45144# VDD.t2718 VDD.t2717 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1615 VSS.t2141 a_22589_40599# a_22537_40625# VSS.t2140 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1616 a_6886_37412# VDAC_Pi.t10 VDD.t2038 VSS.t1790 sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1617 a_6419_46482# a_6165_46155# VSS.t1358 VSS.t1357 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X1618 VSS.t3607 a_768_44030.t11 a_5244_44056# VSS.t3606 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1619 a_n2302_37690# a_n2810_45028.t4 VSS.t2727 VSS.t2726 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1620 VSS.t3238 VDD.t3795 VSS.t3237 VSS.t3190 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1621 VSS.t1899 a_n2946_39072# a_n3565_39304.t4 VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1622 VDD.t973 a_8199_44636# a_8336_45822# VDD.t972 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1623 a_20623_45572# a_20273_45572# a_20528_45572# VDD.t2611 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1624 VSS.t713 a_9396_43370# a_5111_44636# VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1625 a_n2312_39304.t0 a_n1920_47178# VDD.t1174 VDD.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1626 a_20009_46494# a_18819_46122# a_19900_46494# VSS.t2213 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1627 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD.t2492 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1628 a_7309_42852# a_5891_43370.t11 a_7227_42852# VDD.t1877 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1629 a_743_42282.t7 a_13661_43548.t22 VSS.t2904 VSS.t2903 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1630 VSS.t2687 a_n4064_40160.t14 a_n2302_40160# VSS.t2686 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1631 a_22397_42558# a_n913_45002.t17 a_17303_42282# VDD.t2962 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1632 a_12991_43230# a_12545_42858# a_12895_43230# VSS.t1084 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1633 VSS.t2047 a_3905_42865# a_5013_44260# VSS.t2046 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1634 a_22765_42852# a_15743_43084# a_18184_42460.t1 VDD.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1635 a_7705_45326# a_7229_43940# VDD.t2334 VDD.t2333 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1636 VDD.t1019 a_6298_44484# a_4646_46812.t4 VDD.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1637 VSS.t2467 a_10405_44172# a_8016_46348# VSS.t2466 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1638 a_3065_45002# a_1823_45246# VSS.t256 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1639 a_742_44458# a_n443_42852.t8 VSS.t3637 VSS.t3636 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1640 a_310_45028# a_n37_45144# VDD.t2701 VDD.t2700 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1641 VDD.t3037 a_3232_43370.t6 a_2982_43646.t0 VDD.t3036 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1642 VDD.t3479 a_526_44458.t34 a_3905_42558# VDD.t3478 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1643 VSS.t3662 a_18184_42460.t3 a_20256_43172# VSS.t3661 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X1644 VDD.t2276 a_16241_47178# a_16131_47204# VDD.t2275 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1645 a_19466_46812# a_13747_46662.t10 a_19929_45028# VDD.t3090 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1646 VREF.t54 a_n4209_39590.t8 C9_P_btm.t12 VDD.t3072 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1647 a_20850_46482# a_19692_46634.t12 VSS.t1818 VSS.t1817 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1648 VSS.t3615 a_768_44030.t18 a_9028_43914# VSS.t3614 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1649 VDAC_N.t6 a_3422_30871.t7 VCM.t46 VSS.t3509 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1650 a_12089_42308# a_11551_42558# VSS.t686 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1651 a_11173_43940# a_2063_45854.t7 VDD.t1868 VDD.t1867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1652 a_3457_43396# a_1414_42308# VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1653 VDD.t1495 a_5907_46634# a_5894_47026# VDD.t1494 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1654 a_8034_45724# a_8199_44636# VDD.t961 VDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1655 a_5841_46660# a_4651_46660# a_5732_46660# VSS.t2218 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1656 a_22000_46634# a_13507_46334.t12 VSS.t1749 VSS.t1748 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1657 VSS.t2470 a_3699_46348# a_3160_47472# VSS.t2469 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1658 VSS.t1026 a_22223_45036# a_18114_32519.t2 VSS.t1025 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 a_2437_43396# a_1568_43370# VSS.t644 VSS.t643 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VDD.t3329 a_n2104_46634# a_n2312_38680.t0 VDD.t3328 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1661 a_2448_45028# a_2382_45260# a_n2293_45546.t0 VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X1662 C10_P_btm.t19 a_n4315_30879.t11 VREF.t37 VDD.t2071 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1663 a_21167_46155# a_20916_46384# a_20708_46348# VDD.t1054 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1664 a_22725_37990# a_22589_40055# a_22629_37990# VDD.t935 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1665 a_n2438_43548.t28 a_949_44458# VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 a_5205_44484# a_5343_44458# a_5289_44734# VDD.t1262 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1667 a_7499_43078# a_10083_42826# VDD.t917 VDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 a_948_46660# a_33_46660# a_601_46902# VSS.t2471 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1669 VSS.t1050 a_21005_45260# a_19778_44110# VSS.t1049 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1670 VDD.t1151 a_n2302_37690# a_n4209_37414.t3 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1671 VSS.t613 a_13487_47204# a_768_44030.t5 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X1672 a_9241_46436# a_n237_47217.t7 a_8049_45260.t1 VSS.t3031 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1673 a_15015_46420# a_14840_46494# a_15194_46482# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1674 VDD.t132 VSS.t3747 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1675 VSS.t3128 VDD.t3815 VSS.t3127 VSS.t3126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1676 VDD.t2152 a_20567_45036# a_12549_44172.t1 VDD.t2151 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1677 a_21398_44850# a_20640_44752# a_20835_44721# VDD.t2415 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1678 C10_P_btm.t13 a_n4064_40160.t8 VREF_GND.t34 VSS.t2681 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1679 a_1823_45246# a_4704_46090# VSS.t1136 VSS.t1135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1680 a_5527_46155# a_5204_45822# a_5068_46348# VDD.t3483 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1681 a_1606_42308.t2 a_1576_42282# VSS.t100 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1682 VSS.t2460 a_4235_43370# a_4181_43396# VSS.t2459 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 VDD.t939 a_18783_43370# a_18525_43370# VDD.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1684 w_1575_34786.t1 a_n1696_34930.t14 EN_VIN_BSTR_P.t3 w_1575_34786.t0 sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1685 a_n881_46662.t1 a_14495_45572# VDD.t2488 VDD.t2487 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1686 a_21188_45572# a_20107_45572# a_20841_45814# VDD.t2476 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1687 VDD.t78 VSS.t3741 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1688 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS.t2240 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1689 VSS.t3146 VDD.t3821 VSS.t3145 VSS.t3144 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1690 a_22944_39857# a_22613_38993# a_22848_39857# VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1691 VCM.t41 a_5534_30871.t5 C7_N_btm.t1 VSS.t3026 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1692 VSS.t576 a_8270_45546# a_8192_45572# VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1693 VSS.t823 a_6298_44484# a_4646_46812.t27 VSS.t822 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1694 a_5891_43370.t5 a_9127_43156# VSS.t1261 VSS.t1260 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1695 VDD.t699 a_n863_45724# a_3059_42968# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1696 VDD.t2252 a_17609_46634# a_765_45546.t2 VDD.t2251 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1697 VSS.t3383 a_n755_45592.t20 a_3503_45724# VSS.t3382 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 a_19237_31679.t2 a_22959_44484# VSS.t217 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1699 a_12156_46660# a_11813_46116# VDD.t1202 VDD.t1201 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1700 a_n4334_38528# a_n4318_38680.t4 VDD.t2876 VDD.t1983 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1701 a_n901_43156# a_n1076_43230# a_n722_43218# VSS.t1128 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1702 a_n2810_45028.t0 a_n2840_45002# VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1703 VDD.t8 a_949_44458# a_n2438_43548.t5 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1704 a_16333_45814# a_16115_45572# VDD.t540 VDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1705 a_16795_42852# a_n97_42460.t4 a_16877_43172# VSS.t1668 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1706 a_n913_45002.t1 a_526_44458.t8 VDD.t3453 VDD.t2851 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1707 VDD.t1353 a_21188_46660# a_21363_46634# VDD.t1352 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1708 a_6905_45572# a_6151_47436.t5 VSS.t2750 VSS.t2749 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1709 a_14180_45002# a_13059_46348# a_14403_45348# VSS.t1157 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1710 a_16405_45348# a_16375_45002# a_16321_45348# VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1711 VDD.t3688 a_5934_30871.t7 a_8515_42308# VDD.t3687 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1712 VREF.t33 a_19963_31679.t4 C3_N_btm.t2 VDD.t2033 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1713 VDD.t3575 a_3422_30871.t14 a_22315_44484# VDD.t3574 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1714 a_2123_42473# a_n784_42308.t7 VSS.t3532 VSS.t3531 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1715 VSS.t3310 a_n1613_43370.t11 a_n1287_44306# VSS.t3309 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1716 VSS.t1074 a_22223_43948# a_14401_32519.t2 VSS.t1073 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1717 EN_VIN_BSTR_P.t4 a_n1696_34930.t8 w_1575_34786.t3 w_1575_34786.t2 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1718 a_19518_43218# a_16327_47482.t34 VSS.t3296 VSS.t3295 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1719 w_1575_34786.t17 a_n1057_35014.t7 w_1575_34786.t16 w_1575_34786.t10 sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X1720 VSS.t589 a_20075_46420# a_20009_46494# VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1721 VSS.t2593 a_16922_45042# a_16751_45260# VSS.t2592 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1722 VDD.t3041 a_3232_43370.t8 a_11341_43940.t0 VDD.t3040 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X1723 a_1049_43396# a_458_43396# VDD.t2631 VDD.t2630 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1724 VDD.t1204 a_1169_39587# COMP_P.t1 VDD.t1203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1725 VDD.t3467 a_526_44458.t18 a_n913_45002.t0 VDD.t3466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 VDD.t3238 a_n237_47217.t6 a_8270_45546# VDD.t3237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1727 a_1848_45724# a_n237_47217.t12 a_1990_45572# VSS.t3035 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1728 VDD.t1002 a_14539_43914# a_12465_44636# VDD.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1729 VDD.t1784 a_n881_46662.t6 a_7903_47542# VDD.t1783 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1730 VDD.t2947 a_1666_39043.t6 a_1169_39043# VDD.t2946 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1731 VSS.t3482 a_n1696_34930.t15 a_n1057_35014.t0 VSS.t3481 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1732 VDD.t2711 a_n1423_46090# a_n1533_46116# VDD.t2710 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1733 VDD.t1098 a_5111_44636# a_5421_42558# VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1734 a_20623_46660# a_20107_46660# a_20528_46660# VSS.t999 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1735 a_11778_45572# a_10193_42453.t17 a_11688_45572# VSS.t2794 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1736 a_6347_46155# a_6165_46155# VDD.t1566 VDD.t1565 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1737 a_4700_47436# a_n443_46116.t20 a_4842_47570# VSS.t3052 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1738 VDD.t103 VSS.t3737 VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1739 VDD.t2428 a_21359_45002# a_21101_45002# VDD.t2427 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1740 C4_P_btm.t0 a_n3565_38502.t10 VREF.t63 VDD.t3231 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1741 a_14113_42308# a_13575_42558# VSS.t1445 VSS.t1444 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1742 VDD.t2860 a_5755_42308# a_5932_42308.t1 VDD.t2859 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1743 a_10695_43548# a_7499_43078# VDD.t528 VDD.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1744 a_4958_30871.t2 a_17124_42282# VSS.t371 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1745 a_17333_42852# a_16795_42852# VSS.t2124 VSS.t2123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1746 VSS.t1874 a_19339_43156# a_19273_43230# VSS.t1873 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1747 a_8387_43230# a_8037_42858# a_8292_43218# VDD.t1679 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1748 VDD.t2168 a_n2840_44458# a_n4318_40392.t1 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1749 VDD.t534 a_15004_44636# a_14815_43914# VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1750 VSS.t3362 a_16327_47482.t18 a_18861_43218# VSS.t3361 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1751 VSS.t252 a_1823_45246# a_3602_45348# VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VDD.t456 a_18780_47178# a_13661_43548.t1 VDD.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1753 a_n4334_37440# a_n4318_37592.t4 VDD.t3706 VDD.t2043 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1754 VSS.t311 a_8953_45002# a_2324_44458.t26 VSS.t310 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1755 a_2455_43940# a_895_43940# a_2253_43940# VDD.t2250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1756 a_2680_45002# a_3065_45002# a_2809_45028# VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1757 a_13667_43396# a_13661_43548.t6 VDD.t3108 VDD.t3107 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1758 a_21381_43940# a_21115_43940# VSS.t2168 VSS.t2167 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1759 a_380_45546# a_765_45546.t6 a_509_45822# VDD.t3762 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1760 a_15781_43660# a_12549_44172.t9 VDD.t2933 VDD.t2932 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1761 a_16019_45002# a_16147_45260# VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X1762 VDD.t2906 a_3537_45260.t14 a_4558_45348# VDD.t2905 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1763 a_12741_44636.t2 a_6755_46942# a_16789_44484# VSS.t2579 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1764 C9_P_btm.t11 a_n4209_39590.t16 VREF.t60 VDD.t3079 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1765 a_5534_30871.t2 a_12563_42308# VSS.t267 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1766 VSS.t3009 a_2324_44458.t47 a_15682_43940# VSS.t3008 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1767 VDD.t2637 en_comp a_1107_38525# VDD.t2636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1768 VDD.t1452 a_n473_42460# a_n1761_44111# VDD.t1451 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1769 VSS.t1934 a_7754_38470# VSS.t1933 VSS.t1932 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X1770 a_20836_43172# a_20193_45348# VSS.t3449 VSS.t3448 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1771 a_12895_43230# a_12545_42858# a_12800_43218# VDD.t1285 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1772 VSS.t244 a_n2833_47464# CLK_DATA.t6 VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1773 VCM.t54 a_3422_30871.t16 VDAC_N.t0 VSS.t3517 sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X1774 VDD.t1478 a_1123_46634# a_584_46384.t2 VDD.t1477 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 a_726_44056# a_626_44172# a_644_44056# VDD.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1776 a_6655_43762# a_6031_43396# a_6547_43396# VDD.t2435 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1777 DATA[5].t5 a_11459_47204# VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1778 VSS.t416 a_15682_43940# a_11967_42832.t27 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1779 a_2889_44172# a_1414_42308# a_3052_44056# VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1780 VDD.t3039 a_3232_43370.t7 a_3626_43646.t2 VDD.t3038 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1781 a_5700_37509.t19 VDAC_N.t22 a_8912_37509.t30 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1782 a_5343_44458# a_7963_42308# VDD.t1260 VDD.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1783 VSS.t3192 VDD.t3777 VSS.t3191 VSS.t3190 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1784 a_3483_46348.t3 a_4099_45572# VSS.t2444 VSS.t2443 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1785 a_9313_44734.t2 a_5883_43914# a_9241_44734# VDD.t2279 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1786 a_2809_45028# a_1823_45246# VDD.t440 VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1787 VDD.t3608 a_6171_45002.t3 a_11827_44484# VDD.t3607 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1788 w_10694_33990.t9 a_10890_34112.t6 w_10694_33990.t9 w_10694_33990.t7 sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X1789 VDD.t1704 a_9625_46129# a_9569_46155# VDD.t1703 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1790 a_15567_42826# a_15227_44166.t8 VSS.t3589 VSS.t3588 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1791 a_2324_44458.t28 a_8953_45002# VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1792 a_2113_38308# a_2113_38308# a_2113_38308# VSS.t87 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1793 a_7_45899# a_n443_46116.t16 a_n452_45724# VDD.t3252 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1794 a_n2810_45572.t2 a_n2840_45546# VSS.t2324 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1795 a_5732_46660# a_4817_46660# a_5385_46902# VSS.t1019 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1796 a_5708_44484# a_3483_46348.t10 a_5608_44484# VSS.t3077 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X1797 VDD.t256 a_13259_45724.t10 a_22397_42558# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1798 a_11823_42460.t3 a_15051_42282# VDD.t1633 VDD.t1632 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1799 VDD.t1992 a_13507_46334.t3 a_22765_42852# VDD.t1991 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1800 a_13678_32519.t2 a_21855_43396# VSS.t1881 VSS.t1880 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1801 a_5365_45348# a_5111_44636# a_4927_45028# VSS.t907 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1802 a_17021_43396# a_16977_43638# a_16855_43396# VSS.t2397 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1803 VDD.t737 a_7227_47204# DATA[3].t0 VDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1804 VREF_GND.t3 a_n4064_39616.t8 C9_P_btm.t3 VSS.t2844 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1805 a_7989_47542# a_n237_47217.t4 a_7903_47542# VSS.t3030 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1806 a_2324_44458.t16 a_8953_45002# VSS.t316 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1807 a_19332_42282# a_19511_42282# VDD.t2178 VDD.t2177 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1808 VSS.t1987 a_6851_47204# a_7227_47204# VSS.t1986 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1809 a_13607_46688# a_6755_46942# VDD.t2842 VDD.t2841 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1810 a_4880_45572# a_526_44458.t24 a_4808_45572# VSS.t3400 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1811 a_20922_43172# a_10193_42453.t11 a_20836_43172# VSS.t2790 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1812 a_12978_47026# a_11901_46660# a_12816_46660# VDD.t1443 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1813 a_4646_46812.t5 a_6298_44484# VDD.t1007 VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1814 VDD.t1301 a_13720_44458# a_12607_44458# VDD.t1300 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1815 VDD.t665 a_2952_47436# a_2747_46873# VDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1816 a_5147_45002# a_5111_44636# VDD.t1108 VDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1817 VSS.t3236 VDD.t3794 VSS.t3235 VSS.t3234 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1818 VDD.t776 a_14513_46634# a_14543_46987# VDD.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1819 VDD.t1138 a_21259_43561# a_16922_45042# VDD.t1137 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1820 VDD.t1553 a_n4334_38528# a_n4064_38528.t1 VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1821 VSS.t285 a_11459_47204# DATA[5].t6 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1822 VDD.t1752 a_21137_46414# a_21167_46155# VDD.t1751 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1823 C9_N_btm.t6 a_17730_32519.t5 VREF_GND.t8 VSS.t2880 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1824 a_3905_42558# a_1823_45246# VDD.t444 VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1825 VSS.t2318 a_22959_47212# a_22612_30879.t3 VSS.t2317 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1826 a_383_46660# a_33_46660# a_288_46660# VDD.t2727 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1827 VSS.t2581 a_6755_46942# a_13556_45296# VSS.t2580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1828 a_n4209_38216.t4 a_n2302_37984# VSS.t525 VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1829 VSS.t33 a_949_44458# a_n2438_43548.t26 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1830 a_17061_44734# a_11691_44458.t8 a_16979_44734# VDD.t3111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1831 a_4149_42891# a_2382_45260# a_3935_42891# VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X1832 DATA[3].t4 a_7227_47204# VSS.t556 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1833 VDD.t3452 a_n755_45592.t26 a_3318_42354# VDD.t3451 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1834 VDD.t3251 a_n443_46116.t14 a_1427_43646# VDD.t3250 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1835 VDD.t2730 a_5497_46414# a_5527_46155# VDD.t2729 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1836 a_5937_45572.t3 a_5907_45546# VSS.t750 VSS.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1837 a_11323_42473# a_5742_30871.t9 VDD.t2108 VDD.t2107 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1838 VSS.t1508 a_4921_42308# a_5755_42308# VSS.t1507 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1839 a_21076_30879.t0 a_22959_46660# VDD.t945 VDD.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1840 VSS.t3119 VDD.t3812 VSS.t3118 VSS.t3117 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1841 VDD.t2651 a_n2302_38778# a_n4209_38502.t2 VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1842 a_n3565_39304.t6 a_n2946_39072# VSS.t1897 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1843 a_3699_46634# a_3524_46660# a_3878_46660# VSS.t1477 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1844 VDD.t2184 a_17583_46090# a_13259_45724.t0 VDD.t2183 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1845 VSS.t2120 a_3600_43914# a_3499_42826# VSS.t2119 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1846 VSS.t3376 a_n755_45592.t12 a_3318_42354# VSS.t3375 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1847 a_5111_44636# a_9396_43370# VSS.t715 VSS.t714 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1848 a_17595_43084# a_13259_45724.t16 VDD.t252 VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1849 a_13829_44260# a_13059_46348# a_13483_43940# VSS.t1164 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1850 a_18341_45572# a_18175_45572# VSS.t2087 VSS.t2086 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1851 a_9290_44172.t5 a_13635_43156# VSS.t2354 VSS.t2353 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1852 a_12991_46634# a_12816_46660# a_13170_46660# VSS.t3418 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1853 VSS.t932 a_2277_45546# a_2211_45572# VSS.t931 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1854 a_18429_43548# a_18525_43370# VDD.t2520 VDD.t2519 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1855 VSS.t53 a_6453_43914# a_n2661_42282.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1856 a_6773_42558# a_3537_45260.t13 VDD.t2904 VDD.t2903 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1857 a_2253_44260# a_n443_46116.t8 VSS.t3042 VSS.t3041 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1858 C10_N_btm.t7 a_4190_30871.t14 VCM.t9 VSS.t2812 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1859 a_9885_42558# a_7499_43078# a_9803_42558# VDD.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1860 a_16414_43172# a_16137_43396# a_16245_42852# VDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1861 a_21811_47423# SINGLE_ENDED.t0 VDD.t2872 VDD.t2871 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1862 a_2304_45348# a_n863_45724# VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1863 a_3726_37500# a_6886_37412# VSS.t2106 VSS.t2105 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1864 a_13351_46090# a_13507_46334.t6 VDD.t1998 VDD.t1997 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1865 a_n4064_38528.t2 a_n4334_38528# VDD.t1552 VDD.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1866 a_n1435_47204.t1 a_n1605_47204# VSS.t2215 VSS.t2214 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1867 a_n935_46688# a_n1151_42308.t14 a_n1021_46688# VSS.t1661 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1868 VSS.t2703 a_12549_44172.t7 a_17639_46660# VSS.t2702 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X1869 a_6977_45572# a_6598_45938# a_6905_45572# VSS.t2477 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1870 VSS.t2479 a_n23_44458# a_n89_44484# VSS.t2478 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1871 VSS.t2481 a_n1177_43370# a_n1243_43396# VSS.t2480 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1872 VDD.t1671 a_13460_43230# a_13635_43156# VDD.t1670 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1873 VSS.t2729 a_n913_45002.t12 a_n967_45348# VSS.t2728 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1874 VDD.t2603 a_11525_45546# a_11189_46129# VDD.t2602 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1875 VDD.t3440 a_n755_45592.t11 a_626_44172# VDD.t3439 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1876 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1877 VDD.t1842 a_10227_46804.t23 a_10768_47026# VDD.t1841 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1878 a_n755_45592.t3 a_n809_44244# VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1879 a_895_43940# a_644_44056# VSS.t857 VSS.t856 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1880 a_n699_43396# a_n1177_43370# VSS.t2483 VSS.t2482 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1881 a_11136_42852# a_10922_42852# VDD.t2338 VDD.t2337 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1882 VDD.t106 VSS.t3758 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1883 VDD.t2591 a_8568_45546# a_8162_45546# VDD.t2590 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1884 VDD.t1710 a_n4334_37440# a_n4064_37440.t1 VDD.t1709 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1885 a_11551_42558# a_n97_42460.t8 a_11633_42558# VDD.t1897 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_6293_42852# a_5755_42852# VDD.t1416 VDD.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1887 a_n2840_42826# a_n2661_42834.t4 VSS.t1733 VSS.t1732 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1888 a_16131_47204# a_16327_47482.t44 VDD.t3360 VDD.t3359 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1889 a_14033_45572# a_3483_46348.t12 VSS.t3079 VSS.t3078 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1890 a_5289_44734# a_4223_44672.t7 a_5205_44734# VDD.t2898 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1891 VSS.t719 a_n1736_42282# a_n4318_37592.t3 VSS.t718 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1892 VDD.t923 a_10083_42826# a_7499_43078# VDD.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1893 VSS.t3116 VDD.t3811 VSS.t3115 VSS.t3114 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1894 a_768_44030.t4 a_13487_47204# VSS.t609 VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1895 VDD.t2837 a_11415_45002# a_22591_46660# VDD.t2836 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1896 VSS.t673 a_5147_45002# a_5708_44484# VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X1897 VIN_N.t0 EN_VIN_BSTR_N.t8 C8_N_btm.t9 VSS.t2915 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1898 VDD.t243 a_13259_45724.t4 a_14309_45028# VDD.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1899 VSS.t2108 a_6886_37412# a_4338_37500.t6 VSS.t2107 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1900 a_10053_45546# a_10490_45724# a_10210_45822# VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1901 a_n4064_40160.t7 a_n4334_40480# VSS.t2066 VSS.t2065 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1902 VDD.t2182 a_19332_42282# a_4190_30871.t1 VDD.t2181 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1903 a_n998_43396# a_n1613_43370.t10 VSS.t3308 VSS.t3307 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1904 a_3090_45724.t2 a_18911_45144# VDD.t2746 VDD.t2745 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X1905 VSS.t2407 a_18287_44626# a_18248_44752# VSS.t2406 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1906 a_6671_43940# a_6109_44484# a_6453_43914# VDD.t1515 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1907 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD.t2690 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1908 VSS.t851 a_6298_44484# a_4646_46812.t25 VSS.t850 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1909 VDD.t610 a_15682_43940# a_11967_42832.t3 VDD.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1910 VDD.t1154 a_n2302_37690# a_n4209_37414.t2 VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1911 VDD.t1614 a_n2946_37984# a_n3565_38216.t3 VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1912 a_16131_47204# a_15507_47210# a_16023_47582# VDD.t1720 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1913 a_n23_44458# a_n356_44636.t3 VDD.t3655 VDD.t3654 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1914 VSS.t493 a_2779_44458# a_1307_43914.t6 VSS.t492 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1915 a_11750_44172# a_10903_43370.t9 VDD.t3309 VDD.t3308 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1916 a_7845_44172# a_5891_43370.t20 VDD.t1810 VDD.t1809 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1917 VIN_N.t13 EN_VIN_BSTR_N.t21 C1_N_btm.t0 VSS.t2923 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1918 VSS.t3029 a_6123_31319.t6 a_7963_42308# VSS.t1055 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1919 a_5907_46634# a_5732_46660# a_6086_46660# VSS.t1021 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1920 a_8560_45348# a_8746_45002# VSS.t343 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1921 a_19095_43396# a_13661_43548.t18 VSS.t2900 VSS.t2899 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1922 a_21363_46634# a_21188_46660# a_21542_46660# VSS.t1152 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1923 VSS.t1820 a_n4315_30879.t18 a_n4251_40480# VSS.t1819 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1924 VSS.t2847 a_n4064_39616.t10 a_n2302_39866# VSS.t2846 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1925 a_14180_46482# a_14035_46660# VDD.t292 VDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1926 a_n4064_37440.t0 a_n4334_37440# VDD.t1708 VDD.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1927 a_18315_45260# a_18587_45118# a_18545_45144# VDD.t2368 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1928 a_8349_46414# a_8016_46348# VSS.t944 VSS.t943 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1929 a_2537_44260# a_2479_44172# a_2127_44172# VSS.t1877 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1930 C10_N_btm.t24 a_18114_32519.t4 VREF_GND.t16 VSS.t2647 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1931 VSS.t2476 a_3499_42826# a_3445_43172# VSS.t2475 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1932 VDD.t1622 a_3815_47204# a_4007_47204# VDD.t1621 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1933 a_9306_43218# a_n1613_43370.t26 VSS.t3330 VSS.t3329 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1934 VDD.t472 a_6667_45809# a_6598_45938# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1935 a_7230_45938# a_6511_45714# a_6667_45809# VSS.t2494 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1936 VDD.t669 a_2779_44458# a_1307_43914.t3 VDD.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1937 a_8685_43396.t1 a_8147_43396# VSS.t2496 VSS.t2495 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1938 VDD.t1612 a_22400_42852# a_22589_40599# VDD.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1939 VDD.t2059 a_1273_38525.t13 a_1666_39043.t2 VDD.t2056 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1940 VSS.t63 VSS.t61 a_3726_37500# VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X1941 COMP_P.t0 a_1169_39587# VDD.t1206 VDD.t1205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 a_8270_45546# a_n237_47217.t5 VDD.t3236 VDD.t3235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1943 a_15765_45572# a_15599_45572# VSS.t349 VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1944 a_3992_43940# a_768_44030.t14 a_3737_43940# VDD.t3038 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1945 a_3815_47204# a_3785_47178# VSS.t1406 VSS.t1405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1946 a_2063_45854.t3 a_9863_46634# VSS.t2264 VSS.t2263 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1947 VSS.t2577 a_11415_45002# a_22591_46660# VSS.t2576 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1948 a_6755_46942# a_15015_46420# VSS.t616 VSS.t615 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1949 VDD.t2385 a_19431_45546# a_19418_45938# VDD.t2384 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1950 a_11967_42832.t15 a_15682_43940# VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1951 VSS.t2725 a_14021_43940.t2 a_22959_43396# VSS.t1784 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1952 a_19328_44172# a_19478_44306# VSS.t2498 VSS.t2497 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X1953 VSS.t1609 a_10227_46804.t13 a_14537_46482# VSS.t1608 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1954 a_21073_44484# a_16327_47482.t28 VSS.t3369 VSS.t3368 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1955 VDD.t3681 a_768_44030.t10 a_726_44056# VDD.t3680 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1956 VDD.t193 VSS.t3756 VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1957 VDD.t1359 a_13059_46348# a_15297_45822# VDD.t1358 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1958 VSS.t1081 a_12465_44636# a_22223_47212# VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1959 VDD.t2330 a_n1352_43396# a_n1177_43370# VDD.t2329 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1960 VDD.t1655 a_19998_34978# a_21753_35474# VDD.t1654 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1961 VSS.t505 a_n863_45724# a_1067_42314# VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1962 a_19164_43230# a_18083_42858# a_18817_42826# VDD.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1963 a_383_46660# a_n133_46660# a_288_46660# VSS.t1952 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1964 a_3524_46660# a_2443_46660# a_3177_46902# VDD.t2800 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1965 a_13814_43218# a_10227_46804.t11 VSS.t1607 VSS.t1606 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1966 VSS.t1257 a_9127_43156# a_9061_43230# VSS.t1256 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1967 a_11967_42832.t16 a_15682_43940# VSS.t432 VSS.t431 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1968 a_n217_35014# a_n1696_34930.t12 VSS.t3478 VSS.t3477 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1969 VDD.t1295 a_9482_43914# a_10157_44484# VDD.t1294 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1970 VSS.t1536 a_12607_44458# a_12553_44484# VSS.t1535 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1971 VREF.t44 a_n4315_30879.t20 C10_P_btm.t26 VDD.t2080 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1972 VSS.t3095 a_10903_43370.t10 a_11963_45334# VSS.t3094 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1973 VSS.t123 a_17499_43370# a_17433_43396# VSS.t122 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1974 C1_P_btm.t1 a_1606_42308.t5 VCM.t18 VSS.t1728 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1975 VDD.t41 a_12427_45724# a_10490_45724# VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1976 a_13213_44734# a_13259_45724.t8 VDD.t250 VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1977 VSS.t2603 a_14815_43914# a_14761_44260# VSS.t2602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1978 a_12513_46660# a_12469_46902# a_12347_46660# VSS.t1227 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1979 VDD.t404 a_n2302_39072# a_n4209_39304.t2 VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1980 VSS.t2291 a_11323_42473# a_10807_43548# VSS.t2290 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1981 a_18989_43940# a_18451_43940# VDD.t2434 VDD.t2433 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1982 VDD.t6 a_1209_43370# a_n1557_42282# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1983 VSS.t723 a_8667_46634# a_8601_46660# VSS.t722 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1984 VDD.t1084 a_15682_46116# a_11599_46634.t6 VDD.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1985 a_2889_44172# a_2998_44172# VSS.t1107 VSS.t1106 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1986 VSS.t559 a_7281_43914# a_7229_43940# VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VSS.t2316 a_21195_42852# a_21671_42860# VSS.t2315 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1988 a_n2956_38680.t1 a_n2472_46090# VDD.t1733 VDD.t1732 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1989 VSS.t2487 a_n699_43396# a_4743_44484# VSS.t2486 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1990 VDD.t3247 a_n443_46116.t9 a_2437_43646.t1 VDD.t3246 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1991 a_n3565_39590.t6 a_n2946_39866# VSS.t541 VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1992 a_10553_43218# a_10518_42984# a_10083_42826# VSS.t3272 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1993 a_16789_44484# a_14537_43396# VSS.t624 VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1994 VSS.t2356 a_13635_43156# a_13569_43230# VSS.t2355 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1995 a_18834_46812# a_13661_43548.t4 VDD.t3104 VDD.t3103 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1996 a_10405_44172# a_7499_43078# a_10555_44260# VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1997 a_n1151_42308.t3 a_n1329_42308# VSS.t2248 VSS.t2247 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1998 VSS.t240 a_n2833_47464# CLK_DATA.t5 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1999 VSS.t2118 a_18315_45260# a_18189_46348# VSS.t2117 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2000 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS.t2440 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2001 VCM.t4 a_4190_30871.t4 C10_N_btm.t2 VSS.t2801 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2002 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD.t1603 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2003 VDD.t300 a_17499_43370# a_17486_43762# VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2004 VSS.t3168 VDD.t3769 VSS.t3167 VSS.t3166 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2005 VDD.t1438 a_22223_42860# a_22400_42852# VDD.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2006 VDD.t1687 a_3524_46660# a_3699_46634# VDD.t1686 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2007 a_n1059_45260.t2 a_17499_43370# VDD.t306 VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2008 a_5088_37509.t3 VDAC_P.t8 a_8912_37509.t8 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2009 VSS.t2974 a_12861_44030.t15 a_17639_46660# VSS.t2973 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2010 a_10765_43646# a_10695_43548# a_10057_43914# VDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2011 VDD.t2927 a_12549_44172.t5 a_20556_43646# VDD.t2926 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2012 a_15890_42674# a_15803_42450# a_15486_42560# VDD.t2505 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2013 VDD.t1343 a_5815_47464# a_n1613_43370.t3 VDD.t1342 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2014 a_17433_43396# a_16243_43396# a_17324_43396# VSS.t1489 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2015 VCM.t36 a_4958_30871.t10 C9_P_btm.t6 VSS.t2697 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2016 a_11827_44484# a_3232_43370.t10 VDD.t3043 VDD.t3042 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2017 a_1847_42826# a_2351_42308# VSS.t1486 VSS.t1485 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2018 VSS.t2748 a_6151_47436.t4 a_14955_47212# VSS.t2747 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2019 a_20205_31679.t3 a_22223_46124# VSS.t1134 VSS.t1133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2020 VSS.t3603 a_15227_44166.t24 a_15785_43172# VSS.t3602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2021 VDD.t2359 a_1239_47204# a_1431_47204# VDD.t2358 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2022 VDD.t905 a_8667_46634# a_8654_47026# VDD.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2023 VSS.t888 a_15682_46116# a_11599_46634.t27 VSS.t887 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2024 a_n452_45724# a_n443_46116.t12 a_n310_45572# VSS.t3045 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2025 a_700_44734# a_n746_45260# a_327_44734# VDD.t1251 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2026 a_19862_44208# a_13747_46662.t5 VSS.t2862 VSS.t2861 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2027 VREF_GND.t36 a_n4064_40160.t10 C10_P_btm.t10 VSS.t2683 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2028 a_10775_45002# a_9290_44172.t13 VDD.t3266 VDD.t3265 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2029 a_3232_43370.t1 a_526_44458.t16 VDD.t3463 VDD.t3462 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2030 VDD.t394 a_22959_44484# a_19237_31679.t1 VDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2031 a_1115_44172# a_453_43940# a_1443_43940# VDD.t2493 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2032 a_484_44484# a_n863_45724# a_327_44734# VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2033 a_n3690_38528# a_n3674_38680.t4 VDD.t3615 VDD.t2889 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2034 VDD.t2572 a_14543_43071# a_13291_42460# VDD.t2571 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2035 a_2324_44458.t31 a_8953_45002# VSS.t324 VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2036 a_20512_43084# a_11967_42832.t47 VDD.t3150 VDD.t3149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2037 VSS.t2713 a_12549_44172.t21 a_21205_44306# VSS.t2712 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2038 a_20256_43172# a_20202_43084# VSS.t1321 VSS.t1320 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X2039 a_6761_42308# a_n913_45002.t13 a_6773_42558# VDD.t2959 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2040 a_6298_44484# a_2324_44458.t34 VDD.t3205 VDD.t3204 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2041 a_n2840_42282# a_n2661_42282.t2 VSS.t3577 VSS.t3576 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2042 a_n2661_46098# a_1983_46706# a_2162_46660# VSS.t759 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2043 a_5429_46660# a_5385_46902# a_5263_46660# VSS.t997 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2044 VSS.t2504 a_15368_46634# a_15312_46660# VSS.t2503 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2045 VDD.t2868 a_8685_43396.t3 a_14955_43396# VDD.t2867 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2046 VDD.t2349 a_16855_45546# a_16842_45938# VDD.t2348 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2047 VSS.t1144 a_5815_47464# a_n1613_43370.t7 VSS.t1143 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2048 a_11315_46155# a_11133_46155# VDD.t2709 VDD.t2708 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2049 a_16522_42674# a_15803_42450# a_15959_42545# VSS.t2260 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2050 a_1221_42558# a_1184_42692# a_1149_42558# VDD.t2765 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2051 a_20885_46660# a_20841_46902# a_20719_46660# VSS.t2321 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2052 a_20719_45572# a_20273_45572# a_20623_45572# VSS.t2366 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2053 a_1756_43548# a_1307_43914.t18 VSS.t3461 VSS.t3460 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2054 a_14456_42282# a_14635_42282# VSS.t2507 VSS.t2506 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2055 a_n2472_42826# a_n2293_42834.t4 VSS.t1737 VSS.t1736 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2056 a_7276_45260# a_6709_45028# a_7418_45394# VSS.t2429 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2057 VDD.t434 a_1823_45246# a_3232_43370.t2 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2058 a_n4315_30879.t1 a_n2302_40160# VDD.t1372 VDD.t1044 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2059 a_3260_45572# a_3218_45724# a_2957_45546# VSS.t2036 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2060 a_n2497_47436# a_3090_45724.t12 VSS.t1593 VSS.t1592 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2061 VSS.t3506 a_3422_30871.t4 a_22315_44484# VSS.t3505 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2062 C9_N_btm.t16 a_21588_30879.t11 VREF.t11 VDD.t1780 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2063 VDD.t2584 a_10341_42308# a_11554_42852# VDD.t2583 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2064 a_11280_45822# a_2063_45854.t16 a_10907_45822# VDD.t1875 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2065 VDAC_P.t2 a_3422_30871.t10 VCM.t49 VSS.t3512 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2066 a_603_45572# a_310_45028# a_509_45572# VSS.t2468 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2067 a_15002_46116# a_13925_46122# a_14840_46494# VDD.t993 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2068 a_8746_45002# a_7499_43078# VDD.t510 VDD.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2069 a_n906_45572# a_n971_45724.t6 a_n1013_45572# VSS.t1684 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2070 a_11064_45572# a_10903_43370.t5 a_10907_45822# VSS.t3091 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2071 a_21205_44306# a_20935_43940# a_21115_43940# VSS.t2166 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2072 a_2479_44172# a_2905_42968# VDD.t2503 VDD.t2502 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2073 a_12861_44030.t1 a_18143_47464# VDD.t2172 VDD.t2171 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2074 DATA[3].t5 a_7227_47204# VSS.t552 VSS.t551 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2075 VDD.t1408 a_n2840_46090# a_n2956_39304.t1 VDD.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2076 VDD.t2087 a_6945_45028.t4 a_22223_46124# VDD.t2086 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2077 a_11599_46634.t26 a_15682_46116# VSS.t900 VSS.t899 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2078 a_13556_45296# a_6755_46942# VSS.t2583 VSS.t2582 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2079 VREF.t15 a_22612_30879.t7 C10_N_btm.t11 VDD.t1942 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2080 VCM.t22 a_7174_31319.t4 C0_dummy_N_btm.t1 VSS.t1838 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2081 VDD.t969 a_8199_44636# a_9377_42558# VDD.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2082 VREF_GND.t17 a_18114_32519.t11 C10_N_btm.t31 VSS.t2654 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2083 a_n4334_39392# a_n4318_39304.t5 VDD.t1984 VDD.t1983 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2084 a_12710_44260# a_10903_43370.t17 a_12603_44260# VSS.t3099 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2085 a_13777_45326# a_9482_43914# VDD.t1291 VDD.t1290 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2086 a_5088_37509.t5 VDAC_P.t20 a_8912_37509.t10 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2087 a_16522_42674# a_15764_42576# a_15959_42545# VDD.t2479 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2088 a_14205_43396# a_13667_43396# VSS.t2323 VSS.t2322 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X2089 VSS.t25 a_949_44458# a_n2438_43548.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2090 a_8912_37509.t11 VDAC_P.t16 a_5088_37509.t6 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2091 VDD.t1222 a_5732_46660# a_5907_46634# VDD.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2092 a_6419_46155# a_5807_45002# a_6419_46482# VSS.t1281 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2093 VDD.t3581 a_7754_40130.t5 a_8912_37509.t33 VDD.t3580 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2094 a_n2860_39866# a_n2956_39768.t5 a_n2946_39866# VDD.t3093 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2095 VDD.t651 a_13556_45296# a_13857_44734# VDD.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2096 a_18533_44260# a_18326_43940# VSS.t572 VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2097 a_n901_46420# a_n1076_46494# a_n722_46482# VSS.t1251 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2098 a_5066_45546# a_4791_45118.t16 VDD.t2016 VDD.t2015 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2099 a_12861_44030.t5 a_18143_47464# VSS.t1912 VSS.t1911 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2100 VSS.t2955 a_11599_46634.t41 a_18175_45572# VSS.t2954 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2101 VSS.t2352 a_13635_43156# a_9290_44172.t7 VSS.t2351 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2102 VSS.t2947 a_11599_46634.t32 a_18819_46122# VSS.t2946 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2103 a_n3690_37440# a_n3674_37592.t4 VDD.t2894 VDD.t2025 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2104 VSS.t1363 a_n3690_39616# a_n3420_39616.t7 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2105 a_n2442_46660.t3 a_n2472_46634# VSS.t390 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2106 VSS.t1850 a_n1435_47204.t2 a_13487_47204# VSS.t1849 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2107 VDD.t2228 a_3147_46376# a_526_44458.t3 VDD.t2227 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2108 a_8317_43396# a_n755_45592.t9 a_8229_43396# VSS.t3374 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2109 a_n3674_38216.t3 a_n2104_42282# VSS.t141 VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2110 VCM.t45 a_3422_30871.t6 VDAC_N.t4 VSS.t3508 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2111 a_n2312_40392.t3 a_n2288_47178# VSS.t664 VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2112 VDD.t726 a_n1079_45724# a_n1099_45572# VDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2113 VSS.t412 a_22591_44484# a_17730_32519.t3 VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2114 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD.t2774 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2115 a_n97_42460.t0 a_19700_43370# VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2116 VDD.t550 a_n809_44244# a_n755_45592.t1 VDD.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2117 a_3877_44458# a_3699_46634# VSS.t868 VSS.t867 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2118 VDD.t2540 a_22537_40625# a_22725_37990# VDD.t2391 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2119 a_n913_45002.t5 a_1307_43914.t24 VDD.t3530 VDD.t3529 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2120 a_15368_46634# a_15143_45578# VSS.t396 VSS.t395 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2121 a_11206_38545.t0 CAL_N.t4 a_4338_37500.t0 VDD.t3431 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2122 a_4905_42826# a_5379_42460# VSS.t2040 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 VSS.t527 a_10467_46802# a_10428_46928# VSS.t526 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2124 VSS.t1969 a_3147_46376# a_526_44458.t6 VSS.t1968 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2125 a_9313_45822# a_9049_44484# a_9159_45572# VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2126 a_21145_44484# a_20766_44850# a_21073_44484# VSS.t2361 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2127 VDD.t2320 a_n4334_40480# a_n4064_40160.t0 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2128 VSS.t378 a_2680_45002# a_2274_45254# VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2129 VDD.t3211 a_2324_44458.t40 a_15682_43940# VDD.t3210 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2130 VREF_GND.t40 a_n4064_40160.t16 C10_P_btm.t11 VSS.t2689 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2131 a_22613_38993# a_22527_39145# VSS.t482 VSS.t481 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2132 a_10768_47026# a_10554_47026# VDD.t276 VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2133 VSS.t2551 a_21671_42860# a_3422_30871.t2 VSS.t2550 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 a_n785_47204# a_n815_47178# VSS.t3429 VSS.t3428 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 a_5837_45028# a_5807_45002# VDD.t1481 VDD.t1480 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2136 a_5088_37509.t8 VDAC_P.t9 a_8912_37509.t13 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2137 C0_dummy_P_btm.t1 a_7174_31319.t5 VCM.t23 VSS.t1839 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2138 a_14537_43396# a_14358_43442# a_14621_43646# VDD.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2139 a_n3565_38216.t0 a_n2946_37984# VDD.t1613 VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2140 a_n1736_43218# a_n1853_43023# VDD.t587 VDD.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2141 a_6640_46482# a_5257_43370# a_6419_46155# VSS.t1298 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2142 VDD.t1825 a_3090_45724.t20 a_17786_45822# VDD.t1824 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2143 a_n2438_43548.t6 a_949_44458# VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2144 a_15493_43396.t0 a_14955_43396# VDD.t823 VDD.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2145 a_8912_37509.t0 VDAC_P.t22 a_5088_37509.t11 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2146 a_16877_42852# a_n1059_45260.t22 VDD.t2996 VDD.t2995 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2147 a_9823_46482# a_9569_46155# VSS.t1534 VSS.t1533 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X2148 VDD.t2958 a_14021_43940.t3 a_22959_43396# VDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2149 VDD.t2024 a_n3420_38528.t9 a_n2860_38778# VDD.t2023 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2150 VSS.t1603 a_10227_46804.t9 a_12513_46660# VSS.t1602 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2151 VDD.t3293 a_3483_46348.t16 a_17061_44734# VDD.t3292 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2152 VSS.t1483 a_17339_46660# a_19095_43396# VSS.t1482 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2153 a_3699_46348# a_n881_46662.t5 VDD.t1782 VDD.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2154 VSS.t2517 a_10533_42308# a_10723_42308# VSS.t2516 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2155 VSS.t2663 a_3537_45260.t8 a_4223_44672.t3 VSS.t2662 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2156 a_18214_42558# a_n1059_45260.t8 VDD.t2983 VDD.t2982 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2157 VSS.t622 a_14537_43396# a_14180_45002# VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2158 a_16501_45348# a_10193_42453.t9 a_16405_45348# VSS.t2787 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2159 VSS.t652 a_15743_43084# a_15567_42826# VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2160 VSS.t942 a_21259_43561# a_16922_45042# VSS.t941 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2161 VSS.t938 a_n2840_46634# a_n2956_39768.t3 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2162 a_9049_44484# a_8701_44490# VDD.t875 VDD.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2163 VDD.t325 a_2382_45260# a_3737_43940# VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2164 VDD.t2552 a_n967_45348# a_n961_42308# VDD.t2551 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2165 a_19615_44636# a_12861_44030.t10 a_19789_44512# VSS.t2970 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 a_22589_40599# COMP_P.t11 VDD.t1938 VDD.t1937 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2167 a_1273_38525.t1 a_1107_38525# VDD.t2685 VDD.t2684 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2168 VSS.t184 a_1169_39043# comp_n VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2169 a_9863_46634# a_10150_46912# VDD.t2654 VDD.t2653 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2170 VDD.t1796 a_n881_46662.t20 a_n745_45366# VDD.t1795 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2171 VDD.t488 a_8953_45002# a_2324_44458.t2 VDD.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2172 VDD.t2402 a_21496_47436# a_13507_46334.t0 VDD.t2401 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2173 a_n2109_45247# a_n2017_45002.t4 VDD.t3092 VDD.t3091 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2174 VSS.t2519 a_n143_45144# a_n37_45144# VSS.t2518 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2175 SMPL_ON_P.t7 a_n2002_35448# VSS.t2155 VSS.t2154 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2176 a_19418_45938# a_18341_45572# a_19256_45572# VDD.t2344 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2177 VDD.t22 a_949_44458# a_n2438_43548.t14 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2178 VDD.t3742 a_n2438_43548.t38 a_n2433_43396# VDD.t3741 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2179 VDD.t932 a_5907_45546# a_5937_45572.t0 VDD.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X2180 a_11967_42832.t28 a_15682_43940# VSS.t418 VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2181 C5_P_btm.t2 a_n4209_38502.t9 VREF.t52 VDD.t2921 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2182 VSS.t1030 a_n452_44636# a_n2129_44697# VSS.t1029 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2183 a_n2472_42282# a_n2293_42282# VSS.t2521 VSS.t2520 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2184 a_n4318_38680.t3 a_n2472_42826# VSS.t2565 VSS.t2564 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2185 a_5608_44484# a_5111_44636# a_5518_44484# VSS.t915 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X2186 VDD.t975 a_742_44458# a_700_44734# VDD.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2187 VDD.t819 a_n901_43156# a_n443_42852.t2 VDD.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2188 VSS.t3605 a_768_44030.t9 a_13720_44458# VSS.t3604 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2189 VSS.t678 a_7287_43370# a_7221_43396# VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2190 VDD.t2314 a_327_47204# DATA[0].t2 VDD.t2313 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2191 a_2609_46660# a_2443_46660# VDD.t2798 VDD.t2797 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2192 a_n89_44484# a_n467_45028# a_n452_44636# VSS.t2007 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2193 VDD.t3271 a_9290_44172.t21 a_9801_43940# VDD.t3270 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2194 VSS.t3344 a_n1613_43370.t44 a_6809_43396# VSS.t3343 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2195 a_n4064_39616.t5 a_n4334_39616# VSS.t166 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2196 a_556_44484# a_526_44458.t9 a_484_44484# VSS.t3391 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2197 VDD.t784 a_n4334_39392# a_n4064_39072.t2 VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2198 VSS.t2149 a_4007_47204# DATA[2].t6 VSS.t2148 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2199 VDD.t3169 a_2324_44458.t59 a_15682_46116# VDD.t3168 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2200 a_8912_37509.t7 VDAC_P.t11 a_5088_37509.t2 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2201 a_2112_39137# a_1273_38525.t8 VDD.t2055 VDD.t2054 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2202 VSS.t2500 a_19328_44172# a_19279_43940# VSS.t2499 sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2203 VDD.t3432 CAL_N.t5 VDD.t3432 VDD.t1755 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2204 VDD.t3639 a_n3420_37440.t8 a_n2860_37690# VDD.t2887 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2205 a_n3420_38528.t2 a_n3690_38528# VDD.t2524 VDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2206 VSS.t301 a_8953_45002# a_2324_44458.t27 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2207 a_4646_46812.t6 a_6298_44484# VDD.t1021 VDD.t1020 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2208 a_10554_47026# a_10467_46802# a_10150_46912# VDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2209 a_11387_46155# a_n1151_42308.t18 a_11315_46155# VDD.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2210 a_10341_43396.t0 a_9803_43646# VDD.t1550 VDD.t1549 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2211 a_13887_32519.t1 a_22223_43396# VDD.t1561 VDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2212 VSS.t1601 a_10227_46804.t7 a_20885_46660# VSS.t1600 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2213 C0_P_btm.t2 a_n3420_37440.t9 VREF_GND.t45 VSS.t3530 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2214 VIN_P.t15 EN_VIN_BSTR_P.t14 C2_P_btm.t1 VSS.t3566 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2215 VSS.t384 a_16137_43396# a_18548_42308# VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2216 a_n452_45724# a_n743_46660.t3 a_n310_45899# VDD.t3638 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2217 a_11682_45822# a_11652_45724# VDD.t2629 VDD.t2628 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2218 a_n443_42852.t1 a_n901_43156# VDD.t813 VDD.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2219 VDD.t1731 a_n2472_46090# a_n2956_38680.t0 VDD.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2220 VDD.t1080 a_15682_46116# a_11599_46634.t8 VDD.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2221 VDD.t1581 a_11322_45546# a_11280_45822# VDD.t1580 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2222 VSS.t2873 a_13747_46662.t12 a_14495_45572# VSS.t2872 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2223 VDD.t3648 a_10809_44734.t5 a_n2661_42834.t0 VDD.t3647 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2224 C0_dummy_P_btm.t0 EN_VIN_BSTR_P.t17 VIN_P.t12 VSS.t3569 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2225 VSS.t2858 a_n4209_39590.t10 a_n4251_39616# VSS.t1719 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2226 VSS.t2246 a_n1329_42308# a_n1151_42308.t2 VSS.t2245 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2227 a_3381_47502# a_2905_45572# VSS.t2363 VSS.t2362 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2228 VDD.t1595 a_18479_47436# a_13747_46662.t2 VDD.t1594 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2229 VSS.t1046 a_n746_45260# a_261_44278# VSS.t1045 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2230 VDD.t398 a_n2302_39072# a_n4209_39304.t1 VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2231 a_5649_42852.t0 a_5111_42852# VDD.t1560 VDD.t1559 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2232 VSS.t3262 VDD.t3804 VSS.t3261 VSS.t3260 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2233 a_11136_45572# a_3483_46348.t4 a_11064_45572# VSS.t3074 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2234 VSS.t1244 a_13249_42308# a_13904_45546# VSS.t1243 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2235 a_17486_43762# a_16409_43396# a_17324_43396# VDD.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2236 VSS.t2737 a_n913_45002.t24 a_8325_42308# VSS.t2736 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2237 VSS.t3458 a_1307_43914.t16 a_2675_43914# VSS.t3457 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2238 VCM.t17 a_4190_30871.t10 C10_P_btm.t7 VSS.t2808 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2239 a_3699_46634# a_n1613_43370.t28 VDD.t3380 VDD.t3379 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2240 VSS.t71 a_13259_45724.t7 a_14797_45144# VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2241 VSS.t2994 a_2324_44458.t32 a_949_44458# VSS.t2993 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2242 a_20841_45814# a_20623_45572# VDD.t2478 VDD.t2477 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2243 VIN_N.t7 EN_VIN_BSTR_N.t18 C9_N_btm.t8 VSS.t2924 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2244 VDD.t93 VSS.t3731 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2245 a_17639_46660# a_12861_44030.t20 VSS.t2982 VSS.t2981 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2246 a_10341_42308# a_9803_42558# VSS.t2340 VSS.t2339 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2247 a_16327_47482.t0 a_17591_47464# VDD.t2125 VDD.t2124 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2248 a_19998_34978# VDD.t3785 EN_VIN_BSTR_N.t2 VSS.t3211 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X2249 VSS.t2997 a_2324_44458.t36 a_15682_46116# VSS.t1744 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2250 a_1260_45572# a_n755_45592.t18 a_1176_45572# VSS.t3379 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X2251 a_20397_44484# a_20362_44736# a_20159_44458# VSS.t2451 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2252 a_12991_46634# a_10227_46804.t6 VDD.t1830 VDD.t1829 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2253 a_518_46155# a_472_46348# VDD.t1420 VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2254 a_n4064_39072.t0 a_n4334_39392# VDD.t778 VDD.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2255 VDD.t1248 a_20841_45814# a_20731_45938# VDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2256 a_9751_46155# a_9569_46155# VDD.t1748 VDD.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2257 a_1443_43940# a_1414_42308# a_1241_43940# VDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2258 VREF.t14 a_22612_30879.t6 C10_N_btm.t10 VDD.t1941 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X2259 DATA[1].t2 a_1431_47204# VDD.t2117 VDD.t2116 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2260 VDD.t3623 a_11823_42460.t10 a_14033_45822# VDD.t3622 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2261 VSS.t1155 a_n2840_42826# a_n3674_39304.t3 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2262 VSS.t2677 a_3537_45260.t28 a_5365_45348# VSS.t2676 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2263 a_3065_45002# a_3318_42354# VSS.t2345 VSS.t2344 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2264 a_n310_45899# a_n356_45724# VDD.t3513 VDD.t3512 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2265 C8_P_btm.t7 a_n3420_39616.t11 VREF_GND.t29 VSS.t2644 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2266 a_16327_47482.t6 a_17591_47464# VSS.t1867 VSS.t1866 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2267 VDD.t1681 a_22591_46660# a_20820_30879.t1 VDD.t1680 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2268 a_n3420_37440.t2 a_n3690_37440# VDD.t2550 VDD.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2269 a_8337_42558# a_5891_43370.t16 VDD.t1806 VDD.t1805 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2270 VDD.t3127 a_4646_46812.t34 a_7411_46660# VDD.t3126 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2271 a_11186_47026# a_10428_46928# a_10623_46897# VDD.t2294 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2272 a_20273_46660# a_20107_46660# VDD.t1197 VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2273 VSS.t143 a_3877_44458# a_2382_45260# VSS.t142 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2274 VDD.t448 a_n1331_43914# a_n1441_43940# VDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2275 VDD.t2698 a_10835_43094# a_10796_42968# VDD.t2697 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2276 VSS.t168 a_5066_45546# a_9159_45572# VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2277 VSS.t172 a_12883_44458# a_12829_44484# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2278 a_11341_43940.t2 a_10729_43914# a_11257_43940# VDD.t1145 sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2279 VREF.t55 a_n4209_39590.t9 C9_P_btm.t14 VDD.t3073 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2280 VSS.t799 a_564_42282# a_n1794_35082.t2 VSS.t798 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2281 a_12549_44172.t0 a_20567_45036# VDD.t2150 VDD.t2149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2282 VDD.t2771 a_14456_42282# a_5342_30871.t1 VDD.t2770 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2283 a_645_46660# a_601_46902# a_479_46660# VSS.t2001 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2284 VDD.t1866 a_2063_45854.t4 a_10809_44734.t1 VDD.t1865 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2285 VDD.t1162 a_2127_44172# a_n2661_45010# VDD.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2286 VDD.t1856 a_10227_46804.t32 a_16104_42674# VDD.t1855 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2287 a_12861_44030.t3 a_18143_47464# VDD.t2174 VDD.t2173 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2288 a_14513_46634# a_14180_46812# VDD.t2619 VDD.t2618 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2289 a_n2840_46090# a_n2661_46098# VSS.t2502 VSS.t1791 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2290 a_5088_37509.t16 VSS.t3739 VDAC_Ni.t0 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2291 a_21137_46414# a_19692_46634.t3 VDD.t2061 VDD.t2060 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2292 a_1609_45822# a_167_45260# a_1609_45572# VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2293 VREF_GND.t7 a_17730_32519.t6 C9_N_btm.t5 VSS.t2881 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2294 a_14635_42282# a_n913_45002.t26 VSS.t2741 VSS.t2740 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2295 a_10544_45572# a_10490_45724# a_10053_45546# VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X2296 a_10555_44260# a_10949_43914# a_10405_44172# VSS.t859 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X2297 C2_P_btm.t3 a_n3565_38216.t10 VREF.t73 VDD.t3766 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2298 VSS.t1852 a_1431_47204# DATA[1].t6 VSS.t1851 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2299 VDD.t87 VSS.t3723 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2300 a_8952_43230# a_7871_42858# a_8605_42826# VDD.t1674 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2301 a_3067_47026# a_n1613_43370.t36 VDD.t3386 VDD.t3385 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2302 a_9377_42558# a_8685_42308# a_9293_42558# VDD.t2235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2303 a_4190_30871.t2 a_19332_42282# VSS.t1916 VSS.t1915 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2304 VDD.t1214 a_9067_47204# DATA[4].t1 VDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2305 a_15861_45028# a_15595_45028# VDD.t2164 VDD.t2163 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2306 a_15194_46482# a_10227_46804.t4 VSS.t1599 VSS.t1598 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2307 a_6469_45572# a_5907_45546# VSS.t748 VSS.t747 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2308 a_13720_44458# a_9482_43914# a_14112_44734# VDD.t1296 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2309 a_15493_43940# a_14955_43940# VDD.t1734 VDD.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2310 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS.t2075 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2311 a_16245_42852# a_n1059_45260.t9 VDD.t2985 VDD.t2984 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2312 VSS.t1827 a_n357_42282.t5 a_6101_43172# VSS.t1826 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2313 a_20692_30879.t2 a_22959_46124# VSS.t1956 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2314 VSS.t521 a_n2302_37984# a_n4209_38216.t5 VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2315 a_3177_46902# a_2959_46660# VDD.t2784 VDD.t2783 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2316 a_5907_46634# a_n1613_43370.t32 VDD.t3384 VDD.t3383 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2317 a_5497_46414# a_5164_46348# VDD.t362 VDD.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2318 VSS.t928 a_104_43370# a_n971_45724.t3 VSS.t927 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2319 VREF_GND.t21 a_13258_32519.t4 C0_N_btm.t2 VSS.t1673 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2320 VDD.t1315 a_4743_44484# a_4791_45118.t0 VDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2321 a_19700_43370# a_18579_44172# VSS.t2428 VSS.t2427 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2322 a_12861_44030.t7 a_18143_47464# VSS.t1908 VSS.t1907 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2323 a_21363_46634# a_10227_46804.t28 VDD.t1850 VDD.t1849 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2324 VSS.t3649 a_n443_42852.t22 a_15940_43402# VSS.t3648 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X2325 a_12427_45724# a_11823_42460.t22 VDD.t3633 VDD.t3632 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X2326 VSS.t1365 a_n3690_39616# a_n3420_39616.t6 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2327 a_5891_43370.t4 a_9127_43156# VSS.t1253 VSS.t1252 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 a_n1920_47178# a_n1741_47186.t9 VDD.t2110 VDD.t2109 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2329 a_10903_43370.t3 a_13351_46090# VSS.t657 VSS.t656 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2330 a_n955_45028# a_n1059_45260.t20 VDD.t2993 VDD.t2992 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2331 SMPL_ON_P.t6 a_n2002_35448# VSS.t2159 VSS.t2158 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2332 VDD.t2093 a_n357_42282.t11 a_7309_42852# VDD.t2092 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2333 VDD.t2222 a_3147_46376# a_526_44458.t0 VDD.t2221 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2334 a_18596_45572# a_18479_45785# VSS.t2527 VSS.t2526 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2335 a_4185_45028.t2 a_3065_45002# VDD.t563 VDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2336 a_6575_47204# a_6545_47178# VSS.t2193 VSS.t2192 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2337 a_16137_43396# a_15781_43660# VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2338 VCM.t3 a_4190_30871.t5 C10_N_btm.t1 VSS.t2802 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2339 VSS.t1038 a_22775_42308# a_22485_38105# VSS.t1037 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2340 VSS.t388 a_n2472_46634# a_n2442_46660.t2 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2341 a_4649_42852# a_526_44458.t22 VDD.t3473 VDD.t3472 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2342 VSS.t3660 a_2711_45572.t10 a_20107_42308# VSS.t3659 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2343 VSS.t139 a_n2104_42282# a_n3674_38216.t2 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2344 VSS.t618 a_15015_46420# a_14949_46494# VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2345 VSS.t920 a_5691_45260# a_n2109_47186.t1 VSS.t919 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2346 a_17583_46090# a_17715_44484# VSS.t2015 VSS.t2014 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2347 a_17730_32519.t2 a_22591_44484# VSS.t410 VSS.t409 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2348 a_3600_43914# a_1307_43914.t30 VSS.t3470 VSS.t3469 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X2349 VSS.t1941 a_n1550_35448# a_n2002_35448# VSS.t1940 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2350 a_13925_46122# a_13759_46122# VDD.t1625 VDD.t1624 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2351 VDD.t821 a_n901_43156# a_n914_42852# VDD.t820 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2352 a_8191_45002# a_3483_46348.t8 VDD.t3287 VDD.t3286 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2353 VDD.t2212 a_22959_46124# a_20692_30879.t1 VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2354 a_n310_44484# a_n356_44636.t4 VSS.t3581 VSS.t3580 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2355 a_21125_42558# a_18597_46090# VDD.t1398 VDD.t1397 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 VDD.t1208 a_1169_39587# COMP_P.t3 VDD.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2357 a_5932_42308.t0 a_5755_42308# VDD.t2858 VDD.t2857 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2358 VSS.t2329 a_14543_43071# a_13291_42460# VSS.t2328 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2359 VDD.t3553 a_1307_43914.t14 a_n913_45002.t7 VDD.t3552 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2360 VSS.t1973 a_3147_46376# a_526_44458.t7 VSS.t1972 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2361 VDD.t883 a_n2946_38778# a_n3565_38502.t0 VDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2362 VDD.t1388 a_16112_44458# a_14673_44172# VDD.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2363 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD.t1590 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2364 a_3175_45822# a_3316_45546# VDD.t1570 VDD.t1569 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2365 VSS.t707 a_16763_47508# a_5807_45002# VSS.t706 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2366 VREF.t50 a_20447_31679.t4 C5_N_btm.t2 VDD.t2102 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2367 a_14226_46660# a_14180_46812# VSS.t2375 VSS.t2374 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2368 VDD.t2230 a_13348_45260# a_13159_45002# VDD.t2229 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2369 a_4646_46812.t22 a_6298_44484# VSS.t825 VSS.t824 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2370 VDD.t2237 a_6491_46660# a_6851_47204# VDD.t2236 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2371 VSS.t3174 VDD.t3771 VSS.t3173 VSS.t3172 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2372 a_n4209_39590.t3 a_n2302_39866# VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2373 a_6511_45714# a_4646_46812.t40 VDD.t3131 VDD.t3130 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2374 a_n2438_43548.t10 a_949_44458# VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2375 VDD.t1239 a_22775_42308# a_22485_38105# VDD.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2376 a_3422_30871.t3 a_21671_42860# VSS.t2553 VSS.t2552 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2377 VSS.t711 a_16763_47508# a_16697_47582# VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2378 VDD.t1270 a_2889_44172# a_413_45260.t0 VDD.t1269 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X2379 VREF.t22 a_22612_30879.t14 C10_N_btm.t18 VDD.t1949 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2380 VSS.t3652 a_n443_42852.t24 a_1755_42282# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2381 C10_P_btm.t2 a_4190_30871.t8 VCM.t12 VSS.t2805 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2382 a_10405_44172# a_10729_43914# a_10651_43940# VDD.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2383 a_n2840_45546# a_n2661_45546.t3 VDD.t3693 VDD.t2761 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2384 a_14401_32519.t1 a_22223_43948# VDD.t1277 VDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2385 VREF.t3 a_21076_30879.t7 C8_N_btm.t3 VDD.t3557 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2386 a_4558_45348# a_4574_45260# VDD.t2260 VDD.t2259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2387 VDD.t173 VSS.t3745 VDD.t172 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2388 a_5193_42852# a_3905_42865# a_5111_42852# VDD.t2306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2389 a_18143_47464# a_18479_47436# VSS.t1383 VSS.t1382 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2390 a_10533_42308# a_n913_45002.t22 a_10545_42558# VDD.t2964 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2391 VDD.t2266 a_16721_46634# a_16751_46987# VDD.t2265 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2392 a_18909_45814# a_18691_45572# VSS.t3269 VSS.t3268 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2393 a_n2840_45002# a_n2661_45010# VDD.t1164 VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2394 a_948_46660# a_n133_46660# a_601_46902# VDD.t2207 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2395 a_3699_46348# a_3877_44458# a_3873_46454# VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2396 a_117_45144# a_n443_42852.t12 a_45_45144# VDD.t3710 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2397 a_11415_45002# a_13249_42308# VDD.t1449 VDD.t1448 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2398 VSS.t3252 VDD.t3800 VSS.t3251 VSS.t3250 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2399 a_15681_43442# a_12861_44030.t8 VSS.t2967 VSS.t2966 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2400 C10_N_btm.t8 a_22612_30879.t4 VREF.t12 VDD.t1939 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2401 a_n4209_38502.t4 a_n2302_38778# VSS.t2399 VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2402 VREF_GND.t14 a_18114_32519.t9 C10_N_btm.t29 VSS.t2652 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2403 VDD.t3434 CAL_N.t6 VDD.t3433 VDD.t1758 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X2404 VDD.t2989 a_n1059_45260.t16 a_18727_42674# VDD.t2988 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2405 VSS.t3425 a_5013_44260# a_5663_43940# VSS.t3424 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2406 a_9801_43940# a_3483_46348.t7 VDD.t3285 VDD.t3284 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2407 VSS.t2789 a_10193_42453.t10 a_18797_44260# VSS.t2788 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2408 a_n4251_38304# a_n4318_38216.t5 a_n4334_38304# VSS.t1795 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2409 a_2779_44458# a_1423_45028.t4 VDD.t1968 VDD.t1967 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2410 a_19789_44512# a_12549_44172.t27 VSS.t2721 VSS.t2720 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X2411 VDD.t2681 a_1107_38525# a_1273_38525.t2 VDD.t2680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2412 comp_n a_1169_39043# VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2413 VDD.t1311 a_18057_42282# a_n356_44636.t0 VDD.t1310 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X2414 a_13113_42826# a_12895_43230# VDD.t1524 VDD.t1523 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2415 a_16197_42308# a_10227_46804.t22 VSS.t1621 VSS.t1620 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2416 a_11599_46634.t10 a_15682_46116# VDD.t1082 VDD.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2417 VDD.t1493 a_8034_45724# a_n1925_46634.t2 VDD.t1492 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2418 VDD.t3113 a_11691_44458.t9 a_11649_44734# VDD.t3112 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2419 VSS.t3416 a_22581_37893# a_22537_39537# VSS.t753 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2420 VSS.t2157 a_n2002_35448# SMPL_ON_P.t5 VSS.t2156 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2421 a_n3690_39392# a_n3674_39304.t5 VDD.t2890 VDD.t2889 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2422 a_15761_42308# a_15051_42282# VSS.t1422 VSS.t1421 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2423 a_16680_45572# a_15765_45572# a_16333_45814# VSS.t2231 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2424 VSS.t646 a_1568_43370# a_1512_43396# VSS.t645 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2425 VDD.t3060 a_n1794_35082.t8 a_n1696_34930.t0 VDD.t3059 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2426 VDD.t342 a_5066_45546# a_5024_45822# VDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2427 VSS.t361 a_n809_44244# a_n875_44318# VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2428 VDD.t282 a_n2946_37690# a_n3565_37414.t1 VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2429 a_n2267_43396# a_n2433_43396# VDD.t2689 VDD.t2688 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2430 a_10518_42984# a_10796_42968# a_10752_42852# VDD.t3325 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2431 VDD.t1474 a_1123_46634# a_584_46384.t3 VDD.t1473 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2432 a_8189_46660# a_8145_46902# a_8023_46660# VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2433 VDD.t3115 a_13661_43548.t9 a_14976_45028# VDD.t3114 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X2434 a_11691_44458.t2 a_5807_45002# VSS.t1277 VSS.t1276 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2435 VSS.t2860 a_n4064_39072.t10 a_n2302_39072# VSS.t2846 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2436 a_20062_46116# a_18985_46122# a_19900_46494# VDD.t2301 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2437 a_20269_44172# a_20365_43914# VSS.t2418 VSS.t2417 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2438 VSS.t1653 a_5891_43370.t10 a_5837_43396# VSS.t1652 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2439 VSS.t2567 a_n2472_42826# a_n4318_38680.t2 VSS.t2566 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2440 VSS.t1929 a_7754_38470# a_7754_38470# VSS.t1928 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2441 a_18707_42852# a_18083_42858# a_18599_43230# VDD.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2442 VDD.t2312 a_327_47204# DATA[0].t0 VDD.t2311 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2443 a_12638_46436# a_13059_46348# VSS.t1163 VSS.t1162 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2444 VDD.t129 VSS.t3729 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2445 a_n784_42308.t3 a_n961_42308# VSS.t2312 VSS.t2311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2446 a_13157_43218# a_13113_42826# a_12991_43230# VSS.t1317 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2447 VSS.t2145 a_4007_47204# DATA[2].t7 VSS.t2144 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2448 VDD.t800 a_15015_46420# a_15002_46116# VDD.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2449 VDD.t3427 a_16327_47482.t30 a_20159_44458# VDD.t3426 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2450 a_8912_37509.t17 VDAC_N.t9 a_5700_37509.t18 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2451 VSS.t3433 a_n785_47204# a_327_47204# VSS.t3432 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2452 a_18834_46812# a_13661_43548.t8 VSS.t2891 VSS.t2890 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2453 a_n2840_45546# a_n2661_45546.t4 VSS.t3624 VSS.t972 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2454 VSS.t1193 a_21177_47436# a_20990_47178# VSS.t1192 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2455 VSS.t335 a_7499_43078# a_11816_44260# VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2456 a_n3420_38528.t3 a_n3690_38528# VDD.t2523 VDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2457 a_6761_42308# a_3537_45260.t24 VSS.t2674 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2458 a_10623_46897# a_10428_46928# a_10933_46660# VSS.t2038 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2459 a_5263_45724# a_n881_46662.t14 VDD.t1788 VDD.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2460 VDD.t3628 a_11823_42460.t14 a_11322_45546# VDD.t3627 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2461 VSS.t917 a_5111_44636# a_8018_44260# VSS.t916 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2462 a_7903_47542# a_n237_47217.t8 VDD.t3240 VDD.t3239 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2463 VSS.t725 a_8667_46634# a_n237_47217.t3 VSS.t724 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 a_3357_43084.t2 a_4905_42826# VDD.t1557 VDD.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2465 a_n2472_46090# a_n2293_46098.t2 VSS.t2615 VSS.t2614 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2466 VREF.t64 a_19237_31679.t4 C0_N_btm.t0 VDD.t3547 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2467 SMPL_ON_N.t6 a_21753_35474# VSS.t1451 VSS.t1450 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2468 VCM.t24 a_5742_30871.t4 C6_P_btm.t3 VSS.t1843 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2469 VSS.t754 a_22589_40055# a_22527_39145# VSS.t753 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 VDD.t815 a_n901_43156# a_n443_42852.t3 VDD.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2471 VSS.t761 a_22959_46660# a_21076_30879.t3 VSS.t760 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2472 a_10249_46116# a_9823_46155# VDD.t766 VDD.t765 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X2473 VDD.t2426 a_10775_45002# a_10180_45724# VDD.t2425 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X2474 CAL_N.t0 a_22485_38105# VDD.t1244 VDD.t1242 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2475 a_2684_37794# VDAC_Pi.t9 a_2113_38308# VSS.t1789 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2476 VDD.t217 VSS.t3718 VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2477 a_8696_44636.t0 a_16855_45546# VDD.t2347 VDD.t2346 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2478 a_n4209_37414.t6 a_n2302_37690# VSS.t964 VSS.t963 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2479 a_13467_32519.t3 a_21487_43396# VSS.t767 VSS.t766 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2480 a_6633_46155# a_5807_45002# a_6419_46155# VDD.t1489 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2481 a_n2661_42834.t2 a_8975_43940# VDD.t2351 VDD.t2350 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2482 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS.t2439 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2483 a_7274_43762# a_6197_43396# a_7112_43396# VDD.t2331 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2484 a_10922_42852# a_10835_43094# a_10518_42984# VDD.t2699 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2485 DATA[0].t4 a_327_47204# VSS.t2054 VSS.t2053 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2486 VDD.t1488 a_5807_45002# a_11691_44458.t1 VDD.t1487 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2487 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD.t2327 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2488 C10_N_btm.t3 a_4190_30871.t18 VCM.t5 VSS.t2815 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2489 a_n4209_38502.t0 a_n2302_38778# VDD.t2648 VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2490 VSS.t1545 RST_Z.t2 a_14311_47204# VSS.t1544 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2491 a_16327_47482.t3 a_17591_47464# VDD.t2127 VDD.t2126 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2492 a_18285_46348# a_18834_46812# VDD.t2377 VDD.t2376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2493 EN_VIN_BSTR_N.t5 a_18194_34908.t14 w_10694_33990.t11 w_10694_33990.t10 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2494 VREF.t40 a_n4315_30879.t14 C10_P_btm.t22 VDD.t2074 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2495 a_18597_46090# a_19431_45546# VDD.t2387 VDD.t2386 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2496 VSS.t2530 a_18443_44721# a_18374_44850# VSS.t2529 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2497 VSS.t777 a_8199_44636# a_10951_45334# VSS.t776 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2498 a_1176_45572# a_167_45260# VSS.t203 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2499 a_7735_45067# a_6709_45028# a_7276_45260# VDD.t2679 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2500 C8_P_btm.t8 a_5342_30871.t6 VCM.t30 VSS.t2624 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2501 DATA[4].t0 a_9067_47204# VDD.t1212 VDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2502 C10_P_btm.t16 a_n4315_30879.t8 VREF.t34 VDD.t2068 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X2503 a_n3565_39304.t7 a_n2946_39072# VSS.t1898 VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2504 VSS.t2388 a_n2109_45247# en_comp VSS.t2387 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2505 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS.t2514 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2506 DATA[1].t1 a_1431_47204# VDD.t2115 VDD.t2114 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2507 a_13348_45260# a_13556_45296# a_13490_45394# VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2508 C10_P_btm.t8 a_n4064_40160.t17 VREF_GND.t41 VSS.t2690 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2509 a_n2302_40160# a_n2312_40392.t4 VSS.t1647 VSS.t1646 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2510 VSS.t2534 a_21356_42826# a_n357_42282.t3 VSS.t2533 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2511 VDD.t3703 a_11453_44696.t4 a_22959_47212# VDD.t1977 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2512 VSS.t394 a_15037_45618# a_15143_45578# VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2513 VSS.t1714 a_8696_44636.t9 a_8701_44490# VSS.t1713 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2514 a_3878_46660# a_n1613_43370.t16 VSS.t3314 VSS.t3313 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2515 a_2277_45546# a_167_45260# VSS.t207 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2516 a_626_44172# a_n863_45724# VDD.t701 VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2517 a_18479_45785# a_19268_43646# VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2518 a_16327_47482.t7 a_17591_47464# VSS.t1865 VSS.t1864 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2519 a_20273_45572# a_20107_45572# VSS.t2223 VSS.t2222 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2520 a_10555_44260# a_5891_43370.t9 VSS.t1651 VSS.t1650 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2521 a_n3420_37440.t3 a_n3690_37440# VDD.t2548 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2522 VSS.t3639 a_n443_42852.t9 a_742_44458# VSS.t3638 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2523 VSS.t631 a_n901_43156# a_n967_43230# VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2524 a_20820_30879.t0 a_22591_46660# VDD.t1683 VDD.t1682 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2525 VSS.t65 a_13076_44458# a_12883_44458# VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X2526 a_685_42968# a_n443_42852.t16 VSS.t3647 VSS.t3646 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2527 a_17364_32525.t0 a_22959_43396# VDD.t2431 VDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2528 a_13170_46660# a_10227_46804.t20 VSS.t1617 VSS.t1616 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2529 a_11633_42558# a_9290_44172.t19 a_11551_42558# VDD.t3269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2530 VDD.t2008 a_4791_45118.t8 a_6633_46155# VDD.t2007 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2531 a_20731_45938# a_16327_47482.t13 VDD.t3409 VDD.t3408 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2532 a_19700_43370# a_18579_44172# VDD.t2677 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2533 VDD.t3152 a_11599_46634.t34 a_20107_46660# VDD.t3151 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2534 a_16751_45260# a_17023_45118# a_16981_45144# VDD.t2504 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2535 a_2382_45260# a_3877_44458# VSS.t145 VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2536 C9_N_btm.t10 a_21588_30879.t8 VREF.t8 VDD.t1777 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2537 VSS.t607 a_13487_47204# a_768_44030.t7 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2538 a_12829_44484# a_12741_44636.t6 a_n2293_43922.t2 VSS.t1727 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2539 a_11257_43940# a_10807_43548# a_11173_43940# VDD.t1257 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2540 VCM.t43 a_6123_31319.t7 C4_N_btm.t1 VSS.t2678 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2541 VSS.t1412 a_14084_46812# a_14035_46660# VSS.t1411 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2542 VDD.t3564 a_5937_45572.t8 a_8034_45724# VDD.t3563 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2543 a_5342_30871.t0 a_14456_42282# VDD.t2769 VDD.t2768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2544 a_17639_46660# a_12549_44172.t16 VSS.t2710 VSS.t2709 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X2545 a_10809_44734.t0 a_10057_43914# VDD.t310 VDD.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2546 VCM.t56 a_3422_30871.t18 VDAC_P.t5 VSS.t3519 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2547 VDD.t3626 a_11823_42460.t13 a_14853_42852# VDD.t3625 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2548 a_20749_43396# a_20974_43370# VSS.t452 VSS.t451 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2549 VDD.t3146 a_11967_42832.t44 a_16243_43396# VDD.t3145 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2550 a_19511_42282# a_n913_45002.t30 a_21125_42558# VDD.t2968 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2551 VSS.t1854 a_1431_47204# DATA[1].t5 VSS.t1853 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2552 a_1609_45572# a_n443_46116.t22 VSS.t3054 VSS.t3053 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2553 a_17517_44484.t1 a_16979_44734# VSS.t1428 VSS.t1427 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2554 a_20075_46420# a_19900_46494# a_20254_46482# VSS.t2045 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2555 a_n4209_37414.t1 a_n2302_37690# VDD.t1153 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2556 VDD.t915 a_10083_42826# a_7499_43078# VDD.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2557 a_16020_45572# a_15903_45785# VDD.t3506 VDD.t3505 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2558 VSS.t3204 VDD.t3781 VSS.t3203 VSS.t3202 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2559 a_20731_45938# a_20107_45572# a_20623_45572# VDD.t2475 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2560 a_22629_38406# a_22581_37893# CAL_N.t2 VDD.t3480 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2561 VDD.t3031 a_n3420_39072.t8 a_n2860_39072# VDD.t2023 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2562 VSS.t495 a_22731_47423# a_13717_47436.t1 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2563 a_16855_45546# a_16680_45572# a_17034_45572# VSS.t2560 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2564 a_18114_32519.t1 a_22223_45036# VDD.t1229 VDD.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2565 VDD.t616 a_15682_43940# a_11967_42832.t4 VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2566 a_17339_46660# a_12861_44030.t18 VSS.t2978 VSS.t2977 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2567 a_n2472_45546# a_n2293_45546.t4 VDD.t2022 VDD.t2021 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2568 VDD.t622 a_15682_43940# a_11967_42832.t5 VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2569 VSS.t1479 a_18429_43548# a_16823_43084# VSS.t1478 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2570 VSS.t2110 a_n4334_38304# a_n4064_37984.t5 VSS.t1340 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2571 VSS.t2338 a_8325_42308# a_8791_42308# VSS.t2337 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2572 VSS.t3137 VDD.t3818 VSS.t3136 VSS.t3135 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2573 VDD.t1554 a_n4334_38528# a_n4064_38528.t3 VDD.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2574 VSS.t3619 a_768_44030.t22 a_13076_44458# VSS.t3618 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2575 VSS.t2986 a_12861_44030.t24 a_19692_46634.t0 VSS.t2985 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2576 VDD.t2486 a_14495_45572# a_n881_46662.t0 VDD.t2485 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2577 a_18596_45572# a_18479_45785# VDD.t2786 VDD.t2785 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2578 a_n2472_45002# a_n2293_45010# VDD.t3489 VDD.t3488 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2579 VDD.t1792 a_n881_46662.t18 a_6431_45366# VDD.t1791 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2580 a_5326_44056# a_5147_45002# a_5244_44056# VDD.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2581 VSS.t3278 a_22959_42860# a_14097_32519.t3 VSS.t2180 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2582 a_3445_43172# a_3357_43084.t5 a_n2293_42282# VSS.t1798 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2583 a_13003_42852# a_10227_46804.t16 VDD.t1838 VDD.t1837 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2584 VSS.t1259 a_9127_43156# a_5891_43370.t7 VSS.t1258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2585 a_3503_45724# a_3775_45552# VSS.t580 VSS.t579 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2586 C6_N_btm.t2 a_14401_32519.t4 VREF_GND.t19 VSS.t1553 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2587 a_19929_45028# a_19778_44110# VDD.t868 VDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2588 a_3540_43646# a_584_46384.t16 VDD.t3003 VDD.t3002 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2589 VSS.t523 a_n2302_37984# a_n4209_38216.t6 VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2590 DATA[4].t4 a_9067_47204# VSS.t1014 VSS.t1013 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2591 VDD.t184 VSS.t3715 VDD.t183 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2592 VDD.t382 a_167_45260# a_117_45144# VDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2593 a_6086_46660# a_n1613_43370.t15 VSS.t3312 VSS.t3311 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2594 a_3147_46376# a_3483_46348.t6 VDD.t3283 VDD.t3282 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2595 a_n1533_46116# a_n1613_43370.t14 VDD.t3372 VDD.t3371 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2596 VSS.t3696 a_n3565_38216.t9 a_n3607_38304# VSS.t3022 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2597 VSS.t3189 VDD.t3776 VSS.t3188 VSS.t3187 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2598 a_5337_42558# a_5267_42460# a_4905_42826# VDD.t2793 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2599 a_21542_46660# a_10227_46804.t30 VSS.t1625 VSS.t1624 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2600 a_10216_45572# a_10180_45724# VSS.t2416 VSS.t2415 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2601 a_4699_43561# a_3080_42308.t5 VDD.t3429 VDD.t3428 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2602 a_3626_43646.t4 a_3232_43370.t22 a_3457_43396# VSS.t2831 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2603 a_n4064_37984.t4 a_n4334_38304# VSS.t2109 VSS.t1344 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2604 VDD.t2570 a_21613_42308# a_22775_42308# VDD.t2569 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2605 a_16269_42308# a_15890_42674# a_16197_42308# VSS.t2558 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2606 a_1067_42314# a_1184_42692# VSS.t2505 VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2607 VDD.t3561 a_5937_45572.t4 a_6945_45028.t0 VDD.t3560 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2608 COMP_P.t2 a_1169_39587# VDD.t1210 VDD.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2609 a_21356_42826# a_21381_43940# VDD.t2866 VDD.t2865 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2610 VDD.t3699 CLK.t5 a_8953_45002# VDD.t3698 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2611 VDD.t3225 a_2324_44458.t55 a_949_44458# VDD.t3224 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2612 a_4646_46812.t20 a_6298_44484# VSS.t839 VSS.t838 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2613 VDD.t3549 a_1307_43914.t9 a_16237_45028# VDD.t3548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS.t1390 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2615 VSS.t533 a_19862_44208# a_19808_44306# VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2616 VDD.t1814 a_5891_43370.t22 a_8791_43396# VDD.t1813 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2617 VSS.t190 a_n3690_39392# a_n3420_39072.t6 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2618 a_20256_43172# a_18494_42460# VSS.t1109 VSS.t1108 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2619 a_7927_46660# a_7411_46660# a_7832_46660# VSS.t905 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2620 VSS.t3165 VDD.t3768 VSS.t3164 VSS.t3163 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2621 VREF_GND.t33 a_13887_32519.t4 C3_N_btm.t1 VSS.t1802 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2622 a_n3420_39072.t1 a_n3690_39392# VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2623 a_n2472_45546# a_n2293_45546.t5 VSS.t1773 VSS.t1772 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2624 a_17668_45572# a_n881_46662.t7 a_17568_45572# VSS.t1557 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X2625 C9_P_btm.t1 a_n4064_39616.t9 VREF_GND.t1 VSS.t2845 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2626 a_4649_42852# a_1823_45246# VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2627 a_6540_46812# a_3877_44458# a_6682_46660# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2628 VDD.t2752 a_6511_45714# a_6472_45840# VDD.t2751 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2629 VSS.t3039 a_15493_43396.t2 a_19478_44306# VSS.t3038 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2630 a_16664_43396# a_16547_43609# VDD.t2324 VDD.t2323 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2631 VDD.t589 a_5068_46348# a_4955_46873# VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2632 a_9159_44484# a_5883_43914# VSS.t2023 VSS.t2022 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2633 C10_P_btm.t17 a_n4315_30879.t9 VREF.t35 VDD.t2069 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2634 VSS.t1574 a_10341_43396.t2 a_22591_43396# VSS.t1573 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2635 VDD.t1712 a_n4334_37440# a_n4064_37440.t3 VDD.t1711 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2636 VSS.t369 a_17124_42282# a_4958_30871.t3 VSS.t368 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS.t1378 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2638 C8_P_btm.t1 a_n3565_39590.t13 VREF.t69 VDD.t3614 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2639 a_5267_42460# a_4791_45118.t7 VDD.t2006 VDD.t2005 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2640 a_1138_42852# a_791_42968# VDD.t592 VDD.t591 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2641 a_n4318_40392.t0 a_n2840_44458# VDD.t2167 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2642 a_n1644_44306# a_n1761_44111# VSS.t2335 VSS.t2334 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2643 VDD.t3597 a_7754_40130.t12 VDD.t3596 VDD.t3595 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2644 VDD.t388 a_1609_45822# a_n2293_45546.t1 VDD.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2645 a_5267_42460# a_4791_45118.t6 VSS.t1753 VSS.t1752 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2646 VREF_GND.t22 a_17364_32525.t4 C7_N_btm.t4 VSS.t1715 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2647 VDD.t205 VSS.t3726 VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2648 a_2127_44172# a_2675_43914# a_2455_43940# VDD.t2801 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2649 a_11787_45002# a_11823_42460.t8 VDD.t3619 VDD.t3618 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2650 VSS.t841 a_6298_44484# a_4646_46812.t19 VSS.t840 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2651 VDD.t302 a_17499_43370# a_n1059_45260.t0 VDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2652 a_n1057_35014.t3 EN_VIN_BSTR_P.t7 VIN_P.t10 VSS.t3560 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2653 VSS.t1211 a_19333_46634# a_19123_46287# VSS.t1210 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2654 a_11599_46634.t12 a_15682_46116# VDD.t1068 VDD.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2655 a_n2946_37984# a_n2956_38216.t4 VSS.t1552 VSS.t1551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2656 a_3316_45546# a_3537_45260.t9 VDD.t2900 VDD.t2899 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X2657 VSS.t2463 a_13777_45326# a_13711_45394# VSS.t2462 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2658 a_20712_42282# a_n357_42282.t8 VDD.t2089 VDD.t2088 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2659 a_19479_31679.t3 a_22223_45572# VSS.t1230 VSS.t1027 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2660 a_20573_43172# a_20512_43084# a_20256_43172# VSS.t812 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X2661 VSS.t3177 VDD.t3772 VSS.t3176 VSS.t3175 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2662 a_n2293_46634.t0 a_14673_44172# VDD.t1390 VDD.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2663 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS.t2076 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2664 VSS.t3267 VDD.t3807 VSS.t3266 VSS.t3225 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2665 VSS.t3404 a_526_44458.t26 a_5457_43172# VSS.t3403 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2666 a_33_46660# a_n133_46660# VDD.t2209 VDD.t2208 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2667 a_584_46384.t1 a_1123_46634# VDD.t1470 VDD.t1469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 VSS.t902 a_15682_46116# a_11599_46634.t31 VSS.t901 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2669 VDD.t3307 a_10903_43370.t8 a_10849_43646# VDD.t3306 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2670 VDD.t3577 a_7754_40130.t0 a_7754_40130.t1 VDD.t3576 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2671 VSS.t878 a_15682_46116# a_11599_46634.t18 VSS.t877 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2672 a_8495_42852# a_7871_42858# a_8387_43230# VDD.t1677 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2673 VDD.t126 VSS.t3765 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2674 a_5495_43940# a_5244_44056# VSS.t956 VSS.t955 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2675 a_16842_45938# a_15765_45572# a_16680_45572# VDD.t2484 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2676 VDD.t386 a_167_45260# a_2521_46116# VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2677 VDD.t673 a_2779_44458# a_1307_43914.t2 VDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2678 VSS.t2310 a_n961_42308# a_n784_42308.t2 VSS.t2309 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2679 VSS.t73 a_13259_45724.t6 a_17303_42282# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2680 VDD.t3571 a_5937_45572.t17 a_5829_43940# VDD.t2436 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2681 a_17538_32519.t0 a_22959_43948# VDD.t1170 VDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2682 a_21496_47436# a_4883_46098.t2 VSS.t1629 VSS.t1628 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2683 a_11816_44260# a_11750_44172# a_10729_43914# VSS.t2490 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2684 a_9801_43940# a_8199_44636# VDD.t963 VDD.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2685 a_5742_30871.t1 a_10723_42308# VDD.t2414 VDD.t2413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2686 VDD.t1635 a_15051_42282# a_11823_42460.t2 VDD.t1634 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_2123_42473# a_n784_42308.t5 VDD.t3617 VDD.t3616 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2688 a_13565_43940# a_12891_46348# a_13483_43940# VDD.t1643 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2689 a_7227_42852# a_n97_42460.t6 a_7309_43172# VSS.t1669 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2690 a_5257_43370# a_5907_46634# VSS.t1289 VSS.t1288 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2691 VDD.t3089 a_13747_46662.t9 a_13607_46688# VDD.t3088 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2692 a_1667_45002# a_1823_45246# VSS.t248 VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2693 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2694 a_n2293_46098.t0 a_5663_43940# VDD.t2823 VDD.t2822 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2695 a_13003_42852# a_12379_42858# a_12895_43230# VDD.t1667 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2696 a_2711_45572.t3 a_768_44030.t24 VSS.t3621 VSS.t3620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2697 VDD.t171 VSS.t3763 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2698 DATA[0].t5 a_327_47204# VSS.t2060 VSS.t2059 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2699 a_16763_47508# a_16588_47582# a_16942_47570# VSS.t705 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2700 a_4883_46098.t1 a_21363_46634# VSS.t1302 VSS.t1301 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2701 VSS.t568 a_16751_45260# a_6171_45002.t1 VSS.t567 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2702 VDD.t1182 a_20835_44721# a_20766_44850# VDD.t1181 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2703 a_11750_44172# a_10903_43370.t7 VSS.t3093 VSS.t3092 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2704 VSS.t1314 a_15861_45028# a_17668_45572# VSS.t1313 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X2705 a_7845_44172# a_5891_43370.t24 VSS.t1579 VSS.t1578 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2706 a_15597_42852# a_15743_43084# VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2707 a_n4064_39072.t4 a_n4334_39392# VSS.t601 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2708 VSS.t3280 a_9223_42460# a_8953_45546# VSS.t3279 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X2709 VDD.t3135 a_11967_42832.t32 a_18083_42858# VDD.t3134 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2710 a_13487_47204# a_13381_47204# VSS.t605 VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X2711 a_13297_45572# a_13259_45724.t5 VSS.t79 VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X2712 C10_P_btm.t4 a_4190_30871.t20 VCM.t14 VSS.t2817 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2713 C2_N_btm.t1 EN_VIN_BSTR_N.t10 VIN_N.t11 VSS.t2917 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2714 w_10694_33990.t4 a_10890_34112.t7 w_10694_33990.t3 w_10694_33990.t2 sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X2715 C10_N_btm.t33 EN_VIN_BSTR_N.t15 VIN_N.t5 VSS.t2921 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2716 VDD.t3765 a_n3565_38216.t8 a_n3690_38304# VDD.t2956 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2717 a_6101_43172# a_5891_43370.t12 a_5755_42852# VSS.t1654 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2718 a_11901_46660# a_11735_46660# VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2719 a_16979_44734# a_14539_43914# a_17061_44734# VDD.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2720 VSS.t629 a_14955_47212# a_10227_46804.t3 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2721 VDD.t165 VSS.t3740 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2722 a_18443_44721# a_18248_44752# a_18753_44484# VSS.t1944 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2723 VDD.t1564 a_18909_45814# a_18799_45938# VDD.t1563 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2724 VSS.t295 a_8953_45002# a_2324_44458.t29 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2725 a_8912_37509.t28 VDAC_N.t20 a_5700_37509.t15 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2726 a_1431_46436# a_1138_42852# a_1337_46436# VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2727 VREF.t26 a_22612_30879.t18 C10_N_btm.t22 VDD.t1953 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2728 VDD.t3230 a_n4064_37984.t10 a_n2216_37984# VDD.t2027 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2729 a_11967_42832.t6 a_15682_43940# VDD.t608 VDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2730 a_18443_44721# a_18287_44626# a_18588_44850# VDD.t2655 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2731 VDD.t3683 a_768_44030.t12 a_5326_44056# VDD.t3682 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2732 VSS.t1720 a_n4209_39304.t9 a_n4251_39392# VSS.t1719 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2733 a_n357_42282.t2 a_21356_42826# VSS.t2532 VSS.t2531 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2734 VSS.t662 a_n2288_47178# a_n2312_40392.t2 VSS.t661 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2735 a_491_47026# a_n1613_43370.t46 VDD.t3402 VDD.t3401 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2736 a_n901_46420# a_n1613_43370.t42 VDD.t3396 VDD.t3395 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2737 VSS.t3076 a_3483_46348.t5 a_15301_44260# VSS.t3075 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2738 VCM.t19 a_1606_42308.t7 C1_N_btm.t3 VSS.t1731 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2739 VDD.t1727 a_20712_42282# a_10193_42453.t1 VDD.t1726 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2740 VSS.t2350 a_13635_43156# a_9290_44172.t6 VSS.t2349 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2741 a_5068_46348# a_5204_45822# a_5210_46482# VSS.t3417 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2742 a_14033_45822# a_10903_43370.t6 VDD.t3305 VDD.t3304 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2743 VSS.t2957 a_11599_46634.t43 a_20107_45572# VSS.t2956 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2744 a_3537_45260.t3 a_7287_43370# VDD.t858 VDD.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2745 VSS.t2501 a_6761_42308# a_7227_42308# VSS.t1507 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2746 VDD.t3125 a_13661_43548.t24 a_15595_45028# VDD.t3124 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2747 a_9803_42558# a_n97_42460.t5 a_9885_42558# VDD.t1895 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2748 VDD.t1846 a_10227_46804.t26 a_11136_42852# VDD.t1845 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 a_n1177_43370# a_n1613_43370.t30 VDD.t3382 VDD.t3381 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2750 VREF_GND.t28 a_n3420_39616.t10 C8_P_btm.t6 VSS.t2643 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2751 VDD.t2160 a_n2946_39072# a_n3565_39304.t2 VDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2752 a_601_46902# a_383_46660# VDD.t2256 VDD.t2255 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2753 a_5024_45822# a_n443_46116.t24 a_4419_46090# VDD.t3258 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2754 VDAC_Ni.t8 a_3754_38470.t9 a_3726_37500# VSS.t2638 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2755 a_17701_42308# a_17531_42308# VSS.t2122 VSS.t2121 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2756 VSS.t2976 a_12861_44030.t16 a_13487_47204# VSS.t2975 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X2757 a_4808_45572# a_1823_45246# a_4419_46090# VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2758 a_6598_45938# a_6472_45840# a_6194_45824# VSS.t287 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2759 a_n229_43646# a_n2497_47436# a_n447_43370# VDD.t2639 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2760 a_n3607_38304# a_n3674_38216.t5 a_n3690_38304# VSS.t1780 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2761 VSS.t380 a_6969_46634# a_6903_46660# VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2762 a_18214_42558# a_18184_42460.t7 VDD.t3736 VDD.t3735 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2763 a_491_47026# a_n133_46660# a_383_46660# VDD.t2210 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2764 VSS.t1635 a_4883_46098.t9 a_10355_46116# VSS.t1634 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2765 VDD.t3407 a_16327_47482.t12 a_18588_44850# VDD.t3406 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2766 VDD.t3098 a_4646_46812.t32 a_6031_43396# VDD.t3097 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2767 VSS.t3326 a_n1613_43370.t22 a_n1655_43396# VSS.t3325 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2768 a_6812_45938# a_6598_45938# VDD.t2734 VDD.t2733 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2769 a_8147_43396# a_n443_42852.t21 VDD.t3721 VDD.t3720 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2770 VDAC_Ni.t2 VSS.t3736 a_5088_37509.t18 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2771 a_12427_45724# a_12549_44172.t29 VDD.t2952 VDD.t2951 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X2772 C9_N_btm.t7 a_17730_32519.t7 VREF_GND.t9 VSS.t2882 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2773 VDD.t2664 a_19594_46812# a_19551_46910# VDD.t2663 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2774 a_n4318_37592.t2 a_n1736_42282# VSS.t717 VSS.t716 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2775 a_9290_44172.t0 a_13635_43156# VDD.t2601 VDD.t2600 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2776 VSS.t2571 a_2698_46116# a_2804_46116# VSS.t2570 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2777 VDD.t598 a_15682_43940# a_11967_42832.t8 VDD.t597 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2778 a_1414_42308# a_1067_42314# VDD.t787 VDD.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2779 w_1575_34786.t15 a_n1057_35014.t6 w_1575_34786.t15 w_1575_34786.t13 sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X2780 VSS.t1781 a_5649_42852.t2 a_22223_43396# VSS.t1231 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2781 VDD.t239 a_13259_45724.t20 a_14797_45144# VDD.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2782 a_n2288_47178# a_n2109_47186.t3 VDD.t3651 VDD.t3650 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2783 a_4817_46660# a_4651_46660# VDD.t2468 VDD.t2467 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2784 a_8062_46155# a_8016_46348# VDD.t1142 VDD.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2785 a_949_44458# a_2324_44458.t43 VDD.t3215 VDD.t3214 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2786 a_13296_44484# a_12891_46348# VSS.t1435 VSS.t1434 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2787 VDD.t2188 a_20623_43914# a_20365_43914# VDD.t2187 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2788 a_11601_46155# a_11309_47204# a_11387_46155# VDD.t2714 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2789 a_10210_45822# a_8746_45002# VDD.t532 VDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2790 a_18287_44626# a_11967_42832.t34 VSS.t2929 VSS.t2928 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2791 a_8912_37509.t24 VDAC_N.t16 a_5700_37509.t16 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2792 VSS.t2455 a_11189_46129# a_11133_46155# VSS.t2454 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2793 a_n3565_38216.t1 a_n2946_37984# VDD.t1615 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2794 a_6431_45366# a_5937_45572.t14 VDD.t3570 VDD.t3569 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2795 a_6109_44484# a_5518_44484# VSS.t2195 VSS.t2194 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2796 a_14021_43940.t1 a_13483_43940# VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2797 a_17499_43370# a_17324_43396# a_17678_43396# VSS.t2398 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2798 a_3495_45348# a_3429_45260# a_3316_45546# VSS.t1359 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X2799 VDD.t2495 a_1115_44172# a_n2293_45010# VDD.t2494 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2800 VDD.t2796 a_19787_47423# a_19594_46812# VDD.t2795 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2801 a_18707_42852# a_16327_47482.t42 VDD.t3356 VDD.t3355 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2802 a_19787_47423# START.t0 VDD.t2874 VDD.t2873 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2803 a_8667_46634# a_8492_46660# a_8846_46660# VSS.t1895 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2804 a_1208_46090# a_n881_46662.t23 a_1431_46436# VSS.t1572 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2805 a_5431_46482# a_n1151_42308.t5 a_5068_46348# VSS.t1656 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2806 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD.t1317 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2807 a_n2302_39866# a_n2442_46660.t5 VSS.t2884 VSS.t2883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2808 VSS.t3668 a_n2438_43548.t32 a_2443_46660# VSS.t3667 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2809 a_18797_44260# a_13661_43548.t20 a_18451_43940# VSS.t2902 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2810 a_19551_46910# a_19692_46634.t11 VDD.t2067 VDD.t2066 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2811 VDD.t2623 a_8953_45546# a_8049_45260.t0 VDD.t2622 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2812 a_8697_45822# a_3483_46348.t20 VDD.t3299 VDD.t3298 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2813 VDD.t1802 a_10341_43396.t3 a_22591_43396# VDD.t1801 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2814 a_12005_46116# a_2063_45854.t8 VDD.t1870 VDD.t1869 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2815 VSS.t2992 a_12861_44030.t30 a_18911_45144# VSS.t2991 sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2816 a_1241_43940# a_584_46384.t20 VDD.t3007 VDD.t3006 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X2817 VSS.t2591 a_2123_42473# a_1184_42692# VSS.t2590 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2818 a_1273_38525.t5 a_1107_38525# VSS.t2434 VSS.t2389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2819 a_16285_47570# a_16241_47178# a_16119_47582# VSS.t2018 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2820 a_4646_46812.t17 a_6298_44484# VSS.t833 VSS.t832 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2821 a_1423_45028.t2 a_167_45260# VSS.t209 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2822 VDD.t480 a_8953_45002# a_2324_44458.t4 VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2823 VDD.t16 a_949_44458# a_n2438_43548.t12 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2824 a_10617_44484# a_10440_44484# VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2825 C7_P_btm.t0 a_n4064_39072.t9 VREF_GND.t42 VSS.t2859 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2826 VSS.t182 a_1169_39043# comp_n VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2827 VSS.t602 a_961_42354# a_1067_42314# VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2828 VDD.t1335 a_4704_46090# a_1823_45246# VDD.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2829 a_18479_47436# a_20075_46420# VSS.t591 VSS.t590 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2830 a_4646_46812.t31 a_6298_44484# VSS.t821 VSS.t820 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2831 VDD.t2518 a_9313_45822# a_11459_47204# VDD.t2517 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2832 a_n1809_44850# a_n1613_43370.t9 VDD.t3366 VDD.t3365 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2833 VSS.t194 a_n3690_39392# a_n3420_39072.t5 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2834 a_19987_42826# a_10193_42453.t16 a_20573_43172# VSS.t2793 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2835 VSS.t1408 a_3785_47178# a_3815_47204# VSS.t1407 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2836 VDD.t1879 a_5891_43370.t14 a_8375_44464# VDD.t1878 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2837 a_n3420_39072.t0 a_n3690_39392# VDD.t366 VDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2838 VSS.t2266 a_9863_46634# a_2063_45854.t2 VSS.t2265 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X2839 a_7920_46348# a_n1151_42308.t16 a_8062_46155# VDD.t1885 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2840 VDD.t2283 a_22889_38993# a_22581_37893# VDD.t2282 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2841 a_19721_31679.t0 a_22959_45036# VDD.t577 VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2842 a_19808_44306# a_19778_44110# a_19328_44172# VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2843 VDD.t3012 a_10193_42453.t4 a_11633_42558# VDD.t3011 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2844 VDD.t1186 a_15559_46634# a_13059_46348# VDD.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2845 VDD.t2707 a_11189_46129# a_11601_46155# VDD.t2706 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2846 a_5263_45724# a_5257_43370# a_5437_45600# VSS.t1297 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2847 a_12495_44260# a_12429_44172# a_10949_43914# VSS.t858 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X2848 VSS.t115 a_n2840_43370# a_n4318_39304.t3 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2849 a_15037_43396# a_14205_43396# a_14955_43396# VSS.t2512 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2850 VSS.t3682 a_4915_47217.t3 a_12891_46348# VSS.t3681 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 a_14084_46812# a_13885_46660# a_14226_46660# VSS.t2281 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2852 a_6452_43396# a_6293_42852# VDD.t1491 VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2853 VSS.t2431 a_1107_38525# a_1273_38525.t4 VSS.t2430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2854 a_7705_45326# a_7229_43940# VSS.t2080 VSS.t2079 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2855 a_8953_45002# CLK.t6 VSS.t3631 VSS.t3630 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2856 a_16981_45144# a_16922_45042# a_16886_45144# VDD.t2853 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2857 a_1115_44172# a_1307_43914.t22 a_1241_44260# VSS.t3464 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2858 a_19478_44306# a_3090_45724.t10 VSS.t1591 VSS.t1590 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2859 a_11599_46634.t23 a_15682_46116# VSS.t882 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2860 a_4223_44672.t0 a_3537_45260.t18 VDD.t2910 VDD.t2909 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2861 a_7174_31319.t1 a_20107_42308# VDD.t2220 VDD.t2219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2862 VCM.t15 a_4190_30871.t6 C10_P_btm.t5 VSS.t2803 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2863 VDD.t1047 a_n2302_39866# a_n4209_39590.t2 VDD.t1046 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2864 VDD.t1832 a_10227_46804.t8 a_15051_42282# VDD.t1831 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2865 CLK_DATA.t1 a_n2833_47464# VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2866 a_8912_37509.t20 VDAC_N.t12 a_5700_37509.t8 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2867 a_n2833_47464# a_n2497_47436# VSS.t2392 VSS.t2391 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2868 VSS.t1 a_8103_44636# a_7640_43914# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2869 a_15146_44811# a_9482_43914# VDD.t1293 VDD.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2870 a_n4209_39304.t0 a_n2302_39072# VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2871 a_2903_45348# a_n971_45724.t4 a_2809_45348# VSS.t1681 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2872 VSS.t2668 a_3537_45260.t16 a_8103_44636# VSS.t2667 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2873 VSS.t1538 a_21137_46414# a_21071_46482# VSS.t1537 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2874 a_2324_44458.t6 a_8953_45002# VDD.t506 VDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2875 VSS.t473 a_1414_42308# a_2889_44172# VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2876 VDD.t1386 a_1848_45724# a_1799_45572# VDD.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2877 VSS.t2523 a_19279_43940# a_21398_44850# VSS.t2522 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2878 a_1666_39587.t2 a_1273_38525.t11 VDD.t2058 VDD.t2054 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2879 VSS.t400 a_n13_43084# a_n1853_43023# VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2880 a_18479_45785# a_19268_43646# VSS.t215 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2881 VSS.t3122 VDD.t3813 VSS.t3121 VSS.t3120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2882 VSS.t448 a_22485_44484# a_20974_43370# VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2883 VSS.t2630 a_n3420_37984.t8 a_n2946_37984# VSS.t1776 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2884 a_5275_47026# a_n1613_43370.t12 VDD.t3368 VDD.t3367 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2885 a_5841_44260# a_5495_43940# VSS.t2537 VSS.t2536 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2886 C5_N_btm.t0 EN_VIN_BSTR_N.t9 VIN_N.t9 VSS.t2916 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2887 a_n2661_45546.t0 a_4093_43548# VDD.t1426 VDD.t1425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2888 VSS.t2400 a_n2302_38778# a_n4209_38502.t6 VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2889 VSS.t2474 a_5497_46414# a_5431_46482# VSS.t2473 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2890 VSS.t424 a_15682_43940# a_11967_42832.t20 VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2891 VDD.t2137 a_19339_43156# a_19326_42852# VDD.t2136 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2892 VSS.t892 a_15682_46116# a_11599_46634.t30 VSS.t891 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2893 a_8137_45348# a_8049_45260.t6 a_n2293_42834.t1 VSS.t2878 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2894 VDD.t298 a_17499_43370# a_n1059_45260.t1 VDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2895 VDD.t3234 a_6123_31319.t5 a_7963_42308# VDD.t3233 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2896 VDD.t3181 a_12861_44030.t14 a_17339_46660# VDD.t3180 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2897 a_10849_43646# a_10807_43548# a_10765_43646# VDD.t1258 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2898 VSS.t1751 a_13507_46334.t13 a_18997_42308# VSS.t1750 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2899 a_8560_45348# a_3483_46348.t14 a_8488_45348# VSS.t3082 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2900 VDD.t1378 a_n3690_38304# a_n3420_37984.t2 VDD.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2901 a_13249_42308# a_13070_42354# a_13333_42558# VDD.t1271 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2902 a_6969_46634# a_n971_45724.t26 VSS.t1700 VSS.t1699 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2903 a_n2216_37984# a_n2810_45572.t5 a_n2302_37984# VDD.t1761 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2904 VSS.t1132 a_22223_46124# a_20205_31679.t2 VSS.t1131 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2905 a_6194_45824# a_6511_45714# a_6469_45572# VSS.t2493 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2906 a_17613_45144# a_8696_44636.t8 VDD.t1961 VDD.t1960 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2907 a_n229_43646# a_n97_42460.t20 VDD.t1903 VDD.t1902 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2908 VSS.t3328 a_n1613_43370.t24 a_n1379_43218# VSS.t3327 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2909 VDD.t1005 a_6298_44484# a_4646_46812.t15 VDD.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2910 VSS.t2868 a_13747_46662.t11 a_19862_44208# VSS.t2867 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2911 a_17303_42282# a_n913_45002.t16 VSS.t2731 VSS.t2730 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2912 a_8649_43218# a_8605_42826# a_8483_43230# VSS.t1994 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2913 VSS.t2203 a_n901_46420# a_n967_46494# VSS.t2202 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2914 a_15004_44636# a_13556_45296# a_15146_44811# VDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2915 a_11186_47026# a_10467_46802# a_10623_46897# VSS.t529 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2916 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD.t1589 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2917 VSS.t3393 a_526_44458.t12 a_4169_42308# VSS.t3392 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2918 a_n23_45546# a_n356_45724# VDD.t3511 VDD.t3510 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2919 a_3353_43940# a_2998_44172# a_2675_43914# VDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2920 a_11967_42832.t19 a_15682_43940# VSS.t428 VSS.t427 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2921 a_18326_43940# a_18079_43940# VSS.t570 VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2922 a_20922_43172# a_19862_44208# a_20753_42852# VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X2923 a_10334_44484# a_10157_44484# VSS.t1951 VSS.t1950 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2924 VSS.t791 a_742_44458# a_1756_43548# VSS.t790 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2925 C5_P_btm.t1 a_5934_30871.t6 VCM.t63 VSS.t1786 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2926 a_n2017_45002.t3 a_19987_42826# VSS.t231 VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X2927 a_n2956_38216.t1 a_n2472_45546# VDD.t2525 VDD.t1732 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2928 VDD.t3018 a_10193_42453.t8 a_13657_42558# VDD.t3017 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2929 a_13885_46660# a_13607_46688# VDD.t2528 VDD.t2527 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2930 VDD.t2831 a_8191_45002# a_n2293_42834.t2 VDD.t2830 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2931 VSS.t1547 RST_Z.t3 a_7754_39964# VSS.t1546 sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X2932 VSS.t2661 a_4223_44672.t9 a_n2497_47436# VSS.t2660 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2933 a_n217_35014# VDD.t3805 EN_VIN_BSTR_P.t1 VSS.t3263 sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X2934 VDD.t156 VSS.t3749 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2935 a_4699_43561# a_3080_42308.t4 VSS.t3373 VSS.t3372 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2936 a_19511_42282# a_18597_46090# VSS.t1195 VSS.t1194 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2937 a_n1991_46122# a_n2157_46122# VDD.t1587 VDD.t1586 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2938 a_n3420_37984.t4 a_n3690_38304# VSS.t1182 VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2939 VSS.t1814 a_19692_46634.t9 a_743_42282.t3 VSS.t1813 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2940 VDD.t2533 a_22591_43396# a_14209_32519.t1 VDD.t2532 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2941 VDD.t512 a_7499_43078# a_8746_45002# VDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2942 a_n971_45724.t2 a_104_43370# VSS.t930 VSS.t929 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2943 a_22889_38993# a_22400_42852# VDD.t1609 VDD.t1608 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2944 VDD.t780 a_n4334_39392# a_n4064_39072.t1 VDD.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2945 a_20447_31679.t2 a_22959_45572# VSS.t293 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2946 VDD.t1166 a_15493_43940# a_22959_43948# VDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2947 VREF.t38 a_n4315_30879.t12 C10_P_btm.t20 VDD.t2072 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2948 VSS.t962 a_n2302_37690# a_n4209_37414.t5 VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2949 a_18147_46436# a_17339_46660# a_17957_46116# VSS.t1484 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2950 a_8336_45822# a_8270_45546# a_n1925_46634.t0 VDD.t755 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2951 VDD.t1746 a_13527_45546# a_13163_45724# VDD.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X2952 a_n4334_39616# a_n4318_39768.t4 VDD.t1890 VDD.t1889 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2953 a_n2956_39304.t0 a_n2840_46090# VDD.t1406 VDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2954 a_4646_46812.t0 a_6298_44484# VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2955 VDD.t2998 a_584_46384.t9 a_766_43646# VDD.t2997 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2956 w_10694_33990.t13 a_18194_34908.t13 EN_VIN_BSTR_N.t4 w_10694_33990.t12 sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2957 a_11361_45348# a_10907_45822# VSS.t1209 VSS.t1208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2958 VDD.t3160 a_11599_46634.t40 a_11735_46660# VDD.t3159 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2959 a_19431_45546# a_19256_45572# a_19610_45572# VSS.t2371 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2960 VSS.t3069 a_9290_44172.t23 a_12710_44260# VSS.t3068 sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X2961 VDD.t2539 a_11323_42473# a_10807_43548# VDD.t2538 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2962 a_2266_47243# a_n971_45724.t22 VDD.t1924 VDD.t1923 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2963 C10_P_btm.t28 a_n4315_30879.t22 VREF.t46 VDD.t2082 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2964 a_2982_43646.t4 a_2479_44172# a_2896_43646# VDD.t2140 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2965 a_18280_46660# a_12861_44030.t9 VSS.t2969 VSS.t2968 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2966 VDD.t2158 a_8492_46660# a_8667_46634# VDD.t2157 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2967 C1_P_btm.t0 EN_VIN_BSTR_P.t21 VIN_P.t11 VSS.t3569 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2968 VREF_GND.t35 a_n4064_40160.t9 C10_P_btm.t9 VSS.t2682 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2969 VDD.t1456 a_n1076_46494# a_n901_46420# VDD.t1455 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2970 a_n4251_38528# a_n4318_38680.t5 a_n4334_38528# VSS.t1795 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2971 a_4361_42308.t0 a_3823_42558# VDD.t1442 VDD.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2972 VDD.t3139 a_11967_42832.t38 a_12379_42858# VDD.t3138 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2973 VDD.t1053 a_21811_47423# a_20916_46384# VDD.t1052 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2974 VDD.t3158 a_11599_46634.t37 a_13759_46122# VDD.t3157 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2975 a_18985_46122# a_18819_46122# VSS.t2211 VSS.t2210 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2976 VDD.t1916 a_n971_45724.t12 a_3775_45552# VDD.t1915 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2977 VDD.t2030 a_5649_42852.t3 a_22223_43396# VDD.t2029 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2978 VSS.t1058 a_5343_44458# a_8333_44056# VSS.t1057 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2979 VDD.t862 a_7287_43370# a_3537_45260.t1 VDD.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2980 VSS.t3113 VDD.t3810 VSS.t3112 VSS.t3111 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2981 VSS.t1585 a_3090_45724.t7 a_10555_44260# VSS.t1584 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X2982 a_20528_45572# a_19466_46812# VSS.t693 VSS.t692 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2983 a_13487_47204# a_13717_47436.t3 VSS.t2629 VSS.t2628 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2984 VREF_GND.t18 a_13678_32519.t4 C2_N_btm.t2 VSS.t1539 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2985 VDD.t1246 a_22485_38105# a_22581_37893# VDD.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2986 VDD.t3340 a_20269_44172# a_19319_43548# VDD.t3339 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2987 a_5807_45002# a_16763_47508# VSS.t709 VSS.t708 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X2988 VSS.t3302 a_16327_47482.t38 a_16285_47570# VSS.t3301 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2989 a_n23_44458# a_n356_44636.t5 VSS.t3583 VSS.t3582 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2990 VDD.t2987 a_n1059_45260.t14 a_8791_43396# VDD.t2986 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2991 a_1847_42826# a_2351_42308# VDD.t1696 VDD.t1695 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2992 VSS.t3246 VDD.t3798 VSS.t3245 VSS.t3244 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2993 VDD.t612 a_15682_43940# a_11967_42832.t13 VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2994 VSS.t1007 a_1169_39587# COMP_P.t6 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2995 a_19553_46090# a_19335_46494# VDD.t2121 VDD.t2120 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2996 VDD.t2568 a_n2840_45546# a_n2810_45572.t1 VDD.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2997 VSS.t582 a_3503_45724# a_3218_45724# VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2998 a_15037_45618# a_13259_45724.t14 VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2999 a_14537_43646# a_13059_46348# VDD.t1361 VDD.t1360 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3000 VDD.t3532 a_1307_43914.t26 a_n913_45002.t6 VDD.t3531 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3001 a_6671_43940# a_5205_44484# VDD.t3344 VDD.t3343 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3002 a_n1699_43638# a_n1917_43396# VDD.t2422 VDD.t2421 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3003 C6_P_btm.t0 a_n3420_39072.t10 VREF_GND.t4 VSS.t1844 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3004 VDD.t881 a_n2946_38778# a_n3565_38502.t3 VDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3005 VSS.t918 a_5111_44636# a_4905_42826# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3006 VDD.t2035 a_9313_44734.t3 a_22959_42860# VDD.t2034 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3007 a_2124_47436# a_2063_45854.t10 a_2266_47243# VDD.t1871 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3008 VSS.t1494 a_9625_46129# a_9569_46155# VSS.t1493 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3009 a_n4064_37984.t2 a_n4334_38304# VDD.t2360 VDD.t1705 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3010 a_n2438_43548.t13 a_949_44458# VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3011 VDD.t2782 a_19279_43940# a_21398_44850# VDD.t2781 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3012 VDD.t3295 a_3483_46348.t18 a_13565_43940# VDD.t3294 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3013 a_22725_38406# a_22589_40055# a_22629_38406# VDD.t935 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3014 a_6171_42473# a_5932_42308.t7 VSS.t1804 VSS.t1055 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3015 a_17568_45572# a_8696_44636.t3 a_17478_45572# VSS.t1710 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3016 a_18588_44850# a_18374_44850# VDD.t2202 VDD.t2201 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3017 a_18451_43940# a_18579_44172# a_18533_43940# VDD.t2678 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3018 a_22485_38105# a_22775_42308# VSS.t1040 VSS.t1039 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3019 VSS.t2598 a_5755_42308# a_5932_42308.t3 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3020 a_2959_46660# a_2609_46660# a_2864_46660# VDD.t1684 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3021 a_21359_45002# a_21513_45002# VSS.t3290 VSS.t3289 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3022 a_7_47243# a_n746_45260# a_n452_47436# VDD.t1252 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3023 a_15227_46910# a_3090_45724.t18 a_15009_46634# VDD.t1822 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3024 a_14493_46090# a_14275_46494# VSS.t811 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3025 a_19478_44306# a_15493_43396.t3 a_19478_44056# VDD.t3244 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X3026 a_7287_43370# a_7112_43396# a_7466_43396# VSS.t990 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3027 a_12251_46660# a_11901_46660# a_12156_46660# VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3028 a_8495_42852# a_n1613_43370.t40 VDD.t3392 VDD.t3391 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3029 a_n4251_37440# a_n4318_37592.t5 a_n4334_37440# VSS.t3635 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3030 a_11633_42558# a_11823_42460.t24 VDD.t3635 VDD.t3634 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3031 VDD.t3494 a_7276_45260# a_7227_45028# VDD.t3493 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3032 VSS.t1876 a_2479_44172# a_2813_43396# VSS.t1875 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3033 a_15279_43071# a_5342_30871.t8 VDD.t2885 VDD.t2884 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3034 VREF_GND.t20 a_14401_32519.t5 C6_N_btm.t3 VSS.t1554 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3035 VREF.t4 a_21588_30879.t4 C9_N_btm.t9 VDD.t1773 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3036 VDD.t3496 a_n815_47178# a_n785_47204# VDD.t3495 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3037 VDD.t142 VSS.t3754 VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3038 a_1239_47204# a_1209_47178# VSS.t2100 VSS.t2099 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3039 VSS.t3265 VDD.t3806 VSS.t3264 VSS.t3120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3040 VDD.t320 a_3877_44458# a_3699_46348# VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3041 a_9313_45822# a_5937_45572.t6 a_9241_45822# VDD.t3562 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3042 a_20841_45814# a_20623_45572# VSS.t2227 VSS.t2226 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3043 VDD.t1422 a_805_46414# a_835_46155# VDD.t1421 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3044 a_12379_46436# a_12005_46116# a_n1741_47186.t4 VSS.t2113 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3045 VDD.t508 a_8953_45002# a_2324_44458.t14 VDD.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3046 a_6298_44484# a_2324_44458.t42 VSS.t3003 VSS.t3002 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3047 a_4338_37500.t2 a_3754_38470.t10 VDAC_Pi.t4 VSS.t2639 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3048 a_961_42354# a_n1059_45260.t10 VSS.t2760 VSS.t2759 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3049 a_n2956_39768.t2 a_n2840_46634# VSS.t936 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3050 a_n1741_47186.t6 a_12594_46348# VDD.t3502 VDD.t3501 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3051 VDD.t1508 a_5257_43370# a_3905_42865# VDD.t1507 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3052 VSS.t2390 en_comp a_1107_38525# VSS.t2389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3053 VSS.t1249 a_n473_42460# a_n1761_44111# VSS.t1248 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3054 a_13163_45724# a_12549_44172.t19 VDD.t2942 VDD.t2941 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X3055 VDD.t1828 a_10227_46804.t5 a_9863_46634# VDD.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3056 a_10210_45822# a_10586_45546# a_10053_45546# VDD.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3057 comp_n a_1169_39043# VSS.t178 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3058 VSS.t1666 a_4185_45028.t5 a_22959_45036# VSS.t1665 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3059 a_22485_38105# a_22775_42308# VDD.t1241 VDD.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3060 VDD.t3746 a_n2438_43548.t42 a_n2065_43946# VDD.t3745 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3061 VDD.t118 VSS.t3712 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3062 VSS.t2153 a_n2002_35448# SMPL_ON_P.t4 VSS.t2152 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3063 a_5457_43172# a_5111_44636# a_5111_42852# VSS.t910 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3064 VDD.t2615 a_11787_45002# a_11652_45724# VDD.t2614 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3065 a_10695_43548# a_7499_43078# VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3066 VDD.t3056 a_n1794_35082.t5 a_n1696_34930.t3 VDD.t3055 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3067 VDD.t280 a_n2946_37690# a_n3565_37414.t3 VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3068 a_13059_46348# a_15559_46634# VDD.t1188 VDD.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3069 VDD.t2736 a_n23_44458# a_7_44811# VDD.t2735 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3070 a_12891_46348# a_4915_47217.t8 VSS.t3685 VSS.t3684 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3071 a_8023_46660# a_7577_46660# a_7927_46660# VSS.t1506 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3072 VSS.t137 a_10057_43914# a_9672_43914# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3073 a_n237_47217.t2 a_8667_46634# VSS.t727 VSS.t726 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X3074 a_n143_45144# a_n755_45592.t22 VSS.t3385 VSS.t3384 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3075 a_20637_44484# a_20159_44458# VSS.t2423 VSS.t2422 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3076 a_4520_42826# a_4905_42826# a_4649_42852# VDD.t1555 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3077 VSS.t1693 a_n971_45724.t18 a_8423_43396# VSS.t1692 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X3078 VSS.t1549 RST_Z.t4 a_8530_39574# VSS.t1548 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3079 VSS.t1403 a_n2946_37984# a_n3565_38216.t5 VSS.t703 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3080 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS.t1127 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3081 a_8697_45822# a_8199_44636# VDD.t959 VDD.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3082 a_8912_37509.t12 VDAC_P.t13 a_5088_37509.t7 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3083 VDD.t340 a_n4334_39616# a_n4064_39616.t2 VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3084 VSS.t3489 a_3626_43646.t7 a_19647_42308# VSS.t3488 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3085 a_n443_42852.t0 a_n901_43156# VDD.t817 VDD.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3086 VDD.t2355 a_1209_47178# a_1239_47204# VDD.t2354 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3087 a_3094_47243# a_2905_45572# VDD.t2609 VDD.t2608 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3088 a_15051_42282# a_15486_42560# VDD.t2482 VDD.t2481 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3089 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS.t1374 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3090 VDD.t3106 a_13661_43548.t5 a_16241_44734# VDD.t3105 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3091 a_11823_42460.t7 a_15051_42282# VSS.t1420 VSS.t1419 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3092 a_5167_46660# a_4817_46660# a_5072_46660# VDD.t1220 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3093 VSS.t2448 a_10835_43094# a_10796_42968# VSS.t2447 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3094 VDD.t2490 a_20708_46348# a_20411_46873# VDD.t2489 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3095 VSS.t3352 a_16327_47482.t9 a_18005_44484# VSS.t3351 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3096 VSS.t1373 a_16292_46812# a_15811_47375# VSS.t1372 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3097 a_2324_44458.t11 a_8953_45002# VDD.t478 VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3098 a_9482_43914# a_9838_44484# VSS.t1443 VSS.t1442 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3099 a_20623_46660# a_20273_46660# a_20528_46660# VDD.t1350 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3100 VDD.t3504 a_12594_46348# a_n1741_47186.t7 VDD.t3503 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3101 a_18374_44850# a_18287_44626# a_17970_44736# VDD.t2658 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3102 a_16750_47204# a_15673_47210# a_16588_47582# VDD.t2245 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3103 a_6545_47178# a_6419_46155# VSS.t2131 VSS.t2130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3104 a_8783_44734# a_8696_44636.t7 a_8701_44490# VDD.t1959 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3105 a_175_44278# a_n863_45724# VDD.t691 VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3106 VDD.t1611 a_22400_42852# a_22589_40055# VDD.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3107 VDD.t1562 a_22223_43396# a_13887_32519.t0 VDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3108 VSS.t3224 VDD.t3790 VSS.t3223 VSS.t3222 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3109 VSS.t2207 a_n901_46420# a_n443_46116.t7 VSS.t2206 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3110 VDD.t1599 a_18479_47436# a_20935_43940# VDD.t1598 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3111 VSS.t1927 a_7754_38470# VSS.t1926 VSS.t1925 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3112 VSS.t1287 a_5907_46634# a_5841_46660# VSS.t1286 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3113 a_5745_43940# a_5883_43914# a_5829_43940# VDD.t2280 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3114 a_3754_38470.t2 a_7754_38470# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X3115 a_1110_47026# a_33_46660# a_948_46660# VDD.t2728 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3116 a_16434_46987# a_16388_46812# VDD.t657 VDD.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3117 VSS.t3011 a_2324_44458.t51 a_15682_43940# VSS.t3010 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3118 VDD.t1051 a_n2302_39866# a_n4209_39590.t1 VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3119 a_13381_47204# a_12549_44172.t12 VSS.t2706 VSS.t2705 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3120 a_2324_44458.t15 a_8953_45002# VDD.t498 VDD.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3121 a_2998_44172# a_584_46384.t14 VSS.t2779 VSS.t2778 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3122 a_20974_43370# a_22485_44484# VSS.t446 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3123 VDD.t1718 a_4921_42308# a_5755_42308# VDD.t1717 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3124 a_10991_42826# a_10835_43094# a_11136_42852# VDD.t2696 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3125 VDD.t2241 a_6851_47204# a_7227_47204# VDD.t2240 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3126 a_3052_44056# a_2998_44172# VDD.t1305 VDD.t1304 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X3127 VSS.t1341 a_n4334_38528# a_n4064_38528.t4 VSS.t1340 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3128 a_3177_46902# a_2959_46660# VSS.t2525 VSS.t2524 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3129 VSS.t2221 a_1208_46090# a_472_46348# VSS.t2220 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3130 a_9241_44734# a_5937_45572.t13 VDD.t3568 VDD.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3131 a_n1699_43638# a_n1917_43396# VSS.t2170 VSS.t2169 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3132 a_22365_46825# EN_OFFSET_CAL.t0 VDD.t2870 VDD.t2869 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3133 VSS.t880 a_15682_46116# a_11599_46634.t20 VSS.t879 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3134 VSS.t460 a_13163_45724# a_11962_45724# VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3135 a_3055_46660# a_2609_46660# a_2959_46660# VSS.t1475 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3136 a_19326_42852# a_18249_42858# a_19164_43230# VDD.t1121 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3137 a_n443_46116.t4 a_n901_46420# VSS.t2201 VSS.t2200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3138 a_9885_43646# a_8270_45546# a_9803_43646# VDD.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3139 VDD.t1394 a_18597_46090# a_16375_45002# VDD.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3140 a_19431_45546# a_16327_47482.t22 VDD.t3417 VDD.t3416 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3141 VSS.t2181 a_22959_43396# a_17364_32525.t2 VSS.t2180 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3142 w_10694_33990.t8 a_10890_34112.t5 w_10694_33990.t8 w_10694_33990.t7 sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X3143 VDD.t1382 a_n3690_38304# a_n3420_37984.t1 VDD.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3144 a_n4064_39616.t1 a_n4334_39616# VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3145 VSS.t985 a_n1177_44458# a_n1243_44484# VSS.t984 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3146 VREF.t48 a_n4315_30879.t24 C10_P_btm.t30 VDD.t2084 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3147 VSS.t2619 a_n23_45546# a_n89_45572# VSS.t2618 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3148 a_n452_47436# a_n746_45260# a_n310_47570# VSS.t1047 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3149 a_2952_47436# a_n1151_42308.t12 a_3094_47243# VDD.t1884 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3150 VDD.t3485 a_12816_46660# a_12991_46634# VDD.t3484 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3151 VDD.t1029 a_6298_44484# a_4646_46812.t13 VDD.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3152 a_7499_43940# a_7640_43914# VDD.t2146 VDD.t2145 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3153 VSS.t2402 a_n2302_38778# a_n4209_38502.t7 VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3154 a_4235_43370# a_3935_42891# VDD.t2308 VDD.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X3155 a_5105_45348# a_4558_45348# VSS.t2004 VSS.t2003 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3156 a_18051_46116# a_765_45546.t9 a_17957_46116# VDD.t3764 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X3157 a_n1441_43940# a_n1613_43370.t38 VDD.t3390 VDD.t3389 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3158 a_15301_44260# a_15227_44166.t20 a_14955_43940# VSS.t3598 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3159 a_n746_45260# a_n1177_44458# VSS.t983 VSS.t982 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3160 VSS.t3023 a_n3565_38502.t9 a_n3607_38528# VSS.t3022 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3161 a_n2840_43914# a_n2661_43922.t4 VSS.t1543 VSS.t1542 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3162 a_6809_43396# a_6765_43638# a_6643_43396# VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3163 VSS.t176 a_376_46348# a_171_46873# VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3164 a_19443_46116# a_16327_47482.t24 VDD.t3419 VDD.t3418 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3165 VSS.t1166 a_13059_46348# a_15143_45578# VSS.t1165 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3166 VSS.t782 a_8199_44636# a_8701_44490# VSS.t781 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3167 a_7499_43940# a_3090_45724.t14 a_7281_43914# VDD.t1818 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3168 a_9165_43940# a_9290_44172.t17 VDD.t3268 VDD.t3267 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3169 a_453_43940# a_175_44278# VDD.t3519 VDD.t3518 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3170 a_9885_42308# a_7499_43078# VSS.t338 VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3171 a_n3674_39304.t2 a_n2840_42826# VSS.t1156 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3172 a_2959_46660# a_2443_46660# a_2864_46660# VSS.t2541 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3173 a_14543_46987# a_13885_46660# a_14084_46812# VDD.t2529 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3174 VDD.t2105 a_413_45260.t3 a_22959_44484# VDD.t1891 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3175 a_17969_45144# a_16375_45002# a_17896_45144# VDD.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X3176 a_n4064_38528.t5 a_n4334_38528# VSS.t1345 VSS.t1344 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3177 a_16292_46812# a_n743_46660.t8 a_16434_46987# VDD.t3642 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3178 a_21188_46660# a_20107_46660# a_20841_46902# VDD.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3179 a_12251_46660# a_11735_46660# a_12156_46660# VSS.t458 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3180 a_4365_46436# a_4185_45028.t6 a_n1925_42282.t1 VSS.t1667 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3181 a_n998_44484# a_n1613_43370.t18 VSS.t3318 VSS.t3317 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3182 VDD.t2326 a_3177_46902# a_3067_47026# VDD.t2325 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3183 a_7577_46660# a_7411_46660# VDD.t1092 VDD.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3184 VDD.t2526 a_n2472_45546# a_n2956_38216.t0 VDD.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3185 a_14976_45028# a_13059_46348# VDD.t1371 VDD.t1370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3186 a_10835_43094# a_11967_42832.t43 VDD.t3144 VDD.t3011 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3187 a_12638_46436# a_12891_46348# VSS.t1437 VSS.t1436 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3188 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3189 a_n3420_37984.t5 a_n3690_38304# VSS.t1186 VSS.t1185 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3190 VSS.t2898 a_13661_43548.t16 a_743_42282.t5 VSS.t1108 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3191 a_12839_46116# a_12891_46348# a_n1741_47186.t1 VDD.t1645 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3192 VSS.t1597 a_3090_45724.t16 a_4927_45028# VSS.t1596 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3193 VSS.t1066 a_22000_46634# a_15227_44166.t2 VSS.t1065 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3194 VSS.t503 a_n863_45724# a_791_42968# VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3195 a_14209_32519.t0 a_22591_43396# VDD.t2535 VDD.t2534 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3196 a_4646_46812.t12 a_6298_44484# VDD.t1013 VDD.t1012 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3197 VSS.t1496 a_n4334_37440# a_n4064_37440.t7 VSS.t1495 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3198 a_n1613_43370.t0 a_5815_47464# VDD.t1341 VDD.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3199 a_n2661_43922.t0 a_12465_44636# VDD.t1282 VDD.t1281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3200 a_n2012_43396# a_n2129_43609# VSS.t398 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3201 VSS.t3541 a_11823_42460.t20 a_14635_42282# VSS.t3540 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3202 a_19692_46634.t1 a_12549_44172.t13 VSS.t2708 VSS.t2707 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3203 C8_P_btm.t3 a_n3565_39590.t12 VREF.t68 VDD.t3613 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3204 VSS.t1223 a_4520_42826# a_4093_43548# VSS.t1222 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3205 a_5013_44260# a_3905_42865# a_5025_43940# VDD.t2307 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3206 a_8018_44260# a_7499_43078# a_7911_44260# VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X3207 VDD.t3631 a_11823_42460.t18 a_14358_43442# VDD.t3630 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3208 a_167_45260# a_2202_46116# VDD.t1376 VDD.t1127 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3209 a_20254_46482# a_16327_47482.t40 VSS.t3304 VSS.t3303 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3210 VDD.t2722 a_10405_44172# a_8016_46348# VDD.t2721 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X3211 VIN_N.t4 EN_VIN_BSTR_N.t11 C10_N_btm.t32 VSS.t2918 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3212 a_742_44458# a_n443_42852.t25 VDD.t3723 VDD.t3722 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3213 VSS.t1918 a_19332_42282# a_4190_30871.t3 VSS.t1917 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 a_14840_46494# a_13925_46122# a_14493_46090# VSS.t808 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3215 VSS.t469 a_1414_42308# a_3457_43396# VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3216 a_20356_42852# a_18184_42460.t5 a_20256_42852# VDD.t3732 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X3217 a_19006_44850# a_18287_44626# a_18443_44721# VSS.t2408 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3218 a_9420_43940# a_768_44030.t16 a_9165_43940# VDD.t3686 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3219 VDD.t3315 a_10903_43370.t15 a_12005_46116# VDD.t3314 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3220 a_n4209_38216.t7 a_n2302_37984# VSS.t519 VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3221 VSS.t2972 a_12861_44030.t12 a_18280_46660# VSS.t2971 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3222 VSS.t2897 a_13661_43548.t14 a_15685_45394# VSS.t2896 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3223 C4_P_btm.t1 a_6123_31319.t4 VCM.t42 VSS.t1775 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3224 a_13575_42558# a_n97_42460.t14 a_13657_42308# VSS.t1677 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3225 VSS.t958 a_n2302_37690# a_n4209_37414.t4 VSS.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3226 a_8667_46634# a_6151_47436.t2 VDD.t2971 VDD.t2970 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3227 a_n1613_43370.t6 a_5815_47464# VSS.t1142 VSS.t1141 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3228 VDD.t1914 a_n971_45724.t10 a_n229_43646# VDD.t1913 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3229 a_n1057_35014.t1 a_n1696_34930.t13 VSS.t3480 VSS.t3479 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3230 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3231 a_21335_42336# a_16327_47482.t26 VDD.t3423 VDD.t3422 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3232 VSS.t2724 a_n3565_37414.t10 a_n3607_37440# VSS.t2723 sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3233 a_n2946_38778# a_n2956_38680.t5 VSS.t1716 VSS.t1551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3234 VSS.t1255 a_9127_43156# a_5891_43370.t6 VSS.t1254 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3235 VSS.t655 a_13351_46090# a_10903_43370.t2 VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3236 a_14309_45028# a_2711_45572.t11 VDD.t3731 VDD.t3730 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3237 VSS.t1840 a_413_45260.t4 a_22959_44484# VSS.t974 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3238 a_743_42282.t0 a_12549_44172.t10 a_20749_43396# VSS.t2704 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3239 VDD.t316 a_3877_44458# a_4185_45028.t0 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3240 a_13105_45348# a_13017_45260# a_n2661_46634.t1 VSS.t1937 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3241 VSS.t2191 a_6545_47178# a_6575_47204# VSS.t2190 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3242 a_8229_43396# a_7499_43078# a_8147_43396# VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3243 a_19551_46910# a_19466_46812# a_19333_46634# VDD.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3244 a_18280_46660# a_12549_44172.t17 a_17609_46634# VSS.t2711 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3245 VSS.t2127 a_18285_46348# a_18243_46436# VSS.t2126 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X3246 a_6945_45028.t2 a_5205_44484# VDD.t3342 VDD.t3341 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3247 a_3726_37500# a_3754_38470.t8 VDAC_Ni.t7 VSS.t2637 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3248 a_n4064_37440.t6 a_n4334_37440# VSS.t1498 VSS.t1497 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3249 a_20708_46348# a_20916_46384# a_20850_46482# VSS.t866 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3250 a_5167_46660# a_4651_46660# a_5072_46660# VSS.t2219 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3251 VDD.t2720 a_n1352_44484# a_n1177_44458# VDD.t2719 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3252 a_15685_45394# a_15415_45028# a_15595_45028# VSS.t1228 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3253 VDD.t3016 a_10193_42453.t7 a_18214_42558# VDD.t3015 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3254 a_21350_45938# a_20273_45572# a_21188_45572# VDD.t2610 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3255 a_n2002_35448# a_n1550_35448# VSS.t1943 VSS.t1942 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3256 a_7639_45394# a_n1151_42308.t8 a_7276_45260# VSS.t1657 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3257 VSS.t3395 a_526_44458.t14 a_10149_43396# VSS.t3394 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3258 a_7765_42852# a_7227_42852# VSS.t1308 VSS.t1307 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3259 a_501_45348# a_413_45260.t5 a_375_42282# VSS.t1841 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3260 VREF.t16 a_22612_30879.t8 C10_N_btm.t12 VDD.t1943 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3261 COMP_P.t5 a_1169_39587# VSS.t1010 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3262 a_16547_43609# a_16414_43172# VSS.t1242 VSS.t1241 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3263 a_n2438_43548.t7 a_949_44458# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3264 VDD.t3579 a_7754_40130.t4 a_8912_37509.t32 VDD.t3578 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3265 a_n3565_38502.t2 a_n2946_38778# VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3266 a_5891_43370.t3 a_9127_43156# VDD.t1466 VDD.t1465 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3267 a_13857_44734# a_13661_43548.t12 VDD.t3117 VDD.t3116 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3268 a_n2661_46098# a_2107_46812.t3 VDD.t3034 VDD.t3033 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3269 C10_N_btm.t9 a_22612_30879.t5 VREF.t13 VDD.t1940 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3270 VSS.t3356 a_16327_47482.t14 a_18953_45572# VSS.t3355 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3271 VSS.t787 a_742_44458# a_1568_43370# VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3272 a_19273_43230# a_18083_42858# a_19164_43230# VSS.t921 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3273 a_6123_31319.t0 a_7227_42308# VDD.t911 VDD.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3274 a_768_44030.t6 a_13487_47204# VSS.t611 VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3275 a_584_46384.t4 a_1123_46634# VSS.t1270 VSS.t1269 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3276 VDD.t3729 a_2711_45572.t8 a_4099_45572# VDD.t3728 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3277 a_12293_43646# a_9290_44172.t10 VDD.t3262 VDD.t3261 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3278 C8_N_btm.t4 a_5342_30871.t4 VCM.t28 VSS.t2622 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3279 a_8035_47026# a_6151_47436.t12 VDD.t2981 VDD.t2980 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3280 a_10306_45572# a_10193_42453.t6 a_10216_45572# VSS.t2786 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3281 a_18545_45144# a_13259_45724.t18 a_18450_45144# VDD.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X3282 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS.t1122 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3283 a_22629_37990# a_22537_39537# CAL_P.t1 VSS.t2528 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3284 a_n1423_46090# a_n1641_46494# VSS.t3292 VSS.t3291 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3285 a_16977_43638# a_16759_43396# VDD.t992 VDD.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3286 VDD.t2142 a_21855_43396# a_13678_32519.t1 VDD.t2141 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3287 VDD.t2848 a_6540_46812# a_6491_46660# VDD.t2847 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3288 VDD.t1275 a_22223_43948# a_14401_32519.t0 VDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3289 VDD.t683 a_n863_45724# a_n1099_45572# VDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3290 C10_P_btm.t33 EN_VIN_BSTR_P.t18 VIN_P.t4 VSS.t3572 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3291 a_n2946_37690# a_n2956_37592.t5 VSS.t1822 VSS.t1821 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3292 a_5111_42852# a_4905_42826# a_5193_42852# VDD.t1558 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3293 VDD.t1136 a_5263_45724# a_5204_45822# VDD.t1135 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3294 a_n467_45028# a_n745_45366# VSS.t2006 VSS.t2005 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3295 VSS.t3691 a_765_45546.t7 a_1208_46090# VSS.t3690 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3296 VDD.t1303 a_15095_43370# a_14955_43396# VDD.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3297 VDD.t1756 CAL_P.t4 VDD.t1756 VDD.t1755 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X3298 VSS.t2112 a_n4334_38304# a_n4064_37984.t7 VSS.t1342 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3299 VDD.t3487 a_2957_45546# a_2905_45572# VDD.t3486 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3300 a_8855_44734# a_4791_45118.t5 a_8783_44734# VDD.t2004 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3301 a_11963_45334# a_10903_43370.t11 VDD.t3311 VDD.t3310 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3302 a_n2661_44458.t2 a_11453_44696.t5 VDD.t3705 VDD.t3704 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X3303 VDD.t3759 a_4915_47217.t10 a_11415_45002# VDD.t3758 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3304 a_n1741_47186.t2 a_12005_46116# VDD.t2365 VDD.t2364 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3305 a_3600_43914# a_3537_45260.t20 a_3820_44260# VSS.t2670 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3306 a_21588_30879.t2 a_22223_47212# VSS.t2013 VSS.t2012 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3307 a_1848_45724# a_2063_45854.t14 a_1990_45899# VDD.t1872 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3308 a_14537_46482# a_14493_46090# a_14371_46494# VSS.t1894 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3309 a_10425_46660# a_9863_46634# VSS.t2268 VSS.t2267 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3310 a_16241_44734# a_2711_45572.t7 VDD.t3727 VDD.t3726 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3311 a_3905_42865# a_5257_43370# VDD.t1503 VDD.t1502 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3312 a_21811_47423# SINGLE_ENDED.t1 VSS.t2613 VSS.t2612 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3313 a_19365_45572# a_18175_45572# a_19256_45572# VSS.t2089 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3314 VDD.t474 a_22959_45572# a_20447_31679.t0 VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3315 a_3090_45724.t5 a_18911_45144# a_19113_45348# VSS.t2489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3316 DATA[2].t1 a_4007_47204# VDD.t2400 VDD.t2399 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3317 a_13777_45326# a_9482_43914# VSS.t1086 VSS.t1085 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3318 VDD.t3587 a_7754_40130.t8 a_8912_37509.t34 VDD.t3586 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3319 VCM.t62 a_5934_30871.t4 C5_N_btm.t1 VSS.t1774 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3320 a_n3690_39616# a_n3674_39768.t5 VDD.t2919 VDD.t2918 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3321 a_17333_42852# a_16795_42852# VDD.t2375 VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3322 a_11525_45546# a_11962_45724# a_11682_45822# VDD.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3323 VDD.t209 VSS.t3706 VDD.t208 VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3324 a_17595_43084# a_13259_45724.t12 VSS.t81 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3325 a_n13_43084# a_n755_45592.t24 a_133_43172# VSS.t3386 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X3326 a_n1696_34930.t2 a_n1794_35082.t16 VDD.t3067 VDD.t3066 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3327 a_19250_34978# a_18194_34908.t12 VSS.t3704 VSS.t3703 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3328 a_n3565_37414.t0 a_n2946_37690# VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3329 a_n2840_42282# a_n2661_42282.t3 VDD.t3649 VDD.t1981 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3330 a_20193_45348# a_18184_42460.t4 VSS.t3664 VSS.t3663 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3331 a_20719_46660# a_20273_46660# a_20623_46660# VSS.t1150 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3332 a_1756_43548# a_768_44030.t20 VSS.t3617 VSS.t3616 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3333 VSS.t3338 a_n1613_43370.t34 a_n1379_46482# VSS.t3337 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3334 a_n2472_43914# a_n2293_43922.t4 VSS.t2833 VSS.t2832 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3335 a_n2302_39072# a_n2312_39304.t5 VSS.t3474 VSS.t2883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3336 a_14456_42282# a_14635_42282# VDD.t2767 VDD.t2766 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3337 VDD.t768 a_20075_46420# a_20062_46116# VDD.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3338 VSS.t3654 a_2711_45572.t5 a_4099_45572# VSS.t3653 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3339 a_4927_45028# a_5147_45002# a_5105_45348# VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3340 a_21381_43940# a_21115_43940# VDD.t2420 VDD.t2419 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3341 SMPL_ON_N.t5 a_21753_35474# VSS.t1457 VSS.t1456 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 VSS.t1605 a_10227_46804.t10 a_10185_46660# VSS.t1604 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3343 a_n3607_38528# a_n3674_38680.t5 a_n3690_38528# VSS.t1780 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3344 a_4169_42308# a_1823_45246# a_3823_42558# VSS.t250 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3345 CLK_DATA.t4 a_n2833_47464# VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X3346 VDD.t2662 a_20894_47436# a_20843_47204# VDD.t2661 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3347 a_4704_46090# a_4883_46098.t8 VSS.t1633 VSS.t1632 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3348 VSS.t2744 a_n913_45002.t32 a_6761_42308# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3349 VDD.t1284 a_12465_44636# a_22223_47212# VDD.t1283 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3350 VREF.t42 a_n4315_30879.t16 C10_P_btm.t24 VDD.t2076 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3351 VDD.t1637 a_15051_42282# a_11823_42460.t0 VDD.t1636 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3352 VDD.t3515 a_20193_45348# a_20753_42852# VDD.t3514 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3353 VDD.t1078 a_15682_46116# a_11599_46634.t11 VDD.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3354 a_n2438_43548.t23 a_949_44458# VSS.t27 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3355 VDD.t1501 a_5257_43370# a_3357_43084.t0 VDD.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3356 VSS.t721 a_14113_42308# a_16522_42674# VSS.t720 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3357 a_22589_40055# en_comp VDD.t2638 VDD.t1937 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3358 a_2324_44458.t0 a_8953_45002# VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3359 VSS.t1453 a_21753_35474# SMPL_ON_N.t4 VSS.t1452 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3360 a_13460_43230# a_12379_42858# a_13113_42826# VDD.t1666 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3361 a_19240_46482# a_19123_46287# VSS.t1213 VSS.t1212 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3362 a_5829_43940# a_5495_43940# a_5745_43940# VDD.t2794 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3363 a_10227_46804.t2 a_14955_47212# VSS.t627 VSS.t626 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3364 VSS.t765 a_21487_43396# a_13467_32519.t2 VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3365 VDD.t864 a_7287_43370# a_7274_43762# VDD.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3366 VDD.t3187 a_12861_44030.t22 a_18911_45144# VDD.t3186 sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X3367 a_14955_43940# a_14537_43396# a_15037_43940# VDD.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3368 a_15953_42852# a_15227_44166.t16 VDD.t3672 VDD.t3671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3369 a_9114_42852# a_8037_42858# a_8952_43230# VDD.t1678 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3370 a_n4315_30879.t4 a_n2302_40160# VSS.t1176 VSS.t1175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3371 VDD.t1663 a_21753_35474# SMPL_ON_N.t1 VDD.t1662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3372 VSS.t2205 a_n901_46420# a_n443_46116.t6 VSS.t2204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3373 VSS.t309 a_8953_45002# a_2324_44458.t23 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3374 VSS.t780 a_8199_44636# a_8953_45546# VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3375 a_18780_47178# a_18597_46090# VSS.t1197 VSS.t1196 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3376 VDD.t3668 a_15227_44166.t14 a_18285_46348# VDD.t3667 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3377 a_16375_45002# a_18597_46090# VDD.t1400 VDD.t1399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3378 VDD.t3221 a_2324_44458.t49 a_6298_44484# VDD.t3220 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3379 a_15279_43071# a_5342_30871.t7 VSS.t2626 VSS.t2625 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3380 a_10193_42453.t0 a_20712_42282# VDD.t1729 VDD.t1728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3381 a_19335_46494# a_18985_46122# a_19240_46482# VDD.t2302 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3382 VDD.t1031 a_6298_44484# a_4646_46812.t11 VDD.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3383 a_5205_44484# a_5111_44636# VSS.t909 VSS.t908 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3384 C10_N_btm.t20 a_22612_30879.t16 VREF.t24 VDD.t1951 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3385 a_4842_47243# a_4791_45118.t20 VDD.t2020 VDD.t2019 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3386 VSS.t406 a_685_42968# a_791_42968# VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3387 a_11599_46634.t9 a_15682_46116# VDD.t1088 VDD.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3388 VSS.t2031 a_22591_45572# a_19963_31679.t3 VSS.t2030 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3389 C8_N_btm.t2 a_21076_30879.t6 VREF.t2 VDD.t3556 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3390 a_509_45572# a_n1099_45572# VSS.t544 VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3391 VSS.t1369 a_11322_45546# a_12016_45572# VSS.t1368 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X3392 a_n1059_45260.t3 a_17499_43370# VDD.t304 VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3393 a_20753_42852# a_10193_42453.t20 VDD.t3028 VDD.t3027 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3394 DATA[5].t7 a_11459_47204# VSS.t279 VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3395 a_16789_45572# a_15599_45572# a_16680_45572# VSS.t350 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3396 a_20362_44736# a_20640_44752# a_20596_44850# VDD.t2416 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 a_13622_42852# a_12545_42858# a_13460_43230# VDD.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3398 a_n1991_42858# a_n2157_42858# VDD.t1323 VDD.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3399 a_15143_45578# a_11823_42460.t16 VSS.t3538 VSS.t3537 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3400 VSS.t1044 a_n746_45260# a_556_44484# VSS.t1043 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3401 a_8701_44490# a_4791_45118.t14 VSS.t1759 VSS.t1758 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3402 a_n3607_37440# a_n3674_37592.t5 a_n3690_37440# VSS.t2655 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3403 a_10775_45002# a_10951_45334# a_10903_45394# VSS.t2171 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3404 VSS.t554 a_7227_47204# DATA[3].t6 VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3405 VDD.t2973 a_6151_47436.t3 a_14955_47212# VDD.t2972 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3406 a_15673_47210# a_15507_47210# VDD.t1721 VDD.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3407 VDD.t159 VSS.t3707 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3408 VDD.t2390 a_22589_40599# a_22537_40625# VDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3409 a_20679_44626# a_11967_42832.t40 VDD.t3141 VDD.t3140 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3410 VDD.t2162 a_n2946_39072# a_n3565_39304.t1 VDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3411 VDD.t2883 a_10991_42826# a_10922_42852# VDD.t2882 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X3412 a_5815_47464# a_6151_47436.t6 VSS.t2752 VSS.t2751 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X3413 a_8912_37509.t9 VDAC_P.t15 a_5088_37509.t4 VDD.t67 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X3414 a_n2956_37592.t3 a_n2472_45002# VSS.t969 VSS.t968 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3415 a_13667_43396# a_11823_42460.t9 VDD.t3621 VDD.t3620 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X3416 VSS.t979 a_n1920_47178# a_n2312_39304.t3 VSS.t978 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3417 VDD.t2923 a_n4064_40160.t12 a_n2216_40160# VDD.t2922 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3418 a_5164_46348# a_4927_45028# VSS.t1887 VSS.t1886 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X3419 a_949_44458# a_2324_44458.t33 VSS.t2996 VSS.t2995 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3420 a_15940_43402# a_12549_44172.t4 a_15868_43402# VSS.t2701 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3421 VDD.t3132 a_4646_46812.t41 a_4651_46660# VDD.t1592 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3422 a_1427_43646# a_1049_43396# a_1209_43370# VDD.t3507 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3423 a_19164_43230# a_18249_42858# a_18817_42826# VSS.t926 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3424 VDD.t3191 a_12861_44030.t26 a_21845_43940# VDD.t3190 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3425 a_2982_43646.t1 a_3232_43370.t20 VDD.t3049 VDD.t3048 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X3426 w_1575_34786.t9 EN_VIN_BSTR_P.t10 VDD.t3645 w_1575_34786.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3427 VDD.t2372 a_3600_43914# a_3499_42826# VDD.t2371 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3428 a_648_43396# a_526_44458.t30 a_548_43396# VSS.t3409 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3429 a_16409_43396# a_16243_43396# VDD.t1698 VDD.t1697 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3430 VSS.t1637 a_2063_45854.t5 a_11136_45572# VSS.t1636 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3431 VSS.t258 a_1823_45246# a_2202_46116# VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3432 a_10903_45394# a_9290_44172.t8 VSS.t3056 VSS.t3055 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X3433 VDD.t2892 a_n3420_39616.t9 a_n2860_39866# VDD.t2891 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3434 a_18243_46436# a_18189_46348# a_18147_46436# VSS.t998 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X3435 VSS.t1683 a_n971_45724.t5 a_3775_45552# VSS.t1682 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3436 a_9290_44172.t3 a_13635_43156# VDD.t2595 VDD.t2594 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3437 a_4700_47436# a_4915_47217.t4 a_4842_47243# VDD.t3753 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3438 VDD.t52 a_6453_43914# a_n2661_42282.t0 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3439 VSS.t3680 a_n2438_43548.t45 a_n2433_43396# VSS.t3679 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3440 a_11813_46116# a_11387_46155# VSS.t1004 VSS.t1003 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3441 VDD.t3509 a_380_45546# a_n356_45724# VDD.t3508 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3442 VDD.t1130 a_10053_45546# a_9625_46129# VDD.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3443 VDD.t3201 a_12861_44030.t34 a_19615_44636# VDD.t3200 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3444 a_2253_43940# a_n443_46116.t11 VDD.t3249 VDD.t3248 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X3445 VDD.t1526 a_13113_42826# a_13003_42852# VDD.t1525 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3446 a_765_45546.t3 a_17609_46634# VDD.t2254 VDD.t2253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3447 a_3503_45724# a_1823_45246# VSS.t260 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3448 VDD.t2726 a_3699_46348# a_3160_47472# VDD.t2725 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3449 VDD.t1702 a_9625_46129# a_10037_46155# VDD.t1701 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X3450 VDD.t1227 a_22223_45036# a_18114_32519.t0 VDD.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3451 a_18997_42308# a_18727_42674# a_18907_42674# VSS.t1529 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3452 a_5755_42852# a_n97_42460.t18 a_5837_42852# VDD.t1901 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3453 VDAC_Pi.t1 VSS.t3757 a_5700_37509.t1 VDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3454 a_12281_43396# a_n913_45002.t14 a_12293_43646# VDD.t2960 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3455 VDD.t2778 a_10533_42308# a_10723_42308# VDD.t2777 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3456 VSS.t1032 a_9863_47436# a_9804_47204# VSS.t1031 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3457 a_8049_45260.t2 a_n237_47217.t15 VDD.t3243 VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3458 a_11387_46482# a_11133_46155# VSS.t2457 VSS.t2456 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3459 VDD.t1256 a_21005_45260# a_19778_44110# VDD.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3460 VDD.t1404 a_8791_42308# a_5934_30871.t0 VDD.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3461 VDD.t790 a_13487_47204# a_768_44030.t3 VDD.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3462 VSS.t3233 VDD.t3793 VSS.t3232 VSS.t3231 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3463 a_895_43940# a_644_44056# VDD.t1039 VDD.t1038 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3464 VSS.t1777 a_n3420_38528.t10 a_n2946_38778# VSS.t1776 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3465 VDD.t3129 a_4646_46812.t39 a_7871_42858# VDD.t3128 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3466 a_3067_47026# a_2443_46660# a_2959_46660# VDD.t2799 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3467 a_19256_45572# a_18341_45572# a_18909_45814# VSS.t2091 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3468 VDD.t207 VSS.t3742 VDD.t206 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3469 C3_P_btm.t1 a_n4064_37984.t9 VREF_GND.t43 VSS.t1803 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3470 VSS.t1154 a_2713_42308# a_2903_42308# VSS.t1153 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3471 a_9863_47436# a_2063_45854.t6 a_10037_47542# VSS.t1638 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3472 a_15037_45618# a_13259_45724.t17 VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3473 a_3726_37500# CAL_P.t5 a_11206_38545.t4 VDD.t1757 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3474 a_10991_42826# a_10796_42968# a_11301_43218# VSS.t3271 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3475 a_2127_44172# a_1307_43914.t12 a_2253_44260# VSS.t3487 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3476 a_1823_45246# a_4704_46090# VDD.t1337 VDD.t1336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3477 VDD.t3750 a_n2438_43548.t44 a_n2433_44484# VDD.t3749 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3478 a_17678_43396# a_16327_47482.t20 VSS.t3364 VSS.t3363 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3479 a_n452_47436# a_n237_47217.t13 a_n310_47243# VDD.t3242 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3480 VDD.t3313 a_10903_43370.t13 a_12427_45724# VDD.t3312 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X3481 VDD.t112 VSS.t3766 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3482 a_3080_42308.t0 a_2903_42308# VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3483 a_22581_37893# a_22613_38993# VDD.t663 VDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3484 a_18057_42282# a_n1059_45260.t13 a_18310_42308# VSS.t2765 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3485 VSS.t2555 a_n452_45724# a_n1853_46287# VSS.t2554 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3486 a_n3674_39768.t3 a_n2472_43914# VSS.t1959 VSS.t1958 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3487 a_11967_42832.t0 a_15682_43940# VDD.t606 VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3488 a_8846_46660# a_6151_47436.t13 VSS.t2758 VSS.t2757 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3489 a_1307_43914.t4 a_2779_44458# VSS.t491 VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3490 a_22365_46825# EN_OFFSET_CAL.t1 VSS.t2609 VSS.t2608 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3491 VDD.t1760 CAL_P.t6 VDD.t1759 VDD.t1758 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X3492 C10_P_btm.t21 a_n4315_30879.t13 VREF.t39 VDD.t2073 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3493 a_1273_38525.t6 a_1107_38525# VSS.t2436 VSS.t2435 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3494 a_n89_45572# a_n743_46660.t10 a_n452_45724# VSS.t3557 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3495 a_n2472_42282# a_n2293_42282# VDD.t2780 VDD.t1985 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3496 VSS.t83 a_n2840_45002# a_n2810_45028.t2 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3497 a_15928_47570# a_15811_47375# VDD.t1180 VDD.t1179 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3498 a_518_46482# a_472_46348# VSS.t1217 VSS.t1216 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3499 a_15463_44811# a_11691_44458.t7 a_15004_44636# VDD.t3110 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3500 VSS.t801 a_17767_44458# a_17715_44484# VSS.t800 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3501 a_20556_43646# a_19692_46634.t6 a_20301_43646# VDD.t2062 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3502 a_n3420_39616.t1 a_n3690_39616# VDD.t1572 VDD.t1571 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3503 a_14309_45028# a_13059_46348# VDD.t1365 VDD.t1364 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3504 a_16237_45028# a_16375_45002# VDD.t848 VDD.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3505 a_8791_43396# a_3537_45260.t22 VDD.t2912 VDD.t2911 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3506 VDD.t2392 a_22589_40599# a_22725_38406# VDD.t2391 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3507 VDD.t3095 a_n4209_38216.t8 a_n4334_38304# VDD.t3094 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3508 a_9061_43230# a_7871_42858# a_8952_43230# VSS.t1467 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3509 a_1568_43370# a_n863_45724# VSS.t517 VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3510 VDD.t1325 a_n1423_42826# a_n1533_42852# VDD.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3511 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS.t2458 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3512 VSS.t2851 a_n1794_35082.t12 a_n1696_34930.t5 VSS.t2850 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3513 a_13575_42558# a_n97_42460.t7 a_13657_42558# VDD.t1896 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3514 a_6667_45809# a_6511_45714# a_6812_45938# VDD.t2753 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3515 a_3754_39964# a_7754_39964# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X3516 VSS.t3073 a_9290_44172.t27 a_10586_45546# VSS.t3072 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3517 a_16115_45572# a_15765_45572# a_16020_45572# VDD.t2483 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3518 VDD.t2748 a_18911_45144# a_3090_45724.t3 VDD.t2747 sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X3519 a_2725_42558# a_n755_45592.t10 VDD.t3438 VDD.t3437 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3520 a_18504_43218# a_17333_42852# VDD.t2862 VDD.t2861 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3521 VDD.t2732 a_3499_42826# a_n2293_42282# VDD.t2731 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3522 a_16979_44734# a_14539_43914# a_17061_44484# VSS.t815 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3523 a_2253_43940# a_2479_44172# a_2455_43940# VDD.t2138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3524 VDD.t75 VSS.t3751 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3525 VSS.t3468 a_1307_43914.t28 a_3681_42891# VSS.t3467 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3526 a_n310_47243# a_n971_45724.t8 VDD.t1910 VDD.t1909 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3527 a_5025_43940# a_1307_43914.t34 VDD.t3544 VDD.t3543 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3528 VSS.t853 a_626_44172# a_648_43396# VSS.t852 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3529 VSS.t3554 a_n3420_37440.t10 a_n2946_37690# VSS.t3553 sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3530 a_n3420_38528.t4 a_n3690_38528# VSS.t2273 VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3531 a_21356_42826# a_21381_43940# VSS.t2605 VSS.t2604 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3532 a_16877_43172# a_16823_43084# VSS.t1481 VSS.t1480 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3533 a_20841_46902# a_20623_46660# VDD.t2856 VDD.t2855 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3534 VDD.t235 VSS.t3733 VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3535 VDD.t211 VSS.t3724 VDD.t210 VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3536 VSS.t3526 a_6171_45002.t4 a_6125_45348# VSS.t3525 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3537 VSS.t2025 a_17595_43084# a_14539_43914# VSS.t2024 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3538 a_21137_46414# a_19692_46634.t4 VSS.t1810 VSS.t1809 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3539 a_5883_43914# a_8333_44056# VSS.t2020 VSS.t2019 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3540 a_20766_44850# a_20640_44752# a_20362_44736# VSS.t2165 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3541 VSS.t3241 VDD.t3796 VSS.t3240 VSS.t3239 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3542 VSS.t438 a_15682_43940# a_11967_42832.t17 VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3543 a_805_46414# a_472_46348# VDD.t1418 VDD.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3544 a_1176_45822# a_997_45618# VDD.t2589 VDD.t2588 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3545 VSS.t442 a_15682_43940# a_11967_42832.t31 VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3546 a_21887_42336# a_20202_43084# VDD.t1530 VDD.t1529 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3547 VSS.t2933 a_11967_42832.t36 a_18083_42858# VSS.t2932 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3548 DATA[2].t2 a_4007_47204# VDD.t2398 VDD.t2397 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3549 VDD.t442 a_1823_45246# a_3316_45546# VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3550 VDD.t502 a_8953_45002# a_2324_44458.t10 VDD.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3551 a_21513_45002# a_21363_45546# VDD.t1740 VDD.t1739 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3552 a_8704_45028# a_5937_45572.t10 a_8191_45002# VDD.t3565 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3553 a_3232_43370.t5 a_1823_45246# a_3363_44484# VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3554 a_13333_42558# a_13291_42460# a_13249_42558# VDD.t2339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3555 a_13661_43548.t2 a_18780_47178# VSS.t273 VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3556 a_5497_46414# a_5164_46348# VSS.t186 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3557 a_12749_45572# a_12549_44172.t25 a_12649_45572# VSS.t2718 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X3558 VSS.t275 a_n2840_43914# a_n4318_39768.t2 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3559 a_15037_44260# a_13556_45296# VSS.t467 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3560 VSS.t1229 a_22223_45572# a_19479_31679.t2 VSS.t1025 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3561 VDD.t3738 a_n2438_43548.t33 a_n133_46660# VDD.t3737 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3562 VDD.t544 a_n984_44318# a_n809_44244# VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3563 VDD.t2864 a_14815_43914# a_n2293_46634.t2 VDD.t2863 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3564 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS.t2513 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3565 a_8128_46384# a_7903_47542# VSS.t2294 VSS.t2293 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3566 VDD.t743 a_7281_43914# a_7229_43940# VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3567 VDD.t2000 a_13507_46334.t8 a_18907_42674# VDD.t1999 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3568 CLK_DATA.t7 a_n2833_47464# VSS.t242 VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3569 a_479_46660# a_33_46660# a_383_46660# VSS.t2472 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3570 VSS.t289 a_6667_45809# a_6598_45938# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3571 VDD.t2300 a_13904_45546# a_12594_46348# VDD.t2299 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3572 VDD.t1786 a_n881_46662.t13 a_n1021_46688# VDD.t1785 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3573 VDD.t3217 a_2324_44458.t45 a_15682_46116# VDD.t3216 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3574 a_8568_45546# a_8953_45546# a_8697_45822# VDD.t2624 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3575 a_17767_44458# a_17970_44736# VDD.t2200 VDD.t2199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3576 VREF.t70 a_19479_31679.t4 C1_N_btm.t2 VDD.t3663 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3577 VCM.t8 a_4190_30871.t16 C10_N_btm.t6 VSS.t2814 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3578 VDD.t3442 a_n755_45592.t13 a_133_42852# VDD.t3441 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3579 a_16241_44734# a_15227_44166.t12 VDD.t3665 VDD.t3664 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3580 a_10867_43940# a_7499_43078# a_10405_44172# VDD.t518 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3581 C10_N_btm.t16 a_22612_30879.t12 VREF.t20 VDD.t1947 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3582 VDD.t2412 a_10723_42308# a_5742_30871.t0 VDD.t2411 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3583 a_11823_42460.t1 a_15051_42282# VDD.t1631 VDD.t1630 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3584 a_20556_43646# a_20974_43370# VDD.t636 VDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3585 a_n3420_37440.t4 a_n3690_37440# VSS.t2300 VSS.t2299 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3586 a_4574_45260# a_4791_45118.t18 VSS.t1765 VSS.t1764 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3587 a_13483_43940# a_13249_42308# a_13565_43940# VDD.t1450 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3588 VDD.t2672 a_20159_44458# a_19321_45002# VDD.t2671 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X3589 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS.t2239 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3590 a_2583_47243# a_584_46384.t10 a_2124_47436# VDD.t2999 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3591 a_22612_30879.t2 a_22959_47212# VSS.t2320 VSS.t2319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3592 VDD.t1144 a_8349_46414# a_8379_46155# VDD.t1143 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3593 a_11599_46634.t22 a_15682_46116# VSS.t898 VSS.t897 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3594 VSS.t3613 a_768_44030.t17 a_2711_45572.t2 VSS.t3612 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3595 a_n2216_40160# a_n2312_40392.t5 a_n2302_40160# VDD.t1876 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X3596 VSS.t2511 a_14456_42282# a_5342_30871.t3 VSS.t2510 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3597 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD.t1602 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3598 VREF.t17 a_22612_30879.t9 C10_N_btm.t13 VDD.t1944 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3599 a_11608_46482# a_n1151_42308.t10 a_11387_46155# VSS.t1658 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3600 a_5093_45028# a_5111_44636# VDD.t1114 VDD.t1113 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3601 VSS.t303 a_8953_45002# a_2324_44458.t18 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3602 a_19862_44208# a_13747_46662.t4 VDD.t3085 VDD.t3084 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3603 VDD.t3658 a_15227_44166.t5 a_15597_42852# VDD.t3657 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3604 VSS.t21 a_949_44458# a_n2438_43548.t20 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3605 a_19335_46494# a_18819_46122# a_19240_46482# VSS.t2212 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3606 VDD.t3219 a_2324_44458.t48 a_6298_44484# VDD.t3218 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3607 VSS.t3149 VDD.t3822 VSS.t3148 VSS.t3147 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3608 a_8953_45546# a_8685_42308# VSS.t1981 VSS.t1980 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3609 a_n4318_38216.t1 a_n2472_42282# VDD.t2450 VDD.t2449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3610 a_18249_42858# a_18083_42858# VDD.t1120 VDD.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3611 a_12816_46660# a_11735_46660# a_12469_46902# VDD.t641 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3612 a_19268_43646# a_13661_43548.t7 a_19177_43646# VDD.t3109 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X3613 a_13258_32519.t0 a_19647_42308# VDD.t264 VDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3614 a_20256_42852# a_20202_43084# VDD.t1532 VDD.t1531 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X3615 VDD.t2819 a_16680_45572# a_16855_45546# VDD.t2818 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3616 VSS.t2396 a_n447_43370# a_n2129_43609# VSS.t2395 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3617 a_20528_45572# a_19466_46812# VDD.t873 VDD.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3618 a_11525_45546# a_10586_45546# a_11778_45572# VSS.t1079 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3619 VREF.t67 a_n3565_39590.t10 C8_P_btm.t0 VDD.t3610 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3620 a_3537_45260.t2 a_7287_43370# VDD.t860 VDD.t859 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3621 VDD.t3725 a_2711_45572.t4 a_20107_42308# VDD.t3724 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3622 a_16147_45260# a_17478_45572# VSS.t1148 VSS.t1147 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3623 a_n2109_45247# a_n2017_45002.t5 VSS.t2870 VSS.t2869 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3624 a_19610_45572# a_16327_47482.t32 VSS.t3294 VSS.t3293 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3625 a_19963_31679.t2 a_22591_45572# VSS.t2029 VSS.t2028 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3626 a_5837_43172# a_3537_45260.t10 VSS.t2664 VSS.t913 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3627 a_n143_45144# a_n755_45592.t15 VDD.t3445 VDD.t3444 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3628 VDD.t2176 a_18143_47464# a_12861_44030.t0 VDD.t2175 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3629 VDD.t2561 a_22959_47212# a_22612_30879.t1 VDD.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3630 a_n310_45572# a_n356_45724# VSS.t3445 VSS.t3444 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3631 VSS.t3195 VDD.t3778 VSS.t3194 VSS.t3193 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3632 VSS.t550 a_7227_47204# DATA[3].t7 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3633 a_15015_46420# a_10227_46804.t18 VDD.t1840 VDD.t1839 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3634 VSS.t2331 a_7227_45028# a_7230_45938# VSS.t2330 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3635 a_20596_44850# a_20159_44458# VDD.t2674 VDD.t2673 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3636 a_2957_45546# a_3090_45724.t9 VSS.t1589 VSS.t1588 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3637 VSS.t548 a_14579_43548# a_14537_43396# VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3638 VDD.t724 a_n2946_39866# a_n3565_39590.t2 VDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3639 VDD.t3161 a_11599_46634.t42 a_15507_47210# VDD.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3640 VDD.t2979 a_6151_47436.t9 a_6812_45938# VDD.t2978 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3641 VSS.t912 a_5111_44636# a_8333_44056# VSS.t911 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3642 VDD.t856 a_7287_43370# a_3537_45260.t0 VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X3643 a_8912_37509.t22 VDAC_N.t14 a_5700_37509.t7 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3644 VDD.t1648 a_20679_44626# a_20640_44752# VDD.t1647 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3645 a_n3565_39304.t0 a_n2946_39072# VDD.t2159 VDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3646 VDD.t1936 COMP_P.t10 a_n1329_42308# VDD.t1935 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3647 VSS.t1334 a_19321_45002# a_20567_45036# VSS.t1333 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3648 a_n2438_43548.t31 a_949_44458# VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3649 a_14513_46634# a_14180_46812# VSS.t2373 VSS.t2372 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3650 a_10903_43370.t0 a_13351_46090# VDD.t839 VDD.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3651 VSS.t967 a_n2472_45002# a_n2956_37592.t2 VSS.t966 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3652 a_10949_43914# a_10903_43370.t19 VDD.t3321 VDD.t3320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X3653 a_10149_43396# a_5111_44636# a_9803_43646# VSS.t914 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3654 VSS.t2135 a_19431_45546# a_19365_45572# VSS.t2134 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3655 VSS.t2595 a_16922_45042# a_17719_45144# VSS.t2594 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X3656 a_16112_44458# a_14539_43914# a_16241_44734# VDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3657 a_13943_43396# a_11823_42460.t28 a_13837_43396# VSS.t3549 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3658 C8_P_btm.t4 EN_VIN_BSTR_P.t8 VIN_P.t13 VSS.t3561 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3659 VDD.t2693 a_4099_45572# a_3483_46348.t0 VDD.t2692 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3660 a_6197_43396# a_6031_43396# VDD.t2437 VDD.t2436 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3661 VSS.t1910 a_18143_47464# a_12861_44030.t6 VSS.t1909 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3662 a_n2840_46634# a_n2661_46634.t3 VDD.t2040 VDD.t2039 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3663 a_380_45546# a_n357_42282.t4 a_603_45572# VSS.t1825 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3664 a_18533_43940# a_18326_43940# a_18451_43940# VDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3665 a_7309_42852# a_7499_43078# VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3666 VDD.t687 a_n863_45724# a_2448_45028# VDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3667 VSS.t1009 a_1169_39587# COMP_P.t4 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3668 a_5932_42308.t2 a_5755_42308# VSS.t2599 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3669 a_16328_43172# a_n97_42460.t12 VSS.t1675 VSS.t1674 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3670 VSS.t704 a_n2946_38778# a_n3565_38502.t5 VSS.t703 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3671 a_17583_46090# a_17715_44484# VDD.t2272 VDD.t2271 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3672 VDD.t123 VSS.t3767 VDD.t122 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3673 VDD.t2593 a_13635_43156# a_9290_44172.t2 VDD.t2592 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3674 VDD.t980 a_15433_44458# a_15463_44811# VDD.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3675 a_n2267_43396# a_n2433_43396# VSS.t2438 VSS.t2437 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3676 VDD.t3449 a_n755_45592.t21 a_8147_43396# VDD.t3448 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3677 VSS.t2621 a_10991_42826# a_10922_42852# VSS.t2620 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3678 a_5732_46660# a_4651_46660# a_5385_46902# VDD.t2469 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3679 a_19615_44636# a_12549_44172.t8 VDD.t2931 VDD.t2930 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X3680 a_5088_37509.t9 VDAC_P.t19 a_8912_37509.t14 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X3681 VDD.t2154 a_5129_47502# a_5159_47243# VDD.t2153 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3682 a_n2840_46090# a_n2661_46098# VDD.t2762 VDD.t2761 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3683 a_n967_45348# a_n913_45002.t15 a_n955_45028# VDD.t2961 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3684 a_19006_44850# a_18248_44752# a_18443_44721# VDD.t2197 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3685 a_n4209_39590.t6 a_n2302_39866# VSS.t863 VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3686 VDD.t2627 a_18817_42826# a_18707_42852# VDD.t2626 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3687 a_15559_46634# a_13507_46334.t10 VSS.t1745 VSS.t1744 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X3688 a_9803_43646# a_8953_45546# a_9885_43396# VSS.t2377 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3689 VDD.t3046 a_3232_43370.t14 a_9313_44734.t0 VDD.t3045 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3690 VDD.t928 a_n2840_42282# a_n3674_38680.t0 VDD.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3691 a_13460_43230# a_12545_42858# a_13113_42826# VSS.t1083 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3692 a_20362_44736# a_20679_44626# a_20637_44484# VSS.t1438 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3693 a_2713_42308# a_n913_45002.t27 a_2725_42558# VDD.t2966 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3694 a_768_44030.t1 a_13487_47204# VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3695 a_16241_47178# a_16023_47582# VSS.t1514 VSS.t1513 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3696 a_14955_43396# a_14205_43396# VDD.t2772 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3697 VSS.t2746 a_n913_45002.t33 a_10533_42308# VSS.t2745 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3698 a_7466_43396# a_n1613_43370.t19 VSS.t3320 VSS.t3319 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3699 a_n4064_40160.t1 a_n4334_40480# VDD.t2319 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3700 VDD.t2975 a_6151_47436.t7 a_5907_45546# VDD.t2974 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3701 a_16697_47582# a_15507_47210# a_16588_47582# VSS.t1511 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3702 a_n2267_44484# a_n2433_44484# VDD.t1319 VDD.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3703 a_15682_43940# a_2324_44458.t63 VDD.t3175 VDD.t3174 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3704 a_13693_46688# a_6755_46942# a_13607_46688# VSS.t2584 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3705 a_8912_37509.t26 VDAC_N.t18 a_5700_37509.t6 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3706 VDAC_Ni.t6 a_3754_38470.t4 a_3726_37500# VSS.t2633 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3707 a_11967_42832.t14 a_15682_43940# VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3708 VDD.t870 a_19778_44110# a_19741_43940# VDD.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3709 a_2609_46660# a_2443_46660# VSS.t2543 VSS.t2542 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3710 a_5708_44484# a_5257_43370# VSS.t1294 VSS.t1293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X3711 a_18143_47464# a_18479_47436# VDD.t1597 VDD.t1596 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3712 a_5263_46660# a_4817_46660# a_5167_46660# VSS.t1020 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3713 VSS.t1961 a_n2472_43914# a_n3674_39768.t2 VSS.t1960 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3714 VDAC_N.t5 a_3422_30871.t20 VCM.t59 VSS.t3524 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3715 a_12016_45572# a_11962_45724# a_11525_45546# VSS.t1024 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3716 VREF.t6 a_21588_30879.t6 C9_N_btm.t11 VDD.t1775 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3717 VSS.t2433 a_1107_38525# a_1273_38525.t7 VSS.t2432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3718 VSS.t1114 a_18057_42282# a_n356_44636.t1 VSS.t1113 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3719 VDD.t2807 a_21671_42860# a_3422_30871.t0 VDD.t2806 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3720 VDD.t530 a_8746_45002# a_8704_45028# VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3721 C9_N_btm.t1 a_4958_30871.t6 VCM.t33 VSS.t2694 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3722 a_3411_47243# a_3160_47472# a_2952_47436# VDD.t1479 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3723 a_n2840_46634# a_n2661_46634.t4 VSS.t1792 VSS.t1791 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3724 VSS.t2575 a_7705_45326# a_7639_45394# VSS.t2574 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3725 VSS.t201 a_167_45260# a_1423_45028.t3 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3726 a_11967_42832.t18 a_15682_43940# VSS.t422 VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3727 VDD.t895 a_9396_43370# a_5111_44636# VDD.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3728 a_743_42282.t4 a_13661_43548.t15 a_20301_43646# VDD.t3118 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3729 a_n3420_39616.t3 a_n3690_39616# VDD.t1574 VDD.t1573 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3730 a_133_43172# a_n357_42282.t10 VSS.t1833 VSS.t1832 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X3731 VSS.t3259 VDD.t3803 VSS.t3258 VSS.t3105 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3732 C10_N_btm.t17 a_22612_30879.t13 VREF.t21 VDD.t1948 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3733 VSS.t105 a_n2946_37690# a_n3565_37414.t4 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3734 VDD.t998 a_20512_43084# a_19987_42826# VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X3735 a_1891_43646# a_1307_43914.t13 VDD.t3551 VDD.t3550 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X3736 VSS.t3406 a_526_44458.t27 a_2075_43172# VSS.t3405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3737 a_14485_44260# a_5807_45002# a_12465_44636# VSS.t1280 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3738 a_n4318_39304.t2 a_n2840_43370# VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3739 VIN_P.t14 EN_VIN_BSTR_P.t15 C8_P_btm.t5 VSS.t3567 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3740 VSS.t1829 a_n357_42282.t6 a_17141_43172# VSS.t1828 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3741 a_11453_44696.t1 a_17719_45144# VSS.t669 VSS.t668 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X3742 VSS.t2770 a_n1059_45260.t19 a_8945_43396# VSS.t2769 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3743 a_17701_42308# a_17531_42308# VDD.t2374 VDD.t2373 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3744 a_13657_42558# a_11823_42460.t11 a_13575_42558# VDD.t3624 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3745 a_10545_42558# a_7499_43078# VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3746 a_8292_43218# a_7765_42852# VDD.t1519 VDD.t1518 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3747 a_16751_46987# a_5807_45002# a_16292_46812# VDD.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3748 a_10586_45546# a_9290_44172.t12 VSS.t3059 VSS.t3058 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3749 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS.t1121 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3750 VSS.t2092 a_16855_45546# a_16789_45572# VSS.t1711 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3751 a_45_45144# a_n143_45144# a_n37_45144# VDD.t2779 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3752 VDD.t2917 a_3537_45260.t29 a_4223_44672.t1 VDD.t2916 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3753 a_3626_43646.t0 a_1414_42308# a_3540_43646# VDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3754 VSS.t1401 a_n2946_37984# a_n3565_38216.t4 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3755 VDD.t2218 a_20107_42308# a_7174_31319.t0 VDD.t2217 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3756 a_3815_47204# a_3785_47178# VDD.t1620 VDD.t1619 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3757 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD.t2491 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3758 VCM.t29 a_5342_30871.t5 C8_N_btm.t5 VSS.t2623 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3759 a_15567_42826# a_15743_43084# a_15953_42852# VDD.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3760 VSS.t2342 a_10341_42308# a_11554_42852# VSS.t2341 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3761 VSS.t1769 a_4791_45118.t22 a_6640_46482# VSS.t1768 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X3762 a_6755_46942# a_15015_46420# VDD.t802 VDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3763 a_2437_43646.t2 a_1568_43370# VDD.t829 VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3764 VDAC_Pi.t8 a_7754_39632# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X3765 a_n3420_38528.t5 a_n3690_38528# VSS.t2275 VSS.t1185 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3766 a_n4209_39590.t0 a_n2302_39866# VDD.t1045 VDD.t1044 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3767 a_9823_46155# a_9804_47204# a_9823_46482# VSS.t585 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3768 a_1990_45899# a_167_45260# VDD.t378 VDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3769 a_15743_43084# a_19339_43156# VSS.t1872 VSS.t1871 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3770 a_5129_47502# a_4791_45118.t10 VDD.t2010 VDD.t2009 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3771 VDD.t1192 a_5385_46902# a_5275_47026# VDD.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3772 a_9145_43396.t1 a_8791_43396# VSS.t2189 VSS.t2188 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3773 VDD.t2564 a_20841_46902# a_20731_47026# VDD.t2563 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3774 a_n2438_43548.t9 a_949_44458# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3775 VIN_P.t5 EN_VIN_BSTR_P.t9 C10_P_btm.t32 VSS.t3562 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3776 VDD.t3500 a_n785_47204# a_327_47204# VDD.t3499 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3777 a_7276_45260# a_n1151_42308.t7 a_7418_45067# VDD.t1882 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3778 a_8103_44636# a_8375_44464# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3779 VSS.t444 a_15682_43940# a_11967_42832.t21 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3780 a_4915_47217.t1 a_12991_46634# VSS.t2549 VSS.t2548 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3781 VSS.t3159 VDD.t3827 VSS.t3158 VSS.t3129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3782 a_21753_35474# a_19998_34978# VSS.t1447 VSS.t1446 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3783 VDD.t965 a_8199_44636# a_8855_44734# VDD.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3784 VDD.t2929 a_12549_44172.t6 a_21115_43940# VDD.t2928 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3785 VDD.t1514 a_2553_47502# a_2583_47243# VDD.t1513 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3786 a_n327_42558# a_n357_42282.t17 VDD.t2101 VDD.t2100 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3787 a_12800_43218# a_12089_42308# VDD.t2322 VDD.t2321 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3788 VSS.t1924 a_20623_43914# a_20365_43914# VSS.t1923 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3789 VSS.t3559 a_n743_46660.t11 a_16501_45348# VSS.t3558 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3790 VSS.t392 a_22959_45036# a_19721_31679.t2 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3791 VSS.t2935 a_11967_42832.t37 a_16243_43396# VSS.t2934 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3792 VDD.t3583 a_7754_40130.t6 a_11206_38545.t1 VDD.t3582 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3793 a_n4318_38680.t1 a_n2472_42826# VDD.t2825 VDD.t2449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3794 a_3363_44484# a_526_44458.t19 VSS.t3397 VSS.t3396 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3795 a_13483_43940# a_13249_42308# a_13565_44260# VSS.t1247 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3796 a_7754_40130.t2 RST_Z.t5 VDD.t1771 VDD.t1770 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3797 VDD.t2713 a_4235_43370# a_n2661_45546.t2 VDD.t2712 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3798 a_n4209_38502.t5 a_n2302_38778# VSS.t2401 VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3799 a_13249_42558# a_10903_43370.t4 VDD.t3303 VDD.t3302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3800 a_18504_43218# a_17333_42852# VSS.t2601 VSS.t2600 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3801 a_n39_42308# a_n97_42460.t13 a_n473_42460# VSS.t1676 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3802 a_10210_45822# a_10180_45724# VDD.t2666 VDD.t2665 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X3803 VSS.t2937 a_11967_42832.t39 a_20512_43084# VSS.t2936 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3804 VSS.t3047 a_n443_46116.t13 a_2813_43396# VSS.t3046 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3805 VSS.t2911 a_4646_46812.t37 a_7411_46660# VSS.t2910 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3806 a_20273_46660# a_20107_46660# VSS.t1002 VSS.t1001 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3807 VDD.t3656 a_11341_43940.t4 a_22223_43948# VDD.t2029 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3808 a_n2312_38680.t3 a_n2104_46634# VSS.t3276 VSS.t3275 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3809 VDD.t1725 a_12791_45546# a_12427_45724# VDD.t1724 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X3810 a_2324_44458.t19 a_8953_45002# VSS.t305 VSS.t304 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3811 VDD.t1017 a_6298_44484# a_4646_46812.t2 VDD.t1016 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3812 a_19237_31679.t0 a_22959_44484# VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3813 VSS.t3702 a_18194_34908.t10 a_19250_34978# VSS.t3701 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3814 VDD.t2759 a_19328_44172# a_19279_43940# VDD.t2758 sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X3815 VDD.t1934 SMPL_ON_P.t8 a_n1605_47204# VDD.t1933 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3816 VSS.t2939 a_11967_42832.t42 a_12379_42858# VSS.t2938 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3817 VSS.t3597 a_15227_44166.t18 a_17719_45144# VSS.t3596 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3818 VDD.t2370 a_18315_45260# a_18189_46348# VDD.t2369 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X3819 a_10951_45334# a_8199_44636# VDD.t967 VDD.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3820 VREF.t43 a_n4315_30879.t17 C10_P_btm.t25 VDD.t2077 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3821 VDD.t2852 a_2123_42473# a_1184_42692# VDD.t2851 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3822 a_4791_45118.t3 a_4743_44484# VSS.t1118 VSS.t1117 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3823 a_21195_42852# a_20922_43172# VSS.t2314 VSS.t2313 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3824 a_4156_43218# a_3905_42865# a_3935_42891# VSS.t2048 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3825 a_15227_44166.t3 a_22000_46634# VSS.t1064 VSS.t1063 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3826 a_n3420_37440.t5 a_n3690_37440# VSS.t2302 VSS.t2301 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3827 a_n1899_43946# a_n2065_43946# VDD.t1601 VDD.t1600 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3828 VDD.t2131 a_17591_47464# a_16327_47482.t1 VDD.t2130 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3829 a_n743_46660.t1 a_n1021_46688# VSS.t454 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3830 a_n2293_45546.t3 a_2274_45254# VDD.t2776 VDD.t2775 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3831 a_11633_42308# a_9290_44172.t14 VSS.t3061 VSS.t3060 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3832 a_15682_46116# a_2324_44458.t58 VSS.t3021 VSS.t3020 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3833 a_20205_31679.t0 a_22223_46124# VDD.t1331 VDD.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3834 a_n2472_46634# a_n2293_46634.t3 VDD.t2879 VDD.t2878 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3835 a_2698_46116# a_2521_46116# VSS.t2569 VSS.t2568 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3836 a_11599_46634.t24 a_15682_46116# VSS.t894 VSS.t893 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3837 VDD.t3024 a_10193_42453.t14 a_11682_45822# VDD.t3023 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3838 VSS.t3227 VDD.t3791 VSS.t3226 VSS.t3225 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3839 VDD.t190 VSS.t3725 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3840 VDD.t3229 a_n3565_38502.t8 a_n3690_38528# VDD.t3228 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3841 a_5342_30871.t2 a_14456_42282# VSS.t2509 VSS.t2508 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3842 VDD.t2580 a_8325_42308# a_8791_42308# VDD.t2579 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3843 VSS.t31 a_949_44458# a_n2438_43548.t22 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3844 a_548_43396# a_n863_45724# a_458_43396# VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3845 VDD.t334 a_n4334_39616# a_n4064_39616.t0 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3846 VSS.t1902 a_1756_43548# a_1467_44172# VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X3847 a_288_46660# a_171_46873# VDD.t763 VDD.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3848 VSS.t39 a_949_44458# a_n2438_43548.t30 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3849 VDD.t1966 a_17517_44484.t2 a_22591_44484# VDD.t1965 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3850 VSS.t2743 a_n913_45002.t29 a_19511_42282# VSS.t2742 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3851 a_20894_47436# a_20990_47178# VSS.t2411 VSS.t2410 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3852 a_15312_46660# a_14976_45028# a_15009_46634# VSS.t2419 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3853 a_n2472_46090# a_n2293_46098.t3 VDD.t2875 VDD.t2021 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3854 VDD.t3744 a_n2438_43548.t40 a_n2157_46122# VDD.t3743 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3855 VSS.t977 a_22959_43948# a_17538_32519.t2 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3856 a_18194_34908.t2 a_n1794_35082.t18 VDD.t3071 VDD.t3070 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3857 C9_P_btm.t16 EN_VIN_BSTR_P.t11 VIN_P.t0 VSS.t3563 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3858 VDD.t2037 a_n4064_38528.t10 a_n2216_38778# VDD.t2036 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3859 a_8037_42858# a_7871_42858# VDD.t1676 VDD.t1675 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3860 a_n1736_43218# a_n1853_43023# VSS.t402 VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3861 a_n4209_37414.t7 a_n2302_37690# VSS.t960 VSS.t959 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3862 a_13527_45546# a_12861_44030.t32 VDD.t3197 VDD.t3196 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3863 VDD.t2448 a_n2472_42282# a_n4318_38216.t0 VDD.t2447 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3864 a_n2661_43370.t2 a_11415_45002# a_11361_45348# VSS.t2578 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3865 VSS.t1808 a_1273_38525.t12 a_2113_38308# VSS.t1807 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X3866 VDD.t1436 a_22165_42308# a_22223_42860# VDD.t1435 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3867 VDD.t1356 a_n2840_42826# a_n3674_39304.t0 VDD.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3868 VSS.t2589 a_14180_45002# a_13017_45260# VSS.t2588 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3869 a_15681_43442# a_12861_44030.t11 VDD.t3177 VDD.t3176 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3870 VDD.t3603 a_7754_40130.t15 a_8912_37509.t37 VDD.t3602 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3871 C8_N_btm.t0 a_21076_30879.t5 VREF.t0 VDD.t3555 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3872 VSS.t1174 a_n2302_40160# a_n4315_30879.t7 VSS.t1173 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3873 a_8488_45348# a_8199_44636# a_8191_45002# VSS.t783 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X3874 a_16588_47582# a_15673_47210# a_16241_47178# VSS.t1990 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3875 a_18220_42308# a_18184_42460.t8 VSS.t3666 VSS.t3665 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X3876 a_n1423_46090# a_n1641_46494# VDD.t3348 VDD.t3347 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3877 VDD.t3062 a_n1794_35082.t10 a_18194_34908.t1 VDD.t3061 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3878 VSS.t1343 a_n4334_38528# a_n4064_38528.t6 VSS.t1342 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3879 VDD.t2170 a_18143_47464# a_12861_44030.t2 VDD.t2169 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3880 a_17609_46634# a_12549_44172.t23 a_18280_46660# VSS.t2717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3881 a_16115_45572# a_15599_45572# a_16020_45572# VSS.t347 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3882 VSS.t563 a_19700_43370# a_n97_42460.t2 VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3883 VSS.t1504 a_2124_47436# a_1209_47178# VSS.t1503 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3884 VREF_GND.t6 a_17730_32519.t4 C9_N_btm.t4 VSS.t2879 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3885 a_15595_45028# a_15415_45028# VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3886 VDD.t2844 a_6755_46942# a_12741_44636.t1 VDD.t2843 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3887 VSS.t2425 a_19615_44636# a_18579_44172# VSS.t2424 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3888 a_12545_42858# a_12379_42858# VDD.t1669 VDD.t1668 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3889 a_16942_47570# a_16327_47482.t36 VSS.t3298 VSS.t3297 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3890 a_8791_45572# a_7499_43078# a_8697_45572# VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3891 a_14853_42852# a_n913_45002.t23 a_14635_42282# VDD.t2965 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3892 a_n2438_43548.t27 a_949_44458# VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3893 a_8333_44056# a_4223_44672.t8 VSS.t2659 VSS.t2658 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3894 VSS.t2693 a_4958_30871.t5 a_17531_42308# VSS.t2692 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3895 a_6511_45714# a_4646_46812.t36 VSS.t2909 VSS.t2908 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3896 VDD.t1043 a_10949_43914# a_10867_43940# VDD.t1042 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X3897 a_17973_43940# a_17737_43940# VDD.t2381 VDD.t2380 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X3898 a_18494_42460# a_18907_42674# VDD.t1744 VDD.t1743 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3899 a_17061_44734# a_15227_44166.t15 VDD.t3670 VDD.t3669 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3900 a_n2472_46634# a_n2293_46634.t4 VSS.t2617 VSS.t2614 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3901 C2_P_btm.t0 a_3080_42308.t7 VCM.t1 VSS.t2631 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3902 VSS.t2535 a_5267_42460# a_4905_42826# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3903 VSS.t3676 a_n2438_43548.t39 a_n2065_43946# VSS.t3675 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3904 VDD.t3599 a_7754_40130.t13 a_3754_38470.t0 VDD.t3598 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3905 a_22629_38406# a_22537_39537# CAL_N.t1 VSS.t2528 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3906 VDD.t2095 a_n357_42282.t13 a_5837_42852# VDD.t2094 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3907 a_9159_45572# a_5937_45572.t19 VSS.t3502 VSS.t3501 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3908 a_3483_46348.t1 a_4099_45572# VDD.t2695 VDD.t2694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3909 a_8238_44734# a_8199_44636# VDD.t971 VDD.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3910 VSS.t1718 a_17517_44484.t3 a_22591_44484# VSS.t1717 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3911 VDD.t2957 a_n3565_37414.t9 a_n3690_37440# VDD.t2956 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3912 VDD.t2510 a_3381_47502# a_3411_47243# VDD.t2509 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3913 VSS.t2327 a_21613_42308# a_22775_42308# VSS.t2326 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3914 COMP_P.t7 a_1169_39587# VSS.t1008 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3915 a_10150_46912# a_10467_46802# a_10425_46660# VSS.t528 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3916 a_526_44458.t1 a_3147_46376# VDD.t2224 VDD.t2223 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3917 a_n2810_45572.t0 a_n2840_45546# VDD.t2567 VDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3918 a_13675_47204# a_n1435_47204.t3 a_13569_47204# VDD.t2111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X3919 VSS.t174 a_11827_44484# a_22223_45036# VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3920 a_5518_44484# a_3483_46348.t9 VDD.t3289 VDD.t3288 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X3921 VDD.t2028 a_n4064_37440.t10 a_n2216_37690# VDD.t2027 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3922 a_22165_42308# a_21887_42336# VDD.t1148 VDD.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3923 a_n3565_38502.t1 a_n2946_38778# VDD.t885 VDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3924 a_5891_43370.t2 a_9127_43156# VDD.t1464 VDD.t1463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3925 a_13678_32519.t0 a_21855_43396# VDD.t2144 VDD.t2143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3926 a_n2312_40392.t0 a_n2288_47178# VDD.t844 VDD.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3927 VDD.t2249 a_8605_42826# a_8495_42852# VDD.t2248 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3928 a_7499_43078# a_10083_42826# VSS.t738 VSS.t737 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3929 VDD.t3517 a_20193_45348# a_21887_42336# VDD.t3516 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3930 a_18691_45572# a_18341_45572# a_18596_45572# VDD.t2345 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3931 a_13076_44458# a_9482_43914# VSS.t1094 VSS.t1093 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3932 a_3600_43914# a_1307_43914.t23 a_3992_43940# VDD.t3528 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3933 VSS.t1502 a_n4334_37440# a_n4064_37440.t5 VSS.t1501 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3934 a_4743_43172# a_3537_45260.t25 a_4649_43172# VSS.t2675 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3935 a_11387_46155# a_11309_47204# a_11387_46482# VSS.t2461 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3936 a_n755_45592.t5 a_n809_44244# VSS.t363 VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3937 a_15682_43940# a_2324_44458.t50 VDD.t3223 VDD.t3222 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3938 VDD.t2050 a_1666_39587.t4 a_1169_39587# VDD.t2049 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3939 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS.t2465 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3940 a_11554_42852# a_10835_43094# a_10991_42826# VSS.t2445 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3941 VSS.t3131 VDD.t3816 VSS.t3130 VSS.t3129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3942 VDD.t566 a_2680_45002# a_2274_45254# VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3943 C10_N_btm.t4 a_4190_30871.t11 VCM.t6 VSS.t2809 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3944 VSS.t1785 a_9313_44734.t4 a_22959_42860# VSS.t1784 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3945 VSS.t847 a_6298_44484# a_4646_46812.t24 VSS.t846 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3946 VDD.t2740 a_n1177_43370# a_n1190_43762# VDD.t2739 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3947 VDD.t2839 a_6755_46942# a_13556_45296# VDD.t2838 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3948 a_n785_47204# a_n815_47178# VDD.t3498 VDD.t3497 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3949 VDD.t32 a_949_44458# a_n2438_43548.t3 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3950 VDD.t1926 a_n971_45724.t24 a_8147_43396# VDD.t1925 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3951 a_n4251_40480# a_n4318_40392.t5 a_n4334_40480# VSS.t1842 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3952 VSS.t3201 VDD.t3780 VSS.t3200 VSS.t3199 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3953 VDD.t3601 a_7754_40130.t14 a_8912_37509.t36 VDD.t3600 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3954 a_19900_46494# a_18819_46122# a_19553_46090# VDD.t2463 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3955 C9_P_btm.t8 a_n4209_39590.t11 VREF.t56 VDD.t3074 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3956 a_12359_47026# a_10227_46804.t14 VDD.t1836 VDD.t1835 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3957 a_12561_45572# a_11823_42460.t23 VSS.t3545 VSS.t3544 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X3958 a_10083_42826# a_10518_42984# VDD.t3327 VDD.t3326 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3959 VSS.t771 a_10355_46116# a_8199_44636# VSS.t770 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3960 a_3422_30871.t1 a_21671_42860# VDD.t2809 VDD.t2808 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3961 a_5937_45572.t1 a_5907_45546# VDD.t934 VDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3962 a_21005_45260# a_21101_45002# VSS.t2177 VSS.t2176 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X3963 VDD.t3352 a_16327_47482.t35 a_17767_44458# VDD.t3351 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3964 a_12649_45572# a_10903_43370.t22 a_12561_45572# VSS.t3103 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3965 VSS.t1328 a_19321_45002# a_19113_45348# VSS.t1327 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3966 a_5111_44636# a_9396_43370# VDD.t897 VDD.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3967 a_12469_46902# a_12251_46660# VDD.t1428 VDD.t1427 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3968 a_21297_45572# a_20107_45572# a_21188_45572# VSS.t2224 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3969 a_376_46348# a_584_46384.t15 a_518_46482# VSS.t2780 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3970 a_15146_44484# a_9482_43914# VSS.t1100 VSS.t1099 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3971 VIN_P.t1 EN_VIN_BSTR_P.t19 C6_P_btm.t5 VSS.t3573 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3972 a_n1696_34930.t1 a_n1794_35082.t6 VDD.t3058 VDD.t3057 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3973 VDD.t1920 a_n971_45724.t16 a_n327_42558# VDD.t1919 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3974 a_n3565_37414.t2 a_n2946_37690# VDD.t286 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3975 a_14180_45002# a_14537_43396# a_14309_45028# VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3976 VDD.t3026 a_10193_42453.t18 a_16237_45028# VDD.t3025 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3977 a_18681_44484# a_16327_47482.t37 VSS.t3300 VSS.t3299 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3978 VSS.t2333 a_15009_46634# a_14180_46812# VSS.t2332 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3979 a_17829_46910# a_12549_44172.t11 a_765_45546.t0 VDD.t2934 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X3980 a_2304_45348# a_2274_45254# a_2232_45348# VSS.t2515 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3981 VDD.t352 a_1169_39043# comp_n VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3982 a_6598_45938# a_6511_45714# a_6194_45824# VDD.t2754 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3983 VDD.t1072 a_15682_46116# a_11599_46634.t4 VDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3984 a_n3565_38216.t6 a_n2946_37984# VSS.t1402 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3985 a_5745_43940# a_5013_44260# a_5663_43940# VDD.t3492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3986 VDD.t3014 a_10193_42453.t5 a_18533_43940# VDD.t3013 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3987 SMPL_ON_P.t2 a_n2002_35448# VDD.t2406 VDD.t2405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3988 a_5742_30871.t2 a_10723_42308# VSS.t2161 VSS.t2160 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3989 VDD.t1060 a_15682_46116# a_11599_46634.t3 VDD.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3990 a_19478_44056# a_3090_45724.t17 VDD.t1821 VDD.t1820 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3991 a_10890_34112.t0 EN_VIN_BSTR_N.t16 VIN_N.t2 VSS.t2922 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3992 VSS.t1426 a_15051_42282# a_11823_42460.t5 VSS.t1425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3993 a_10185_46660# a_10150_46912# a_9863_46634# VSS.t2405 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3994 a_8192_45572# a_8199_44636# VSS.t773 VSS.t772 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3995 a_15890_42674# a_15764_42576# a_15486_42560# VSS.t2229 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3996 a_10835_43094# a_11967_42832.t49 VSS.t2945 VSS.t2944 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3997 VSS.t414 a_15682_43940# a_11967_42832.t26 VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3998 a_n699_43396# a_n1177_43370# VDD.t2738 VDD.t2737 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3999 a_14033_45822# a_3483_46348.t11 VDD.t3291 VDD.t3290 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4000 VSS.t3221 VDD.t3789 VSS.t3220 VSS.t3219 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4001 a_6101_44260# a_1307_43914.t35 a_5663_43940# VSS.t3471 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4002 a_7927_46660# a_7577_46660# a_7832_46660# VDD.t1715 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4003 a_21496_47436# a_4883_46098.t6 VDD.t1862 VDD.t1861 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X4004 a_16721_46634# a_16388_46812# VDD.t659 VDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4005 a_5826_44734# a_5147_45002# a_5518_44484# VDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X4006 VDD.t893 a_16763_47508# a_16750_47204# VDD.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4007 VSS.t827 a_6298_44484# a_4646_46812.t26 VSS.t826 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4008 VDD.t1254 a_n746_45260# a_175_44278# VDD.t1253 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4009 a_n443_46116.t5 a_n901_46420# VSS.t2209 VSS.t2208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4010 a_2813_43396# a_3232_43370.t16 a_2982_43646.t2 VSS.t2827 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4011 a_6171_42473# a_5932_42308.t5 VDD.t2053 VDD.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4012 VDD.t2258 a_601_46902# a_491_47026# VDD.t2257 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4013 VSS.t2907 a_4646_46812.t35 a_6031_43396# VSS.t2906 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4014 VDD.t84 VSS.t3710 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4015 VDD.t1476 a_1123_46634# a_1110_47026# VDD.t1475 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4016 VSS.t1168 a_13059_46348# a_12638_46436# VSS.t1167 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4017 C10_N_btm.t26 a_18114_32519.t6 VREF_GND.t15 VSS.t2649 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4018 a_11787_45002# a_11963_45334# a_11915_45394# VSS.t2368 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4019 VSS.t2785 a_584_46384.t23 a_2998_44172# VSS.t2784 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4020 a_8292_43218# a_7765_42852# VSS.t1310 VSS.t1309 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4021 VDD.t2824 a_n2472_42826# a_n4318_38680.t0 VDD.t2447 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4022 a_1667_45002# a_1823_45246# VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X4023 VDD.t2522 a_n3690_38528# a_n3420_38528.t1 VDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4024 a_20731_47026# a_10227_46804.t12 VDD.t1834 VDD.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4025 a_8062_46482# a_8016_46348# VSS.t946 VSS.t945 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4026 VDD.t1035 a_6298_44484# a_4646_46812.t7 VDD.t1034 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4027 a_n2216_38778# a_n2312_38680.t5 a_n2302_38778# VDD.t2877 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4028 VSS.t2963 a_11599_46634.t49 a_20107_46660# VSS.t2962 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4029 a_13925_46122# a_13759_46122# VSS.t1414 VSS.t1413 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 VSS.t3625 CLK.t0 a_8953_45002# VSS.t1077 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4031 VSS.t3274 a_n2104_46634# a_n2312_38680.t2 VSS.t3273 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4032 a_5385_46902# a_5167_46660# VDD.t1190 VDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4033 a_n1177_44458# a_n1613_43370.t41 VDD.t3394 VDD.t3393 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4034 VDD.t524 a_7499_43078# a_10729_43914# VDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4035 a_9803_43646# a_8953_45546# a_9885_43646# VDD.t2625 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4036 VDD.t2617 a_19256_45572# a_19431_45546# VDD.t2616 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4037 a_7911_44260# a_7845_44172# a_7542_44172# VSS.t2561 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X4038 VDD.t1102 a_5111_44636# a_7542_44172# VDD.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4039 VDD.t2760 a_6761_42308# a_7227_42308# VDD.t1877 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4040 VDD.t2123 a_19553_46090# a_19443_46116# VDD.t2122 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4041 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS.t1126 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4042 a_5205_44484# a_5343_44458# VSS.t1060 VSS.t1059 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4043 a_22400_42852# a_22223_42860# VSS.t1236 VSS.t1235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4044 a_12603_44260# a_12549_44172.t26 a_12495_44260# VSS.t2719 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X4045 a_3638_45822# a_1823_45246# VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X4046 a_17324_43396# a_16243_43396# a_16977_43638# VDD.t1700 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4047 a_19452_47524# a_19386_47436# a_13747_46662.t1 VSS.t1335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4048 a_5275_47026# a_4651_46660# a_5167_46660# VDD.t2470 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4049 VSS.t2056 a_327_47204# DATA[0].t6 VSS.t2055 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4050 a_11915_45394# a_11823_42460.t25 VSS.t3547 VSS.t3546 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X4051 a_14447_46660# a_n1151_42308.t15 a_14084_46812# VSS.t1662 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4052 a_20731_47026# a_20107_46660# a_20623_46660# VDD.t1198 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4053 VSS.t3334 a_n1613_43370.t31 a_n1655_44484# VSS.t3333 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4054 a_12800_43218# a_12089_42308# VSS.t2070 VSS.t2069 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4055 VDD.t490 a_8953_45002# a_2324_44458.t7 VDD.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4056 VDAC_N.t7 a_3422_30871.t8 VCM.t47 VSS.t3510 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4057 VSS.t1519 a_20712_42282# a_10193_42453.t3 VSS.t1518 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4058 a_15720_42674# a_15051_42282# VDD.t1629 VDD.t1628 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4059 VSS.t3651 a_n443_42852.t23 a_421_43172# VSS.t3650 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4060 a_14493_46090# a_14275_46494# VDD.t996 VDD.t995 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4061 VDD.t3167 a_11599_46634.t48 a_15599_45572# VDD.t3166 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4062 a_n659_45366# a_n746_45260# a_n745_45366# VSS.t1048 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4063 a_15682_46116# a_2324_44458.t60 VSS.t2965 VSS.t2964 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4064 a_n881_46662.t2 a_14495_45572# VSS.t2234 VSS.t2233 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4065 a_8685_43396.t0 a_8147_43396# VDD.t2756 VDD.t2755 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4066 C7_P_btm.t2 a_n4209_39304.t8 VREF.t30 VDD.t1969 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4067 a_765_45546.t4 a_17609_46634# a_17639_46660# VSS.t1997 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4068 a_8912_37509.t23 VDAC_N.t15 a_5700_37509.t5 VDD.t67 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X4069 a_11554_42852# a_10796_42968# a_10991_42826# VDD.t3324 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4070 a_19386_47436# a_19321_45002# VSS.t1332 VSS.t1331 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4071 a_8492_46660# a_7411_46660# a_8145_46902# VDD.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4072 a_2063_45854.t1 a_9863_46634# VDD.t2516 VDD.t2515 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4073 VDD.t2507 a_15803_42450# a_15764_42576# VDD.t2506 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4074 a_1337_46436# a_1176_45822# VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4075 VSS.t23 a_949_44458# a_n2438_43548.t16 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4076 VSS.t2137 a_4419_46090# a_4365_46436# VSS.t2136 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4077 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4078 VDD.t1218 a_9067_47204# DATA[4].t2 VDD.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4079 VSS.t1939 a_6575_47204# a_9067_47204# VSS.t1938 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4080 a_n1331_43914# a_n1549_44318# VSS.t262 VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4081 VDD.t2902 a_3537_45260.t12 a_5093_45028# VDD.t2901 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4082 VSS.t2453 a_11189_46129# a_11608_46482# VSS.t2452 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4083 a_20835_44721# a_20640_44752# a_21145_44484# VSS.t2164 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X4084 w_10694_33990.t6 a_10890_34112.t4 w_10694_33990.t5 w_10694_33990.t2 sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X4085 a_n327_42558# a_n97_42460.t22 a_n473_42460# VDD.t1905 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X4086 a_8147_43396# a_7499_43078# VDD.t514 VDD.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X4087 VDD.t2549 a_n3690_37440# a_n3420_37440.t1 VDD.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4088 a_19431_46494# a_18985_46122# a_19335_46494# VSS.t2043 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4089 VDD.t1750 a_12607_44458# a_n2661_43922.t2 VDD.t1749 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4090 VDD.t2647 a_17324_43396# a_17499_43370# VDD.t2646 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4091 a_8685_42308# a_8515_42308# VSS.t1979 VSS.t1978 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4092 a_1414_42308# a_1067_42314# VSS.t603 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4093 VDD.t1864 a_4883_46098.t7 a_10355_46116# VDD.t1863 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4094 a_n2216_37690# a_n2810_45028.t5 a_n2302_37690# VDD.t1761 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4095 VDD.t3020 a_10193_42453.t12 a_9885_42558# VDD.t3019 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4096 VDD.t2790 a_21356_42826# a_n357_42282.t0 VDD.t2789 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4097 a_16977_43638# a_16759_43396# VSS.t807 VSS.t806 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4098 VSS.t2064 a_n4334_40480# a_n4064_40160.t4 VSS.t2063 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4099 VSS.t3033 a_n237_47217.t9 a_8270_45546# VSS.t3032 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4100 a_10555_43940# a_5891_43370.t18 VDD.t1808 VDD.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4101 a_1049_43396# a_458_43396# VSS.t2384 VSS.t2383 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4102 VSS.t1036 a_22775_42308# a_22485_38105# VSS.t1035 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4103 VDD.t3708 a_n443_42852.t10 a_742_44458# VDD.t3707 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4104 a_8145_46902# a_7927_46660# VSS.t235 VSS.t234 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4105 a_21613_42308# a_21335_42336# VDD.t2291 VDD.t2290 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4106 VDD.t2881 a_n23_45546# a_7_45899# VDD.t2880 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4107 VSS.t57 a_16019_45002# a_15903_45785# VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X4108 VCM.t31 a_5342_30871.t9 C8_P_btm.t9 VSS.t2627 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4109 VDD.t2829 a_2698_46116# a_2804_46116# VDD.t2828 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4110 a_20935_43940# a_18479_47436# VSS.t1385 VSS.t1384 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4111 a_18194_34908.t0 a_n1794_35082.t17 VDD.t3069 VDD.t3068 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4112 a_2713_42308# a_n755_45592.t27 VSS.t3390 VSS.t3389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4113 VDD.t2744 a_n699_43396# a_4743_44484# VDD.t2743 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4114 DATA[1].t4 a_1431_47204# VSS.t1856 VSS.t1855 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4115 a_17591_47464# a_10227_46804.t21 VSS.t1619 VSS.t1618 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4116 a_9223_42460# a_5891_43370.t21 VDD.t1812 VDD.t1811 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4117 a_12741_44636.t0 a_14537_43396# VDD.t806 VDD.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4118 a_2684_37794# a_1666_39587.t5 a_1666_39043.t0 VSS.t1801 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4119 VDD.t1534 a_20202_43084# a_21335_42336# VDD.t1533 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4120 a_564_42282# a_743_42282.t8 VSS.t3473 VSS.t3472 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4121 a_15367_44484# a_13556_45296# a_15004_44636# VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4122 VSS.t1170 a_n2302_40160# a_n4315_30879.t6 VSS.t1169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4123 VSS.t1337 a_n452_47436# a_n815_47178# VSS.t1336 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4124 VDD.t1874 a_2063_45854.t15 a_9863_47436# VDD.t1873 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4125 a_2981_46116# a_2804_46116# VSS.t3282 VSS.t3281 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4126 VSS.t2492 a_6511_45714# a_6472_45840# VSS.t2491 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4127 VSS.t1977 a_13159_45002# a_13105_45348# VSS.t1976 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4128 a_11967_42832.t1 a_15682_43940# VDD.t604 VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4129 EN_VIN_BSTR_P.t5 a_n1696_34930.t9 w_1575_34786.t5 w_1575_34786.t4 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4130 a_9223_42460# a_5891_43370.t19 VSS.t1577 VSS.t1576 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4131 VSS.t229 a_19987_42826# a_n2017_45002.t2 VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X4132 a_20692_30879.t0 a_22959_46124# VDD.t2211 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4133 a_21188_45572# a_20273_45572# a_20841_45814# VSS.t2367 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4134 a_9028_43914# a_9482_43914# VSS.t1092 VSS.t1091 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4135 VDD.t2274 a_17715_44484# a_17737_43940# VDD.t2273 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4136 VSS.t1904 a_n2840_44458# a_n4318_40392.t2 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4137 VSS.t346 a_15004_44636# a_14815_43914# VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4138 a_16759_43396# a_16243_43396# a_16664_43396# VSS.t1490 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4139 a_4574_45260# a_4791_45118.t19 VDD.t2018 VDD.t2017 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4140 a_17829_46910# a_12861_44030.t13 VDD.t3179 VDD.t3178 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4141 VSS.t3049 a_n443_46116.t15 a_4880_45572# VSS.t3048 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X4142 a_n4064_38528.t0 a_n4334_38528# VDD.t1551 VDD.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4143 VDD.t941 a_1799_45572# a_1983_46706# VDD.t940 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4144 VDD.t1738 a_21363_45546# a_21350_45938# VDD.t1737 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4145 SMPL_ON_P.t1 a_n2002_35448# VDD.t2408 VDD.t2407 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4146 a_n4064_40160.t6 a_n4334_40480# VSS.t2068 VSS.t2067 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X4147 VDD.t1235 a_22775_42308# a_22485_38105# VDD.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4148 a_13259_45724.t2 a_17583_46090# VSS.t1920 VSS.t1919 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4149 w_1575_34786.t14 a_n1057_35014.t5 w_1575_34786.t14 w_1575_34786.t13 sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X4150 VDAC_P.t0 a_3422_30871.t5 VCM.t44 VSS.t3507 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4151 C1_P_btm.t3 a_n4064_37440.t9 VREF_GND.t25 VSS.t1728 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4152 VIN_P.t6 EN_VIN_BSTR_P.t22 C4_P_btm.t2 VSS.t3575 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4153 a_6575_47204# a_6545_47178# VDD.t2442 VDD.t2441 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4154 VSS.t3695 a_765_45546.t11 a_380_45546# VSS.t3694 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4155 VSS.t2283 a_327_44734# a_501_45348# VSS.t2282 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4156 a_104_43370# a_n699_43396# VSS.t2485 VSS.t2484 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4157 VDD.t3335 a_22959_42860# a_14097_32519.t0 VDD.t3334 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4158 a_n2293_42282# a_3357_43084.t6 VDD.t2048 VDD.t2047 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4159 VSS.t2039 a_6171_42473# a_5379_42460# VSS.t1055 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4160 a_3935_42891# a_2382_45260# a_3935_43218# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4161 VSS.t1016 a_9067_47204# DATA[4].t5 VSS.t1015 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD.t414 a_8145_46902# a_8035_47026# VDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4163 VDD.t695 a_n863_45724# a_327_44734# VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4164 C10_P_btm.t27 a_n4315_30879.t21 VREF.t45 VDD.t2081 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4165 a_17141_43172# a_n1059_45260.t23 a_16795_42852# VSS.t2771 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4166 VDD.t1458 a_9127_43156# a_5891_43370.t0 VDD.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4167 a_15433_44458# a_9482_43914# VDD.t1288 VDD.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4168 VSS.t2792 a_10193_42453.t15 a_11897_42308# VSS.t2791 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4169 VSS.t1757 a_4791_45118.t13 a_5066_45546# VSS.t1756 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4170 VDD.t1116 a_5691_45260# a_n2109_47186.t0 VDD.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4171 VDD.t2196 a_n1550_35448# a_n2002_35448# VDD.t2195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4172 VSS.t3152 VDD.t3823 VSS.t3151 VSS.t3150 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4173 VDD.t943 a_1983_46706# a_n2661_46098# VDD.t942 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4174 a_15227_46910# a_15368_46634# VDD.t2764 VDD.t2763 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4175 a_18753_44484# a_18374_44850# a_18681_44484# VSS.t1947 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4176 a_15486_42560# a_15803_42450# a_15761_42308# VSS.t2259 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X4177 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD.t2773 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4178 a_6682_46987# a_n971_45724.t28 VDD.t1932 VDD.t1931 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4179 a_n1079_45724# a_n755_45592.t17 VDD.t3447 VDD.t3446 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4180 a_12429_44172# a_12861_44030.t23 VSS.t2984 VSS.t2983 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X4181 a_1568_43370# a_1847_42826# VSS.t2250 VSS.t2249 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4182 VSS.t3198 VDD.t3779 VSS.t3197 VSS.t3196 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4183 VSS.t2857 a_n1794_35082.t19 a_n1696_34930.t4 VSS.t2856 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4184 VSS.t3162 VDD.t3767 VSS.t3161 VSS.t3160 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4185 a_10890_34112.t3 a_18194_34908.t9 VSS.t3700 VSS.t3699 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4186 VDD.t913 a_7227_42308# a_6123_31319.t1 VDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4187 VSS.t1264 a_1123_46634# a_584_46384.t7 VSS.t1263 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4188 a_3457_43396# a_3232_43370.t21 a_3626_43646.t3 VSS.t2830 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4189 a_7174_31319.t2 a_20107_42308# VSS.t1965 VSS.t1964 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4190 a_8952_43230# a_8037_42858# a_8605_42826# VSS.t1469 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4191 VSS.t205 a_167_45260# a_n37_45144# VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4192 a_13490_45067# a_9482_43914# VDD.t1299 VDD.t1298 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4193 a_4181_44734# a_3090_45724.t21 a_n2497_47436# VDD.t1826 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4194 VSS.t3528 a_6171_45002.t5 a_11909_44484# VSS.t3527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4195 VSS.t860 a_n2302_39866# a_n4209_39590.t5 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4196 a_33_46660# a_n133_46660# VSS.t1954 VSS.t1953 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4197 a_16388_46812# a_17957_46116# VSS.t3453 VSS.t3452 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X4198 VDD.t2293 a_3218_45724# a_3175_45822# VDD.t2292 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4199 a_8283_46482# a_n1151_42308.t19 a_7920_46348# VSS.t1663 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4200 a_8953_45002# CLK.t7 VDD.t3701 VDD.t3700 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4201 VSS.t357 a_n809_44244# a_n755_45592.t7 VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4202 VDD.t730 a_15279_43071# a_14579_43548# VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4203 VDD.t891 a_16763_47508# a_5807_45002# VDD.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 VDD.t2724 a_310_45028# a_509_45822# VDD.t2723 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4205 a_n23_47502# a_n971_45724.t20 VDD.t1922 VDD.t1921 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4206 a_n1099_45572# a_n971_45724.t25 VDD.t1928 VDD.t1927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X4207 VDD.t3317 a_10903_43370.t16 a_10907_45822# VDD.t3316 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4208 a_3935_43218# a_3681_42891# VSS.t497 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4209 a_14949_46494# a_13759_46122# a_14840_46494# VSS.t1416 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4210 a_11599_46634.t1 a_15682_46116# VDD.t1086 VDD.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4211 a_6851_47204# a_6491_46660# VSS.t1985 VSS.t1984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4212 a_13556_45296# a_6755_46942# VDD.t2846 VDD.t2845 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4213 VDD.t2079 a_n4315_30879.t19 a_n4334_40480# VDD.t2078 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4214 VSS.t3591 a_15227_44166.t10 a_14539_43914# VSS.t3590 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X4215 a_19987_42826# a_18494_42460# a_20356_42852# VDD.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X4216 a_n2833_47464# a_n2497_47436# VDD.t2641 VDD.t2640 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4217 a_3524_46660# a_2609_46660# a_3177_46902# VSS.t1476 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4218 a_n4209_39304.t7 a_n2302_39072# VSS.t223 VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4219 VSS.t2011 a_22223_47212# a_21588_30879.t3 VSS.t2010 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4220 VSS.t2754 a_6151_47436.t10 a_6229_45572# VSS.t2753 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X4221 a_18533_43940# a_13661_43548.t17 VDD.t3120 VDD.t3119 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4222 a_14205_43396# a_13667_43396# VDD.t2566 VDD.t2565 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4223 VREF.t66 a_n3565_39590.t9 C8_P_btm.t2 VDD.t3609 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4224 VCM.t51 a_3422_30871.t12 VDAC_N.t2 VSS.t3514 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4225 VDD.t30 a_949_44458# a_n2438_43548.t1 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4226 a_n4064_37440.t2 a_n4334_37440# VDD.t1706 VDD.t1705 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4227 a_16377_45572# a_16333_45814# a_16211_45572# VSS.t2559 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4228 a_4646_46812.t28 a_6298_44484# VSS.t829 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X4229 a_10044_46482# a_n743_46660.t5 a_9823_46155# VSS.t3555 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4230 a_19113_45348# a_18911_45144# a_3090_45724.t4 VSS.t2488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4231 VSS.t1102 a_13720_44458# a_12607_44458# VSS.t1101 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4232 a_n2860_37984# a_n2956_38216.t5 a_n2946_37984# VDD.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4233 a_2266_47570# a_n971_45724.t19 VSS.t1695 VSS.t1694 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4234 a_5837_43396# a_5111_44636# a_5147_45002# VSS.t913 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4235 a_5934_30871.t1 a_8791_42308# VDD.t1402 VDD.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4236 a_10861_46660# a_10227_46804.t17 VSS.t1613 VSS.t1612 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4237 VSS.t660 a_7920_46348# a_7715_46873# VSS.t659 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4238 a_14383_46116# a_10227_46804.t24 VDD.t1844 VDD.t1843 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4239 a_2809_45348# a_526_44458.t23 VSS.t3399 VSS.t3398 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4240 a_2905_42968# a_742_44458# VSS.t793 VSS.t792 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4241 a_6540_46812# a_6755_46942# a_6682_46987# VDD.t2840 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4242 a_6709_45028# a_6431_45366# VSS.t1072 VSS.t1071 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4243 a_8953_45002# CLK.t4 VSS.t3629 VSS.t3628 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4244 VSS.t1112 a_18494_42460# a_20193_45348# VSS.t1111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4245 a_n2442_46660.t0 a_n2472_46634# VDD.t574 VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4246 C7_P_btm.t4 EN_VIN_BSTR_P.t12 VIN_P.t3 VSS.t3564 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4247 a_13249_42308# a_13070_42354# VSS.t1070 VSS.t1069 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4248 a_n1991_42858# a_n2157_42858# VSS.t1124 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4249 VDD.t153 VSS.t3734 VDD.t152 VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4250 VDD.t1090 a_15682_46116# a_11599_46634.t7 VDD.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4251 a_13348_45260# a_12891_46348# a_13490_45067# VDD.t1640 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4252 VREF_GND.t2 a_n4064_39616.t13 C9_P_btm.t2 VSS.t2849 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4253 a_17061_44484# a_11691_44458.t5 VSS.t2887 VSS.t2886 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4254 comp_n a_1169_39043# VDD.t358 VDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4255 VDD.t146 VSS.t3760 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4256 VDD.t2788 a_18443_44721# a_18374_44850# VDD.t2787 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4257 VDD.t139 VSS.t3720 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4258 a_1512_43396# a_n443_46116.t17 a_1209_43370# VSS.t3050 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4259 VDD.t3605 a_n3565_39304.t10 a_n3690_39392# VDD.t3228 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4260 VDD.t596 a_22591_44484# a_17730_32519.t0 VDD.t595 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4261 VDD.t3482 a_22581_37893# a_22537_39537# VDD.t3481 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4262 VDD.t2410 a_n2002_35448# SMPL_ON_P.t0 VDD.t2409 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4263 VSS.t2258 a_15803_42450# a_15764_42576# VSS.t2257 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4264 a_11901_46660# a_11735_46660# VSS.t457 VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4265 a_21076_30879.t2 a_22959_46660# VSS.t763 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4266 a_3877_44458# a_3699_46634# VDD.t1058 VDD.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4267 VDD.t3081 a_n4064_39072.t8 a_n2216_39072# VDD.t2036 sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4268 a_11599_46634.t19 a_15682_46116# VSS.t874 VSS.t873 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4269 a_11691_44458.t0 a_5807_45002# VDD.t1485 VDD.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4270 a_15368_46634# a_15143_45578# VDD.t581 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X4271 VSS.t3423 a_9028_43914# a_8975_43940# VSS.t3422 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4272 a_2813_43396# a_n443_46116.t10 VSS.t3044 VSS.t3043 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X4273 C8_N_btm.t7 a_17538_32519.t5 VREF_GND.t31 VSS.t2646 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4274 a_5093_45028# a_4558_45348# a_5009_45028# VDD.t2261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4275 VSS.t2799 a_10193_42453.t22 a_13921_42308# VSS.t2798 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4276 a_15597_42852# a_15567_42826# a_15095_43370# VDD.t2652 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X4277 a_2553_47502# a_n971_45724.t14 VDD.t1918 VDD.t1917 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4278 VDD.t1369 a_13059_46348# a_12839_46116# VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4279 C10_N_btm.t14 a_22612_30879.t10 VREF.t18 VDD.t1945 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4280 a_3823_42558# a_3065_45002# a_3905_42308# VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4281 VDD.t3475 a_526_44458.t28 a_5193_42852# VDD.t3474 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4282 VSS.t501 a_1667_45002# a_n863_45724# VSS.t500 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4283 a_1307_43914.t0 a_2779_44458# VDD.t671 VDD.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4284 VDD.t2521 a_n3690_38528# a_n3420_38528.t0 VDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4285 VDD.t1392 a_21177_47436# a_20990_47178# VDD.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4286 a_16855_45546# a_16327_47482.t39 VDD.t3354 VDD.t3353 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4287 a_5495_43940# a_5244_44056# VDD.t1150 VDD.t1149 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4288 VDD.t1339 a_5815_47464# a_n1613_43370.t1 VDD.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4289 VSS.t2539 a_19787_47423# a_19594_46812# VSS.t2538 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4290 VDD.t1528 a_22365_46825# a_20202_43084# VDD.t1527 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4291 a_5063_47570# a_4915_47217.t11 a_4700_47436# VSS.t3689 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4292 a_n1736_46482# a_n1853_46287# VSS.t2098 VSS.t2097 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4293 VDD.t462 a_11459_47204# DATA[5].t1 VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4294 a_11322_45546# a_11823_42460.t12 VSS.t3534 VSS.t3533 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4295 a_19787_47423# START.t1 VSS.t2611 VSS.t2610 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4296 a_3754_39466# a_7754_39632# VSS.t564 sky130_fd_pr__res_high_po_0p35 l=18
X4297 a_n4251_39616# a_n4318_39768.t5 a_n4334_39616# VSS.t1664 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4298 VDD.t1462 a_9127_43156# a_9114_42852# VDD.t1461 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4299 a_10384_47026# a_9863_46634# VDD.t2514 VDD.t2513 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4300 VSS.t3218 VDD.t3788 VSS.t3217 VSS.t3216 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4301 VSS.t2360 a_11525_45546# a_11189_46129# VSS.t2359 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4302 SMPL_ON_N.t2 a_21753_35474# VDD.t1665 VDD.t1664 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4303 VSS.t3257 VDD.t3802 VSS.t3256 VSS.t3255 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4304 a_10729_43914# a_11750_44172# VDD.t2750 VDD.t2749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4305 a_4921_42308# a_n913_45002.t28 a_4933_42558# VDD.t2967 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4306 VSS.t2289 a_n23_47502# a_n89_47570# VSS.t2288 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4307 a_20528_46660# a_20411_46873# VSS.t2033 VSS.t2032 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4308 VSS.t2348 a_8568_45546# a_8162_45546# VSS.t2347 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4309 a_13657_42558# a_13259_45724.t23 VDD.t241 VDD.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4310 VDD.t96 VSS.t3753 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4311 VSS.t2657 a_4223_44672.t6 a_5205_44484# VSS.t2656 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4312 a_18005_44484# a_17970_44736# a_17767_44458# VSS.t1946 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4313 a_13837_43396# a_13259_45724.t22 a_13749_43396# VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4314 a_19177_43646# a_17339_46660# VDD.t1692 VDD.t1691 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X4315 a_196_42282# a_375_42282# VSS.t1949 VSS.t1948 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4316 a_791_42968# a_n1059_45260.t12 VSS.t2764 VSS.t2763 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4317 VSS.t2058 a_327_47204# DATA[0].t7 VSS.t2057 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4318 a_11309_47204# a_11031_47542# VSS.t2298 VSS.t2297 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4319 VSS.t2913 a_4646_46812.t38 a_7871_42858# VSS.t2912 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4320 VSS.t1146 a_5815_47464# a_n1613_43370.t4 VSS.t1145 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4321 a_n23_45546# a_n356_45724# VSS.t3443 VSS.t3442 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4322 a_18691_45572# a_18175_45572# a_18596_45572# VSS.t2088 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4323 a_9885_42558# a_9290_44172.t11 VDD.t3264 VDD.t3263 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4324 VSS.t1381 a_4700_47436# a_3785_47178# VSS.t1380 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4325 a_5700_37509.t10 VDAC_N.t19 a_8912_37509.t27 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4326 a_4361_42308.t1 a_3823_42558# VSS.t1238 VSS.t1237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4327 VDD.t1132 a_n2840_46634# a_n2956_39768.t0 VDD.t1131 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4328 a_4817_46660# a_4651_46660# VSS.t2217 VSS.t2216 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4329 VDD.t2597 a_13635_43156# a_13622_42852# VDD.t2596 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4330 VDD.t3748 a_n2438_43548.t43 a_n2157_42858# VDD.t3747 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4331 a_8415_44056# a_5343_44458# a_8333_44056# VDD.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4332 a_8912_37509.t1 VDAC_P.t12 a_5088_37509.t12 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4333 VSS.t3466 a_1307_43914.t25 a_4156_43218# VSS.t3465 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4334 a_n1699_44726# a_n1917_44484# VDD.t330 VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4335 a_1525_44260# a_1467_44172# a_1115_44172# VSS.t3456 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4336 VDD.t718 a_n2946_39866# a_n3565_39590.t0 VDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4337 a_14976_45028# a_14797_45144# a_15060_45348# VSS.t2464 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X4338 VSS.t3143 VDD.t3820 VSS.t3142 VSS.t3141 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4339 a_2324_44458.t30 a_8953_45002# VSS.t318 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4340 VSS.t3183 VDD.t3774 VSS.t3182 VSS.t3181 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4341 a_n3565_39304.t3 a_n2946_39072# VDD.t2161 VDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4342 VSS.t2557 a_15959_42545# a_15890_42674# VSS.t2556 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4343 a_n2312_39304.t2 a_n1920_47178# VSS.t981 VSS.t980 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4344 VDD.t600 a_15682_43940# a_11967_42832.t7 VDD.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4345 VIN_N.t12 EN_VIN_BSTR_N.t12 C7_N_btm.t0 VSS.t2919 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4346 VDD.t2052 a_1666_39587.t6 a_1666_39043.t1 VDD.t2051 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X4347 VDD.t2547 a_n3690_37440# a_n3420_37440.t0 VDD.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4348 VSS.t1526 a_21363_45546# a_21297_45572# VSS.t1525 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4349 VDD.t1231 a_n452_44636# a_n2129_44697# VDD.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4350 a_19443_46116# a_18819_46122# a_19335_46494# VDD.t2464 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4351 VDD.t1184 a_7112_43396# a_7287_43370# VDD.t1183 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4352 a_310_45028# a_n37_45144# VSS.t2450 VSS.t2449 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4353 VDD.t1100 a_5111_44636# a_5518_44484# VDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X4354 a_17719_45144# a_17613_45144# VSS.t3455 VSS.t3454 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4355 a_17499_43370# a_16327_47482.t11 VDD.t3405 VDD.t3404 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4356 VDD.t452 a_12563_42308# a_5534_30871.t0 VDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4357 VSS.t2866 a_13747_46662.t8 a_19466_46812# VSS.t2865 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4358 a_14112_44734# a_768_44030.t19 a_13857_44734# VDD.t3689 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4359 VSS.t702 a_n2946_38778# a_n3565_38502.t4 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 a_n357_42282.t1 a_21356_42826# VDD.t2792 VDD.t2791 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4361 VDD.t199 VSS.t3708 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4362 VDD.t3301 a_3483_46348.t22 a_15037_43940# VDD.t3300 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4363 VCM.t11 a_4190_30871.t12 C10_P_btm.t1 VSS.t2810 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4364 a_5700_37509.t11 VDAC_N.t23 a_8912_37509.t31 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4365 VDD.t2599 a_13635_43156# a_9290_44172.t1 VDD.t2598 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4366 VDD.t794 a_13487_47204# a_768_44030.t0 VDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4367 a_14097_32519.t2 a_22959_42860# VSS.t3277 VSS.t2178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4368 a_3094_47570# a_2905_45572# VSS.t2365 VSS.t2364 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4369 a_8270_45546# a_n237_47217.t14 VSS.t3037 VSS.t3036 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 a_8781_46436# a_8199_44636# a_8034_45724# VSS.t784 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4371 VDD.t220 VSS.t3722 VDD.t219 VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4372 VSS.t2824 a_3232_43370.t12 a_11541_44484# VSS.t2823 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4373 DATA[4].t7 a_9067_47204# VSS.t1012 VSS.t1011 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4374 a_20841_46902# a_20623_46660# VSS.t2597 VSS.t2596 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4375 a_13527_45546# a_12861_44030.t28 VSS.t2990 VSS.t2989 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4376 a_10533_42308# a_7499_43078# VSS.t340 VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 a_17896_45144# a_16922_45042# a_17801_45144# VDD.t2854 sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X4378 DATA[1].t7 a_1431_47204# VSS.t1858 VSS.t1857 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4379 a_18817_42826# a_18599_43230# VSS.t2296 VSS.t2295 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4380 a_104_43370# a_n699_43396# VDD.t2742 VDD.t2741 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4381 C10_P_btm.t18 a_n4315_30879.t10 VREF.t36 VDD.t2070 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4382 a_16211_45572# a_15765_45572# a_16115_45572# VSS.t2232 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4383 VDD.t2897 a_4223_44672.t5 a_4181_44734# VDD.t2896 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4384 VSS.t989 a_20835_44721# a_20766_44850# VSS.t988 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4385 a_19741_43940# a_19478_44306# a_19328_44172# VDD.t2757 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4386 VDD.t3087 a_13747_46662.t6 a_14495_45572# VDD.t3086 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4387 a_2487_47570# a_2063_45854.t17 a_2124_47436# VSS.t1645 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4388 VSS.t3571 a_10809_44734.t6 a_22959_46124# VSS.t1725 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4389 a_11967_42832.t12 a_15682_43940# VDD.t626 VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 C10_N_btm.t30 a_18114_32519.t10 VREF_GND.t12 VSS.t2653 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4391 VSS.t1936 a_7754_38470# a_6886_37412# VSS.t1935 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4392 VSS.t1891 a_20567_45036# a_12549_44172.t3 VSS.t1890 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4393 a_21359_45002# a_21513_45002# VDD.t3346 VDD.t3345 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4394 a_18451_43940# a_18579_44172# a_18533_44260# VSS.t2426 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4395 a_13904_45546# a_13249_42308# a_14033_45822# VDD.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X4396 VSS.t2893 a_13661_43548.t10 a_18587_45118# VSS.t2892 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4397 a_6547_43396# a_6031_43396# a_6452_43396# VSS.t2186 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
R0 a_13259_45724.n20 a_13259_45724.n19 589.152
R1 a_13259_45724.t18 a_13259_45724.t11 378.255
R2 a_13259_45724.n13 a_13259_45724.t21 334.723
R3 a_13259_45724.n7 a_13259_45724.t9 334.723
R4 a_13259_45724.n4 a_13259_45724.t18 332.308
R5 a_13259_45724.n19 a_13259_45724.n0 289.462
R6 a_13259_45724.n6 a_13259_45724.t23 256.716
R7 a_13259_45724.n10 a_13259_45724.t8 241.536
R8 a_13259_45724.n9 a_13259_45724.t4 241.536
R9 a_13259_45724.n1 a_13259_45724.t10 231.835
R10 a_13259_45724.n3 a_13259_45724.n1 206.881
R11 a_13259_45724.n13 a_13259_45724.t5 206.19
R12 a_13259_45724.n7 a_13259_45724.t22 206.19
R13 a_13259_45724.n2 a_13259_45724.t16 201.369
R14 a_13259_45724.n11 a_13259_45724.n9 193.643
R15 a_13259_45724.n8 a_13259_45724.n6 192.037
R16 a_13259_45724.n17 a_13259_45724.n5 179.357
R17 a_13259_45724.n3 a_13259_45724.n2 179.332
R18 a_13259_45724.n14 a_13259_45724.n13 177.531
R19 a_13259_45724.n8 a_13259_45724.n7 172.637
R20 a_13259_45724.n11 a_13259_45724.n10 170.416
R21 a_13259_45724.n10 a_13259_45724.t13 169.237
R22 a_13259_45724.n9 a_13259_45724.t15 169.237
R23 a_13259_45724.n16 a_13259_45724.n15 167.631
R24 a_13259_45724.n6 a_13259_45724.t19 161.275
R25 a_13259_45724.n1 a_13259_45724.t6 157.07
R26 a_13259_45724.n5 a_13259_45724.t20 142.994
R27 a_13259_45724.n15 a_13259_45724.t14 137.177
R28 a_13259_45724.n2 a_13259_45724.t12 132.282
R29 a_13259_45724.n5 a_13259_45724.t7 126.927
R30 a_13259_45724.n15 a_13259_45724.t17 121.109
R31 a_13259_45724.n0 a_13259_45724.t3 38.5719
R32 a_13259_45724.n0 a_13259_45724.t2 38.5719
R33 a_13259_45724.t0 a_13259_45724.n20 26.5955
R34 a_13259_45724.n20 a_13259_45724.t1 26.5955
R35 a_13259_45724.n18 a_13259_45724.n17 17.4579
R36 a_13259_45724.n19 a_13259_45724.n18 17.2128
R37 a_13259_45724.n12 a_13259_45724.n8 11.7999
R38 a_13259_45724.n4 a_13259_45724.n3 9.27935
R39 a_13259_45724.n16 a_13259_45724.n14 9.1023
R40 a_13259_45724.n17 a_13259_45724.n16 4.97577
R41 a_13259_45724.n12 a_13259_45724.n11 4.5005
R42 a_13259_45724.n14 a_13259_45724.n12 4.4222
R43 a_13259_45724.n18 a_13259_45724.n4 1.99363
R44 VSS.n4892 VSS.t1452 1.14713e+06
R45 VSS.n4111 VSS.t963 1.03856e+06
R46 VSS.n3994 VSS.n3993 461132
R47 VSS.n4299 VSS.n3874 39462.7
R48 VSS.n4168 VSS.n4167 30027
R49 VSS.n3989 VSS.n3970 27875.5
R50 VSS.n3871 VSS.n3815 27875.5
R51 VSS.n3989 VSS.n3971 27736.4
R52 VSS.n3815 VSS.n3814 27736.4
R53 VSS.n3977 VSS.n3970 27701.7
R54 VSS.n3871 VSS.n3817 27701.7
R55 VSS.n3977 VSS.n3971 27562.6
R56 VSS.n3817 VSS.n3814 27562.6
R57 VSS.n4817 VSS.n4801 22537
R58 VSS.n4206 VSS.n4203 19062.6
R59 VSS.n4280 VSS.n4203 19062.6
R60 VSS.n4279 VSS.n4206 19062.6
R61 VSS.n4280 VSS.n4279 19062.6
R62 VSS.n3990 VSS.n3969 18180.1
R63 VSS.n4801 VSS.n4800 15727.3
R64 VSS.n3993 VSS.t3153 15408.2
R65 VSS.n3840 VSS.n3839 11539.6
R66 VSS.n4228 VSS.n1774 8128.61
R67 VSS.n4300 VSS.n4299 7785.2
R68 VSS.n4226 VSS.n4222 6361.94
R69 VSS.n4222 VSS.n4215 6361.94
R70 VSS.n3996 VSS.t2389 5807.56
R71 VSS.t1548 VSS.t1925 5523.02
R72 VSS.n4231 VSS.n4226 5446.47
R73 VSS.n4217 VSS.n4215 5446.47
R74 VSS.n3993 VSS.n3992 5420.59
R75 VSS.n4255 VSS.n4252 5419.2
R76 VSS.n4298 VSS.n3875 5342.18
R77 VSS.n4298 VSS.n3877 5342.18
R78 VSS.n3876 VSS.n3875 5342.18
R79 VSS.n3877 VSS.n3876 5342.18
R80 VSS.n4800 VSS.n4799 5197.83
R81 VSS.n4229 VSS.n4228 4819.77
R82 VSS.n4035 VSS.t96 4752.56
R83 VSS.n4881 VSS.n1732 4345.59
R84 VSS.n1734 VSS.n1732 4345.59
R85 VSS.n4868 VSS.n1743 4345.59
R86 VSS.n1748 VSS.n1743 4345.59
R87 VSS.n4025 VSS.n3954 4345.59
R88 VSS.n4025 VSS.n4024 4345.59
R89 VSS.n4146 VSS.n3950 4345.59
R90 VSS.n4050 VSS.n3950 4345.59
R91 VSS.n4799 VSS.t1842 4286.04
R92 VSS.n4173 VSS.n3915 4154.38
R93 VSS.n4196 VSS.n3915 4154.38
R94 VSS.n4266 VSS.n4257 3743
R95 VSS.n4268 VSS.n4257 3743
R96 VSS.n4282 VSS.n3908 3743
R97 VSS.n4282 VSS.n3909 3743
R98 VSS.n4275 VSS.n4208 3685.06
R99 VSS.n4251 VSS.n4208 3685.06
R100 VSS.n4275 VSS.n4209 3685.06
R101 VSS.n4251 VSS.n4209 3685.06
R102 VSS.t3234 VSS.n4913 3683.8
R103 VSS.n3992 VSS.n3969 3578.95
R104 VSS.n3874 VSS.n1755 3235.7
R105 VSS.n4228 VSS.t1932 3221.17
R106 VSS.n1744 VSS.n1739 3128.82
R107 VSS.n1744 VSS.n1738 3128.82
R108 VSS.n4878 VSS.n1733 3128.82
R109 VSS.n4878 VSS.n1735 3128.82
R110 VSS.n4042 VSS.n3949 3128.82
R111 VSS.n4042 VSS.n3951 3128.82
R112 VSS.n4039 VSS.n4038 3128.82
R113 VSS.n4038 VSS.n3953 3128.82
R114 VSS.n4857 VSS.n1755 3082.34
R115 VSS.n4859 VSS.n1755 3082.34
R116 VSS.n4015 VSS.n3966 3082.34
R117 VSS.n4018 VSS.n3966 3082.34
R118 VSS.t3244 VSS.t2293 2948.87
R119 VSS.n4200 VSS.n3911 2914.44
R120 VSS.t3683 VSS.t3150 2902.25
R121 VSS.t3150 VSS.t1638 2902.25
R122 VSS.n4170 VSS.n4169 2885.47
R123 VSS.n4200 VSS.n3910 2885.47
R124 VSS.n4170 VSS.n3933 2821.74
R125 VSS.n492 VSS.t3216 2714.18
R126 VSS.t3684 VSS.t3260 2704.11
R127 VSS.t1335 VSS.t1196 2698.28
R128 VSS.t1938 VSS.t3244 2698.28
R129 VSS.t2412 VSS.t3184 2692.45
R130 VSS.n4864 VSS.n1750 2690.47
R131 VSS.n4864 VSS.n1749 2690.47
R132 VSS.n4032 VSS.n3962 2690.47
R133 VSS.n3962 VSS.n3959 2690.47
R134 VSS.n3832 VSS.n3827 2549.41
R135 VSS.n3832 VSS.n1725 2549.41
R136 VSS.n3837 VSS.n1723 2549.41
R137 VSS.n4894 VSS.n1723 2549.41
R138 VSS.t1397 VSS.t481 2438.55
R139 VSS.t3184 VSS.n265 2412.72
R140 VSS.n4913 VSS.n4912 2402.01
R141 VSS.n4912 VSS.n4911 2402.01
R142 VSS.n4911 VSS.n4910 2402.01
R143 VSS.t542 VSS.t3166 2377.01
R144 VSS.t1427 VSS.t800 2360.15
R145 VSS.t3196 VSS.t3108 2326.44
R146 VSS.n4821 VSS.n4819 2192
R147 VSS.n3843 VSS.n3822 2192
R148 VSS.t2192 VSS.t2751 2185.43
R149 VSS.n4802 VSS.n1773 2174.6
R150 VSS.n3825 VSS.n3824 2174.6
R151 VSS.t2950 VSS.t628 2173.77
R152 VSS.t1080 VSS.t2612 2167.95
R153 VSS.t3114 VSS.t3428 2167.95
R154 VSS.t1458 VSS.t2069 2149.43
R155 VSS.t2447 VSS.t2341 2149.43
R156 VSS.t903 VSS.t2385 2149.43
R157 VSS.n4910 VSS.n4909 2136.38
R158 VSS.n4230 VSS.n4216 2126.44
R159 VSS.n4236 VSS.n4216 2126.44
R160 VSS.t1111 VSS.t692 2115.71
R161 VSS.t118 VSS.t2499 2115.71
R162 VSS.t461 VSS.t2832 2115.71
R163 VSS.t181 VSS.t1799 2065.13
R164 VSS.n3839 VSS.n1719 2019.64
R165 VSS.t3070 VSS.t3155 1989.27
R166 VSS.n4262 VSS.n4259 1970
R167 VSS.n4262 VSS.n4258 1970
R168 VSS.t3129 VSS.t290 1963.98
R169 VSS.n1444 VSS.t2441 1963.98
R170 VSS.t84 VSS.t3190 1963.98
R171 VSS.t2180 VSS.t3135 1963.98
R172 VSS.t112 VSS.t3105 1963.98
R173 VSS.t218 VSS.t3225 1963.98
R174 VSS.t276 VSS.t3144 1963.98
R175 VSS.t3228 VSS.t760 1963.98
R176 VSS.t935 VSS.t3120 1963.98
R177 VSS.t3219 VSS.t173 1955.56
R178 VSS.t3193 VSS.t1280 1955.56
R179 VSS.t3166 VSS.t3196 1938.7
R180 VSS.t1041 VSS.t753 1930.27
R181 VSS.t3030 VSS.t553 1888.21
R182 VSS.n4184 VSS.n3923 1877.29
R183 VSS.t3260 VSS.n199 1876.56
R184 VSS.n1758 VSS.n1757 1857.31
R185 VSS.n1757 VSS.n1754 1857.31
R186 VSS.n3967 VSS.n3961 1857.31
R187 VSS.n3968 VSS.n3967 1857.31
R188 VSS.n4299 VSS.t1548 1849.37
R189 VSS.t2079 VSS.t1285 1829.12
R190 VSS.t3642 VSS.t3231 1786.97
R191 VSS.n4184 VSS.n3924 1784.59
R192 VSS.t1478 VSS.t922 1778.54
R193 VSS.n4266 VSS.n4259 1773
R194 VSS.n4259 VSS.n3908 1773
R195 VSS.n4268 VSS.n4258 1773
R196 VSS.n4258 VSS.n3909 1773
R197 VSS.t1524 VSS.t1527 1753.26
R198 VSS.t1152 VSS.t1301 1753.26
R199 VSS.t1895 VSS.t726 1753.26
R200 VSS.t1477 VSS.t867 1753.26
R201 VSS.t703 VSS.t1540 1744.83
R202 VSS.t2883 VSS.t534 1744.83
R203 VSS.t1780 VSS.t1342 1677.39
R204 VSS.t159 VSS.t2640 1677.39
R205 VSS.t272 VSS.t1382 1643.44
R206 VSS.t171 VSS.t64 1626.82
R207 VSS.t3126 VSS.t1762 1620.13
R208 VSS.t2214 VSS.t3114 1620.13
R209 VSS.t332 VSS.t1465 1618.39
R210 VSS.t2095 VSS.t3092 1618.39
R211 VSS.t2778 VSS.t2662 1618.39
R212 VSS.t1413 VSS.t1411 1618.39
R213 VSS.t1925 VSS.n3875 1615.98
R214 VSS.t1932 VSS.n3877 1615.98
R215 VSS.t919 VSS.t1886 1609.96
R216 VSS.t2486 VSS.t2784 1609.96
R217 VSS.t511 VSS.t377 1601.53
R218 VSS.t3584 VSS.t2936 1601.53
R219 VSS.t1091 VSS.t120 1601.53
R220 VSS.t1665 VSS.t2030 1593.1
R221 VSS.t2172 VSS.t1077 1593.1
R222 VSS.t968 VSS.t972 1593.1
R223 VSS.t2286 VSS.t1784 1593.1
R224 VSS.t1231 VSS.t1882 1593.1
R225 VSS.t1222 VSS.t2051 1593.1
R226 VSS.t2564 VSS.t1732 1593.1
R227 VSS.t411 VSS.t974 1593.1
R228 VSS.t1104 VSS.t1723 1593.1
R229 VSS.t1958 VSS.t1542 1593.1
R230 VSS.t1725 VSS.t1473 1593.1
R231 VSS.t1198 VSS.t2125 1593.1
R232 VSS.t389 VSS.t1791 1593.1
R233 VSS.t1682 VSS.t3653 1584.67
R234 VSS.t579 VSS.t1682 1584.67
R235 VSS.t2387 VSS.t1772 1584.67
R236 VSS.t2934 VSS.t4 1584.67
R237 VSS.t3272 VSS.t739 1584.67
R238 VSS.t913 VSS.t1292 1584.67
R239 VSS.t3669 VSS.t1736 1584.67
R240 VSS.t867 VSS.t1667 1584.67
R241 VSS.t3671 VSS.t2614 1584.67
R242 VSS.t2704 VSS.t2793 1576.25
R243 VSS.t3141 VSS.t1063 1576.25
R244 VSS.t1274 VSS.t2132 1567.82
R245 VSS.t3108 VSS.t2869 1567.82
R246 VSS.n4242 VSS.n4213 1564.22
R247 VSS.n4242 VSS.n4214 1564.22
R248 VSS.n4244 VSS.n4214 1564.22
R249 VSS.n4244 VSS.n4213 1564.22
R250 VSS.t2948 VSS.t3594 1550.96
R251 VSS.t3636 VSS.t6 1550.96
R252 VSS.n548 VSS.t1265 1550.96
R253 VSS.t3422 VSS.t3492 1542.53
R254 VSS.t2045 VSS.t2032 1542.53
R255 VSS.t3175 VSS.t2979 1534.1
R256 VSS.t1654 VSS.t1652 1517.24
R257 VSS.t3471 VSS.t1293 1517.24
R258 VSS.n3816 VSS.n1774 1497.06
R259 VSS.n3976 VSS.n1774 1495.7
R260 VSS.n3833 VSS.n3828 1494.88
R261 VSS.n3833 VSS.n1724 1494.88
R262 VSS.t986 VSS.t1509 1486.09
R263 VSS.n4912 VSS.t3129 1483.52
R264 VSS.n5376 VSS.t3190 1483.52
R265 VSS.n4910 VSS.t3135 1483.52
R266 VSS.n5376 VSS.t3105 1483.52
R267 VSS.n4911 VSS.t3225 1483.52
R268 VSS.n5376 VSS.t3144 1483.52
R269 VSS.n4913 VSS.t3228 1483.52
R270 VSS.t3120 VSS.n5376 1483.52
R271 VSS.n2337 VSS.t858 1466.67
R272 VSS.n4255 VSS.n4254 1447.27
R273 VSS.t2574 VSS.t2079 1416.09
R274 VSS.t2478 VSS.t3582 1416.09
R275 VSS.t379 VSS.t1699 1416.09
R276 VSS.n3874 VSS.n3873 1413.27
R277 VSS.n3992 VSS.n3991 1413.27
R278 VSS.t3271 VSS.t2083 1399.23
R279 VSS.t158 VSS.t2240 1399.23
R280 VSS.t101 VSS.t2038 1399.23
R281 VSS.t2568 VSS.t565 1399.23
R282 VSS.t3250 VSS.t282 1398.68
R283 VSS.n178 VSS.t1015 1398.68
R284 VSS.t1139 VSS.t3126 1398.68
R285 VSS.t3169 VSS.t2055 1398.68
R286 VSS.t3160 VSS.t237 1398.68
R287 VSS.t2071 VSS.t385 1390.8
R288 VSS.n4193 VSS.n3916 1390.59
R289 VSS.n4193 VSS.n3917 1390.59
R290 VSS.n4173 VSS.n3933 1390.59
R291 VSS.n4196 VSS.n3911 1390.59
R292 VSS.n3925 VSS.n3919 1390.59
R293 VSS.n3925 VSS.n3920 1390.59
R294 VSS.n4178 VSS.n3929 1390.59
R295 VSS.n4178 VSS.n4177 1390.59
R296 VSS.t1405 VSS.t2362 1375.36
R297 VSS.t3432 VSS.t1697 1369.54
R298 VSS.n157 VSS.t1982 1363.71
R299 VSS.t484 VSS.t1686 1363.71
R300 VSS.t2099 VSS.t3169 1363.71
R301 VSS.t2317 VSS.t3234 1357.88
R302 VSS.t2269 VSS.t2297 1357.88
R303 VSS.t3199 VSS.t232 1352.05
R304 VSS.n3844 VSS.n1774 1348.8
R305 VSS.n4818 VSS.n1774 1348.64
R306 VSS.t3436 VSS.t1900 1340.23
R307 VSS.t1283 VSS.t1214 1340.23
R308 VSS.t2890 VSS.t1212 1340.23
R309 VSS.t1632 VSS.t1463 1340.23
R310 VSS.t2097 VSS.t1738 1340.23
R311 VSS.t532 VSS.n2205 1323.37
R312 VSS.t583 VSS.t3163 1323.37
R313 VSS.t1320 VSS.t228 1306.51
R314 VSS.t2150 VSS.t1740 1305.43
R315 VSS.t864 VSS.t1628 1299.6
R316 VSS.t1113 VSS.t2121 1299.46
R317 VSS.n1719 VSS.t1397 1298.8
R318 VSS.t755 VSS.t925 1289.66
R319 VSS.t939 VSS.t674 1281.23
R320 VSS.t737 VSS.t2377 1281.23
R321 VSS.t2822 VSS.t949 1281.23
R322 VSS.t1089 VSS.t136 1281.23
R323 VSS.t3046 VSS.t3484 1272.8
R324 VSS.t520 VSS.n4732 1272.8
R325 VSS.n4732 VSS.t224 1272.8
R326 VSS.n4733 VSS.t1183 1264.37
R327 VSS.t193 VSS.n4798 1264.37
R328 VSS.t1962 VSS.t1516 1259.07
R329 VSS.t2134 VSS.t3293 1255.94
R330 VSS.t747 VSS.t2753 1255.94
R331 VSS.t1360 VSS.t1359 1255.94
R332 VSS.t3295 VSS.t1873 1255.94
R333 VSS.t3329 VSS.t1256 1255.94
R334 VSS.t3345 VSS.t630 1255.94
R335 VSS.t2422 VSS.t3353 1255.94
R336 VSS.t1299 VSS.t1624 1255.94
R337 VSS.t617 VSS.t1598 1255.94
R338 VSS.t1604 VSS.t2267 1255.94
R339 VSS.t2892 VSS.t1356 1247.51
R340 VSS.t619 VSS.t2740 1247.51
R341 VSS.n4909 VSS.t3239 1245.01
R342 VSS.n4205 VSS.n3905 1239.46
R343 VSS.n4859 VSS.n1754 1238.21
R344 VSS.n4857 VSS.n1758 1238.21
R345 VSS.n4015 VSS.n3961 1238.21
R346 VSS.n4018 VSS.n3968 1238.21
R347 VSS.t3181 VSS.t1317 1230.65
R348 VSS.t1177 VSS.t3667 1230.65
R349 VSS.n4881 VSS.n1733 1216.76
R350 VSS.n4872 VSS.n1733 1216.76
R351 VSS.n4872 VSS.n1739 1216.76
R352 VSS.n4868 VSS.n1739 1216.76
R353 VSS.n1735 VSS.n1734 1216.76
R354 VSS.n4874 VSS.n1735 1216.76
R355 VSS.n4874 VSS.n1738 1216.76
R356 VSS.n1748 VSS.n1738 1216.76
R357 VSS.n4039 VSS.n3954 1216.76
R358 VSS.n4040 VSS.n4039 1216.76
R359 VSS.n4040 VSS.n3949 1216.76
R360 VSS.n4146 VSS.n3949 1216.76
R361 VSS.n4024 VSS.n3953 1216.76
R362 VSS.n4045 VSS.n3953 1216.76
R363 VSS.n4045 VSS.n3951 1216.76
R364 VSS.n4050 VSS.n3951 1216.76
R365 VSS.t3032 VSS.t1493 1213.79
R366 VSS.t2136 VSS.n519 1213.79
R367 VSS.t708 VSS.t705 1212.19
R368 VSS.t2034 VSS.t1324 1211.94
R369 VSS.n4231 VSS.n4230 1210.97
R370 VSS.n4236 VSS.n4217 1210.97
R371 VSS.n5375 VSS.n5374 1198.25
R372 VSS.n5313 VSS.n117 1198.25
R373 VSS.n5265 VSS.n138 1198.25
R374 VSS.n5218 VSS.n157 1198.25
R375 VSS.n5169 VSS.n178 1198.25
R376 VSS.n5117 VSS.n199 1198.25
R377 VSS.n5074 VSS.n221 1198.25
R378 VSS.n5031 VSS.n241 1198.25
R379 VSS.n4991 VSS.n265 1198.25
R380 VSS.n4915 VSS.n4914 1198.25
R381 VSS.n903 VSS.n340 1198.25
R382 VSS.n855 VSS.n368 1198.25
R383 VSS.n811 VSS.n408 1198.25
R384 VSS.n466 VSS.n439 1198.25
R385 VSS.n638 VSS.n519 1198.25
R386 VSS.n588 VSS.n548 1198.25
R387 VSS.n5449 VSS.n5377 1198.25
R388 VSS.n957 VSS.n956 1198.25
R389 VSS.n2205 VSS.n2204 1198.25
R390 VSS.n2338 VSS.n2337 1198.25
R391 VSS.n2475 VSS.n2474 1198.25
R392 VSS.n2473 VSS.n1970 1198.25
R393 VSS.n2636 VSS.n2635 1198.25
R394 VSS.n2083 VSS.n2061 1198.25
R395 VSS.n2891 VSS.n2890 1198.25
R396 VSS.n2941 VSS.n2915 1198.25
R397 VSS.n3108 VSS.n3011 1198.25
R398 VSS.n3010 VSS.n2988 1198.25
R399 VSS.n3293 VSS.n3292 1198.25
R400 VSS.n3295 VSS.n3294 1198.25
R401 VSS.n3054 VSS.n3033 1198.25
R402 VSS.n1329 VSS.n1328 1198.25
R403 VSS.n1444 VSS.n1443 1198.25
R404 VSS.n1446 VSS.n1445 1198.25
R405 VSS.n1567 VSS.n1566 1198.25
R406 VSS.n1569 VSS.n1568 1198.25
R407 VSS.n1627 VSS.n1626 1198.25
R408 VSS.n1675 VSS.n1004 1198.25
R409 VSS.n1718 VSS.n1717 1198.25
R410 VSS.n4012 VSS.n4011 1198.25
R411 VSS.n4110 VSS.n4109 1198.25
R412 VSS.n4520 VSS.n3605 1198.25
R413 VSS.n4473 VSS.n3628 1198.25
R414 VSS.n3667 VSS.n3646 1198.25
R415 VSS.n4390 VSS.n3668 1198.25
R416 VSS.n3717 VSS.n3716 1198.25
R417 VSS.n4908 VSS.n4907 1198.25
R418 VSS.n3728 VSS.n3727 1198.25
R419 VSS.n4301 VSS.n3689 1198.25
R420 VSS.n4303 VSS.n4302 1198.25
R421 VSS.n3812 VSS.n3811 1198.25
R422 VSS.n4611 VSS.n3569 1198.25
R423 VSS.n4731 VSS.n4730 1198.25
R424 VSS.n4563 VSS.n3586 1198.25
R425 VSS.n2336 VSS.n2335 1198.01
R426 VSS.n2207 VSS.n2206 1197.79
R427 VSS.n2892 VSS.n2765 1197.79
R428 VSS.n3997 VSS.t179 1196.93
R429 VSS.n726 VSS.n467 1196.63
R430 VSS.n681 VSS.n492 1194.5
R431 VSS.n2634 VSS.n2633 1194.5
R432 VSS.n2472 VSS.n2471 1194.5
R433 VSS.n3354 VSS.n2942 1194.5
R434 VSS.n3457 VSS.n2893 1194.5
R435 VSS.n1327 VSS.n1326 1194.5
R436 VSS.n1625 VSS.n1624 1194.5
R437 VSS.n1718 VSS.t1025 1188.51
R438 VSS.n3033 VSS.t1233 1188.51
R439 VSS.n1004 VSS.t2956 1180.08
R440 VSS.n1626 VSS.t2093 1180.08
R441 VSS.n1568 VSS.t41 1180.08
R442 VSS.n1568 VSS.t3094 1180.08
R443 VSS.t2049 VSS.t3202 1180.08
R444 VSS.n2061 VSS.t1988 1180.08
R445 VSS.n2205 VSS.t2420 1180.08
R446 VSS.n2336 VSS.t345 1180.08
R447 VSS.n957 VSS.t2608 1180.08
R448 VSS.n368 VSS.t1919 1180.08
R449 VSS.n519 VSS.t2875 1180.08
R450 VSS.t3673 VSS.t2206 1180.08
R451 VSS.n4733 VSS.t1551 1180.08
R452 VSS.n4798 VSS.t1734 1180.08
R453 VSS.n4254 VSS.t1507 1171.78
R454 VSS.t3172 VSS.t3219 1163.22
R455 VSS.t1097 VSS.t1522 1163.22
R456 VSS.n3839 VSS.n3838 1163.22
R457 VSS.t2466 VSS.t1950 1154.79
R458 VSS.t1907 VSS.t1618 1148.08
R459 VSS.t2024 VSS.t122 1146.36
R460 VSS.n3844 VSS.n3840 1133.58
R461 VSS.n4818 VSS.n4817 1133.58
R462 VSS.t1754 VSS.t1288 1129.5
R463 VSS.t2381 VSS.t2359 1121.07
R464 VSS.t1742 VSS.t2584 1121.07
R465 VSS.n4800 VSS.t1795 1121.07
R466 VSS.n4799 VSS.t1664 1121.07
R467 VSS.t1544 VSS.t612 1118.94
R468 VSS.t1984 VSS.t2190 1118.94
R469 VSS.t1409 VSS.t1407 1113.11
R470 VSS.t2103 VSS.t2101 1113.11
R471 VSS.t3355 VSS.t3268 1112.64
R472 VSS.t2749 VSS.t288 1112.64
R473 VSS.t1614 VSS.t1315 1112.64
R474 VSS.t1622 VSS.t2620 1112.64
R475 VSS.t1992 VSS.t3331 1112.64
R476 VSS.t1392 VSS.t3343 1112.64
R477 VSS.t3291 VSS.t3337 1112.64
R478 VSS.t2705 VSS.t3681 1107.28
R479 VSS.t2391 VSS.t663 1107.28
R480 VSS.t3578 VSS.t980 1101.46
R481 VSS.t1994 VSS.t1692 1095.79
R482 VSS.t3503 VSS.t3633 1095.63
R483 VSS.t1192 VSS.t2410 1095.63
R484 VSS.t2538 VSS.t1331 1095.63
R485 VSS.t604 VSS.t2705 1095.63
R486 VSS.t1847 VSS.t1703 1095.63
R487 VSS.n221 VSS.t3199 1072.32
R488 VSS.n199 VSS.t3250 1072.32
R489 VSS.t1031 VSS.n178 1072.32
R490 VSS.t2462 VSS.t2041 1070.5
R491 VSS.n3828 VSS.n3827 1054.53
R492 VSS.n3837 VSS.n3828 1054.53
R493 VSS.n4894 VSS.n1724 1054.53
R494 VSS.n1725 VSS.n1724 1054.53
R495 VSS.t463 VSS.t1431 1053.64
R496 VSS.t3035 VSS.t1644 1053.64
R497 VSS.t2048 VSS.t149 1053.64
R498 VSS.t150 VSS.t254 1036.78
R499 VSS.t3417 VSS.t997 1036.78
R500 VSS.t2235 VSS.t70 1028.35
R501 VSS.t1475 VSS.t1966 1028.35
R502 VSS.n5376 VSS.t3160 1025.7
R503 VSS.t560 VSS.t1870 1019.92
R504 VSS.t132 VSS.t1610 1019.92
R505 VSS.t355 VSS.t1029 1011.49
R506 VSS.t2043 VSS.t690 1011.49
R507 VSS.t3418 VSS.t656 1011.49
R508 VSS.t3038 VSS.t2424 1003.07
R509 VSS.t2016 VSS.t2128 1003.07
R510 VSS.t2014 VSS.t2709 1003.07
R511 VSS.t1239 VSS.t2114 1003.07
R512 VSS.t2174 VSS.t3357 994.636
R513 VSS.t1557 VSS.t1313 994.636
R514 VSS.t3202 VSS.t1348 994.636
R515 VSS.n3933 VSS.n3924 979.207
R516 VSS.t1762 VSS.t1892 979.073
R517 VSS.t2362 VSS.t2261 979.073
R518 VSS.t1686 VSS.t1303 979.073
R519 VSS.t1697 VSS.t2288 979.073
R520 VSS.t1311 VSS.t2560 977.779
R521 VSS.t636 VSS.n2891 977.779
R522 VSS.n5377 VSS.t2200 977.779
R523 VSS.t1181 VSS.t3022 969.35
R524 VSS.t1344 VSS.t2679 969.35
R525 VSS.t3521 VSS.t191 969.35
R526 VSS.t1719 VSS.t163 969.35
R527 VSS.t2018 VSS.t1991 967.418
R528 VSS.n3923 VSS.n3917 961.823
R529 VSS.n4177 VSS.n3924 961.823
R530 VSS.t286 VSS.t3497 960.92
R531 VSS.t1600 VSS.t3587 960.92
R532 VSS.t915 VSS.t955 952.49
R533 VSS.t3132 VSS.t2078 944.062
R534 VSS.t3222 VSS.t1378 944.062
R535 VSS.t516 VSS.t645 935.633
R536 VSS.t3283 VSS.t2420 935.633
R537 VSS.t3459 VSS.t2232 927.203
R538 VSS.t2359 VSS.t2578 927.203
R539 VSS.t2367 VSS.t2224 918.774
R540 VSS.t197 VSS.t1187 918.774
R541 VSS.t3444 VSS.t2554 918.774
R542 VSS.t1083 VSS.t1461 918.774
R543 VSS.t2409 VSS.t1945 918.774
R544 VSS.t1247 VSS.t1101 918.774
R545 VSS.t1151 VSS.t1000 918.774
R546 VSS.t2237 VSS.t1817 918.774
R547 VSS.t2044 VSS.t2213 918.774
R548 VSS.t2452 VSS.t1003 918.774
R549 VSS.t1019 VSS.t2218 918.774
R550 VSS.t1377 VSS.t1379 918.774
R551 VSS.n3916 VSS.n3910 915.471
R552 VSS.n4189 VSS.n3916 915.471
R553 VSS.n4189 VSS.n3919 915.471
R554 VSS.n4182 VSS.n3919 915.471
R555 VSS.n4182 VSS.n3929 915.471
R556 VSS.n4169 VSS.n3929 915.471
R557 VSS.n4188 VSS.n3917 915.471
R558 VSS.n4188 VSS.n3920 915.471
R559 VSS.n3928 VSS.n3920 915.471
R560 VSS.n4177 VSS.n3928 915.471
R561 VSS.n4232 VSS.n4231 915.471
R562 VSS.n4232 VSS.n4217 915.471
R563 VSS.t567 VSS.t2231 910.346
R564 VSS.t1366 VSS.t1636 910.346
R565 VSS.t575 VSS.t772 910.346
R566 VSS.t3048 VSS.t3400 910.346
R567 VSS.t230 VSS.t2427 910.346
R568 VSS.t2403 VSS.t640 910.346
R569 VSS.t1678 VSS.t2484 910.346
R570 VSS.t951 VSS.t1584 910.346
R571 VSS.t908 VSS.t2046 910.346
R572 VSS.t3391 VSS.t1043 910.346
R573 VSS.t1045 VSS.t3450 910.346
R574 VSS.t2469 VSS.t1558 910.346
R575 VSS.t453 VSS.t1562 910.346
R576 VSS.t2464 VSS.t2895 901.917
R577 VSS.t2346 VSS.t3379 901.917
R578 VSS.n3870 VSS.n3869 894.395
R579 VSS.n3980 VSS.n3979 894.212
R580 VSS.t1550 VSS.t1103 893.487
R581 VSS.t1240 VSS.t1436 893.487
R582 VSS.t2473 VSS.t995 893.487
R583 VSS.n3923 VSS.n3911 886.5
R584 VSS.t931 VSS.t152 885.058
R585 VSS.t2313 VSS.t451 885.058
R586 VSS.t2825 VSS.t751 876.629
R587 VSS.t653 VSS.t2966 876.629
R588 VSS.t325 VSS.t859 876.629
R589 VSS.t486 VSS.t2544 876.629
R590 VSS.t456 VSS.t1639 876.629
R591 VSS.n3865 VSS.n3819 871.289
R592 VSS.n3978 VSS.n3973 871.111
R593 VSS.n4285 VSS.n3905 870.4
R594 VSS.t3297 VSS.t710 868.345
R595 VSS.n3981 VSS.n3972 867.322
R596 VSS.n3863 VSS.n3818 867.322
R597 VSS.t1864 VSS.n241 862.518
R598 VSS.n241 VSS.t706 862.518
R599 VSS.n138 VSS.t2148 862.518
R600 VSS.n117 VSS.t1851 862.518
R601 VSS.t3053 VSS.t200 859.77
R602 VSS.t2942 VSS.t2985 859.77
R603 VSS.t1439 VSS.t2867 859.77
R604 VSS.t2019 VSS.t1713 859.77
R605 VSS.t1608 VSS.t2372 859.77
R606 VSS.t2378 VSS.t3036 859.77
R607 VSS.t2257 VSS.t720 858.456
R608 VSS.t6 VSS.t407 851.341
R609 VSS.t3247 VSS.t1434 851.341
R610 VSS.t3089 VSS.t2540 851.341
R611 VSS.t1787 VSS.t524 851.341
R612 VSS.t1776 VSS.t697 851.341
R613 VSS.t222 VSS.t2846 851.341
R614 VSS.t540 VSS.t2641 851.341
R615 VSS.n3988 VSS.n3987 850.336
R616 VSS.n3866 VSS.n3864 850.336
R617 VSS.n4891 VSS.t1448 850.068
R618 VSS.t3102 VSS.t2716 842.913
R619 VSS.t459 VSS.t78 842.913
R620 VSS.t3103 VSS.t2718 842.913
R621 VSS.t749 VSS.t1278 842.913
R622 VSS.t3440 VSS.t2449 842.913
R623 VSS.t3661 VSS.t1320 842.913
R624 VSS.t1489 VSS.t2123 842.913
R625 VSS.t4 VSS.t651 842.913
R626 VSS.t2512 VSS.t3540 842.913
R627 VSS.t1834 VSS.t336 842.913
R628 VSS.t3403 VSS.t910 842.913
R629 VSS.t3409 VSS.t506 842.913
R630 VSS.t2902 VSS.t2788 842.913
R631 VSS.t3351 VSS.t1129 842.913
R632 VSS.t3080 VSS.t3599 842.913
R633 VSS.t1164 VSS.t3085 842.913
R634 VSS.t3077 VSS.t915 842.913
R635 VSS.t668 VSS.t2954 834.484
R636 VSS.t926 VSS.t2295 834.484
R637 VSS.t1315 VSS.t1083 834.484
R638 VSS.t2077 VSS.t1392 834.484
R639 VSS.t399 VSS.t1671 834.484
R640 VSS.t988 VSS.t2165 834.484
R641 VSS.t2239 VSS.t156 834.484
R642 VSS.t1859 VSS.t2044 834.484
R643 VSS.t810 VSS.t808 834.484
R644 VSS.t2037 VSS.t381 834.484
R645 VSS.t234 VSS.t1505 834.484
R646 VSS.t2471 VSS.t1999 834.484
R647 VSS.t1379 VSS.t3291 834.484
R648 VSS.n4277 VSS.n4207 834.412
R649 VSS.n1754 VSS.n1750 833.155
R650 VSS.n1758 VSS.n1749 833.155
R651 VSS.n4032 VSS.n3961 833.155
R652 VSS.n3968 VSS.n3959 833.155
R653 VSS.t3430 VSS.n5375 827.551
R654 VSS.t3055 VSS.t2172 826.054
R655 VSS.t941 VSS.t2313 826.054
R656 VSS.t2295 VSS.t647 826.054
R657 VSS.t3414 VSS.t3616 826.054
R658 VSS.t781 VSS.t694 826.054
R659 VSS.t3163 VSS.t1953 826.054
R660 VSS.n4914 VSS.t2010 821.722
R661 VSS.t1986 VSS.n157 821.722
R662 VSS.t2117 VSS.t3592 817.625
R663 VSS.t395 VSS.t1165 817.625
R664 VSS.t2449 VSS.t204 817.625
R665 VSS.t3380 VSS.t509 817.625
R666 VSS.t80 VSS.t3590 817.625
R667 VSS.t3542 VSS.t1160 817.625
R668 VSS.t1798 VSS.t2827 817.625
R669 VSS.t2451 VSS.t3283 817.625
R670 VSS.t955 VSS.t3606 817.625
R671 VSS.t1592 VSS.t3469 817.625
R672 VSS.t3608 VSS.t856 817.625
R673 VSS.t1370 VSS.t2456 817.625
R674 VSS.t757 VSS.t2819 817.625
R675 VSS.n4914 VSS.t494 815.894
R676 VSS.n265 VSS.t2610 815.894
R677 VSS.t2747 VSS.n221 815.894
R678 VSS.t1380 VSS.n138 815.894
R679 VSS.t1503 VSS.n117 815.894
R680 VSS.n5375 VSS.t1336 815.894
R681 VSS.t2224 VSS.t1525 809.196
R682 VSS.t2088 VSS.t2090 809.196
R683 VSS.t1711 VSS.t350 809.196
R684 VSS.t1900 VSS.t348 809.196
R685 VSS.t74 VSS.t1157 809.196
R686 VSS.t2979 VSS.t1937 809.196
R687 VSS.t778 VSS.t296 809.196
R688 VSS.t341 VSS.t778 809.196
R689 VSS.t2081 VSS.t2429 809.196
R690 VSS.t249 VSS.t372 809.196
R691 VSS.t3694 VSS.t1825 809.196
R692 VSS.t1825 VSS.t2468 809.196
R693 VSS.t2618 VSS.t3557 809.196
R694 VSS.t3045 VSS.t3444 809.196
R695 VSS.t925 VSS.t924 809.196
R696 VSS.t804 VSS.t1490 809.196
R697 VSS.t3549 VSS.t3066 809.196
R698 VSS.t1461 VSS.t2355 809.196
R699 VSS.t1460 VSS.t1084 809.196
R700 VSS.t2734 VSS.t2938 809.196
R701 VSS.t2078 VSS.t2186 809.196
R702 VSS.t1348 VSS.t246 809.196
R703 VSS.t2051 VSS.t2459 809.196
R704 VSS.t2074 VSS.t2440 809.196
R705 VSS.t2885 VSS.t1099 809.196
R706 VSS.t3686 VSS.t1191 809.196
R707 VSS.t2888 VSS.t2823 809.196
R708 VSS.t2007 VSS.t2478 809.196
R709 VSS.t360 VSS.t1391 809.196
R710 VSS.t353 VSS.t1390 809.196
R711 VSS.t1748 VSS.t1823 809.196
R712 VSS.t999 VSS.t1150 809.196
R713 VSS.t2210 VSS.t2890 809.196
R714 VSS.t615 VSS.t993 809.196
R715 VSS.t2456 VSS.t2461 809.196
R716 VSS.t2038 VSS.t529 809.196
R717 VSS.t3555 VSS.t1491 809.196
R718 VSS.t906 VSS.t722 809.196
R719 VSS.t1663 VSS.t947 809.196
R720 VSS.t945 VSS.t658 809.196
R721 VSS.t2585 VSS.t379 809.196
R722 VSS.t1357 VSS.t1281 809.196
R723 VSS.t2540 VSS.t869 809.196
R724 VSS.t1572 VSS.t642 809.196
R725 VSS.t1267 VSS.t1955 809.196
R726 VSS.t1220 VSS.t3556 809.196
R727 VSS.t2780 VSS.t1216 809.196
R728 VSS.t1378 VSS.t1374 809.196
R729 VSS.n4839 VSS.t1446 802.178
R730 VSS.t292 VSS.t1665 800.766
R731 VSS.t2028 VSS.t1796 800.766
R732 VSS.t173 VSS.t1027 800.766
R733 VSS.t692 VSS.t2225 800.766
R734 VSS.n1626 VSS.t1710 800.766
R735 VSS.t247 VSS.t500 800.766
R736 VSS.t1772 VSS.t966 800.766
R737 VSS.t972 VSS.t82 800.766
R738 VSS.t1784 VSS.t2178 800.766
R739 VSS.t1235 VSS.t1231 800.766
R740 VSS.t1880 VSS.t1793 800.766
R741 VSS.t2552 VSS.t2315 800.766
R742 VSS.t766 VSS.t1782 800.766
R743 VSS.t2604 VSS.t2533 800.766
R744 VSS.t2349 VSS.t3542 800.766
R745 VSS.t2069 VSS.t1460 800.766
R746 VSS.t2341 VSS.t2445 800.766
R747 VSS.t2186 VSS.t1283 800.766
R748 VSS.t2782 VSS.t852 800.766
R749 VSS.t1732 VSS.t114 800.766
R750 VSS.t974 VSS.t216 800.766
R751 VSS.t2522 VSS.t1441 800.766
R752 VSS.t2408 VSS.t118 800.766
R753 VSS.t2490 VSS.t2888 800.766
R754 VSS.t1950 VSS.t1089 800.766
R755 VSS.t1117 VSS.t2486 800.766
R756 VSS.t1542 VSS.t274 800.766
R757 VSS.t762 VSS.t1725 800.766
R758 VSS.t1471 VSS.t2576 800.766
R759 VSS.t1065 VSS.t1748 800.766
R760 VSS.t1212 VSS.t2212 800.766
R761 VSS.t2503 VSS.t615 800.766
R762 VSS.t1005 VSS.t458 800.766
R763 VSS.t2385 VSS.t905 800.766
R764 VSS.t1137 VSS.t1632 800.766
R765 VSS.t257 VSS.t1177 800.766
R766 VSS.t1952 VSS.t583 800.766
R767 VSS.t1374 VSS.t2097 800.766
R768 VSS.t1738 VSS.t3273 800.766
R769 VSS.t2614 VSS.t387 800.766
R770 VSS.t1791 VSS.t937 800.766
R771 VSS.n4892 VSS.t2842 792.418
R772 VSS.t2840 VSS.n4111 792.418
R773 VSS.t1527 VSS.t3172 792.337
R774 VSS.t3078 VSS.t3539 792.337
R775 VSS.t3398 VSS.t1681 792.337
R776 VSS.t2169 VSS.t2513 792.337
R777 VSS.t1717 VSS.t445 792.337
R778 VSS.t3063 VSS.t3083 792.337
R779 VSS.t998 VSS.t2126 792.337
R780 VSS.t3094 VSS.t1368 783.909
R781 VSS.t2562 VSS.t3490 783.909
R782 VSS.t2544 VSS.t3004 783.909
R783 VSS.t953 VSS.t2730 781.025
R784 VSS.t2093 VSS.t1311 775.48
R785 VSS.t1278 VSS.t919 775.48
R786 VSS.t2005 VSS.n1327 775.48
R787 VSS.t1573 VSS.t649 775.48
R788 VSS.t2427 VSS.t1871 775.48
R789 VSS.t640 VSS.t2625 775.48
R790 VSS.t1214 VSS.t1826 775.48
R791 VSS.t1832 VSS.t399 775.48
R792 VSS.t3505 VSS.t3584 775.48
R793 VSS.t3604 VSS.t1095 775.48
R794 VSS.t3618 VSS.t1093 775.48
R795 VSS.t3469 VSS.t3622 775.48
R796 VSS.t1823 VSS.t1318 775.48
R797 VSS.t3434 VSS.t1240 775.48
R798 VSS.t1513 VSS.t3301 769.271
R799 VSS.t2753 VSS.t2343 767.051
R800 VSS.t1841 VSS.t3440 767.051
R801 VSS.t1610 VSS.t3272 767.051
R802 VSS.t965 VSS.t3329 767.051
R803 VSS.t990 VSS.t3319 767.051
R804 VSS.t1946 VSS.t3351 767.051
R805 VSS.t2826 VSS.t1091 767.051
R806 VSS.t1624 VSS.t1152 767.051
R807 VSS.t2709 VSS.t2702 767.051
R808 VSS.t2548 VSS.t1742 767.051
R809 VSS.t3311 VSS.t1021 767.051
R810 VSS.t1251 VSS.t3321 767.051
R811 VSS.t2508 VSS.t1444 760.519
R812 VSS.t2290 VSS.t2162 760.519
R813 VSS.t3289 VSS.t1524 758.621
R814 VSS.t2794 VSS.t2381 758.621
R815 VSS.t1416 VSS.t2332 758.621
R816 VSS.t1662 VSS.t1894 758.621
R817 VSS.t1493 VSS.n467 758.621
R818 VSS.t2218 VSS.t1770 758.621
R819 VSS.t2742 VSS.t3367 754.093
R820 VSS.t1147 VSS.t668 750.192
R821 VSS.t407 VSS.t2383 750.192
R822 VSS.t64 VSS.t3247 750.192
R823 VSS.t1968 VSS.t1476 750.192
R824 VSS.t2542 VSS.t2568 750.192
R825 VSS.t3544 VSS.t3103 741.763
R826 VSS.t2869 VSS.t2387 741.763
R827 VSS.t2806 VSS.t941 741.763
R828 VSS.t1103 VSS.t2512 741.763
R829 VSS.t1648 VSS.t2187 741.763
R830 VSS.t1580 VSS.t2019 741.763
R831 VSS.t3490 VSS.t2194 741.763
R832 VSS.t169 VSS.t1596 733.333
R833 VSS.t846 VSS.t327 733.333
R834 VSS.t3689 VSS.t3052 728.477
R835 VSS.t1660 VSS.t1273 728.477
R836 VSS.t1645 VSS.t2781 728.477
R837 VSS.t3034 VSS.t1047 728.477
R838 VSS.t3098 VSS.t3657 724.904
R839 VSS.t3630 VSS.t3626 724.904
R840 VSS.t313 VSS.t310 724.904
R841 VSS.t317 VSS.t294 724.904
R842 VSS.t294 VSS.t298 724.904
R843 VSS.t298 VSS.t306 724.904
R844 VSS.t315 VSS.t308 724.904
R845 VSS.t167 VSS.t323 724.904
R846 VSS.t304 VSS.t167 724.904
R847 VSS.t300 VSS.t304 724.904
R848 VSS.t296 VSS.t300 724.904
R849 VSS.t2036 VSS.t1360 724.904
R850 VSS.t1811 VSS.t1108 724.904
R851 VSS.t1108 VSS.t2903 724.904
R852 VSS.t2271 VSS.t2600 724.904
R853 VSS.t910 VSS.t1290 724.904
R854 VSS.t2831 VSS.t2772 724.904
R855 VSS.t468 VSS.t470 724.904
R856 VSS.t470 VSS.t2774 724.904
R857 VSS.t2827 VSS.t2829 724.904
R858 VSS.t1878 VSS.t3046 724.904
R859 VSS.t645 VSS.t3050 724.904
R860 VSS.t1671 VSS.t1685 724.904
R861 VSS.t441 VSS.t431 724.904
R862 VSS.t431 VSS.t425 724.904
R863 VSS.t421 VSS.t433 724.904
R864 VSS.t433 VSS.t439 724.904
R865 VSS.t415 VSS.t435 724.904
R866 VSS.t413 VSS.t427 724.904
R867 VSS.t3018 VSS.t3010 724.904
R868 VSS.t3010 VSS.t3016 724.904
R869 VSS.t2894 VSS.t3604 724.904
R870 VSS.t76 VSS.t3618 724.904
R871 VSS.t1434 VSS.t76 724.904
R872 VSS.t859 VSS.t1643 724.904
R873 VSS.t573 VSS.t3062 724.904
R874 VSS.t842 VSS.t824 724.904
R875 VSS.t838 VSS.t842 724.904
R876 VSS.t828 VSS.t830 724.904
R877 VSS.t834 VSS.t850 724.904
R878 VSS.t850 VSS.t844 724.904
R879 VSS.t844 VSS.t840 724.904
R880 VSS.t832 VSS.t3012 724.904
R881 VSS.t3002 VSS.t3000 724.904
R882 VSS.t3000 VSS.t3006 724.904
R883 VSS.t2670 VSS.t150 724.904
R884 VSS.t492 VSS.t486 724.904
R885 VSS.t2995 VSS.t2993 724.904
R886 VSS.t2993 VSS.t2998 724.904
R887 VSS.t16 VSS.t10 724.904
R888 VSS.t18 VSS.t16 724.904
R889 VSS.t32 VSS.t18 724.904
R890 VSS.t24 VSS.t12 724.904
R891 VSS.t36 VSS.t30 724.904
R892 VSS.t26 VSS.t22 724.904
R893 VSS.t3582 VSS.t507 724.904
R894 VSS.t883 VSS.t877 724.904
R895 VSS.t871 VSS.t883 724.904
R896 VSS.t881 VSS.t871 724.904
R897 VSS.t889 VSS.t881 724.904
R898 VSS.t887 VSS.t897 724.904
R899 VSS.t873 VSS.t885 724.904
R900 VSS.t875 VSS.t891 724.904
R901 VSS.t879 VSS.t875 724.904
R902 VSS.t3014 VSS.t899 724.904
R903 VSS.t3020 VSS.t3014 724.904
R904 VSS.t1744 VSS.t3020 724.904
R905 VSS.t2964 VSS.t1744 724.904
R906 VSS.t2419 VSS.t2503 724.904
R907 VSS.t1183 VSS.t1185 724.904
R908 VSS.t1185 VSS.t1179 724.904
R909 VSS.t1179 VSS.t1181 724.904
R910 VSS.t1342 VSS.t1346 724.904
R911 VSS.t1346 VSS.t1340 724.904
R912 VSS.t1340 VSS.t1344 724.904
R913 VSS.t195 VSS.t193 724.904
R914 VSS.t189 VSS.t195 724.904
R915 VSS.t191 VSS.t189 724.904
R916 VSS.t165 VSS.t159 724.904
R917 VSS.t161 VSS.t165 724.904
R918 VSS.t163 VSS.t161 724.904
R919 VSS.t308 VSS.t319 716.476
R920 VSS.t1588 VSS.t2036 716.476
R921 VSS.t385 VSS.t2766 716.476
R922 VSS.t401 VSS.t2074 716.476
R923 VSS.t429 VSS.t415 716.476
R924 VSS.t3317 VSS.t261 716.476
R925 VSS.t2220 VSS.t1267 716.476
R926 VSS.t290 VSS.t292 708.047
R927 VSS.t1027 VSS.t1025 708.047
R928 VSS.t1888 VSS.t1890 708.047
R929 VSS.t687 VSS.t2865 708.047
R930 VSS.t2488 VSS.t1327 708.047
R931 VSS.t3592 VSS.t66 708.047
R932 VSS.t2954 VSS.t2086 708.047
R933 VSS.t665 VSS.t3596 708.047
R934 VSS.t2594 VSS.t665 708.047
R935 VSS.t2592 VSS.t1711 708.047
R936 VSS.t1165 VSS.t3537 708.047
R937 VSS.t3537 VSS.t393 708.047
R938 VSS.t2233 VSS.t2235 708.047
R939 VSS.t1243 VSS.t74 708.047
R940 VSS.t78 VSS.t1974 708.047
R941 VSS.t1937 VSS.t1976 708.047
R942 VSS.t3533 VSS.t3535 708.047
R943 VSS.t2578 VSS.t1208 708.047
R944 VSS.t2330 VSS.t2081 708.047
R945 VSS.t751 VSS.t749 708.047
R946 VSS.t245 VSS.t2671 708.047
R947 VSS.t2671 VSS.t2002 708.047
R948 VSS.t2443 VSS.t2441 708.047
R949 VSS.t374 VSS.t148 708.047
R950 VSS.t1681 VSS.t3419 708.047
R951 VSS.t3620 VSS.t3612 708.047
R952 VSS.t500 VSS.t498 708.047
R953 VSS.t199 VSS.t3053 708.047
R954 VSS.t200 VSS.t208 708.047
R955 VSS.t3644 VSS.t2518 708.047
R956 VSS.t1568 VSS.t1048 708.047
R957 VSS.t966 VSS.t968 708.047
R958 VSS.t82 VSS.t84 708.047
R959 VSS.t2178 VSS.t2180 708.047
R960 VSS.t1233 VSS.t1235 708.047
R961 VSS.t1882 VSS.t1880 708.047
R962 VSS.t2550 VSS.t2552 708.047
R963 VSS.t764 VSS.t766 708.047
R964 VSS.t2533 VSS.t2531 708.047
R965 VSS.t562 VSS.t560 708.047
R966 VSS.t2899 VSS.t1482 708.047
R967 VSS.t128 VSS.t130 708.047
R968 VSS.t130 VSS.t124 708.047
R969 VSS.t806 VSS.t2771 708.047
R970 VSS.t2353 VSS.t2349 708.047
R971 VSS.t2357 VSS.t2351 708.047
R972 VSS.t2355 VSS.t2901 708.047
R973 VSS.t2938 VSS.t1458 708.047
R974 VSS.t2944 VSS.t2447 708.047
R975 VSS.t1254 VSS.t1252 708.047
R976 VSS.t712 VSS.t714 708.047
R977 VSS.t2188 VSS.t1467 708.047
R978 VSS.t675 VSS.t681 708.047
R979 VSS.t2184 VSS.t2906 708.047
R980 VSS.t1292 VSS.t1350 708.047
R981 VSS.t1290 VSS.t1295 708.047
R982 VSS.t1022 VSS.t3407 708.047
R983 VSS.t2475 VSS.t1798 708.047
R984 VSS.t513 VSS.t792 708.047
R985 VSS.t3484 VSS.t3462 708.047
R986 VSS.t3462 VSS.t3463 708.047
R987 VSS.t3410 VSS.t3405 708.047
R988 VSS.t3405 VSS.t3401 708.047
R989 VSS.t3401 VSS.t3414 708.047
R990 VSS.t790 VSS.t3460 708.047
R991 VSS.t2249 VSS.t786 708.047
R992 VSS.t786 VSS.t516 708.047
R993 VSS.t502 VSS.t2763 708.047
R994 VSS.t2763 VSS.t405 708.047
R995 VSS.t927 VSS.t929 708.047
R996 VSS.t634 VSS.t632 708.047
R997 VSS.t2437 VSS.t3679 708.047
R998 VSS.t2566 VSS.t2564 708.047
R999 VSS.t114 VSS.t112 708.047
R1000 VSS.t216 VSS.t218 708.047
R1001 VSS.t1073 VSS.t1075 708.047
R1002 VSS.t2936 VSS.t2942 708.047
R1003 VSS.t2985 VSS.t2707 708.047
R1004 VSS.t2940 VSS.t1439 708.047
R1005 VSS.t2867 VSS.t2861 708.047
R1006 VSS.t1590 VSS.t3038 708.047
R1007 VSS.t2406 VSS.t2928 708.047
R1008 VSS.t1191 VSS.t2602 708.047
R1009 VSS.t1245 VSS.t3686 708.047
R1010 VSS.t1280 VSS.t818 708.047
R1011 VSS.t3099 VSS.t3068 708.047
R1012 VSS.t3570 VSS.t2095 708.047
R1013 VSS.t3527 VSS.t2828 708.047
R1014 VSS.t334 VSS.t2490 708.047
R1015 VSS.t2823 VSS.t3632 708.047
R1016 VSS.t949 VSS.t1051 708.047
R1017 VSS.t1051 VSS.t1641 708.047
R1018 VSS.t330 VSS.t325 708.047
R1019 VSS.t1758 VSS.t781 708.047
R1020 VSS.t1713 VSS.t1758 708.047
R1021 VSS.t2658 VSS.t911 708.047
R1022 VSS.t1057 VSS.t2658 708.047
R1023 VSS.t2667 VSS.t2 708.047
R1024 VSS.t774 VSS.t2667 708.047
R1025 VSS.t327 VSS.t916 708.047
R1026 VSS.t830 VSS.t1586 708.047
R1027 VSS.t2656 VSS.t908 708.047
R1028 VSS.t2046 VSS.t3485 708.047
R1029 VSS.t1115 VSS.t1117 708.047
R1030 VSS.t2662 VSS.t2665 708.047
R1031 VSS.t2660 VSS.t1592 708.047
R1032 VSS.t142 VSS.t144 708.047
R1033 VSS.t253 VSS.t3396 708.047
R1034 VSS.t3396 VSS.t3412 708.047
R1035 VSS.t3457 VSS.t1104 708.047
R1036 VSS.t856 VSS.t26 708.047
R1037 VSS.t507 VSS.t1045 708.047
R1038 VSS.t358 VSS.t364 708.047
R1039 VSS.t1119 VSS.t3677 708.047
R1040 VSS.t1960 VSS.t1958 708.047
R1041 VSS.t274 VSS.t276 708.047
R1042 VSS.t760 VSS.t762 708.047
R1043 VSS.t1133 VSS.t1131 708.047
R1044 VSS.t1063 VSS.t1065 708.047
R1045 VSS.t588 VSS.t2962 708.047
R1046 VSS.t1200 VSS.t1198 708.047
R1047 VSS.t2717 VSS.t2711 708.047
R1048 VSS.t2968 VSS.t2717 708.047
R1049 VSS.t2977 VSS.t2987 708.047
R1050 VSS.t993 VSS.t991 708.047
R1051 VSS.t2584 VSS.t2863 708.047
R1052 VSS.t656 VSS.t654 708.047
R1053 VSS.t1639 VSS.t3104 708.047
R1054 VSS.t2960 VSS.t456 708.047
R1055 VSS.t768 VSS.t770 708.047
R1056 VSS.t3036 VSS.t3032 708.047
R1057 VSS.t3031 VSS.t2378 708.047
R1058 VSS.t726 VSS.t724 708.047
R1059 VSS.t722 VSS.t784 708.047
R1060 VSS.t2910 VSS.t903 708.047
R1061 VSS.t2819 VSS.t759 708.047
R1062 VSS.t1265 VSS.t1271 708.047
R1063 VSS.t1271 VSS.t1263 708.047
R1064 VSS.t1953 VSS.t3673 708.047
R1065 VSS.t2206 VSS.t2208 708.047
R1066 VSS.t2204 VSS.t2200 708.047
R1067 VSS.t387 VSS.t389 708.047
R1068 VSS.t937 VSS.t935 708.047
R1069 VSS.t177 VSS.t181 708.047
R1070 VSS.t183 VSS.t177 708.047
R1071 VSS.t179 VSS.t183 708.047
R1072 VSS.t518 VSS.t520 708.047
R1073 VSS.t522 VSS.t518 708.047
R1074 VSS.t524 VSS.t522 708.047
R1075 VSS.t1540 VSS.t1787 708.047
R1076 VSS.t699 VSS.t703 708.047
R1077 VSS.t701 VSS.t699 708.047
R1078 VSS.t697 VSS.t701 708.047
R1079 VSS.t1551 VSS.t1776 708.047
R1080 VSS.t224 VSS.t226 708.047
R1081 VSS.t226 VSS.t220 708.047
R1082 VSS.t220 VSS.t222 708.047
R1083 VSS.t2846 VSS.t2883 708.047
R1084 VSS.t534 VSS.t536 708.047
R1085 VSS.t536 VSS.t538 708.047
R1086 VSS.t538 VSS.t540 708.047
R1087 VSS.t2641 VSS.t1734 708.047
R1088 VSS.n3718 VSS.n3717 708.047
R1089 VSS.t2026 VSS.t483 708.047
R1090 VSS.t1399 VSS.t1041 708.047
R1091 VSS.t2231 VSS.t3558 699.617
R1092 VSS.t3539 VSS.t2588 699.617
R1093 VSS.t3091 VSS.t2171 699.617
R1094 VSS.t451 VSS.t530 699.617
R1095 VSS.t805 VSS.t1828 699.617
R1096 VSS.t51 VSS.t653 699.617
R1097 VSS.t409 VSS.t447 699.617
R1098 VSS.t1945 VSS.t571 699.617
R1099 VSS.t2022 VSS.t3614 699.617
R1100 VSS.t848 VSS.t1884 699.617
R1101 VSS.t820 VSS.t557 699.617
R1102 VSS.t22 VSS.t2243 699.617
R1103 VSS.t2946 VSS.t3600 699.617
R1104 VSS.t455 VSS.t1429 699.617
R1105 VSS.t1634 VSS.t528 699.617
R1106 VSS.t1135 VSS.t2216 699.617
R1107 VSS.t1375 VSS.t3275 699.617
R1108 VSS.t2089 VSS.t1329 691.188
R1109 VSS.t449 VSS.t2790 691.188
R1110 VSS.t2722 VSS.t3448 691.188
R1111 VSS.t545 VSS.t1550 691.188
R1112 VSS.t2776 VSS.t28 691.188
R1113 VSS.t1079 VSS.t2369 682.76
R1114 VSS.t2284 VSS.t1746 682.76
R1115 VSS.t1487 VSS.t1674 682.76
R1116 VSS.t3319 VSS.t1669 682.76
R1117 VSS.t1875 VSS.t2251 682.76
R1118 VSS.t852 VSS.t3646 682.76
R1119 VSS.t1250 VSS.t401 682.76
R1120 VSS.t802 VSS.t569 682.76
R1121 VSS.t464 VSS.t102 682.76
R1122 VSS.t672 VSS.t3424 682.76
R1123 VSS.t3487 VSS.t20 682.76
R1124 VSS.t1167 VSS.t3418 682.76
R1125 VSS.t3663 VSS.t2222 674.331
R1126 VSS.t3454 VSS.t1582 674.331
R1127 VSS.t351 VSS.t2787 674.331
R1128 VSS.t772 VSS.t783 674.331
R1129 VSS.t372 VSS.t1588 674.331
R1130 VSS.t213 VSS.t921 674.331
R1131 VSS.t2966 VSS.t2403 674.331
R1132 VSS.t3638 VSS.t3438 674.331
R1133 VSS.t2484 VSS.t3386 674.331
R1134 VSS.t982 VSS.t360 674.331
R1135 VSS.t3064 VSS.t268 668.768
R1136 VSS.t3359 VSS.t1049 665.9
R1137 VSS.t1158 VSS.n1625 665.9
R1138 VSS.t1157 VSS.t2872 665.9
R1139 VSS.t3087 VSS.t342 665.9
R1140 VSS.t2572 VSS.t575 665.9
R1141 VSS.t1101 VSS.t1164 665.9
R1142 VSS.n2634 VSS.t38 665.9
R1143 VSS.t1815 VSS.t1859 665.9
R1144 VSS.t3435 VSS.t1225 665.9
R1145 VSS.t3313 VSS.t147 665.9
R1146 VSS.t264 VSS.n3667 660.612
R1147 VSS.t2896 VSS.t1228 657.471
R1148 VSS.t621 VSS.t2233 657.471
R1149 VSS.t2368 VSS.t3546 657.471
R1150 VSS.t2171 VSS.t3055 657.471
R1151 VSS.t696 VSS.t315 657.471
R1152 VSS.t3372 VSS.t2675 657.471
R1153 VSS.t3307 VSS.t2514 657.471
R1154 VSS.t2712 VSS.t2166 657.471
R1155 VSS.t2240 VSS.t1388 657.471
R1156 VSS.t2596 VSS.t1537 657.471
R1157 VSS.t381 VSS.t3058 657.471
R1158 VSS.n467 VSS.t1533 657.471
R1159 VSS.t1286 VSS.t1756 657.471
R1160 VSS.t3667 VSS.t210 657.471
R1161 VSS.t2226 VSS.t2176 649.043
R1162 VSS.t2253 VSS.t3043 649.043
R1163 VSS.t2465 VSS.t354 649.043
R1164 VSS.t1830 VSS.t1194 646.366
R1165 VSS.t3501 VSS.t302 640.614
R1166 VSS.t3525 VSS.t2825 640.614
R1167 VSS.t2282 VSS.t543 640.614
R1168 VSS.t1668 VSS.t1480 640.614
R1169 VSS.t2377 VSS.t577 640.614
R1170 VSS.n2942 VSS.t1258 640.614
R1171 VSS.t1680 VSS.t913 640.614
R1172 VSS.t1352 VSS.t2049 640.614
R1173 VSS.t3650 VSS.t1678 640.614
R1174 VSS.t1384 VSS.t988 640.614
R1175 VSS.t815 VSS.t2886 640.614
R1176 VSS.t623 VSS.t429 640.614
R1177 VSS.t625 VSS.t345 640.614
R1178 VSS.t1432 VSS.t1247 640.614
R1179 VSS.t809 VSS.t1662 640.614
R1180 VSS.t1162 VSS.t1616 640.614
R1181 VSS.t1970 VSS.t2524 640.614
R1182 VSS.t1915 VSS.t1530 636.266
R1183 VSS.t2767 VSS.t383 636.266
R1184 VSS.t370 VSS.t2930 636.266
R1185 VSS.t1511 VSS.t1990 635.232
R1186 VSS.t1766 VSS.t1380 635.232
R1187 VSS.t2364 VSS.t484 635.232
R1188 VSS.t1694 VSS.t1503 635.232
R1189 VSS.t1701 VSS.t1336 635.232
R1190 VSS.t3488 VSS.t1913 632.9
R1191 VSS.t1529 VSS.t2767 632.9
R1192 VSS.t1636 VSS.t776 632.184
R1193 VSS.n1567 VSS.t319 632.184
R1194 VSS.t2429 VSS.t2491 632.184
R1195 VSS.t1260 VSS.t712 632.184
R1196 VSS.t427 VSS.t2580 632.184
R1197 VSS.n2474 VSS.t822 632.184
R1198 VSS.t2958 VSS.t2452 632.184
R1199 VSS.t2297 VSS.t1564 629.404
R1200 VSS.t1560 VSS.t1031 629.404
R1201 VSS.t2293 VSS.t1566 629.404
R1202 VSS.t2115 VSS.t2088 623.755
R1203 VSS.t2625 VSS.t2606 623.755
R1204 VSS.t2440 VSS.t1123 623.755
R1205 VSS.t1325 VSS.t1438 623.755
R1206 VSS.t2579 VSS.t423 623.755
R1207 VSS.t901 VSS.t1282 623.755
R1208 VSS.t1021 VSS.t1754 623.755
R1209 VSS.t3281 VSS.t1475 623.755
R1210 VSS.t610 VSS.t2975 617.749
R1211 VSS.t1849 VSS.t604 617.749
R1212 VSS.t287 VSS.t1570 615.327
R1213 VSS.t3008 VSS.t2582 615.327
R1214 VSS.t1727 VSS.t2983 615.327
R1215 VSS.t1535 VSS.t3099 615.327
R1216 VSS.t3012 VSS.t52 615.327
R1217 VSS.t2973 VSS.t998 615.327
R1218 VSS.t2546 VSS.t1162 615.327
R1219 VSS.t2570 VSS.t2541 615.327
R1220 VSS.t1042 VSS.t3359 606.898
R1221 VSS.t2560 VSS.t2255 606.898
R1222 VSS.t2718 VSS.t1515 606.898
R1223 VSS.t1368 VSS.t1024 606.898
R1224 VSS.t3074 VSS.t3091 606.898
R1225 VSS.t1077 VSS.t40 606.898
R1226 VSS.t783 VSS.t3082 606.898
R1227 VSS.t1555 VSS.t907 606.898
R1228 VSS.t674 VSS.t2003 606.898
R1229 VSS.t212 VSS.t2515 606.898
R1230 VSS.t3231 VSS.t3694 606.898
R1231 VSS.t3361 VSS.t2380 606.898
R1232 VSS.t3349 VSS.t2397 606.898
R1233 VSS.t1490 VSS.t1241 606.898
R1234 VSS.t1317 VSS.t1614 606.898
R1235 VSS.t3117 VSS.t3271 606.898
R1236 VSS.t2083 VSS.t1622 606.898
R1237 VSS.t2669 VSS.t1575 606.898
R1238 VSS.t683 VSS.t1834 606.898
R1239 VSS.t3343 VSS.t1394 606.898
R1240 VSS.n2891 VSS.t1128 606.898
R1241 VSS.t1127 VSS.t2169 606.898
R1242 VSS.t2361 VSS.t3368 606.898
R1243 VSS.t3299 VSS.t1947 606.898
R1244 VSS.t2426 VSS.t3299 606.898
R1245 VSS.t136 VSS.t1442 606.898
R1246 VSS.t2021 VSS.t2536 606.898
R1247 VSS.t1995 VSS.t1877 606.898
R1248 VSS.t3464 VSS.t24 606.898
R1249 VSS.t515 VSS.t3391 606.898
R1250 VSS.t1001 VSS.t2045 606.898
R1251 VSS.t3498 VSS.t1895 606.898
R1252 VSS.t236 VSS.t2755 606.898
R1253 VSS.t3339 VSS.t2001 606.898
R1254 VSS.n5377 VSS.t1251 606.898
R1255 VSS.t3337 VSS.t2458 606.898
R1256 VSS.t3022 VSS.t1780 606.898
R1257 VSS.t2679 VSS.t1795 606.898
R1258 VSS.t2640 VSS.t3521 606.898
R1259 VSS.t1664 VSS.t1719 606.898
R1260 VSS.n4798 VSS.n4797 599.125
R1261 VSS.n4762 VSS.n4733 599.125
R1262 VSS.t3384 VSS.t3045 598.467
R1263 VSS.t813 VSS.t3363 598.467
R1264 VSS.t2701 VSS.t3602 598.467
R1265 VSS.t3465 VSS.t1224 598.467
R1266 VSS.t2514 VSS.t2480 598.467
R1267 VSS.t816 VSS.t437 598.467
R1268 VSS.t785 VSS.t1721 598.467
R1269 VSS.t1106 VSS.t490 598.467
R1270 VSS.t3041 VSS.t14 598.467
R1271 VSS.n2635 VSS.t3323 598.467
R1272 VSS.t2454 VSS.t1370 598.467
R1273 VSS.t1756 VSS.t3311 598.467
R1274 VSS.n3812 VSS.t1705 590.73
R1275 VSS.t1333 VSS.t2366 590.038
R1276 VSS.t2347 VSS.t3495 590.038
R1277 VSS.t2494 VSS.t3426 590.038
R1278 VSS.n1445 VSS.t2494 590.038
R1279 VSS.t1468 VSS.t3374 590.038
R1280 VSS.t2167 VSS.t2164 590.038
R1281 VSS.t1944 VSS.t2182 590.038
R1282 VSS.t590 VSS.t999 590.038
R1283 VSS.t2971 VSS.t3452 590.038
R1284 VSS.t458 VSS.n466 590.038
R1285 VSS.t1533 VSS.t2263 590.038
R1286 VSS.t659 VSS.t1506 590.038
R1287 VSS.t1656 VSS.t3315 590.038
R1288 VSS.t2472 VSS.t175 590.038
R1289 VSS.t933 VSS.t317 581.61
R1290 VSS.n1328 VSS.t3035 581.61
R1291 VSS.t1813 VSS.t812 581.61
R1292 VSS.t2861 VSS.t2522 581.61
R1293 VSS.t472 VSS.t488 581.61
R1294 VSS.t474 VSS.t8 581.61
R1295 VSS.t3323 VSS.t982 581.61
R1296 VSS.t1997 VSS.t2014 581.61
R1297 VSS.t1990 VSS.t1513 576.955
R1298 VSS.t344 VSS.t3628 573.181
R1299 VSS.t1870 VSS.t214 573.181
R1300 VSS.t2397 VSS.t1668 573.181
R1301 VSS.t3648 VSS.t3588 573.181
R1302 VSS.t77 VSS.t1462 573.181
R1303 VSS.t1669 VSS.t677 573.181
R1304 VSS.t1128 VSS.t2482 573.181
R1305 VSS.t1061 VSS.t2439 573.181
R1306 VSS.t1029 VSS.t362 573.181
R1307 VSS.t984 VSS.t3309 573.181
R1308 VSS.t1210 VSS.t2043 573.181
R1309 VSS.t1331 VSS.t1386 565.298
R1310 VSS.t1382 VSS.t1909 565.298
R1311 VSS.t1618 VSS.t1862 565.298
R1312 VSS.t280 VSS.t2269 565.298
R1313 VSS.t1011 VSS.t1938 565.298
R1314 VSS.t551 VSS.t1986 565.298
R1315 VSS.t2751 VSS.t1145 565.298
R1316 VSS.t2142 VSS.t1409 565.298
R1317 VSS.t1857 VSS.t2103 565.298
R1318 VSS.t2059 VSS.t3432 565.298
R1319 VSS.t239 VSS.t2391 565.298
R1320 VSS.t1087 VSS.t1532 564.751
R1321 VSS.t2620 VSS.t328 564.751
R1322 VSS.t2128 VSS.t1946 564.751
R1323 VSS.t822 VSS.t558 564.751
R1324 VSS.t254 VSS.t2119 564.751
R1325 VSS.t3104 VSS.t1005 564.751
R1326 VSS.t2265 VSS.t3555 564.751
R1327 VSS.t146 VSS.t2130 564.751
R1328 VSS.t2586 VSS.t1298 564.751
R1329 VSS.t710 VSS.t1511 559.471
R1330 VSS.t1991 VSS.t1512 559.471
R1331 VSS.t1892 VSS.t3689 559.471
R1332 VSS.t3052 VSS.t1766 559.471
R1333 VSS.t2261 VSS.t1660 559.471
R1334 VSS.t1273 VSS.t2364 559.471
R1335 VSS.t1303 VSS.t1645 559.471
R1336 VSS.t2781 VSS.t1694 559.471
R1337 VSS.t2288 VSS.t3034 559.471
R1338 VSS.t1047 VSS.t1701 559.471
R1339 VSS.t2228 VSS.t2558 558.837
R1340 VSS.n3901 VSS.t3711 557.02
R1341 VSS.n3896 VSS.t3717 557.013
R1342 VSS.n3901 VSS.t3743 556.54
R1343 VSS.n3899 VSS.t3739 556.54
R1344 VSS.n3900 VSS.t3738 556.54
R1345 VSS.n3898 VSS.t3748 556.54
R1346 VSS.n3897 VSS.t3736 556.54
R1347 VSS.n3896 VSS.t3757 556.54
R1348 VSS.t347 VSS.t56 556.322
R1349 VSS.t508 VSS.t3642 556.322
R1350 VSS.t1048 VSS.t3380 556.322
R1351 VSS.t466 VSS.t3598 556.322
R1352 VSS.t824 VSS.t2561 556.322
R1353 VSS.t1122 VSS.t3675 556.322
R1354 VSS.t596 VSS.t1608 556.322
R1355 VSS.t403 VSS.t2219 556.322
R1356 VSS.t3633 VSS.t2319 553.643
R1357 VSS.t2012 VSS.t1080 553.643
R1358 VSS.t1628 VSS.t2150 553.643
R1359 VSS.t1740 VSS.t1192 553.643
R1360 VSS.t2410 VSS.t2412 553.643
R1361 VSS.t1196 VSS.t270 553.643
R1362 VSS.t1512 VSS.t986 553.643
R1363 VSS.t626 VSS.t2747 553.643
R1364 VSS.t978 VSS.t1847 553.643
R1365 VSS.t661 VSS.t3578 553.643
R1366 VSS.t3475 VSS.t3207 550.402
R1367 VSS.t3305 VSS.t2592 547.894
R1368 VSS.t2901 VSS.t1606 547.894
R1369 VSS.t3270 VSS.t3096 547.894
R1370 VSS.t2769 VSS.t1469 547.894
R1371 VSS.t689 VSS.t2970 547.894
R1372 VSS.t2497 VSS.t2720 547.894
R1373 VSS.t263 VSS.t2239 547.894
R1374 VSS.t2962 VSS.t3303 547.894
R1375 VSS.t3213 VSS.t879 547.894
R1376 VSS.t784 VSS.t2757 547.894
R1377 VSS.t288 VSS.t1071 539.465
R1378 VSS.t3590 VSS.t2398 539.465
R1379 VSS.t1258 VSS.t1630 539.465
R1380 VSS.t681 VSS.t1307 539.465
R1381 VSS.t2439 VSS.t3327 539.465
R1382 VSS.t970 VSS.t38 539.465
R1383 VSS.t261 VSS.t984 539.465
R1384 VSS.t895 VSS.t476 539.465
R1385 VSS.t2863 VSS.t2952 539.465
R1386 VSS.t2405 VSS.t586 539.465
R1387 VSS.t3335 VSS.t2220 539.465
R1388 VSS.t2202 VSS.t1661 539.465
R1389 VSS.t3714 VSS.n1849 538.312
R1390 VSS.n4205 VSS.n4204 538.28
R1391 VSS.t66 VSS.t2526 531.034
R1392 VSS.t43 VSS.t347 531.034
R1393 VSS.t152 VSS.t206 531.034
R1394 VSS.t1309 VSS.t332 531.034
R1395 VSS.t397 VSS.t3669 531.034
R1396 VSS.t1411 VSS.t116 531.034
R1397 VSS.t526 VSS.t1658 531.034
R1398 VSS.t705 VSS.t3297 530.332
R1399 VSS.n3891 VSS.t58 526.735
R1400 VSS.n3816 VSS.t2925 526.693
R1401 VSS.n3976 VSS.t3574 526.693
R1402 VSS.n3895 VSS.t61 526.552
R1403 VSS.t1276 VSS.t2371 522.606
R1404 VSS.t2989 VSS.t2462 522.606
R1405 VSS.t2908 VSS.t2574 522.606
R1406 VSS.t3382 VSS.t1690 522.606
R1407 VSS.t581 VSS.t2673 522.606
R1408 VSS.t794 VSS.t3075 522.606
R1409 VSS.t94 VSS.t1650 522.606
R1410 VSS.t2461 VSS.t526 522.606
R1411 VSS.t995 VSS.t185 522.606
R1412 VSS.t2489 VSS.t2091 514.177
R1413 VSS.t68 VSS.t1158 514.177
R1414 VSS.t509 VSS.t2728 514.177
R1415 VSS.t1684 VSS.t2761 514.177
R1416 VSS.t3586 VSS.t419 514.177
R1417 VSS.t3333 VSS.t2334 514.177
R1418 VSS.t2321 VSS.t866 514.177
R1419 VSS.t2981 VSS.t1484 514.177
R1420 VSS.t494 VSS.t3503 512.848
R1421 VSS.t2612 VSS.t864 512.848
R1422 VSS.t2610 VSS.t2538 512.848
R1423 VSS.t232 VSS.t1544 512.848
R1424 VSS.t1703 VSS.t2214 512.848
R1425 VSS.t1297 VSS.t2676 505.748
R1426 VSS.t1338 VSS.t731 505.748
R1427 VSS.t1470 VSS.t3641 505.748
R1428 VSS.t2076 VSS.t1125 505.748
R1429 VSS.t2166 VSS.t2361 505.748
R1430 VSS.t2529 VSS.t2426 505.748
R1431 VSS.t1067 VSS.t492 505.748
R1432 VSS.t1452 VSS.t1450 502.858
R1433 VSS.t1450 VSS.t1454 502.858
R1434 VSS.t1454 VSS.t1456 502.858
R1435 VSS.t1446 VSS.t1448 502.858
R1436 VSS.t1909 VSS.t1911 501.192
R1437 VSS.t1911 VSS.t1905 501.192
R1438 VSS.t1905 VSS.t1907 501.192
R1439 VSS.t1862 VSS.t1866 501.192
R1440 VSS.t1866 VSS.t1868 501.192
R1441 VSS.t1868 VSS.t1864 501.192
R1442 VSS.t282 VSS.t278 501.192
R1443 VSS.t278 VSS.t284 501.192
R1444 VSS.t284 VSS.t280 501.192
R1445 VSS.t1015 VSS.t1013 501.192
R1446 VSS.t1013 VSS.t1017 501.192
R1447 VSS.t1017 VSS.t1011 501.192
R1448 VSS.t553 VSS.t555 501.192
R1449 VSS.t555 VSS.t549 501.192
R1450 VSS.t549 VSS.t551 501.192
R1451 VSS.t1145 VSS.t1141 501.192
R1452 VSS.t1141 VSS.t1143 501.192
R1453 VSS.t1143 VSS.t1139 501.192
R1454 VSS.t2148 VSS.t2146 501.192
R1455 VSS.t2146 VSS.t2144 501.192
R1456 VSS.t2144 VSS.t2142 501.192
R1457 VSS.t1851 VSS.t1855 501.192
R1458 VSS.t1855 VSS.t1853 501.192
R1459 VSS.t1853 VSS.t1857 501.192
R1460 VSS.t2055 VSS.t2053 501.192
R1461 VSS.t2053 VSS.t2057 501.192
R1462 VSS.t2057 VSS.t2059 501.192
R1463 VSS.t241 VSS.t239 501.192
R1464 VSS.t243 VSS.t241 501.192
R1465 VSS.t237 VSS.t243 501.192
R1466 VSS.t3400 VSS.t1764 497.318
R1467 VSS.t3598 VSS.t2885 497.318
R1468 VSS.t0 VSS.t1578 497.318
R1469 VSS.t1059 VSS.t670 497.318
R1470 VSS.t2241 VSS.t32 497.318
R1471 VSS.t1204 VSS.t3279 491.382
R1472 VSS.t2319 VSS.t2317 489.536
R1473 VSS.t2010 VSS.t2012 489.536
R1474 VSS.t1386 VSS.t1335 489.536
R1475 VSS.t270 VSS.t272 489.536
R1476 VSS.t706 VSS.t708 489.536
R1477 VSS.t1509 VSS.t2950 489.536
R1478 VSS.t628 VSS.t626 489.536
R1479 VSS.t612 VSS.t608 489.536
R1480 VSS.t608 VSS.t606 489.536
R1481 VSS.t606 VSS.t610 489.536
R1482 VSS.t2975 VSS.t2628 489.536
R1483 VSS.t2628 VSS.t1849 489.536
R1484 VSS.t3681 VSS.t3684 489.536
R1485 VSS.t1564 VSS.t3683 489.536
R1486 VSS.t1638 VSS.t1560 489.536
R1487 VSS.t1566 VSS.t3030 489.536
R1488 VSS.t1982 VSS.t1984 489.536
R1489 VSS.t2190 VSS.t2192 489.536
R1490 VSS.t1407 VSS.t1405 489.536
R1491 VSS.t2101 VSS.t2099 489.536
R1492 VSS.t3428 VSS.t3430 489.536
R1493 VSS.t980 VSS.t978 489.536
R1494 VSS.t663 VSS.t661 489.536
R1495 VSS.t3550 VSS.t1069 489.342
R1496 VSS.t393 VSS.t2464 488.889
R1497 VSS.t1085 VSS.t3078 488.889
R1498 VSS.t632 VSS.t2395 488.889
R1499 VSS.t3325 VSS.t1126 488.889
R1500 VSS.t3353 VSS.t2417 488.889
R1501 VSS.t858 VSS.t1082 488.889
R1502 VSS.t333 VSS.t134 488.889
R1503 VSS.t840 VSS.t3287 488.889
R1504 VSS.t836 VSS.t3500 488.889
R1505 VSS.t854 VSS.t788 488.889
R1506 VSS.t1809 VSS.t1299 488.889
R1507 VSS.t1998 VSS.t1921 488.889
R1508 VSS.t3552 VSS.t893 488.889
R1509 VSS.t1594 VSS.t614 488.889
R1510 VSS.t585 VSS.t2265 488.889
R1511 VSS.t2130 VSS.t2585 488.889
R1512 VSS.t1281 VSS.t2586 488.889
R1513 VSS.t743 VSS.t3123 482.221
R1514 VSS.t1890 VSS.t1042 480.461
R1515 VSS.n2941 VSS.t2077 480.461
R1516 VSS.t2830 VSS.t496 480.461
R1517 VSS.t826 VSS.t1305 480.461
R1518 VSS.t808 VSS.n408 480.461
R1519 VSS.n4302 VSS.t88 474.675
R1520 VSS.n3668 VSS.t2506 473.031
R1521 VSS.n3667 VSS.t685 473.031
R1522 VSS.t2559 VSS.t3459 472.031
R1523 VSS.t321 VSS.t2415 472.031
R1524 VSS.t208 VSS.t2346 472.031
R1525 VSS.t122 VSS.n3010 472.031
R1526 VSS.t2322 VSS.t2353 472.031
R1527 VSS.t1053 VSS.t733 472.031
R1528 VSS.t3407 VSS.n2893 472.031
R1529 VSS.t3463 VSS.t3051 472.031
R1530 VSS.t3483 VSS.t643 472.031
R1531 VSS.t3368 VSS.t1384 472.031
R1532 VSS.t417 VSS.t1189 472.031
R1533 VSS.n2472 VSS.t3083 472.031
R1534 VSS.t3456 VSS.t34 472.031
R1535 VSS.n340 VSS.t588 472.031
R1536 VSS.t3341 VSS.t1970 472.031
R1537 VSS.t1262 VSS.t54 472.031
R1538 VSS.n4302 VSS.t3659 471.308
R1539 VSS.t2692 VSS.n4301 471.308
R1540 VSS.n4301 VSS.t366 471.308
R1541 VSS.t1708 VSS.t1557 463.603
R1542 VSS.t2878 VSS.t1149 463.603
R1543 VSS.t3467 VSS.t468 463.603
R1544 VSS.t1505 VSS.t943 463.603
R1545 VSS.t1218 VSS.t2471 463.603
R1546 VSS.t45 VSS.t1706 458.776
R1547 VSS.t3557 VSS.t3384 455.173
R1548 VSS.t3066 VSS.t2357 455.173
R1549 VSS.t1394 VSS.t3132 455.173
R1550 VSS.t3058 VSS.t1612 455.173
R1551 VSS.t943 VSS.t906 455.173
R1552 VSS.t1688 VSS.t1768 455.173
R1553 VSS.t1269 VSS.t1572 455.173
R1554 VSS.t1955 VSS.t1218 455.173
R1555 VSS.t2208 VSS.t3208 455.173
R1556 VSS.t2458 VSS.t3222 455.173
R1557 VSS.t3665 VSS.t1113 447.743
R1558 VSS.t1049 VSS.t2226 446.743
R1559 VSS.t3387 VSS.t202 446.743
R1560 VSS.t2772 VSS.t3467 446.743
R1561 VSS.t356 VSS.t1659 446.743
R1562 VSS.t3370 VSS.t1815 446.743
R1563 VSS.t1602 VSS.t3435 446.743
R1564 VSS.t187 VSS.t1020 446.743
R1565 VSS.t1790 VSS.n4239 445.438
R1566 VSS.t3348 VSS.n4207 445.438
R1567 VSS.t1620 VSS.t2556 444.377
R1568 VSS.t2787 VSS.t3365 438.315
R1569 VSS.t3628 VSS.t2786 438.315
R1570 VSS.t3497 VSS.t2477 438.315
R1571 VSS.t228 VSS.n3011 438.315
R1572 VSS.t3394 VSS.t735 438.315
R1573 VSS.t2187 VSS.n2941 438.315
R1574 VSS.t2602 VSS.n2336 438.315
R1575 VSS.t478 VSS.t889 438.315
R1576 VSS.n408 VSS.t1416 438.315
R1577 VSS.t506 VSS.t3650 429.885
R1578 VSS.t1923 VSS.t2422 429.885
R1579 VSS.t2905 VSS.t443 429.885
R1580 VSS.t3016 VSS.t1097 429.885
R1581 VSS.t92 VSS.t2466 429.885
R1582 VSS.t2491 VSS.t1657 421.457
R1583 VSS.t1082 VSS.t2719 421.457
R1584 VSS.t134 VSS.t951 421.457
R1585 VSS.t1043 VSS.t854 421.457
R1586 VSS.t2987 VSS.n368 421.457
R1587 VSS.t3301 VSS.t2018 419.603
R1588 VSS.t259 VSS.t251 413.027
R1589 VSS.t1129 VSS.t802 413.027
R1590 VSS.t1095 VSS.t3193 413.027
R1591 VSS.t2702 VSS.t3692 413.027
R1592 VSS.t2281 VSS.t809 413.027
R1593 VSS.t2374 VSS.t1415 413.027
R1594 VSS.t3479 VSS.t1940 405.053
R1595 VSS.t1796 VSS.n1718 404.599
R1596 VSS.t2865 VSS.n1004 404.599
R1597 VSS.t2493 VSS.t3494 404.599
R1598 VSS.t3494 VSS.t747 404.599
R1599 VSS.t2554 VSS.t2005 404.599
R1600 VSS.n3033 VSS.t1573 404.599
R1601 VSS.t2771 VSS.t3349 404.599
R1602 VSS.t3155 VSS.t2944 404.599
R1603 VSS.t735 VSS.t914 404.599
R1604 VSS.t577 VSS.t1254 404.599
R1605 VSS.n2061 VSS.t1717 404.599
R1606 VSS.n2206 VSS.t3080 404.599
R1607 VSS.n2337 VSS.t3570 404.599
R1608 VSS.t3632 VSS.t2822 404.599
R1609 VSS.t2576 VSS.n957 404.599
R1610 VSS.t2008 VSS.t887 404.599
R1611 VSS.n548 VSS.t757 404.599
R1612 VSS.n3717 VSS.t2026 404.599
R1613 VSS.t2765 VSS.t2797 403.979
R1614 VSS.t1930 VSS.t1928 401.39
R1615 VSS.t1925 VSS.t1930 401.39
R1616 VSS.t1928 VSS.t1935 401.39
R1617 VSS.t1932 VSS.t1935 401.39
R1618 VSS.t1110 VSS.t2765 397.247
R1619 VSS.t2002 VSS.n1444 396.17
R1620 VSS.t1685 VSS.t638 396.17
R1621 VSS.t1415 VSS.t2281 396.17
R1622 VSS.t2114 VSS.t1227 396.17
R1623 VSS.t339 VSS.t2339 391.474
R1624 VSS.t3442 VSS.t3644 387.74
R1625 VSS.t2761 VSS.t542 387.74
R1626 VSS.t2393 VSS.t634 387.74
R1627 VSS.t690 VSS.t1861 387.74
R1628 VSS.t116 VSS.t2374 387.74
R1629 VSS.t2736 VSS.t3610 383.673
R1630 VSS.t1978 VSS.t2337 383.515
R1631 VSS.t2230 VSS.t1417 383.318
R1632 VSS.t75 VSS.t1677 383.318
R1633 VSS.t3548 VSS.t1679 383.318
R1634 VSS.t3060 VSS.t1845 383.318
R1635 VSS.t2516 VSS.t2745 383.318
R1636 VSS.t3057 VSS.t1670 383.318
R1637 VSS.t1576 VSS.n3628 381.279
R1638 VSS.n4144 VSS.t2850 380.635
R1639 VSS.t1710 VSS.t1708 379.31
R1640 VSS.t1359 VSS.t581 379.31
R1641 VSS.t206 VSS.t511 379.31
R1642 VSS.t3327 VSS.t2075 379.31
R1643 VSS.t1438 VSS.t1923 379.31
R1644 VSS.t1372 VSS.t895 379.31
R1645 VSS.t1491 VSS.t2405 379.31
R1646 VSS.t1419 VSS.n3668 375.163
R1647 VSS.t3207 VSS.n3960 372.932
R1648 VSS.t3365 VSS.t667 370.882
R1649 VSS.t2600 VSS.t1478 370.882
R1650 VSS.t126 VSS.t2932 370.882
R1651 VSS.t2740 VSS.n3293 370.882
R1652 VSS.t547 VSS.t3027 370.882
R1653 VSS.t2328 VSS.t547 370.882
R1654 VSS.n3294 VSS.t2734 370.882
R1655 VSS.t3096 VSS.t2446 370.882
R1656 VSS.t1467 VSS.t2769 370.882
R1657 VSS.t679 VSS.t2912 370.882
R1658 VSS.t1947 VSS.t2902 370.882
R1659 VSS.n2206 VSS.t1427 370.882
R1660 VSS.t1121 VSS.t263 370.882
R1661 VSS.t2952 VSS.t2279 370.882
R1662 VSS.t1667 VSS.t3178 370.882
R1663 VSS.t1966 VSS.t2073 370.882
R1664 VSS.n4220 VSS.n4219 369.245
R1665 VSS.t72 VSS.t2140 365.563
R1666 VSS.t3446 VSS.t953 363.582
R1667 VSS.t1322 VSS.t2034 363.582
R1668 VSS.t2030 VSS.t3111 362.452
R1669 VSS.n2893 VSS.t1222 362.452
R1670 VSS.t2424 VSS.t2497 362.452
R1671 VSS.t443 VSS.t3655 362.452
R1672 VSS.t3655 VSS.t417 362.452
R1673 VSS.t120 VSS.n2472 362.452
R1674 VSS.t3580 VSS.t356 362.452
R1675 VSS.t1473 VSS.t3255 362.452
R1676 VSS.t1020 VSS.t3417 362.452
R1677 VSS.t2219 VSS.t187 362.452
R1678 VSS.t3389 VSS.t1485 357.058
R1679 VSS.n4860 VSS.n1753 356.894
R1680 VSS.n4019 VSS.n3965 356.894
R1681 VSS.t3616 VSS.n2892 354.024
R1682 VSS.n2892 VSS.t790 354.024
R1683 VSS.t2784 VSS.n2473 354.024
R1684 VSS.n2473 VSS.t2778 354.024
R1685 VSS.t3072 VSS.t101 354.024
R1686 VSS.t1768 VSS.t146 354.024
R1687 VSS.t1298 VSS.t1688 354.024
R1688 VSS.t2073 VSS.t1972 354.024
R1689 VSS.t1263 VSS.t3690 354.024
R1690 VSS.t3690 VSS.t1269 354.024
R1691 VSS.t3138 VSS.t3576 353.904
R1692 VSS.n4225 VSS.n4221 353.882
R1693 VSS.n4234 VSS.n4220 353.882
R1694 VSS.n2966 VSS.n2963 352
R1695 VSS.t1153 VSS.t2738 349.62
R1696 VSS.t1729 VSS.t3531 349.62
R1697 VSS.n4297 VSS.n4296 347.404
R1698 VSS.n4297 VSS.n3878 347.3
R1699 VSS.t1456 VSS.n4891 347.212
R1700 VSS.t3111 VSS.t2028 345.594
R1701 VSS.t2041 VSS.t1085 345.594
R1702 VSS.t362 VSS.t3580 345.594
R1703 VSS.t3255 VSS.t1471 345.594
R1704 VSS.t891 VSS.t1372 345.594
R1705 VSS.n4276 VSS.t62 338.784
R1706 VSS.n4252 VSS.t59 338.784
R1707 VSS.t1356 VSS.t2991 337.166
R1708 VSS.t3285 VSS.t2749 337.166
R1709 VSS.t922 VSS.t126 337.166
R1710 VSS.t2932 VSS.t128 337.166
R1711 VSS.n3010 VSS.t1489 337.166
R1712 VSS.n3293 VSS.t3540 337.166
R1713 VSS.t3027 VSS.t619 337.166
R1714 VSS.t1160 VSS.t2328 337.166
R1715 VSS.n3294 VSS.t3070 337.166
R1716 VSS.t2446 VSS.t1053 337.166
R1717 VSS.t1465 VSS.t679 337.166
R1718 VSS.t2912 VSS.t675 337.166
R1719 VSS.t2213 VSS.n340 337.166
R1720 VSS.t2279 VSS.t1413 337.166
R1721 VSS.t3178 VSS.t2136 337.166
R1722 VSS.n4856 VSS.n1753 333.628
R1723 VSS.n4014 VSS.n3965 333.628
R1724 VSS.t2556 VSS.t2229 333.283
R1725 VSS.n5376 VSS.t2061 331.171
R1726 VSS.t1530 VSS.t1750 329.916
R1727 VSS.t2369 VSS.t2794 328.736
R1728 VSS.t149 VSS.t2830 328.736
R1729 VSS.t1861 VSS.t2414 328.736
R1730 VSS.t1227 VSS.t2113 328.736
R1731 VSS.t1506 VSS.t945 328.736
R1732 VSS.t1216 VSS.t2472 328.736
R1733 VSS.t2260 VSS.t2228 323.183
R1734 VSS.t3268 VSS.t2489 320.307
R1735 VSS.t3082 VSS.t2347 320.307
R1736 VSS.t204 VSS.t3442 320.307
R1737 VSS.t2518 VSS.t2618 320.307
R1738 VSS.t1462 VSS.t3549 320.307
R1739 VSS.t638 VSS.t2393 320.307
R1740 VSS.t2513 VSS.t3325 320.307
R1741 VSS.t1578 VSS.t774 320.307
R1742 VSS.t916 VSS.t0 320.307
R1743 VSS.t1000 VSS.t1809 320.307
R1744 VSS.t893 VSS.t2008 320.307
R1745 VSS.t759 VSS.t257 320.307
R1746 VSS.t642 VSS.t1262 320.307
R1747 VSS.t1518 VSS.t1830 319.817
R1748 VSS.t3659 VSS.t1964 319.817
R1749 VSS.t90 VSS.t3488 319.817
R1750 VSS.t1913 VSS.t1917 319.817
R1751 VSS.t366 VSS.t368 319.817
R1752 VSS.t720 VSS.t2260 319.817
R1753 VSS.t1037 VSS.t3239 318.553
R1754 VSS.t2229 VSS.t2259 315.173
R1755 VSS.n4863 VSS.n4862 312.094
R1756 VSS.n4022 VSS.n4021 312.094
R1757 VSS.t3646 VSS.t3409 311.877
R1758 VSS.t3424 VSS.t3077 311.877
R1759 VSS.t185 VSS.t1019 311.877
R1760 VSS.t1948 VSS.t796 308.572
R1761 VSS.t3377 VSS.t594 308.572
R1762 VSS.n228 VSS.t987 307.536
R1763 VSS.n909 VSS.t2033 307.536
R1764 VSS.n350 VSS.t1213 307.536
R1765 VSS.n798 VSS.t117 307.536
R1766 VSS.n765 VSS.t1006 307.536
R1767 VSS.n756 VSS.t1371 307.536
R1768 VSS.n514 VSS.t1464 307.536
R1769 VSS.n538 VSS.t566 307.536
R1770 VSS.n5392 VSS.t2098 307.536
R1771 VSS.n2052 VSS.t2523 307.536
R1772 VSS.n2188 VSS.t119 307.536
R1773 VSS.n2681 VSS.t2335 307.536
R1774 VSS.n2650 VSS.t462 307.536
R1775 VSS.n2801 VSS.t398 307.536
R1776 VSS.n2832 VSS.t402 307.536
R1777 VSS.n3424 VSS.t1284 307.536
R1778 VSS.n2925 VSS.t1310 307.536
R1779 VSS.n3141 VSS.t2601 307.536
R1780 VSS.n1452 VSS.t2331 307.536
R1781 VSS.n1078 VSS.t3437 307.536
R1782 VSS.n1017 VSS.t2527 307.536
R1783 VSS.n1682 VSS.t693 307.536
R1784 VSS.n3683 VSS.t721 307.536
R1785 VSS.n486 VSS.t2386 306.988
R1786 VSS.t3472 VSS.t2759 306.94
R1787 VSS.t1696 VSS.t1676 306.94
R1788 VSS.t2245 VSS.t2307 306.94
R1789 VSS.t2924 VSS.t3517 304.856
R1790 VSS.t3516 VSS.t3563 304.856
R1791 VSS.n5469 VSS.t584 304.238
R1792 VSS.n3311 VSS.t2342 304.238
R1793 VSS.n2983 VSS.t2072 304.238
R1794 VSS.n3251 VSS.t2070 304.238
R1795 VSS.n1756 VSS.t3154 303.978
R1796 VSS.t1421 VSS.t1626 303.8
R1797 VSS.t1570 VSS.t2493 303.449
R1798 VSS.t907 VSS.t939 303.449
R1799 VSS.t914 VSS.t737 303.449
R1800 VSS.t3331 VSS.t2495 303.449
R1801 VSS.t2495 VSS.t1994 303.449
R1802 VSS.t1692 VSS.t1470 303.449
R1803 VSS.t3641 VSS.t1468 303.449
R1804 VSS.t630 VSS.t2076 303.449
R1805 VSS.t869 VSS.t2469 303.449
R1806 VSS.t2797 VSS.t3665 302.985
R1807 VSS.n4865 VSS.t3211 299.248
R1808 VSS.n1756 VSS.t3211 299.248
R1809 VSS.t2121 VSS.t2692 296.252
R1810 VSS.n4278 VSS.n4277 296.18
R1811 VSS.t1071 VSS.t287 295.019
R1812 VSS.t251 VSS.t3382 295.019
R1813 VSS.t2673 VSS.t259 295.019
R1814 VSS.t2165 VSS.t1325 295.019
R1815 VSS.t419 VSS.t2905 295.019
R1816 VSS.t3068 VSS.t1727 295.019
R1817 VSS.t1817 VSS.t2321 295.019
R1818 VSS.t3692 VSS.t2981 295.019
R1819 VSS.t54 VSS.t3335 295.019
R1820 VSS.n4061 VSS.t962 294.036
R1821 VSS.n1824 VSS.t1174 294.036
R1822 VSS.n4233 VSS.n4232 292.5
R1823 VSS.n4232 VSS.t1546 292.5
R1824 VSS.n4218 VSS.n4216 292.5
R1825 VSS.n4216 VSS.t1546 292.5
R1826 VSS.n4223 VSS.n4222 292.5
R1827 VSS.n4222 VSS.t1546 292.5
R1828 VSS.n4188 VSS.n4187 292.5
R1829 VSS.t1801 VSS.n4188 292.5
R1830 VSS.n3928 VSS.n3922 292.5
R1831 VSS.t2715 VSS.n3928 292.5
R1832 VSS.n3912 VSS.n3910 292.5
R1833 VSS.n3910 VSS.t1807 292.5
R1834 VSS.n4190 VSS.n4189 292.5
R1835 VSS.n4189 VSS.t1801 292.5
R1836 VSS.n4182 VSS.n4181 292.5
R1837 VSS.t2715 VSS.n4182 292.5
R1838 VSS.n4169 VSS.n3930 292.5
R1839 VSS.n4169 VSS.t1805 292.5
R1840 VSS.n1761 VSS.t1453 292.252
R1841 VSS.n4117 VSS.t2159 292.252
R1842 VSS.n4224 VSS.n3890 290.296
R1843 VSS.n3117 VSS.t215 290.289
R1844 VSS.n4836 VSS.t2843 289.26
R1845 VSS.n4140 VSS.t2841 289.188
R1846 VSS.t1431 VSS.t2989 286.591
R1847 VSS.t2786 VSS.t321 286.591
R1848 VSS.t1657 VSS.t2908 286.591
R1849 VSS.t647 VSS.t3361 286.591
R1850 VSS.t3075 VSS.t466 286.591
R1851 VSS.t2719 VSS.t1535 286.591
R1852 VSS.t1584 VSS.t94 286.591
R1853 VSS.t1390 VSS.t3333 286.591
R1854 VSS.t897 VSS.t478 286.591
R1855 VSS.t1288 VSS.t1357 286.591
R1856 VSS.n4004 VSS.t1009 286.433
R1857 VSS.n4004 VSS.t182 286.433
R1858 VSS.n862 VSS.t2710 286.426
R1859 VSS.t1802 VSS.t2678 285.803
R1860 VSS.t1539 VSS.t1802 285.803
R1861 VSS.t1731 VSS.t1539 285.803
R1862 VSS.t1673 VSS.t1731 285.803
R1863 VSS.t1838 VSS.t1673 285.803
R1864 VSS.t2915 VSS.t1838 285.803
R1865 VSS.t2916 VSS.t2920 285.803
R1866 VSS.t2926 VSS.t2916 285.803
R1867 VSS.t2917 VSS.t2926 285.803
R1868 VSS.t3566 VSS.t3575 285.803
R1869 VSS.t3575 VSS.t3565 285.803
R1870 VSS.t3565 VSS.t3573 285.803
R1871 VSS.t3561 VSS.t1839 285.803
R1872 VSS.t1839 VSS.t3530 285.803
R1873 VSS.t3530 VSS.t1728 285.803
R1874 VSS.t1728 VSS.t2631 285.803
R1875 VSS.t2631 VSS.t1803 285.803
R1876 VSS.t1803 VSS.t1775 285.803
R1877 VSS.n4010 VSS.t1010 285.481
R1878 VSS.n4010 VSS.t180 285.481
R1879 VSS.t337 VSS.n3628 285.45
R1880 VSS.t1715 VSS.t2918 284.442
R1881 VSS.t3572 VSS.t2859 284.442
R1882 VSS.n3353 VSS.t1255 283.214
R1883 VSS.n785 VSS.t1168 283.175
R1884 VSS.n778 VSS.t1437 283.175
R1885 VSS.n1860 VSS.t2062 283.175
R1886 VSS.n4748 VSS.t1343 283.175
R1887 VSS.n4748 VSS.t2112 283.175
R1888 VSS.n4761 VSS.t2274 283.175
R1889 VSS.n4761 VSS.t1184 283.175
R1890 VSS.n4108 VSS.t2304 283.175
R1891 VSS.n4097 VSS.t1502 283.175
R1892 VSS.n4783 VSS.t160 283.175
R1893 VSS.n4783 VSS.t598 283.175
R1894 VSS.n1777 VSS.t1365 283.175
R1895 VSS.n1777 VSS.t194 283.175
R1896 VSS.t1554 VSS.t3026 283.082
R1897 VSS.t2678 VSS.t1774 283.082
R1898 VSS.t2920 VSS.t2919 283.082
R1899 VSS.t2923 VSS.t2917 283.082
R1900 VSS.t3569 VSS.t3566 283.082
R1901 VSS.t3573 VSS.t3564 283.082
R1902 VSS.t1775 VSS.t1786 283.082
R1903 VSS.t1844 VSS.t3025 283.082
R1904 VSS.t1324 VSS.t3446 282.786
R1905 VSS.t3367 VSS.t1322 282.786
R1906 VSS.t1194 VSS.t2742 282.786
R1907 VSS.t1516 VSS.t1518 282.786
R1908 VSS.t1964 VSS.t1962 282.786
R1909 VSS.t88 VSS.t90 282.786
R1910 VSS.t1917 VSS.t1915 282.786
R1911 VSS.t368 VSS.t370 282.786
R1912 VSS.t2930 VSS.t2257 282.786
R1913 VSS.n1897 VSS.t521 282.565
R1914 VSS.n1897 VSS.t2400 282.565
R1915 VSS.n1906 VSS.t1403 282.565
R1916 VSS.n1906 VSS.t704 282.565
R1917 VSS.n4069 VSS.t105 282.565
R1918 VSS.n1803 VSS.t1896 282.565
R1919 VSS.n1803 VSS.t535 282.565
R1920 VSS.n1792 VSS.t225 282.565
R1921 VSS.n1792 VSS.t860 282.565
R1922 VSS.n1747 VSS.n1746 282.353
R1923 VSS.n1736 VSS.n1730 282.353
R1924 VSS.n4049 VSS.n4048 282.353
R1925 VSS.n4026 VSS.n4023 282.353
R1926 VSS.n1726 VSS.t1457 282.327
R1927 VSS.n4120 VSS.t2157 282.327
R1928 VSS.n214 VSS.t613 282.147
R1929 VSS.n4225 VSS.n4224 281.771
R1930 VSS.n3093 VSS.t1814 281.25
R1931 VSS.n4843 VSS.t2855 281.13
R1932 VSS.n4137 VSS.t2851 281.13
R1933 VSS.n5461 VSS.t2207 280.945
R1934 VSS.n549 VSS.t1266 280.822
R1935 VSS.n2715 VSS.t365 280.822
R1936 VSS.n2876 VSS.t639 280.822
R1937 VSS.n3385 VSS.t680 280.822
R1938 VSS.n3347 VSS.t738 280.822
R1939 VSS.n3143 VSS.t127 280.822
R1940 VSS.n3224 VSS.t2350 280.822
R1941 VSS.n3670 VSS.t1420 280.822
R1942 VSS.t2232 VSS.t43 278.161
R1943 VSS.t776 VSS.t3074 278.161
R1944 VSS.t1886 VSS.t1297 278.161
R1945 VSS.t2417 VSS.t2451 278.161
R1946 VSS.t1099 VSS.t625 278.161
R1947 VSS.t1650 VSS.t92 278.161
R1948 VSS.t2414 VSS.t3370 278.161
R1949 VSS.t1598 VSS.t1594 278.161
R1950 VSS.t2113 VSS.t1602 278.161
R1951 VSS.n1831 VSS.t1647 276.098
R1952 VSS.n1905 VSS.t2616 276.098
R1953 VSS.n1905 VSS.t1541 276.098
R1954 VSS.n1918 VSS.t1716 276.098
R1955 VSS.n1918 VSS.t1552 276.098
R1956 VSS.n4068 VSS.t2727 276.098
R1957 VSS.n4083 VSS.t1822 276.098
R1958 VSS.n1776 VSS.t2871 276.098
R1959 VSS.n1776 VSS.t1735 276.098
R1960 VSS.n1785 VSS.t2884 276.098
R1961 VSS.n1785 VSS.t3474 276.098
R1962 VSS.n2525 VSS.t909 275.293
R1963 VSS.n2760 VSS.t517 275.293
R1964 VSS.n2977 VSS.t652 275.293
R1965 VSS.n3716 VSS.t2027 274.296
R1966 VSS.n4171 VSS.n4168 270.63
R1967 VSS.t2991 VSS.t3355 269.733
R1968 VSS.t2477 VSS.t3285 269.733
R1969 VSS.n3011 VSS.t230 269.733
R1970 VSS.t328 VSS.t3270 269.733
R1971 VSS.t731 VSS.t3394 269.733
R1972 VSS.t1391 VSS.t2465 269.733
R1973 VSS.t1661 VSS.t1377 269.733
R1974 VSS.n290 VSS.t3762 262.784
R1975 VSS.n291 VSS.t3719 262.784
R1976 VSS.n5404 VSS.t3715 262.784
R1977 VSS.n5405 VSS.t3749 262.784
R1978 VSS.n2066 VSS.t3724 262.784
R1979 VSS.n2067 VSS.t3767 262.784
R1980 VSS.n2659 VSS.t3721 262.784
R1981 VSS.n2660 VSS.t3744 262.784
R1982 VSS.n3038 VSS.t3731 262.784
R1983 VSS.n3039 VSS.t3745 262.784
R1984 VSS.n2808 VSS.t3752 262.784
R1985 VSS.n2809 VSS.t3716 262.784
R1986 VSS.n985 VSS.t3751 262.784
R1987 VSS.n964 VSS.t3742 262.784
R1988 VSS.n965 VSS.t3725 262.784
R1989 VSS.n1262 VSS.t3761 262.784
R1990 VSS.n1279 VSS.t3727 262.784
R1991 VSS.n1280 VSS.t3741 262.784
R1992 VSS.n3239 VSS.t3755 262.719
R1993 VSS.t1750 VSS.t1529 262.587
R1994 VSS.n3904 VSS.n3903 262.551
R1995 VSS.t1525 VSS.t2174 261.303
R1996 VSS.t3379 VSS.t3387 261.303
R1997 VSS.t202 VSS.t508 261.303
R1998 VSS.t1125 VSS.t3307 261.303
R1999 VSS.t3450 VSS.t515 261.303
R2000 VSS.t1659 VSS.t358 261.303
R2001 VSS.t658 VSS.t236 261.303
R2002 VSS.t2001 VSS.t2780 261.303
R2003 VSS.t2590 VSS.n3569 260.356
R2004 VSS.n3547 VSS.t3647 259.51
R2005 VSS.n3205 VSS.t2967 259.51
R2006 VSS.n1180 VSS.t3385 259.51
R2007 VSS.n1365 VSS.t1683 259.51
R2008 VSS.n1015 VSS.t2893 259.51
R2009 VSS.n4630 VSS.t2760 259.51
R2010 VSS.n44 VSS.t3720 259.082
R2011 VSS.n5332 VSS.t3728 259.082
R2012 VSS.n5245 VSS.t3737 259.082
R2013 VSS.n5120 VSS.t3718 259.082
R2014 VSS.n5078 VSS.t3710 259.082
R2015 VSS.n4924 VSS.t3758 259.082
R2016 VSS.n306 VSS.t3722 259.082
R2017 VSS.n633 VSS.t3759 259.082
R2018 VSS.n2323 VSS.t3766 259.082
R2019 VSS.n3448 VSS.t3707 259.082
R2020 VSS.n3302 VSS.t3709 259.082
R2021 VSS.n980 VSS.t3754 259.082
R2022 VSS.n1836 VSS.t3747 259.082
R2023 VSS.n3796 VSS.t3713 259.082
R2024 VSS.n4688 VSS.t3706 259.082
R2025 VSS.n1052 VSS.t1312 258.892
R2026 VSS.t2854 VSS.n4839 258.289
R2027 VSS.n5103 VSS.t2706 256.065
R2028 VSS.n2449 VSS.t1581 255.326
R2029 VSS.n1094 VSS.t69 255.326
R2030 VSS.t2415 VSS.t313 252.875
R2031 VSS.t1189 VSS.t413 252.875
R2032 VSS.t1522 VSS.t794 252.875
R2033 VSS.t12 VSS.t3456 252.875
R2034 VSS.t2372 VSS.t810 252.875
R2035 VSS.t1612 VSS.t3072 252.875
R2036 VSS.t1972 VSS.t3341 252.875
R2037 VSS.t3208 VSS.t2204 252.875
R2038 VSS.n1975 VSS.t671 246.506
R2039 VSS.n1960 VSS.t473 246.506
R2040 VSS.t3293 VSS.t1276 244.445
R2041 VSS.t56 VSS.t3436 244.445
R2042 VSS.t1532 VSS.t463 244.445
R2043 VSS.t3495 VSS.t3087 244.445
R2044 VSS.t1149 VSS.t2572 244.445
R2045 VSS.t714 VSS.t965 244.445
R2046 VSS.t496 VSS.t2831 244.445
R2047 VSS.t2928 VSS.t1590 244.445
R2048 VSS.t1305 VSS.t832 244.445
R2049 VSS.t3675 VSS.t461 244.445
R2050 VSS.t2126 VSS.t2971 244.445
R2051 VSS.t1463 VSS.t403 244.445
R2052 VSS.n4265 VSS.n4248 243.306
R2053 VSS.n41 VSS.t238 243.286
R2054 VSS.n101 VSS.t2056 243.286
R2055 VSS.n115 VSS.t1852 243.286
R2056 VSS.n136 VSS.t2149 243.286
R2057 VSS.n146 VSS.t1140 243.286
R2058 VSS.n162 VSS.t554 243.286
R2059 VSS.n176 VSS.t1016 243.286
R2060 VSS.n5125 VSS.t283 243.286
R2061 VSS.n5030 VSS.t1865 243.286
R2062 VSS.n247 VSS.t1908 243.286
R2063 VSS.n536 VSS.t1967 243.286
R2064 VSS.n2575 VSS.t487 243.286
R2065 VSS.n3793 VSS.t1038 243.286
R2066 VSS.n1022 VSS.t3455 242.965
R2067 VSS.n4897 VSS.t2292 242.945
R2068 VSS.n1628 VSS.t1709 242.395
R2069 VSS.t383 VSS.t1110 242.387
R2070 VSS.t2558 VSS.t1620 242.387
R2071 VSS.n854 VSS.t878 242.067
R2072 VSS.n2208 VSS.t442 242.067
R2073 VSS.n2435 VSS.t847 242.067
R2074 VSS.n2611 VSS.t27 242.067
R2075 VSS.n1479 VSS.t297 242.067
R2076 VSS.n1938 VSS.t855 241.971
R2077 VSS.n4897 VSS.t2139 241.695
R2078 VSS.n3101 VSS.t2904 241.054
R2079 VSS.n824 VSS.t2965 240.948
R2080 VSS.n1536 VSS.t777 240.575
R2081 VSS.n1118 VSS.t3095 240.575
R2082 VSS.n4323 VSS.t2768 240.575
R2083 VSS.n4201 VSS.t1807 240.221
R2084 VSS.t2715 VSS.n3927 240.221
R2085 VSS.n4247 VSS.n4210 239.843
R2086 VSS.n4274 VSS.n4210 239.435
R2087 VSS.n856 VSS.t1920 238.856
R2088 VSS.n823 VSS.t994 238.856
R2089 VSS.n786 VSS.t657 238.856
R2090 VSS.n741 VSS.t771 238.856
R2091 VSS.n2528 VSS.t1116 238.856
R2092 VSS.n1208 VSS.t499 238.856
R2093 VSS.n1029 VSS.t2236 238.856
R2094 VSS.n4723 VSS.t2246 238.856
R2095 VSS.t3475 VSS.n3957 238.794
R2096 VSS.n4037 VSS.t3477 238.794
R2097 VSS.n4037 VSS.t3568 238.794
R2098 VSS.t3479 VSS.n4144 238.794
R2099 VSS.n1104 VSS.t2990 238.311
R2100 VSS.n5032 VSS.t707 238.083
R2101 VSS.n727 VSS.t2264 238.083
R2102 VSS.n719 VSS.t725 238.083
R2103 VSS.n1420 VSS.t750 238.083
R2104 VSS.n2021 VSS.t3017 237.381
R2105 VSS.n1983 VSS.t3007 237.381
R2106 VSS.n2578 VSS.t3005 237.381
R2107 VSS.n1544 VSS.t3625 237.381
R2108 VSS.n2203 VSS.t533 237.332
R2109 VSS.n2113 VSS.t1385 237.327
R2110 VSS.n1085 VSS.t3595 237.327
R2111 VSS.t667 VSS.t2559 236.016
R2112 VSS.t2343 VSS.t3525 236.016
R2113 VSS.t2903 VSS.t3661 236.016
R2114 VSS.t2351 VSS.t2322 236.016
R2115 VSS.t733 VSS.t132 236.016
R2116 VSS.t3051 VSS.t3483 236.016
R2117 VSS.t643 VSS.t3410 236.016
R2118 VSS.t2480 VSS.t1061 236.016
R2119 VSS.t2164 VSS.t2712 236.016
R2120 VSS.t3287 VSS.t836 236.016
R2121 VSS.t3500 VSS.t826 236.016
R2122 VSS.t1723 VSS.t472 236.016
R2123 VSS.t3309 VSS.t1121 236.016
R2124 VSS.t2212 VSS.t1210 236.016
R2125 VSS.n2430 VSS.t1885 234.239
R2126 VSS.n2862 VSS.t1672 234.239
R2127 VSS.n3092 VSS.t3449 234.239
R2128 VSS.n3192 VSS.t1675 234.239
R2129 VSS.n1156 VSS.t1361 234.239
R2130 VSS.n4195 VSS.n4194 232.619
R2131 VSS.n207 VSS.t605 231.744
R2132 VSS.n1350 VSS.t373 231.613
R2133 VSS.n2223 VSS.t817 230.977
R2134 VSS.n1999 VSS.t137 230.977
R2135 VSS.n1126 VSS.t2376 230.977
R2136 VSS.n1613 VSS.t1244 230.977
R2137 VSS.n897 VSS.t1816 230.488
R2138 VSS.n399 VSS.t2504 230.488
R2139 VSS.n1987 VSS.t3288 230.488
R2140 VSS.n3518 VSS.t646 230.488
R2141 VSS.t2309 VSS.n4731 230.204
R2142 VSS.t1805 VSS.t87 229.578
R2143 VSS.n4731 VSS.t1248 228.571
R2144 VSS.n1581 VSS.t2980 228.052
R2145 VSS.t1039 VSS.t1035 227.815
R2146 VSS.n864 VSS.t3693 227.68
R2147 VSS.n581 VSS.t3691 227.68
R2148 VSS.n3447 VSS.t1349 227.68
R2149 VSS.n1196 VSS.t3695 227.68
R2150 VSS.n1619 VSS.t622 227.68
R2151 VSS.n1328 VSS.t197 227.587
R2152 VSS.t124 VSS.t80 227.587
R2153 VSS.t2075 VSS.t1127 227.587
R2154 VSS.t8 VSS.t2241 227.587
R2155 VSS.t885 VSS.t3552 227.587
R2156 VSS.t614 VSS.t2419 227.587
R2157 VSS.t586 VSS.t1604 227.587
R2158 VSS.n238 VSS.t709 226.882
R2159 VSS.n910 VSS.t591 226.882
R2160 VSS.n787 VSS.t2549 226.882
R2161 VSS.n464 VSS.t2266 226.882
R2162 VSS.n473 VSS.t727 226.882
R2163 VSS.n524 VSS.t868 226.882
R2164 VSS.n2130 VSS.t2421 226.882
R2165 VSS.n2856 VSS.t2483 226.882
R2166 VSS.n3007 VSS.t1872 226.882
R2167 VSS.n1389 VSS.t752 226.882
R2168 VSS.n1052 VSS.t2094 226.882
R2169 VSS.t1801 VSS.t86 226.538
R2170 VSS.n4909 VSS.n4908 226.296
R2171 VSS.n667 VSS.t1289 225.448
R2172 VSS.n990 VSS.t1528 224.214
R2173 VSS.n4172 VSS.n4171 223.498
R2174 VSS.n822 VSS.t616 223.315
R2175 VSS.n2163 VSS.t801 223.315
R2176 VSS.n2702 VSS.t983 223.315
R2177 VSS.n1006 VSS.t2133 223.315
R2178 VSS.n1821 VSS.n1820 221.894
R2179 VSS.n1893 VSS.n1891 221.894
R2180 VSS.n1893 VSS.n1892 221.894
R2181 VSS.n1885 VSS.n1883 221.894
R2182 VSS.n1885 VSS.n1884 221.894
R2183 VSS.n4058 VSS.n4057 221.894
R2184 VSS.n4078 VSS.n4077 221.894
R2185 VSS.n1810 VSS.n1779 221.894
R2186 VSS.n1810 VSS.n1780 221.894
R2187 VSS.n1797 VSS.n1787 221.894
R2188 VSS.n1797 VSS.n1788 221.894
R2189 VSS.t3123 VSS.t3147 221.45
R2190 VSS.t2654 VSS.n3813 220.476
R2191 VSS.t2685 VSS.n3990 220.476
R2192 VSS.t2225 VSS.t1333 219.157
R2193 VSS.n1445 VSS.t286 219.157
R2194 VSS.t2395 VSS.t636 219.157
R2195 VSS.t1441 VSS.t2167 219.157
R2196 VSS.t2182 VSS.t2408 219.157
R2197 VSS.t1643 VSS.t333 219.157
R2198 VSS.t490 VSS.t1067 219.157
R2199 VSS.t788 VSS.t3608 219.157
R2200 VSS.t1921 VSS.t1997 219.157
R2201 VSS.t1919 VSS.t1998 219.157
R2202 VSS.n466 VSS.t1239 219.157
R2203 VSS.t2263 VSS.t585 219.157
R2204 VSS.t905 VSS.t659 219.157
R2205 VSS.t3315 VSS.t2473 219.157
R2206 VSS.t175 VSS.t1952 219.157
R2207 VSS.n79 VSS.t3756 218.308
R2208 VSS.n5454 VSS.t3753 218.308
R2209 VSS.n392 VSS.t3735 218.308
R2210 VSS.n15 VSS.t3765 218.308
R2211 VSS.n2295 VSS.t3705 218.308
R2212 VSS.n1229 VSS.t3733 218.308
R2213 VSS.n1112 VSS.t3740 218.308
R2214 VSS.n4509 VSS.t3764 218.308
R2215 VSS.n2289 VSS.n2281 218
R2216 VSS.n4036 VSS.t3568 216.954
R2217 VSS.n4861 VSS.n1752 216.847
R2218 VSS.n4020 VSS.n3964 216.847
R2219 VSS.n4035 VSS.n3569 215.724
R2220 VSS.n988 VSS.t3173 215.407
R2221 VSS.n1312 VSS.t3197 215.407
R2222 VSS.n1867 VSS.n1850 214.956
R2223 VSS.n1760 VSS.n1752 214.589
R2224 VSS.n4863 VSS.n1751 214.589
R2225 VSS.n3964 VSS.n3963 214.589
R2226 VSS.n4030 VSS.n4022 214.589
R2227 VSS.n196 VSS.t3252 214.456
R2228 VSS.n5119 VSS.t3251 214.456
R2229 VSS.n5144 VSS.t3151 214.456
R2230 VSS.n184 VSS.t3152 214.456
R2231 VSS.n5182 VSS.t3245 214.456
R2232 VSS.n166 VSS.t3246 214.456
R2233 VSS.n5246 VSS.t3128 214.456
R2234 VSS.n5243 VSS.t3127 214.456
R2235 VSS.n5333 VSS.t3171 214.456
R2236 VSS.n5330 VSS.t3170 214.456
R2237 VSS.n78 VSS.t3116 214.456
R2238 VSS.n29 VSS.t3115 214.456
R2239 VSS.n43 VSS.t3162 214.456
R2240 VSS.n46 VSS.t3161 214.456
R2241 VSS.n4975 VSS.t3185 214.456
R2242 VSS.n266 VSS.t3186 214.456
R2243 VSS.n5077 VSS.t3201 214.456
R2244 VSS.n5076 VSS.t3200 214.456
R2245 VSS.n5111 VSS.t3261 214.456
R2246 VSS.n200 VSS.t3262 214.456
R2247 VSS.n4922 VSS.t3236 214.456
R2248 VSS.n4923 VSS.t3235 214.456
R2249 VSS.n304 VSS.t3257 214.456
R2250 VSS.n302 VSS.t3256 214.456
R2251 VSS.n290 VSS.t3230 214.456
R2252 VSS.n290 VSS.t3229 214.456
R2253 VSS.n291 VSS.t3243 214.456
R2254 VSS.n291 VSS.t3242 214.456
R2255 VSS.n5427 VSS.t3224 214.456
R2256 VSS.n5385 VSS.t3223 214.456
R2257 VSS.n5453 VSS.t3210 214.456
R2258 VSS.n20 VSS.t3209 214.456
R2259 VSS.n16 VSS.t3165 214.456
R2260 VSS.n5470 VSS.t3164 214.456
R2261 VSS.n632 VSS.t3180 214.456
R2262 VSS.n523 VSS.t3179 214.456
R2263 VSS.n490 VSS.t3218 214.456
R2264 VSS.n687 VSS.t3217 214.456
R2265 VSS.n393 VSS.t3215 214.456
R2266 VSS.n833 VSS.t3214 214.456
R2267 VSS.n324 VSS.t3143 214.456
R2268 VSS.n316 VSS.t3142 214.456
R2269 VSS.n5404 VSS.t3265 214.456
R2270 VSS.n5404 VSS.t3264 214.456
R2271 VSS.n5405 VSS.t3122 214.456
R2272 VSS.n5405 VSS.t3121 214.456
R2273 VSS.n2066 VSS.t3267 214.456
R2274 VSS.n2066 VSS.t3266 214.456
R2275 VSS.n2067 VSS.t3227 214.456
R2276 VSS.n2067 VSS.t3226 214.456
R2277 VSS.n2294 VSS.t3249 214.456
R2278 VSS.n2276 VSS.t3248 214.456
R2279 VSS.n2322 VSS.t3195 214.456
R2280 VSS.n2268 VSS.t3194 214.456
R2281 VSS.n2659 VSS.t3254 214.456
R2282 VSS.n2659 VSS.t3253 214.456
R2283 VSS.n2660 VSS.t3146 214.456
R2284 VSS.n2660 VSS.t3145 214.456
R2285 VSS.n3038 VSS.t3206 214.456
R2286 VSS.n3038 VSS.t3205 214.456
R2287 VSS.n3039 VSS.t3137 214.456
R2288 VSS.n3039 VSS.t3136 214.456
R2289 VSS.n3303 VSS.t3157 214.456
R2290 VSS.n3300 VSS.t3156 214.456
R2291 VSS.n3309 VSS.t3118 214.456
R2292 VSS.n2958 VSS.t3119 214.456
R2293 VSS.n3407 VSS.t3133 214.456
R2294 VSS.n2909 VSS.t3134 214.456
R2295 VSS.n3446 VSS.t3204 214.456
R2296 VSS.n3445 VSS.t3203 214.456
R2297 VSS.n2808 VSS.t3259 214.456
R2298 VSS.n2808 VSS.t3258 214.456
R2299 VSS.n2809 VSS.t3107 214.456
R2300 VSS.n2809 VSS.t3106 214.456
R2301 VSS.n3241 VSS.t3183 214.456
R2302 VSS.n3234 VSS.t3182 214.456
R2303 VSS.n1230 VSS.t3233 214.456
R2304 VSS.n1220 VSS.t3232 214.456
R2305 VSS.n1114 VSS.t3177 214.456
R2306 VSS.n1580 VSS.t3176 214.456
R2307 VSS.n985 VSS.t3221 214.456
R2308 VSS.n985 VSS.t3220 214.456
R2309 VSS.n987 VSS.t3174 214.456
R2310 VSS.n978 VSS.t3113 214.456
R2311 VSS.n976 VSS.t3112 214.456
R2312 VSS.n964 VSS.t3131 214.456
R2313 VSS.n964 VSS.t3130 214.456
R2314 VSS.n965 VSS.t3159 214.456
R2315 VSS.n965 VSS.t3158 214.456
R2316 VSS.n1296 VSS.t3110 214.456
R2317 VSS.n1263 VSS.t3109 214.456
R2318 VSS.n1265 VSS.t3198 214.456
R2319 VSS.n1262 VSS.t3168 214.456
R2320 VSS.n1262 VSS.t3167 214.456
R2321 VSS.n1279 VSS.t3192 214.456
R2322 VSS.n1279 VSS.t3191 214.456
R2323 VSS.n1280 VSS.t3238 214.456
R2324 VSS.n1280 VSS.t3237 214.456
R2325 VSS.n1837 VSS.t3140 214.456
R2326 VSS.n1818 VSS.t3139 214.456
R2327 VSS.n1839 VSS.t3148 214.456
R2328 VSS.n1853 VSS.t3149 214.456
R2329 VSS.n3610 VSS.t3189 214.456
R2330 VSS.n4507 VSS.t3188 214.456
R2331 VSS.n3798 VSS.t3241 214.456
R2332 VSS.n3795 VSS.t3240 214.456
R2333 VSS.n4687 VSS.t3125 214.456
R2334 VSS.n4686 VSS.t3124 214.456
R2335 VSS.t2730 VSS.t72 214.351
R2336 VSS.n320 VSS.t1302 214.197
R2337 VSS.n1964 VSS.n1963 211.242
R2338 VSS.t2366 VSS.t1888 210.728
R2339 VSS.t3426 VSS.t2330 210.728
R2340 VSS.t3374 VSS.t1309 210.728
R2341 VSS.t1224 VSS.t2048 210.728
R2342 VSS.t437 VSS.t3586 210.728
R2343 VSS.t1721 VSS.t3063 210.728
R2344 VSS.t3606 VSS.t1059 210.728
R2345 VSS.t670 VSS.t2656 210.728
R2346 VSS.t2032 VSS.t590 210.728
R2347 VSS.n3480 VSS.n2782 210.721
R2348 VSS.n2518 VSS.n2517 210.601
R2349 VSS.n2569 VSS.n2568 210.601
R2350 VSS.n2610 VSS.n2605 210.601
R2351 VSS.n3888 VSS.t1549 209.686
R2352 VSS.n236 VSS.n235 209.254
R2353 VSS.n930 VSS.n325 209.254
R2354 VSS.n339 VSS.n338 209.254
R2355 VSS.n735 VSS.n461 209.254
R2356 VSS.n476 VSS.n475 209.254
R2357 VSS.n661 VSS.n504 209.254
R2358 VSS.n573 VSS.n557 209.254
R2359 VSS.n2122 VSS.n2121 209.254
R2360 VSS.n2170 VSS.n2154 209.254
R2361 VSS.n2695 VSS.n2641 209.254
R2362 VSS.n2796 VSS.n2795 209.254
R2363 VSS.n2855 VSS.n2854 209.254
R2364 VSS.n3400 VSS.n2917 209.254
R2365 VSS.n2935 VSS.n2934 209.254
R2366 VSS.n2952 VSS.n2951 209.254
R2367 VSS.n3005 VSS.n3004 209.254
R2368 VSS.n3162 VSS.n3161 209.254
R2369 VSS.n3232 VSS.n3231 209.254
R2370 VSS.n1392 VSS.n1391 209.254
R2371 VSS.n1058 VSS.n1048 209.254
R2372 VSS.n1010 VSS.n1009 209.254
R2373 VSS.n1703 VSS.n1701 209.254
R2374 VSS.n3676 VSS.n3675 209.254
R2375 VSS.n2358 VSS.n2008 208.719
R2376 VSS.n1825 VSS.n1823 208.719
R2377 VSS.n1899 VSS.n1895 208.719
R2378 VSS.n1899 VSS.n1896 208.719
R2379 VSS.n1912 VSS.n1887 208.719
R2380 VSS.n1912 VSS.n1888 208.719
R2381 VSS.n4062 VSS.n4060 208.719
R2382 VSS.n4075 VSS.n4054 208.719
R2383 VSS.n1783 VSS.n1781 208.719
R2384 VSS.n1783 VSS.n1782 208.719
R2385 VSS.n1791 VSS.n1789 208.719
R2386 VSS.n1791 VSS.n1790 208.719
R2387 VSS.n3366 VSS.n2933 208.553
R2388 VSS.n5090 VSS.n213 207.965
R2389 VSS.n5456 VSS.n22 207.965
R2390 VSS.n357 VSS.n356 207.965
R2391 VSS.n363 VSS.n362 207.965
R2392 VSS.n582 VSS.n551 207.965
R2393 VSS.n1948 VSS.n1947 207.965
R2394 VSS.n2879 VSS.n2878 207.965
R2395 VSS.n2922 VSS.n2921 207.965
R2396 VSS.n3355 VSS.n2940 207.965
R2397 VSS.n3345 VSS.n2946 207.965
R2398 VSS.n3148 VSS.n2992 207.965
R2399 VSS.n3279 VSS.n3226 207.965
R2400 VSS.n4384 VSS.n3672 207.965
R2401 VSS.n1763 VSS.n1762 207.213
R2402 VSS.n4837 VSS.n4835 207.213
R2403 VSS.n2373 VSS.n2372 207.213
R2404 VSS.n2784 VSS.n2783 207.213
R2405 VSS.n3487 VSS.n2777 207.213
R2406 VSS.n3505 VSS.n2767 207.213
R2407 VSS.n2769 VSS.n2768 207.213
R2408 VSS.n2774 VSS.n2773 207.213
R2409 VSS.n3002 VSS.n3001 207.213
R2410 VSS.n4001 VSS.n3999 207.213
R2411 VSS.n4001 VSS.n4000 207.213
R2412 VSS.n4141 VSS.n4113 207.213
R2413 VSS.n4116 VSS.n4115 207.213
R2414 VSS.n826 VSS.n394 206.909
R2415 VSS.n2498 VSS.n2497 206.909
R2416 VSS.n1955 VSS.n1954 206.909
R2417 VSS.n2585 VSS.n2584 206.909
R2418 VSS.n1502 VSS.n1501 206.909
R2419 VSS.n1549 VSS.n1504 206.909
R2420 VSS.n2509 VSS.n1980 206.619
R2421 VSS.n2751 VSS.n2750 206.619
R2422 VSS.n1633 VSS.n1023 206.619
R2423 VSS.n3938 VSS.n3937 206.333
R2424 VSS.n379 VSS.n378 205.899
R2425 VSS.n840 VSS.n381 205.899
R2426 VSS.n2222 VSS.n2221 205.899
R2427 VSS.n2032 VSS.n2031 205.899
R2428 VSS.n1994 VSS.n1993 205.899
R2429 VSS.n1991 VSS.n1990 205.899
R2430 VSS.n2628 VSS.n2593 205.899
R2431 VSS.n1120 VSS.n1119 205.899
R2432 VSS.n1565 VSS.n1496 205.899
R2433 VSS.n1664 VSS.n1011 205.707
R2434 VSS.n374 VSS.n373 205.481
R2435 VSS.n2035 VSS.n2034 205.481
R2436 VSS.n2429 VSS.n2416 205.481
R2437 VSS.n2621 VSS.n2598 205.481
R2438 VSS.n2601 VSS.n2600 205.481
R2439 VSS.n1491 VSS.n1490 205.481
R2440 VSS.n53 VSS.n52 205.078
R2441 VSS.n5351 VSS.n100 205.078
R2442 VSS.n5318 VSS.n114 205.078
R2443 VSS.n5270 VSS.n135 205.078
R2444 VSS.n5237 VSS.n148 205.078
R2445 VSS.n5212 VSS.n161 205.078
R2446 VSS.n5175 VSS.n175 205.078
R2447 VSS.n194 VSS.n193 205.078
R2448 VSS.n244 VSS.n243 205.078
R2449 VSS.n5018 VSS.n249 205.078
R2450 VSS.n2571 VSS.n2570 205.078
R2451 VSS.n3804 VSS.n3791 205.078
R2452 VSS.n852 VSS.n372 204.692
R2453 VSS.n2038 VSS.n2037 204.692
R2454 VSS.n2229 VSS.n2228 204.692
R2455 VSS.n2414 VSS.n2413 204.692
R2456 VSS.n2486 VSS.n2485 204.692
R2457 VSS.n2588 VSS.n2587 204.692
R2458 VSS.n2615 VSS.n2604 204.692
R2459 VSS.n1484 VSS.n1483 204.692
R2460 VSS.n1559 VSS.n1558 204.692
R2461 VSS.n5200 VSS.n5199 204.457
R2462 VSS.n5163 VSS.n5162 204.457
R2463 VSS.n5137 VSS.n189 204.457
R2464 VSS.n1942 VSS.n1941 204.457
R2465 VSS.n1428 VSS.n1382 204.457
R2466 VSS.n1395 VSS.n1394 204.457
R2467 VSS.n3770 VSS.n3769 204.457
R2468 VSS.n3734 VSS.n3733 204.457
R2469 VSS.n1857 VSS.n1856 204.435
R2470 VSS.n4094 VSS.n4093 204.435
R2471 VSS.n2138 VSS.n2137 204.083
R2472 VSS.t2798 VSS.t75 203.893
R2473 VSS.t2791 VSS.t3548 203.893
R2474 VSS.t2795 VSS.t3057 203.893
R2475 VSS.n39 VSS.n38 203.619
R2476 VSS.n5353 VSS.n98 203.619
R2477 VSS.n112 VSS.n111 203.619
R2478 VSS.n133 VSS.n132 203.619
R2479 VSS.n150 VSS.n149 203.619
R2480 VSS.n159 VSS.n158 203.619
R2481 VSS.n5177 VSS.n173 203.619
R2482 VSS.n5131 VSS.n192 203.619
R2483 VSS.n5024 VSS.n246 203.619
R2484 VSS.n251 VSS.n250 203.619
R2485 VSS.n365 VSS.n364 203.619
R2486 VSS.n825 VSS.n395 203.619
R2487 VSS.n427 VSS.n426 203.619
R2488 VSS.n459 VSS.n458 203.619
R2489 VSS.n532 VSS.n531 203.619
R2490 VSS.n2532 VSS.n1973 203.619
R2491 VSS.n2566 VSS.n1961 203.619
R2492 VSS.n1206 VSS.n1205 203.619
R2493 VSS.n1041 VSS.n1040 203.619
R2494 VSS.n3806 VSS.n3790 203.619
R2495 VSS.n4672 VSS.n4671 203.619
R2496 VSS.n404 VSS.n403 203.526
R2497 VSS.n431 VSS.n430 203.526
R2498 VSS.n530 VSS.n529 203.526
R2499 VSS.n5382 VSS.n5381 203.526
R2500 VSS.n2703 VSS.n2638 203.526
R2501 VSS.n2215 VSS.n2214 203.519
R2502 VSS.n4877 VSS.n4876 203.294
R2503 VSS.n1741 VSS.n1737 203.294
R2504 VSS.n3955 VSS.n3952 203.294
R2505 VSS.n4047 VSS.n3947 203.294
R2506 VSS.n846 VSS.n377 203.262
R2507 VSS.n2119 VSS.n2118 203.016
R2508 VSS.n3131 VSS.n3130 203.016
R2509 VSS.n1703 VSS.n1702 203.016
R2510 VSS.n391 VSS.n390 202.724
R2511 VSS.n2025 VSS.n2024 202.724
R2512 VSS.n2243 VSS.n2023 202.724
R2513 VSS.n2489 VSS.n2488 202.724
R2514 VSS.n2418 VSS.n2417 202.463
R2515 VSS.n4998 VSS.n260 202.349
R2516 VSS.n884 VSS.n352 202.349
R2517 VSS.n589 VSS.n545 202.349
R2518 VSS.n2345 VSS.n2344 202.349
R2519 VSS.n1199 VSS.n1198 202.349
R2520 VSS.n1376 VSS.n1375 202.349
R2521 VSS.t2676 VSS.t1555 202.299
R2522 VSS.t2445 VSS.t3117 202.299
R2523 VSS.t739 VSS.t1338 202.299
R2524 VSS.t1442 VSS.t785 202.299
R2525 VSS.t877 VSS.t2977 202.299
R2526 VSS.t529 VSS.t2454 202.299
R2527 VSS.n2511 VSS.n2510 202.067
R2528 VSS.n2623 VSS.n2597 201.458
R2529 VSS.n1486 VSS.n1125 201.129
R2530 VSS.n4877 VSS.n1731 201.036
R2531 VSS.n4870 VSS.n1741 201.036
R2532 VSS.n1746 VSS.n1742 201.036
R2533 VSS.n4883 VSS.n1730 201.036
R2534 VSS.n4027 VSS.n3955 201.036
R2535 VSS.n4148 VSS.n3947 201.036
R2536 VSS.n4048 VSS.n3948 201.036
R2537 VSS.n4029 VSS.n4026 201.036
R2538 VSS.n613 VSS.n535 200.812
R2539 VSS.t2105 VSS.t62 200.761
R2540 VSS.t59 VSS.t2107 200.761
R2541 VSS.n5155 VSS.n5154 200.692
R2542 VSS.n5193 VSS.n5192 200.692
R2543 VSS.n4986 VSS.n4985 200.692
R2544 VSS.n5429 VSS.n5428 200.692
R2545 VSS.n936 VSS.n322 200.692
R2546 VSS.n3321 VSS.n3320 200.692
R2547 VSS.n3419 VSS.n3418 200.692
R2548 VSS.n1298 VSS.n1297 200.692
R2549 VSS.n5097 VSS.n209 200.516
R2550 VSS.n574 VSS.n556 200.516
R2551 VSS.n2402 VSS.n2401 200.516
R2552 VSS.n2406 VSS.n2405 200.516
R2553 VSS.n2442 VSS.n2408 200.516
R2554 VSS.n2589 VSS.n2586 200.516
R2555 VSS.n2616 VSS.n2603 200.516
R2556 VSS.n3533 VSS.n2754 200.516
R2557 VSS.n2765 VSS.n2764 200.516
R2558 VSS.n3488 VSS.n2776 200.516
R2559 VSS.n1242 VSS.n1188 200.516
R2560 VSS.n1164 VSS.n1163 200.516
R2561 VSS.n1384 VSS.n1383 200.516
R2562 VSS.n1529 VSS.n1514 200.516
R2563 VSS.n1606 VSS.n1605 200.516
R2564 VSS.n1612 VSS.n1611 200.516
R2565 VSS.n1032 VSS.n1031 200.516
R2566 VSS.n1057 VSS.n1049 200.516
R2567 VSS.n1635 VSS.n1634 200.516
R2568 VSS.n1649 VSS.n1648 200.516
R2569 VSS.n4334 VSS.n3694 200.516
R2570 VSS.n4625 VSS.n4624 200.516
R2571 VSS.n4164 VSS.n3936 200.516
R2572 VSS.n386 VSS.n385 200.508
R2573 VSS.n832 VSS.n387 200.508
R2574 VSS.n2234 VSS.n2027 200.508
R2575 VSS.n2480 VSS.n1989 200.508
R2576 VSS.n1952 VSS.n1951 200.508
R2577 VSS.n1555 VSS.n1500 200.508
R2578 VSS.n2106 VSS.n2105 200.231
R2579 VSS.n1542 VSS.n1508 200.231
R2580 VSS.n1524 VSS.n1518 200.231
R2581 VSS.n1079 VSS.n1038 200.231
R2582 VSS.n4317 VSS.n3702 200.231
R2583 VSS.n2521 VSS.n2520 200.127
R2584 VSS.n3334 VSS.n2954 200.127
R2585 VSS.n3159 VSS.n3158 200.127
R2586 VSS.n3200 VSS.n3199 200.127
R2587 VSS.n3591 VSS.n3590 200.127
R2588 VSS.n4481 VSS.n4480 200.127
R2589 VSS.n3655 VSS.n3654 200.127
R2590 VSS.n4578 VSS.n4577 200.127
R2591 VSS.n425 VSS.n422 200.105
R2592 VSS.n527 VSS.n526 200.105
R2593 VSS.n5379 VSS.n5378 200.105
R2594 VSS.n1176 VSS.n1175 200.105
R2595 VSS.n2129 VSS.n2128 199.966
R2596 VSS.n2152 VSS.n2151 199.966
R2597 VSS.n2997 VSS.n2996 199.966
R2598 VSS.n3194 VSS.n2979 199.917
R2599 VSS.n36 VSS.n35 199.739
R2600 VSS.n33 VSS.n32 199.739
R2601 VSS.n73 VSS.n72 199.739
R2602 VSS.n92 VSS.n91 199.739
R2603 VSS.n5311 VSS.n119 199.739
R2604 VSS.n5294 VSS.n125 199.739
R2605 VSS.n5263 VSS.n140 199.739
R2606 VSS.n5084 VSS.n217 199.739
R2607 VSS.n223 VSS.n222 199.739
R2608 VSS.n5062 VSS.n227 199.739
R2609 VSS.n5049 VSS.n232 199.739
R2610 VSS.n255 VSS.n254 199.739
R2611 VSS.n4993 VSS.n263 199.739
R2612 VSS.n279 VSS.n278 199.739
R2613 VSS.n4943 VSS.n283 199.739
R2614 VSS.n4936 VSS.n4917 199.739
R2615 VSS.n4931 VSS.n4920 199.739
R2616 VSS.n289 VSS.n287 199.739
R2617 VSS.n289 VSS.n288 199.739
R2618 VSS.n952 VSS.n311 199.739
R2619 VSS.n951 VSS.n312 199.739
R2620 VSS.n329 VSS.n328 199.739
R2621 VSS.n915 VSS.n332 199.739
R2622 VSS.n336 VSS.n335 199.739
R2623 VSS.n883 VSS.n353 199.739
R2624 VSS.n799 VSS.n418 199.739
R2625 VSS.n438 VSS.n437 199.739
R2626 VSS.n763 VSS.n443 199.739
R2627 VSS.n762 VSS.n446 199.739
R2628 VSS.n448 VSS.n447 199.739
R2629 VSS.n733 VSS.n463 199.739
R2630 VSS.n699 VSS.n480 199.739
R2631 VSS.n693 VSS.n483 199.739
R2632 VSS.n674 VSS.n496 199.739
R2633 VSS.n498 VSS.n497 199.739
R2634 VSS.n646 VSS.n513 199.739
R2635 VSS.n641 VSS.n516 199.739
R2636 VSS.n640 VSS.n517 199.739
R2637 VSS.n596 VSS.n540 199.739
R2638 VSS.n562 VSS.n561 199.739
R2639 VSS.n11 VSS.n10 199.739
R2640 VSS.n5422 VSS.n5394 199.739
R2641 VSS.n5421 VSS.n5395 199.739
R2642 VSS.n5399 VSS.n5397 199.739
R2643 VSS.n5399 VSS.n5398 199.739
R2644 VSS.n5403 VSS.n5401 199.739
R2645 VSS.n5403 VSS.n5402 199.739
R2646 VSS.n2060 VSS.n2059 199.739
R2647 VSS.n2065 VSS.n2063 199.739
R2648 VSS.n2065 VSS.n2064 199.739
R2649 VSS.n2086 VSS.n2085 199.739
R2650 VSS.n2057 VSS.n2056 199.739
R2651 VSS.n2098 VSS.n2097 199.739
R2652 VSS.n2150 VSS.n2149 199.739
R2653 VSS.n2709 VSS.n1949 199.739
R2654 VSS.n2693 VSS.n2642 199.739
R2655 VSS.n2686 VSS.n2645 199.739
R2656 VSS.n2679 VSS.n2649 199.739
R2657 VSS.n2665 VSS.n2656 199.739
R2658 VSS.n2665 VSS.n2657 199.739
R2659 VSS.n3032 VSS.n3031 199.739
R2660 VSS.n3037 VSS.n3035 199.739
R2661 VSS.n3037 VSS.n3036 199.739
R2662 VSS.n2816 VSS.n2814 199.739
R2663 VSS.n2816 VSS.n2815 199.739
R2664 VSS.n2830 VSS.n2829 199.739
R2665 VSS.n2839 VSS.n2838 199.739
R2666 VSS.n2846 VSS.n2845 199.739
R2667 VSS.n2869 VSS.n2865 199.739
R2668 VSS.n3454 VSS.n2895 199.739
R2669 VSS.n2906 VSS.n2905 199.739
R2670 VSS.n3372 VSS.n2930 199.739
R2671 VSS.n2938 VSS.n2937 199.739
R2672 VSS.n3029 VSS.n3027 199.739
R2673 VSS.n3029 VSS.n3028 199.739
R2674 VSS.n3025 VSS.n3024 199.739
R2675 VSS.n3068 VSS.n3067 199.739
R2676 VSS.n3022 VSS.n3021 199.739
R2677 VSS.n3074 VSS.n3073 199.739
R2678 VSS.n3077 VSS.n3076 199.739
R2679 VSS.n3014 VSS.n3013 199.739
R2680 VSS.n3111 VSS.n3110 199.739
R2681 VSS.n3129 VSS.n3128 199.739
R2682 VSS.n3171 VSS.n3170 199.739
R2683 VSS.n2981 VSS.n2980 199.739
R2684 VSS.n2973 VSS.n2972 199.739
R2685 VSS.n1255 VSS.n1179 199.739
R2686 VSS.n1174 VSS.n1173 199.739
R2687 VSS.n1369 VSS.n1148 199.739
R2688 VSS.n1451 VSS.n1450 199.739
R2689 VSS.n1140 VSS.n1139 199.739
R2690 VSS.n1573 VSS.n1116 199.739
R2691 VSS.n1594 VSS.n1593 199.739
R2692 VSS.n1080 VSS.n1037 199.739
R2693 VSS.n1066 VSS.n1065 199.739
R2694 VSS.n1642 VSS.n1641 199.739
R2695 VSS.n1678 VSS.n1677 199.739
R2696 VSS.n999 VSS.n998 199.739
R2697 VSS.n1712 VSS.n1710 199.739
R2698 VSS.n1712 VSS.n1711 199.739
R2699 VSS.n963 VSS.n961 199.739
R2700 VSS.n963 VSS.n962 199.739
R2701 VSS.n1291 VSS.n1273 199.739
R2702 VSS.n1291 VSS.n1274 199.739
R2703 VSS.n1278 VSS.n1276 199.739
R2704 VSS.n1278 VSS.n1277 199.739
R2705 VSS.n4540 VSS.n3596 199.739
R2706 VSS.n4534 VSS.n3599 199.739
R2707 VSS.n3608 VSS.n3607 199.739
R2708 VSS.n4502 VSS.n3614 199.739
R2709 VSS.n4494 VSS.n3618 199.739
R2710 VSS.n4489 VSS.n3621 199.739
R2711 VSS.n3636 VSS.n3635 199.739
R2712 VSS.n4447 VSS.n3640 199.739
R2713 VSS.n3649 VSS.n3648 199.739
R2714 VSS.n3665 VSS.n3664 199.739
R2715 VSS.n4366 VSS.n3680 199.739
R2716 VSS.n4353 VSS.n3685 199.739
R2717 VSS.n4347 VSS.n3688 199.739
R2718 VSS.n4341 VSS.n3691 199.739
R2719 VSS.n3705 VSS.n3704 199.739
R2720 VSS.n4308 VSS.n3707 199.739
R2721 VSS.n3745 VSS.n3744 199.739
R2722 VSS.n3757 VSS.n3756 199.739
R2723 VSS.n4593 VSS.n4592 199.739
R2724 VSS.n3572 VSS.n3571 199.739
R2725 VSS.n4607 VSS.n4606 199.739
R2726 VSS.n3566 VSS.n3565 199.739
R2727 VSS.n4633 VSS.n4632 199.739
R2728 VSS.n4650 VSS.n4649 199.739
R2729 VSS.n4669 VSS.n4668 199.739
R2730 VSS.n4675 VSS.n4674 199.739
R2731 VSS.n4678 VSS.n4677 199.739
R2732 VSS.n4681 VSS.n4680 199.739
R2733 VSS.n4684 VSS.n4683 199.739
R2734 VSS.n1618 VSS.n1098 199.662
R2735 VSS.n3327 VSS.n3326 199.541
R2736 VSS.n1248 VSS.n1184 199.352
R2737 VSS.n2411 VSS.n2410 199.052
R2738 VSS.n1321 VSS.n1259 199.052
R2739 VSS.n1155 VSS.n1152 199.052
R2740 VSS.n1028 VSS.n1027 199.052
R2741 VSS.n4202 VSS.t49 198.987
R2742 VSS.n2158 VSS.n2157 198.986
R2743 VSS.n2142 VSS.n2140 198.974
R2744 VSS.n2183 VSS.n2146 198.964
R2745 VSS.n2207 VSS.n2041 198.964
R2746 VSS.n2251 VSS.n2250 198.964
R2747 VSS.n2270 VSS.n2269 198.964
R2748 VSS.n2351 VSS.n2350 198.964
R2749 VSS.n2466 VSS.n2395 198.964
R2750 VSS.n2397 VSS.n2396 198.964
R2751 VSS.n2546 VSS.n2545 198.964
R2752 VSS.n2871 VSS.n2864 198.964
R2753 VSS.n3436 VSS.n2902 198.964
R2754 VSS.n3425 VSS.n2908 198.964
R2755 VSS.n3344 VSS.n2947 198.964
R2756 VSS.n3169 VSS.n3168 198.964
R2757 VSS.n1421 VSS.n1387 198.964
R2758 VSS.n1134 VSS.n1133 198.964
R2759 VSS.n1855 VSS.n1854 198.964
R2760 VSS.n4742 VSS.n4740 198.964
R2761 VSS.n4742 VSS.n4741 198.964
R2762 VSS.n4746 VSS.n4744 198.964
R2763 VSS.n4746 VSS.n4745 198.964
R2764 VSS.n4755 VSS.n4753 198.964
R2765 VSS.n4755 VSS.n4754 198.964
R2766 VSS.n4736 VSS.n4734 198.964
R2767 VSS.n4736 VSS.n4735 198.964
R2768 VSS.n4087 VSS.n4086 198.964
R2769 VSS.n4102 VSS.n4089 198.964
R2770 VSS.n4095 VSS.n4092 198.964
R2771 VSS.n4776 VSS.n4774 198.964
R2772 VSS.n4776 VSS.n4775 198.964
R2773 VSS.n4779 VSS.n4777 198.964
R2774 VSS.n4779 VSS.n4778 198.964
R2775 VSS.n4771 VSS.n4769 198.964
R2776 VSS.n4771 VSS.n4770 198.964
R2777 VSS.n4792 VSS.n4790 198.964
R2778 VSS.n4792 VSS.n4791 198.964
R2779 VSS.n4465 VSS.n3631 198.964
R2780 VSS.n4436 VSS.n3645 198.964
R2781 VSS.n4403 VSS.n3660 198.964
R2782 VSS.n3583 VSS.n3582 198.964
R2783 VSS.n4663 VSS.n4662 198.964
R2784 VSS.n2576 VSS.n1957 198.77
R2785 VSS.n2595 VSS.n2594 198.77
R2786 VSS.n1435 VSS.n1379 198.77
R2787 VSS.n1301 VSS.n1267 198.696
R2788 VSS.n3531 VSS.n2756 198.654
R2789 VSS.n1186 VSS.n1185 198.654
R2790 VSS.n1358 VSS.n1357 198.654
R2791 VSS.n1046 VSS.n1045 198.654
R2792 VSS.n1644 VSS.n1643 198.654
R2793 VSS.n3563 VSS.n3562 198.654
R2794 VSS.n211 VSS.n210 198.475
R2795 VSS.n2455 VSS.n2399 198.475
R2796 VSS.n3486 VSS.n2779 198.475
R2797 VSS.n1020 VSS.n1019 198.475
R2798 VSS.n2142 VSS.n2141 198.248
R2799 VSS.t3100 VSS.t3064 197.776
R2800 VSS.t779 VSS.t1576 197.776
R2801 VSS.n3087 VSS.n3018 197.488
R2802 VSS.n4908 VSS.n1719 197.37
R2803 VSS.n872 VSS.n359 197.219
R2804 VSS.n2029 VSS.n2028 197.219
R2805 VSS.n1996 VSS.n1995 197.219
R2806 VSS.n2503 VSS.n1982 197.219
R2807 VSS.n3456 VSS.n2894 197.219
R2808 VSS.n1154 VSS.n1153 197.219
R2809 VSS.n1132 VSS.n1131 197.219
R2810 VSS.n1556 VSS.n1499 197.219
R2811 VSS.n3512 VSS.n2762 196.831
R2812 VSS.n3220 VSS.n3219 196.831
R2813 VSS.n1694 VSS.n994 196.619
R2814 VSS.t2520 VSS.t2198 196.613
R2815 VSS.t3576 VSS.t745 196.613
R2816 VSS.n305 VSS.n303 196.442
R2817 VSS.n317 VSS.n315 196.442
R2818 VSS.n896 VSS.n343 196.442
R2819 VSS.n383 VSS.n382 196.442
R2820 VSS.n414 VSS.n413 196.442
R2821 VSS.n424 VSS.n423 196.442
R2822 VSS.n455 VSS.n454 196.442
R2823 VSS.n488 VSS.n487 196.442
R2824 VSS.n653 VSS.n510 196.442
R2825 VSS.n614 VSS.n534 196.442
R2826 VSS.n5437 VSS.n5386 196.442
R2827 VSS.n2112 VSS.n2049 196.442
R2828 VSS.n2259 VSS.n2257 196.442
R2829 VSS.n2370 VSS.n2003 196.442
R2830 VSS.n2672 VSS.n2652 196.442
R2831 VSS.n2671 VSS.n2653 196.442
R2832 VSS.n3287 VSS.n3222 196.442
R2833 VSS.n2823 VSS.n2803 196.442
R2834 VSS.n2822 VSS.n2804 196.442
R2835 VSS.n3462 VSS.n2788 196.442
R2836 VSS.n3409 VSS.n2914 196.442
R2837 VSS.n3387 VSS.n2924 196.442
R2838 VSS.n2994 VSS.n2993 196.442
R2839 VSS.n3262 VSS.n3236 196.442
R2840 VSS.n1269 VSS.n1268 196.442
R2841 VSS.n1403 VSS.n1397 196.442
R2842 VSS.n1109 VSS.n1108 196.442
R2843 VSS.n1658 VSS.n1014 196.442
R2844 VSS.n996 VSS.n995 196.442
R2845 VSS.n979 VSS.n977 196.442
R2846 VSS.n2320 VSS.n2319 196.192
R2847 VSS.t2326 VSS.t1395 196.026
R2848 VSS.n2440 VSS.n2409 195.752
R2849 VSS.n1087 VSS.n1034 195.752
R2850 VSS.t2259 VSS.t1421 195.738
R2851 VSS.n780 VSS.n433 195.667
R2852 VSS.n2303 VSS.n2275 195.667
R2853 VSS.n2607 VSS.n2606 195.667
R2854 VSS.n3392 VSS.n2920 195.667
R2855 VSS.n1167 VSS.n1166 195.667
R2856 VSS.n1436 VSS.n1378 195.667
R2857 VSS.n1129 VSS.n1128 195.667
R2858 VSS.n1123 VSS.n1122 195.667
R2859 VSS.n1535 VSS.n1511 195.667
R2860 VSS.n2447 VSS.n2404 195.612
R2861 VSS.n3511 VSS.n2763 195.612
R2862 VSS.n4143 VSS.n4142 195
R2863 VSS.n4841 VSS.n4840 195
R2864 VSS.t2091 VSS.t2488 193.87
R2865 VSS.t2895 VSS.t68 193.87
R2866 VSS.t1024 VSS.t2368 193.87
R2867 VSS.t2728 VSS.t1684 193.87
R2868 VSS.t214 VSS.t3295 193.87
R2869 VSS.t1241 VSS.t2071 193.87
R2870 VSS.t1606 VSS.t77 193.87
R2871 VSS.t2482 VSS.t3345 193.87
R2872 VSS.t1484 VSS.t2973 193.87
R2873 VSS.t2506 VSS.t2510 193.698
R2874 VSS.t266 VSS.t264 193.698
R2875 VSS.t2160 VSS.t2516 193.698
R2876 VSS.t2337 VSS.t1202 193.698
R2877 VSS.n4838 VSS.t3697 191.613
R2878 VSS.t3699 VSS.n4879 191.613
R2879 VSS.n4879 VSS.t2927 191.613
R2880 VSS.n1745 VSS.t2922 191.613
R2881 VSS.t3701 VSS.n1745 191.613
R2882 VSS.t3703 VSS.n4866 191.613
R2883 VSS.n4278 VSS.t564 191.417
R2884 VSS.n5153 VSS.n5152 190.399
R2885 VSS.n5191 VSS.n5190 190.399
R2886 VSS.n4984 VSS.n4983 190.399
R2887 VSS.n5391 VSS.n5389 190.399
R2888 VSS.n938 VSS.n937 190.399
R2889 VSS.n3319 VSS.n3318 190.399
R2890 VSS.n3417 VSS.n3416 190.399
R2891 VSS.n19 VSS.n18 189.481
R2892 VSS.n3244 VSS.n3243 189.481
R2893 VSS.n2966 VSS.n2965 189.201
R2894 VSS.t1444 VSS.t2798 187.582
R2895 VSS.t685 VSS.t2791 187.582
R2896 VSS.t2339 VSS.t2795 187.582
R2897 VSS.t1626 VSS.t2230 185.542
R2898 VSS.t2176 VSS.t2367 185.441
R2899 VSS.t2371 VSS.t1274 185.441
R2900 VSS.t1690 VSS.t579 185.441
R2901 VSS.t1480 VSS.t804 185.441
R2902 VSS.t2788 VSS.t1944 185.441
R2903 VSS.t800 VSS.t2016 185.441
R2904 VSS.t14 VSS.t970 185.441
R2905 VSS.t1150 VSS.t2237 185.441
R2906 VSS.t476 VSS.t901 185.441
R2907 VSS.t2755 VSS.t1663 185.441
R2908 VSS.t2541 VSS.t3281 185.441
R2909 VSS.t565 VSS.t2570 185.441
R2910 VSS.t3556 VSS.t3339 185.441
R2911 VSS.n5362 VSS.n5361 185
R2912 VSS.n5360 VSS.n5359 185
R2913 VSS.n5304 VSS.n5303 185
R2914 VSS.n5302 VSS.n5301 185
R2915 VSS.n5287 VSS.n5286 185
R2916 VSS.n5285 VSS.n5284 185
R2917 VSS.n5256 VSS.n5255 185
R2918 VSS.n5254 VSS.n5253 185
R2919 VSS.n4969 VSS.n4968 185
R2920 VSS.n4961 VSS.n4960 185
R2921 VSS.n276 VSS.n275 185
R2922 VSS.n924 VSS.n923 185
R2923 VSS.n922 VSS.n326 185
R2924 VSS.n349 VSS.n348 185
R2925 VSS.n347 VSS.n346 185
R2926 VSS.n407 VSS.n406 185
R2927 VSS.n405 VSS.n401 185
R2928 VSS.n753 VSS.n752 185
R2929 VSS.n755 VSS.n754 185
R2930 VSS.n703 VSS.n702 185
R2931 VSS.n701 VSS.n478 185
R2932 VSS.n605 VSS.n604 185
R2933 VSS.n598 VSS.n597 185
R2934 VSS.n544 VSS.n543 185
R2935 VSS.n565 VSS.n564 185
R2936 VSS.n567 VSS.n566 185
R2937 VSS.n2197 VSS.n2196 185
R2938 VSS.n2195 VSS.n2139 185
R2939 VSS.n2311 VSS.n2310 185
R2940 VSS.n2313 VSS.n2312 185
R2941 VSS.n2375 VSS.n2374 185
R2942 VSS.n2383 VSS.n2382 185
R2943 VSS.n2390 VSS.n2389 185
R2944 VSS.n2458 VSS.n2457 185
R2945 VSS.n2460 VSS.n2459 185
R2946 VSS.n2422 VSS.n2421 185
R2947 VSS.n2424 VSS.n2423 185
R2948 VSS.n2490 VSS.n1985 185
R2949 VSS.n2492 VSS.n2491 185
R2950 VSS.n2555 VSS.n2554 185
R2951 VSS.n2553 VSS.n2552 185
R2952 VSS.n2719 VSS.n2718 185
R2953 VSS.n2717 VSS.n1943 185
R2954 VSS.n2881 VSS.n2880 185
R2955 VSS.n2883 VSS.n2882 185
R2956 VSS.n3523 VSS.n3522 185
R2957 VSS.n3525 VSS.n3524 185
R2958 VSS.n3474 VSS.n3473 185
R2959 VSS.n3472 VSS.n3471 185
R2960 VSS.n3085 VSS.n3084 185
R2961 VSS.n3083 VSS.n3082 185
R2962 VSS.n3100 VSS.n3099 185
R2963 VSS.n3186 VSS.n3185 185
R2964 VSS.n3184 VSS.n3183 185
R2965 VSS.n1162 VSS.n1161 185
R2966 VSS.n1160 VSS.n1158 185
R2967 VSS.n1459 VSS.n1458 185
R2968 VSS.n1461 VSS.n1460 185
R2969 VSS.n1602 VSS.n1601 185
R2970 VSS.n1604 VSS.n1603 185
R2971 VSS.t2726 VSS.t104 184.785
R2972 VSS.n4229 VSS.t1546 184.208
R2973 VSS.n4237 VSS.t1546 184.208
R2974 VSS.n4241 VSS.n4240 183.341
R2975 VSS.n4241 VSS.n4211 183.341
R2976 VSS.t3610 VSS.t1978 179.593
R2977 VSS.t1845 VSS.t2290 179.425
R2978 VSS.t2655 VSS.t1501 177.643
R2979 VSS.t2526 VSS.t2115 177.012
R2980 VSS.t1596 VSS.t3048 177.012
R2981 VSS.t1644 VSS.t212 177.012
R2982 VSS.t3043 VSS.t513 177.012
R2983 VSS.t1123 VSS.t397 177.012
R2984 VSS.t1537 VSS.t1151 177.012
R2985 VSS.t899 VSS.t3213 177.012
R2986 VSS.t1658 VSS.t2958 177.012
R2987 VSS.t3321 VSS.t453 177.012
R2988 VSS.t47 VSS.t1153 176.669
R2989 VSS.t716 VSS.t1173 175.917
R2990 VSS.n4017 VSS.t3263 175.411
R2991 VSS.t1173 VSS.t1171 173.849
R2992 VSS.t2686 VSS.t1646 173.849
R2993 VSS.t2198 VSS.t2196 173.849
R2994 VSS.t745 VSS.t743 173.849
R2995 VSS.n4295 VSS.n4294 172.139
R2996 VSS.t1417 VSS.t1423 171.27
R2997 VSS.t1425 VSS.t1419 171.27
R2998 VSS.t2510 VSS.t2508 171.27
R2999 VSS.t1069 VSS.t2084 171.27
R3000 VSS.t2084 VSS.t3100 171.27
R3001 VSS.t268 VSS.t266 171.27
R3002 VSS.t2162 VSS.t2160 171.27
R3003 VSS.t2745 VSS.t339 171.27
R3004 VSS.t1980 VSS.t779 171.27
R3005 VSS.t3279 VSS.t1980 171.27
R3006 VSS.t1202 VSS.t1204 171.27
R3007 VSS.t2398 VSS.t813 168.583
R3008 VSS.t1084 VSS.t3181 168.583
R3009 VSS.t1630 VSS.t1260 168.583
R3010 VSS.t1575 VSS.t1992 168.583
R3011 VSS.t1307 VSS.t683 168.583
R3012 VSS.t2561 VSS.t846 168.583
R3013 VSS.n2635 VSS.t355 168.583
R3014 VSS.t1562 VSS.t2202 168.583
R3015 VSS.n4903 VSS.t482 166.978
R3016 VSS.n3831 VSS.n3830 165.648
R3017 VSS.n3831 VSS.n3829 165.648
R3018 VSS.n3836 VSS.n1721 165.648
R3019 VSS.n4243 VSS.t1790 165.209
R3020 VSS.n4243 VSS.t3348 165.209
R3021 VSS.n2709 VSS.t363 164.097
R3022 VSS.n2938 VSS.t1261 164.097
R3023 VSS.n4271 VSS.n4270 163.742
R3024 VSS.t1485 VSS.t1729 163.653
R3025 VSS.t3531 VSS.t2590 163.653
R3026 VSS.t1836 VSS.t1696 163.266
R3027 VSS.n86 VSS.t3429 162.471
R3028 VSS.n109 VSS.t2100 162.471
R3029 VSS.n5278 VSS.t1406 162.471
R3030 VSS.n152 VSS.t2193 162.471
R3031 VSS.n155 VSS.t1983 162.471
R3032 VSS.n5106 VSS.t3685 162.471
R3033 VSS.n877 VSS.t1201 162.471
R3034 VSS.n470 VSS.t3033 162.471
R3035 VSS.n659 VSS.t1771 162.471
R3036 VSS.n2091 VSS.t2937 162.471
R3037 VSS.n2099 VSS.t2868 162.471
R3038 VSS.n2364 VSS.t326 162.471
R3039 VSS.n2534 VSS.t2785 162.471
R3040 VSS.n2539 VSS.t2663 162.471
R3041 VSS.n1966 VSS.t145 162.471
R3042 VSS.n3519 VSS.t3639 162.471
R3043 VSS.n3442 VSS.t1296 162.471
R3044 VSS.n1344 VSS.t3613 162.471
R3045 VSS.n1115 VSS.t3534 162.471
R3046 VSS.n1670 VSS.t1275 162.471
R3047 VSS.n3721 VSS.t2141 161.968
R3048 VSS.n23 VSS.t2201 161.744
R3049 VSS.n2359 VSS.t1642 161.302
R3050 VSS.n855 VSS.t2988 161.042
R3051 VSS.n1202 VSS.t201 160.8
R3052 VSS.n554 VSS.t1270 160.8
R3053 VSS.n2889 VSS.t637 160.8
R3054 VSS.n3394 VSS.t684 160.8
R3055 VSS.n2949 VSS.t740 160.8
R3056 VSS.n3152 VSS.t125 160.8
R3057 VSS.n3229 VSS.t2358 160.8
R3058 VSS.n4378 VSS.t1418 160.8
R3059 VSS.t961 VSS.t2156 160.701
R3060 VSS.t959 VSS.t2154 160.701
R3061 VSS.t957 VSS.t2152 160.701
R3062 VSS.t963 VSS.t2158 160.701
R3063 VSS.t2255 VSS.t3305 160.154
R3064 VSS.t2970 VSS.t532 160.154
R3065 VSS.t2720 VSS.t689 160.154
R3066 VSS.t3303 VSS.t1001 160.154
R3067 VSS.t2757 VSS.t3498 160.154
R3068 VSS.n25 VSS.t3431 160.017
R3069 VSS.n5324 VSS.t2102 160.017
R3070 VSS.n5276 VSS.t1408 160.017
R3071 VSS.n5225 VSS.t2191 160.017
R3072 VSS.n5224 VSS.t1985 160.017
R3073 VSS.n5104 VSS.t3682 160.017
R3074 VSS.n354 VSS.t1199 160.017
R3075 VSS.n746 VSS.t3073 160.017
R3076 VSS.n662 VSS.t1757 160.017
R3077 VSS.n2103 VSS.t2862 160.017
R3078 VSS.n2538 VSS.t2779 160.017
R3079 VSS.n1968 VSS.t2666 160.017
R3080 VSS.n1213 VSS.t209 160.017
R3081 VSS.n1574 VSS.t3536 160.017
R3082 VSS.n1007 VSS.t1277 160.017
R3083 VSS.n853 VSS.t2978 160.017
R3084 VSS.n2360 VSS.t331 160.017
R3085 VSS.n2900 VSS.t1291 160.017
R3086 VSS.n1340 VSS.t3621 160.017
R3087 VSS.n4183 VSS.t3347 159.642
R3088 VSS.n1656 VSS.t2992 159.45
R3089 VSS.n2054 VSS.t2943 159.315
R3090 VSS.t3263 VSS.n3958 159.224
R3091 VSS.n720 VSS.t3037 158.796
R3092 VSS.n2060 VSS.t446 158.583
R3093 VSS.n2546 VSS.t143 158.583
R3094 VSS.n4002 VSS.t2714 158.361
R3095 VSS.n4002 VSS.t1800 158.361
R3096 VSS.n3713 VSS.t3416 158.361
R3097 VSS.n3713 VSS.t754 158.361
R3098 VSS.n4902 VSS.t1398 158.361
R3099 VSS.n870 VSS.t2974 157.993
R3100 VSS.n2241 VSS.t2583 157.291
R3101 VSS.n1728 VSS.t1449 157.291
R3102 VSS.n457 VSS.t3059 157.291
R3103 VSS.n2078 VSS.t448 157.291
R3104 VSS.n4125 VSS.t1943 157.291
R3105 VSS.n2544 VSS.t1593 156.915
R3106 VSS.n2969 VSS.t2735 156.915
R3107 VSS.n3588 VSS.t2733 156.915
R3108 VSS.n3600 VSS.t2732 156.915
R3109 VSS.n3603 VSS.t2744 156.915
R3110 VSS.n3616 VSS.t2737 156.915
R3111 VSS.n4459 VSS.t2746 156.915
R3112 VSS.n3763 VSS.t2743 156.915
R3113 VSS.n3783 VSS.t2731 156.915
R3114 VSS.n3574 VSS.t2739 156.915
R3115 VSS.n2562 VSS.t1105 156.915
R3116 VSS.n3291 VSS.t2741 156.915
R3117 VSS.n1001 VSS.t1112 156.915
R3118 VSS.t3207 VSS.n3958 156.745
R3119 VSS.t49 VSS.t47 156.214
R3120 VSS.t2738 VSS.t3389 156.214
R3121 VSS.n1675 VSS.t2866 156.133
R3122 VSS.n2098 VSS.t2708 155.679
R3123 VSS.n3032 VSS.t650 155.679
R3124 VSS.n2505 VSS.t2195 155.51
R3125 VSS.n3532 VSS.t2384 155.51
R3126 VSS.n1636 VSS.t1148 155.51
R3127 VSS.n4885 VSS.t1447 155.286
R3128 VSS.n3521 VSS.t3637 155.286
R3129 VSS.n4127 VSS.t1941 155.286
R3130 VSS.n2236 VSS.t2581 155.286
R3131 VSS.t798 VSS.t3472 155.102
R3132 VSS.t592 VSS.t1948 155.102
R3133 VSS.t2307 VSS.t2311 155.102
R3134 VSS.t1706 VSS.t2247 155.102
R3135 VSS.t718 VSS.t45 155.102
R3136 VSS.t1677 VSS.t3550 154.958
R3137 VSS.t1679 VSS.t3060 154.958
R3138 VSS.t1670 VSS.t337 154.958
R3139 VSS.n59 VSS.t664 154.561
R3140 VSS.n65 VSS.t981 154.561
R3141 VSS.n5068 VSS.t629 154.561
R3142 VSS.n5011 VSS.t273 154.561
R3143 VSS.n4941 VSS.t2011 154.561
R3144 VSS.n4929 VSS.t2318 154.561
R3145 VSS.n294 VSS.t1957 154.561
R3146 VSS.n294 VSS.t761 154.561
R3147 VSS.n285 VSS.t1132 154.561
R3148 VSS.n639 VSS.t1136 154.561
R3149 VSS.n5420 VSS.t3276 154.561
R3150 VSS.n5414 VSS.t1521 154.561
R3151 VSS.n5414 VSS.t390 154.561
R3152 VSS.n5408 VSS.t1207 154.561
R3153 VSS.n5408 VSS.t936 154.561
R3154 VSS.n2070 VSS.t977 154.561
R3155 VSS.n2070 VSS.t219 154.561
R3156 VSS.n2084 VSS.t1074 154.561
R3157 VSS.n2654 VSS.t1959 154.561
R3158 VSS.n2658 VSS.t277 154.561
R3159 VSS.n2658 VSS.t1903 154.561
R3160 VSS.n3042 VSS.t3278 154.561
R3161 VSS.n3042 VSS.t2181 154.561
R3162 VSS.n2807 VSS.t1156 154.561
R3163 VSS.n2807 VSS.t113 154.561
R3164 VSS.n2805 VSS.t2565 154.561
R3165 VSS.n3361 VSS.t715 154.561
R3166 VSS.n3055 VSS.t1234 154.561
R3167 VSS.n3055 VSS.t1354 154.561
R3168 VSS.n3061 VSS.t1883 154.561
R3169 VSS.n3115 VSS.t561 154.561
R3170 VSS.n1371 VSS.t2442 154.561
R3171 VSS.n1689 VSS.t1891 154.561
R3172 VSS.n958 VSS.t1026 154.561
R3173 VSS.n958 VSS.t1229 154.561
R3174 VSS.n968 VSS.t392 154.561
R3175 VSS.n968 VSS.t291 154.561
R3176 VSS.n1289 VSS.t969 154.561
R3177 VSS.n1289 VSS.t2278 154.561
R3178 VSS.n1283 VSS.t85 154.561
R3179 VSS.n1283 VSS.t2324 154.561
R3180 VSS.n3597 VSS.t2598 154.561
R3181 VSS.n4514 VSS.t730 154.561
R3182 VSS.n4487 VSS.t1205 154.561
R3183 VSS.n4453 VSS.t2163 154.561
R3184 VSS.n4423 VSS.t269 154.561
R3185 VSS.n4397 VSS.t2509 154.561
R3186 VSS.n3686 VSS.t371 154.561
R3187 VSS.n4315 VSS.t1916 154.561
R3188 VSS.n3709 VSS.t89 154.561
R3189 VSS.n3749 VSS.t1963 154.561
R3190 VSS.n3741 VSS.t1517 154.561
R3191 VSS.n3576 VSS.t50 154.561
R3192 VSS.n4618 VSS.t100 154.561
R3193 VSS.n4647 VSS.t797 154.561
R3194 VSS.n4654 VSS.t595 154.561
R3195 VSS.n4729 VSS.t2310 154.561
R3196 VSS.n4711 VSS.t717 154.561
R3197 VSS.n4705 VSS.t141 154.561
R3198 VSS.n4699 VSS.t2197 154.561
R3199 VSS.n4693 VSS.t744 154.561
R3200 VSS.n2054 VSS.t2986 154.131
R3201 VSS.n1972 VSS.t3486 154.131
R3202 VSS.n2540 VSS.t2661 154.131
R3203 VSS.n1964 VSS.t3458 154.131
R3204 VSS.n2967 VSS.t3071 154.131
R3205 VSS.n2970 VSS.t3541 154.131
R3206 VSS.n1260 VSS.t2762 154.131
R3207 VSS.n1676 VSS.t3664 154.131
R3208 VSS.n4558 VSS.t1761 154.131
R3209 VSS.n4528 VSS.t3652 154.131
R3210 VSS.n4527 VSS.t2674 154.131
R3211 VSS.n4500 VSS.t1655 154.131
R3212 VSS.n3633 VSS.t340 154.131
R3213 VSS.n3739 VSS.t1195 154.131
R3214 VSS.n3729 VSS.t73 154.131
R3215 VSS.n4599 VSS.t3390 154.131
R3216 VSS.n2871 VSS.t930 153.673
R3217 VSS.n3025 VSS.t2551 153.673
R3218 VSS.n3068 VSS.t765 153.673
R3219 VSS.n3077 VSS.t2532 153.673
R3220 VSS.t2850 VSS.t2836 152.791
R3221 VSS.t2856 VSS.t2840 152.791
R3222 VSS.t2838 VSS.t2842 152.791
R3223 VSS.t2852 VSS.t2854 152.791
R3224 VSS.n2526 VSS.t2047 152.381
R3225 VSS.n1320 VSS.t2729 152.381
R3226 VSS.n5192 VSS.n168 152
R3227 VSS.n5154 VSS.n183 152
R3228 VSS.n4985 VSS.n268 152
R3229 VSS.n936 VSS.n935 152
R3230 VSS.n5430 VSS.n5429 152
R3231 VSS.n3418 VSS.n2911 152
R3232 VSS.n3320 VSS.n2960 152
R3233 VSS.n1299 VSS.n1298 152
R3234 VSS.n1867 VSS.n1866 152
R3235 VSS.n1870 VSS.n1869 152
R3236 VSS.n1849 VSS.n1846 152
R3237 VSS.t2090 VSS.t2892 151.725
R3238 VSS.n1625 VSS.t70 151.725
R3239 VSS.t3626 VSS.t344 151.725
R3240 VSS.t2468 VSS.t2282 151.725
R3241 VSS.t1295 VSS.t1352 151.725
R3242 VSS.t246 VSS.t3372 151.725
R3243 VSS.t558 VSS.t828 151.725
R3244 VSS.t1388 VSS.t1122 151.725
R3245 VSS.t3587 VSS.t2596 151.725
R3246 VSS.n764 VSS.t1640 150.922
R3247 VSS.n720 VSS.t2379 150.922
R3248 VSS.n713 VSS.t3499 150.922
R3249 VSS.n2220 VSS.t624 150.922
R3250 VSS.n2335 VSS.t2603 150.922
R3251 VSS.n2330 VSS.t819 150.922
R3252 VSS.n2329 VSS.t1246 150.922
R3253 VSS.n2279 VSS.t172 150.922
R3254 VSS.n2287 VSS.t1536 150.922
R3255 VSS.n2342 VSS.t2096 150.922
R3256 VSS.n2343 VSS.t3528 150.922
R3257 VSS.n3480 VSS.t2476 150.922
R3258 VSS.n3437 VSS.t1351 150.922
R3259 VSS.n3430 VSS.t1653 150.922
R3260 VSS.n1189 VSS.t2283 150.922
R3261 VSS.n1214 VSS.t3388 150.922
R3262 VSS.n1202 VSS.t3054 150.922
R3263 VSS.n1147 VSS.t375 150.922
R3264 VSS.n1468 VSS.t2573 150.922
R3265 VSS.n3719 VSS.t1396 150.922
R3266 VSS.n3715 VSS.t1400 150.922
R3267 VSS.n300 VSS.t1474 150.376
R3268 VSS.n944 VSS.t1064 150.376
R3269 VSS.n2076 VSS.t412 150.376
R3270 VSS.n3048 VSS.t2287 150.376
R3271 VSS.n974 VSS.t2031 150.376
R3272 VSS.n3049 VSS.t1747 150.101
R3273 VSS.n1671 VSS.t688 150.101
R3274 VSS.n3934 VSS.t2431 149.762
R3275 VSS.n1064 VSS.t3559 149.395
R3276 VSS.n1519 VSS.t1369 149.02
R3277 VSS.n3698 VSS.t384 149.02
R3278 VSS.n3109 VSS.t231 148.536
R3279 VSS.n3967 VSS.n3958 147.942
R3280 VSS.n3926 VSS.t1789 147.478
R3281 VSS.n521 VSS.t2137 147.411
R3282 VSS.n2004 VSS.t135 147.411
R3283 VSS.n3499 VSS.t644 147.411
R3284 VSS.n3464 VSS.t2460 147.411
R3285 VSS.n1398 VSS.t3286 147.411
R3286 VSS.n1512 VSS.t1209 147.411
R3287 VSS.n1588 VSS.t1977 147.411
R3288 VSS.n3960 VSS.n3957 147.405
R3289 VSS.n4253 VSS.t564 147.288
R3290 VSS.n3874 VSS.t3212 146.667
R3291 VSS.n4050 VSS.n4049 146.25
R3292 VSS.n4051 VSS.n4050 146.25
R3293 VSS.n4046 VSS.n4045 146.25
R3294 VSS.n4045 VSS.n4044 146.25
R3295 VSS.n4024 VSS.n4023 146.25
R3296 VSS.n4024 VSS.n3956 146.25
R3297 VSS.n4028 VSS.n3954 146.25
R3298 VSS.n4034 VSS.n3954 146.25
R3299 VSS.n4040 VSS.n3946 146.25
R3300 VSS.n4041 VSS.n4040 146.25
R3301 VSS.n4147 VSS.n4146 146.25
R3302 VSS.n4146 VSS.n4145 146.25
R3303 VSS.n4895 VSS.n4894 146.25
R3304 VSS.n4894 VSS.n4893 146.25
R3305 VSS.n3830 VSS.n1725 146.25
R3306 VSS.n4893 VSS.n1725 146.25
R3307 VSS.n3829 VSS.n3827 146.25
R3308 VSS.n3838 VSS.n3827 146.25
R3309 VSS.n3837 VSS.n3836 146.25
R3310 VSS.n3838 VSS.n3837 146.25
R3311 VSS.n1748 VSS.n1747 146.25
R3312 VSS.n4867 VSS.n1748 146.25
R3313 VSS.n4875 VSS.n4874 146.25
R3314 VSS.n4874 VSS.n4873 146.25
R3315 VSS.n1736 VSS.n1734 146.25
R3316 VSS.n4880 VSS.n1734 146.25
R3317 VSS.n4882 VSS.n4881 146.25
R3318 VSS.n4881 VSS.n4880 146.25
R3319 VSS.n4872 VSS.n4871 146.25
R3320 VSS.n4873 VSS.n4872 146.25
R3321 VSS.n4869 VSS.n4868 146.25
R3322 VSS.n4868 VSS.n4867 146.25
R3323 VSS.n4236 VSS.n4235 146.25
R3324 VSS.n4237 VSS.n4236 146.25
R3325 VSS.n4230 VSS.n4227 146.25
R3326 VSS.n4230 VSS.n4229 146.25
R3327 VSS.n4240 VSS.n4213 146.25
R3328 VSS.n4239 VSS.n4213 146.25
R3329 VSS.n4214 VSS.n4211 146.25
R3330 VSS.n4214 VSS.n4207 146.25
R3331 VSS.n1505 VSS.t1078 145.724
R3332 VSS.n2215 VSS.t2887 145.212
R3333 VSS.n3353 VSS.t578 145.212
R3334 VSS.n4472 VSS.t338 145.212
R3335 VSS.n3641 VSS.t3061 145.212
R3336 VSS.n4410 VSS.t3551 145.212
R3337 VSS.n4575 VSS.t155 145.212
R3338 VSS.n4655 VSS.t3378 145.212
R3339 VSS.n2176 VSS.t572 145.212
R3340 VSS.n3548 VSS.t3651 145.212
R3341 VSS.n2903 VSS.t2664 145.212
R3342 VSS.n3402 VSS.t1649 145.212
R3343 VSS.n3178 VSS.t1481 145.212
R3344 VSS.n1414 VSS.t3526 145.212
R3345 VSS.n3206 VSS.t2404 144.886
R3346 VSS.t140 VSS.t2686 144.874
R3347 VSS.n3443 VSS.t2050 144.365
R3348 VSS.t2872 VSS.t621 143.296
R3349 VSS.t3546 VSS.t1079 143.296
R3350 VSS.t310 VSS.t933 143.296
R3351 VSS.t1285 VSS.t2878 143.296
R3352 VSS.t812 VSS.t1811 143.296
R3353 VSS.t2119 VSS.t253 143.296
R3354 VSS.n2258 VSS.t467 142.821
R3355 VSS.n2274 VSS.t1433 142.821
R3356 VSS.n4861 VSS.n4860 141.554
R3357 VSS.n4020 VSS.n4019 141.554
R3358 VSS.n3838 VSS.t2138 141.261
R3359 VSS.n4893 VSS.t2528 141.261
R3360 VSS.n4858 VSS.t3154 140.754
R3361 VSS.n4858 VSS.t3212 140.754
R3362 VSS.n3888 VSS.n3887 139.548
R3363 VSS.n4199 VSS.n3912 139.06
R3364 VSS.n4227 VSS.n4218 138.166
R3365 VSS.n4235 VSS.n4218 138.166
R3366 VSS.t796 VSS.t798 137.143
R3367 VSS.t594 VSS.t592 137.143
R3368 VSS.t2311 VSS.t2309 137.143
R3369 VSS.t2247 VSS.t2245 137.143
R3370 VSS.n4732 VSS.t716 136.595
R3371 VSS.n3728 VSS.t1033 135.1
R3372 VSS.t3558 VSS.t351 134.867
R3373 VSS.n1327 VSS.t1568 134.867
R3374 VSS.t1873 VSS.t213 134.867
R3375 VSS.t1828 VSS.t806 134.867
R3376 VSS.t651 VSS.t3648 134.867
R3377 VSS.t336 VSS.t990 134.867
R3378 VSS.t571 VSS.t2529 134.867
R3379 VSS.t34 VSS.t474 134.867
R3380 VSS.n4300 VSS.t1425 134.57
R3381 VSS.n4110 VSS.t2303 133.901
R3382 VSS.n3931 VSS.n3930 133.026
R3383 VSS.t2834 VSS.t1169 132.456
R3384 VSS.n4036 VSS.t1248 132.245
R3385 VSS.t2156 VSS.n1919 131.276
R3386 VSS.t2651 VSS.t2654 130.654
R3387 VSS.t2648 VSS.t2651 130.654
R3388 VSS.t2649 VSS.t2648 130.654
R3389 VSS.t2652 VSS.t2649 130.654
R3390 VSS.t2647 VSS.t2650 130.654
R3391 VSS.t2650 VSS.t2653 130.654
R3392 VSS.t2653 VSS.t2879 130.654
R3393 VSS.t2879 VSS.t2882 130.654
R3394 VSS.t2882 VSS.t2881 130.654
R3395 VSS.t2881 VSS.t2880 130.654
R3396 VSS.t2880 VSS.t2645 130.654
R3397 VSS.t2645 VSS.t2646 130.654
R3398 VSS.t2646 VSS.t1715 130.654
R3399 VSS.t2918 VSS.t2921 130.654
R3400 VSS.t2921 VSS.t2924 130.654
R3401 VSS.t3517 VSS.t3513 130.654
R3402 VSS.t3513 VSS.t3514 130.654
R3403 VSS.t3514 VSS.t3524 130.654
R3404 VSS.t3524 VSS.t3508 130.654
R3405 VSS.t3508 VSS.t3509 130.654
R3406 VSS.t3509 VSS.t3515 130.654
R3407 VSS.t3515 VSS.t3510 130.654
R3408 VSS.t3510 VSS.t2814 130.654
R3409 VSS.t2814 VSS.t2815 130.654
R3410 VSS.t2815 VSS.t2801 130.654
R3411 VSS.t2801 VSS.t2804 130.654
R3412 VSS.t2804 VSS.t2813 130.654
R3413 VSS.t2813 VSS.t2809 130.654
R3414 VSS.t2809 VSS.t2802 130.654
R3415 VSS.t2802 VSS.t2812 130.654
R3416 VSS.t2812 VSS.t2699 130.654
R3417 VSS.t2699 VSS.t2691 130.654
R3418 VSS.t2691 VSS.t2700 130.654
R3419 VSS.t2623 VSS.t2694 130.654
R3420 VSS.t2622 VSS.t2623 130.654
R3421 VSS.t3026 VSS.t2622 130.654
R3422 VSS.t1553 VSS.t1554 130.654
R3423 VSS.t1774 VSS.t1553 130.654
R3424 VSS.t2914 VSS.t2915 130.654
R3425 VSS.t2919 VSS.t2914 130.654
R3426 VSS.t3564 VSS.t3567 130.654
R3427 VSS.t3567 VSS.t3561 130.654
R3428 VSS.t1786 VSS.t1843 130.654
R3429 VSS.t1843 VSS.t1844 130.654
R3430 VSS.t3025 VSS.t2627 130.654
R3431 VSS.t2627 VSS.t2624 130.654
R3432 VSS.t2624 VSS.t2697 130.654
R3433 VSS.t2698 VSS.t2695 130.654
R3434 VSS.t2695 VSS.t2696 130.654
R3435 VSS.t2696 VSS.t2803 130.654
R3436 VSS.t2803 VSS.t2805 130.654
R3437 VSS.t2805 VSS.t2811 130.654
R3438 VSS.t2811 VSS.t2816 130.654
R3439 VSS.t2816 VSS.t2810 130.654
R3440 VSS.t2810 VSS.t2817 130.654
R3441 VSS.t2817 VSS.t2808 130.654
R3442 VSS.t2808 VSS.t2818 130.654
R3443 VSS.t2818 VSS.t3523 130.654
R3444 VSS.t3523 VSS.t3518 130.654
R3445 VSS.t3518 VSS.t3520 130.654
R3446 VSS.t3520 VSS.t3507 130.654
R3447 VSS.t3507 VSS.t3519 130.654
R3448 VSS.t3519 VSS.t3512 130.654
R3449 VSS.t3512 VSS.t3511 130.654
R3450 VSS.t3511 VSS.t3516 130.654
R3451 VSS.t3563 VSS.t3562 130.654
R3452 VSS.t3562 VSS.t3572 130.654
R3453 VSS.t2859 VSS.t2643 130.654
R3454 VSS.t2643 VSS.t2644 130.654
R3455 VSS.t2644 VSS.t2844 130.654
R3456 VSS.t2844 VSS.t2848 130.654
R3457 VSS.t2848 VSS.t2849 130.654
R3458 VSS.t2849 VSS.t2845 130.654
R3459 VSS.t2845 VSS.t2689 130.654
R3460 VSS.t2689 VSS.t2681 130.654
R3461 VSS.t2681 VSS.t2688 130.654
R3462 VSS.t2684 VSS.t2682 130.654
R3463 VSS.t2682 VSS.t2690 130.654
R3464 VSS.t2690 VSS.t2683 130.654
R3465 VSS.t2683 VSS.t2685 130.654
R3466 VSS.n4121 VSS.n1919 130
R3467 VSS.n4891 VSS.n4890 130
R3468 VSS.n4296 VSS.n4295 129.748
R3469 VSS.n3887 VSS.n3878 129.385
R3470 VSS.t3477 VSS.n4036 129.317
R3471 VSS.n4270 VSS.n4248 128.982
R3472 VSS.n4732 VSS.t1942 128.25
R3473 VSS.n4264 VSS.n4263 128
R3474 VSS.n4263 VSS.n4249 128
R3475 VSS.t3263 VSS.n4016 127.18
R3476 VSS.t1313 VSS.t3454 126.438
R3477 VSS.t342 VSS.t341 126.438
R3478 VSS.t3386 VSS.t927 126.438
R3479 VSS.t569 VSS.t2409 126.438
R3480 VSS.t435 VSS.t816 126.438
R3481 VSS.t2536 VSS.t672 126.438
R3482 VSS.t488 VSS.t1106 126.438
R3483 VSS.t20 VSS.t3041 126.438
R3484 VSS.n4271 VSS.n4247 126.291
R3485 VSS.t3153 VSS.n3969 125.293
R3486 VSS.t1821 VSS.n4110 124.975
R3487 VSS.n4274 VSS.n4273 124.236
R3488 VSS.t1676 VSS.t3377 124.082
R3489 VSS.n200 VSS.t3723 121.927
R3490 VSS.n490 VSS.t3708 121.927
R3491 VSS.n987 VSS.t3729 121.927
R3492 VSS.n4801 VSS.t3635 118.727
R3493 VSS.n4866 VSS.n4865 118.281
R3494 VSS.t1329 VSS.t2134 118.008
R3495 VSS.t3535 VSS.t3544 118.008
R3496 VSS.t40 VSS.t3630 118.008
R3497 VSS.t3612 VSS.t3398 118.008
R3498 VSS.t2606 VSS.t545 118.008
R3499 VSS.t3460 VSS.t2249 118.008
R3500 VSS.t1126 VSS.t1250 118.008
R3501 VSS.t28 VSS.t3464 118.008
R3502 VSS.t354 VSS.t3317 118.008
R3503 VSS.t3452 VSS.t2968 118.008
R3504 VSS.t947 VSS.t234 118.008
R3505 VSS.t1999 VSS.t1220 118.008
R3506 VSS.n5463 VSS.n19 117.334
R3507 VSS.n3245 VSS.n3244 117.334
R3508 VSS.n1581 VSS.n1110 117.334
R3509 VSS.n4021 VSS.n3959 117.001
R3510 VSS.t3207 VSS.n3959 117.001
R3511 VSS.n4032 VSS.n4031 117.001
R3512 VSS.t3207 VSS.n4032 117.001
R3513 VSS.n3834 VSS.n3833 117.001
R3514 VSS.n3833 VSS.t480 117.001
R3515 VSS.n3832 VSS.n3831 117.001
R3516 VSS.t480 VSS.n3832 117.001
R3517 VSS.n1723 VSS.n1721 117.001
R3518 VSS.t480 VSS.n1723 117.001
R3519 VSS.n1759 VSS.n1749 117.001
R3520 VSS.n1749 VSS.t3211 117.001
R3521 VSS.n4862 VSS.n1750 117.001
R3522 VSS.n1750 VSS.t3211 117.001
R3523 VSS.n4179 VSS.n4178 117.001
R3524 VSS.n4178 VSS.n3927 117.001
R3525 VSS.n3925 VSS.n3921 117.001
R3526 VSS.n3926 VSS.n3925 117.001
R3527 VSS.n4193 VSS.n4192 117.001
R3528 VSS.n4194 VSS.n4193 117.001
R3529 VSS.n4174 VSS.n4173 117.001
R3530 VSS.n4173 VSS.n4172 117.001
R3531 VSS.n4197 VSS.n4196 117.001
R3532 VSS.n4196 VSS.n4195 117.001
R3533 VSS.n4265 VSS.n4264 115.201
R3534 VSS.n4264 VSS.n3906 115.201
R3535 VSS.n3374 VSS.n2929 114.376
R3536 VSS.n3208 VSS.n3207 114.376
R3537 VSS.n3278 VSS.n3227 114.376
R3538 VSS.n2196 VSS.n2195 111.43
R3539 VSS.n2956 VSS.n2955 111.15
R3540 VSS.n3285 VSS.n3223 111.15
R3541 VSS.n4546 VSS.n3593 111.15
R3542 VSS.n4478 VSS.n3625 111.15
R3543 VSS.n4417 VSS.n3653 111.15
R3544 VSS.n4585 VSS.n4584 111.15
R3545 VSS.n4043 VSS.n4042 111.001
R3546 VSS.n4239 VSS.n4238 110.838
R3547 VSS.n4256 VSS.t2639 109.695
R3548 VSS.t138 VSS.t1175 109.691
R3549 VSS.t2588 VSS.t3098 109.579
R3550 VSS.t1764 VSS.t245 109.579
R3551 VSS.t1482 VSS.t926 109.579
R3552 VSS.t2380 VSS.t755 109.579
R3553 VSS.t3363 VSS.t2024 109.579
R3554 VSS.t3588 VSS.t2701 109.579
R3555 VSS.t2459 VSS.t3465 109.579
R3556 VSS.t2582 VSS.t3018 109.579
R3557 VSS.t52 VSS.t3002 109.579
R3558 VSS.t1429 VSS.t2546 109.579
R3559 VSS.t770 VSS.t2037 109.579
R3560 VSS.t2267 VSS.t1634 109.579
R3561 VSS.n4284 VSS.n3906 108.8
R3562 VSS.n2929 VSS.t1693 108.505
R3563 VSS.n3207 VSS.t2607 108.505
R3564 VSS.n3227 VSS.t3067 108.505
R3565 VSS.t2759 VSS.t98 108.121
R3566 VSS.n3151 VSS.n3150 107.853
R3567 VSS.n3873 VSS.t2647 107.516
R3568 VSS.n3991 VSS.t2688 107.516
R3569 VSS.t2638 VSS.t2344 103.602
R3570 VSS.t2299 VSS.t2723 102.659
R3571 VSS.t1497 VSS.t3687 102.659
R3572 VSS.n4291 VSS.t2336 102.332
R3573 VSS.n2933 VSS.t2770 101.43
R3574 VSS.t3419 VSS.t249 101.15
R3575 VSS.t921 VSS.t2899 101.15
R3576 VSS.t1256 VSS.t2188 101.15
R3577 VSS.t2906 VSS.t1654 101.15
R3578 VSS.t405 VSS.t2782 101.15
R3579 VSS.t439 VSS.t2579 101.15
R3580 VSS.t818 VSS.t1245 101.15
R3581 VSS.t1282 VSS.t873 101.15
R3582 VSS.t528 VSS.t768 101.15
R3583 VSS.t724 VSS.t3031 101.15
R3584 VSS.t147 VSS.t1477 101.15
R3585 VSS.t483 VSS.t1399 101.15
R3586 VSS.n4250 VSS.t2105 100.38
R3587 VSS.t2107 VSS.n4250 100.38
R3588 VSS.n4043 VSS.t3481 100.368
R3589 VSS.t3560 VSS.n4043 100.368
R3590 VSS.n235 VSS.t3298 100.001
R3591 VSS.n325 VSS.t1625 100.001
R3592 VSS.n338 VSS.t3304 100.001
R3593 VSS.n403 VSS.t1599 100.001
R3594 VSS.n430 VSS.t1617 100.001
R3595 VSS.n461 VSS.t1605 100.001
R3596 VSS.n475 VSS.t2758 100.001
R3597 VSS.n504 VSS.t3312 100.001
R3598 VSS.n529 VSS.t3314 100.001
R3599 VSS.n557 VSS.t3336 100.001
R3600 VSS.n5381 VSS.t3322 100.001
R3601 VSS.n2121 VSS.t3354 100.001
R3602 VSS.n2154 VSS.t3352 100.001
R3603 VSS.n2638 VSS.t3324 100.001
R3604 VSS.n2641 VSS.t3318 100.001
R3605 VSS.n2795 VSS.t3308 100.001
R3606 VSS.n2854 VSS.t3346 100.001
R3607 VSS.n2917 VSS.t3320 100.001
R3608 VSS.n2934 VSS.t3330 100.001
R3609 VSS.n2951 VSS.t1611 100.001
R3610 VSS.n3004 VSS.t3296 100.001
R3611 VSS.n3161 VSS.t3364 100.001
R3612 VSS.n3231 VSS.t1607 100.001
R3613 VSS.n1391 VSS.t2754 100.001
R3614 VSS.n1048 VSS.t3306 100.001
R3615 VSS.n1009 VSS.t3294 100.001
R3616 VSS.n1701 VSS.t3358 100.001
R3617 VSS.n3675 VSS.t1627 100.001
R3618 VSS.n376 VSS.t2009 99.9005
R3619 VSS.n412 VSS.t597 99.9005
R3620 VSS.n469 VSS.t1534 99.9005
R3621 VSS.n493 VSS.t380 99.9005
R3622 VSS.n501 VSS.t1358 99.9005
R3623 VSS.n508 VSS.t2474 99.9005
R3624 VSS.n2020 VSS.t795 99.9005
R3625 VSS.n1182 VSS.t2619 99.9005
R3626 VSS.n1169 VSS.t932 99.9005
R3627 VSS.n1306 VSS.t3760 99.7825
R3628 VSS.n4143 VSS.t2856 98.2229
R3629 VSS.n4840 VSS.t2838 98.2229
R3630 VSS.n4839 VSS.n4838 98.1726
R3631 VSS.n4242 VSS.n4241 97.5005
R3632 VSS.n4243 VSS.n4242 97.5005
R3633 VSS.n4245 VSS.n4244 97.5005
R3634 VSS.n4244 VSS.n4243 97.5005
R3635 VSS.n5255 VSS.n5254 97.1434
R3636 VSS.n5286 VSS.n5285 97.1434
R3637 VSS.n5303 VSS.n5302 97.1434
R3638 VSS.n5361 VSS.n5360 97.1434
R3639 VSS.n566 VSS.n565 97.1434
R3640 VSS.n702 VSS.n701 97.1434
R3641 VSS.n754 VSS.n753 97.1434
R3642 VSS.n923 VSS.n922 97.1434
R3643 VSS.n2718 VSS.n2717 97.1434
R3644 VSS.n3473 VSS.n3472 97.1434
R3645 VSS.n1460 VSS.n1459 97.1434
R3646 VSS.n1603 VSS.n1602 97.1434
R3647 VSS.n3835 VSS.n3834 97.1299
R3648 VSS.n3834 VSS.n1722 97.1299
R3649 VSS.n3872 VSS.t2694 96.629
R3650 VSS.t2697 VSS.n3975 96.629
R3651 VSS.n4862 VSS.n4861 95.2476
R3652 VSS.n4021 VSS.n4020 95.2476
R3653 VSS.t2435 VSS.t2430 93.4991
R3654 VSS.t2389 VSS.t2432 93.4991
R3655 VSS.t1801 VSS.t1789 92.7441
R3656 VSS.t2086 VSS.t2117 92.7208
R3657 VSS.t1582 VSS.t2594 92.7208
R3658 VSS.t306 VSS.n1567 92.7208
R3659 VSS.t2774 VSS.t2475 92.7208
R3660 VSS.t2580 VSS.t3008 92.7208
R3661 VSS.t3085 VSS.t464 92.7208
R3662 VSS.t2983 VSS.t171 92.7208
R3663 VSS.n2474 VSS.t834 92.7208
R3664 VSS.t1877 VSS.t2995 92.7208
R3665 VSS.t2334 VSS.t158 92.7208
R3666 VSS.t866 VSS.t1600 92.7208
R3667 VSS.t1035 VSS.n3728 92.7157
R3668 VSS.n4224 VSS.n4223 90.9607
R3669 VSS.n4192 VSS.n4191 90.3534
R3670 VSS.n4192 VSS.n3913 90.3534
R3671 VSS.n3921 VSS.n3918 90.3534
R3672 VSS.n4186 VSS.n3921 90.3534
R3673 VSS.n4180 VSS.n4179 90.3534
R3674 VSS.n4179 VSS.n4176 90.3534
R3675 VSS.t108 VSS.t3553 90.1608
R3676 VSS.n4277 VSS.n4276 89.9245
R3677 VSS.t1940 VSS.t1942 89.7746
R3678 VSS.t1033 VSS.n3718 87.4177
R3679 VSS.t3375 VSS.n4202 87.3505
R3680 VSS.n2141 VSS.t1591 85.7148
R3681 VSS.n4254 VSS.t2736 85.7148
R3682 VSS.n4896 VSS.n1721 85.0829
R3683 VSS.n846 VSS.n376 84.6851
R3684 VSS.n726 VSS.n469 84.6851
R3685 VSS.n667 VSS.n501 84.6851
R3686 VSS.n1248 VSS.n1182 84.6851
R3687 VSS.t3657 VSS.t1243 84.2917
R3688 VSS.t323 VSS.t3501 84.2917
R3689 VSS.t2675 VSS.t1022 84.2917
R3690 VSS.t3599 VSS.t441 84.2917
R3691 VSS.t423 VSS.t623 84.2917
R3692 VSS.t911 VSS.t1580 84.2917
R3693 VSS.t2 VSS.t1057 84.2917
R3694 VSS.t2665 VSS.t2660 84.2917
R3695 VSS.t364 VSS.t2007 84.2917
R3696 VSS.t1616 VSS.t1167 84.2917
R3697 VSS.t2524 VSS.t1968 84.2917
R3698 VSS.n2979 VSS.t3649 83.899
R3699 VSS.t480 VSS.t2138 83.7104
R3700 VSS.t480 VSS.t2528 83.7104
R3701 VSS.n3909 VSS.n3907 83.5719
R3702 VSS.n4260 VSS.n3909 83.5719
R3703 VSS.n4269 VSS.n4268 83.5719
R3704 VSS.n4268 VSS.n4267 83.5719
R3705 VSS.n4266 VSS.n4265 83.5719
R3706 VSS.n4267 VSS.n4266 83.5719
R3707 VSS.n3908 VSS.n3906 83.5719
R3708 VSS.n4260 VSS.n3908 83.5719
R3709 VSS.n4272 VSS.n4209 83.5719
R3710 VSS.n4250 VSS.n4209 83.5719
R3711 VSS.n4210 VSS.n4208 83.5719
R3712 VSS.n4250 VSS.n4208 83.5719
R3713 VSS.n4199 VSS.n4198 83.1211
R3714 VSS.n415 VSS.n412 82.5518
R3715 VSS.n680 VSS.n493 82.5518
R3716 VSS.n509 VSS.n508 82.5518
R3717 VSS.n2248 VSS.n2020 82.5518
R3718 VSS.n1170 VSS.n1169 82.5518
R3719 VSS.n4856 VSS.n4855 81.9205
R3720 VSS.n4014 VSS.n4013 81.9205
R3721 VSS.n2297 VSS.n2278 81.4574
R3722 VSS.n1759 VSS.n1751 80.9605
R3723 VSS.n1760 VSS.n1759 80.9605
R3724 VSS.n4031 VSS.n3963 80.9605
R3725 VSS.n4031 VSS.n4030 80.9605
R3726 VSS.n4896 VSS.n4895 80.5652
R3727 VSS.t504 VSS.t98 79.915
R3728 VSS.n4202 VSS.n4201 79.0606
R3729 VSS.n4876 VSS.n1736 79.0593
R3730 VSS.n4876 VSS.n4875 79.0593
R3731 VSS.n4875 VSS.n1737 79.0593
R3732 VSS.n1747 VSS.n1737 79.0593
R3733 VSS.n4023 VSS.n3952 79.0593
R3734 VSS.n4046 VSS.n3952 79.0593
R3735 VSS.n4047 VSS.n4046 79.0593
R3736 VSS.n4049 VSS.n4047 79.0593
R3737 VSS.n4227 VSS.n4221 78.6829
R3738 VSS.n4235 VSS.n4234 78.6829
R3739 VSS.n4175 VSS.n3931 77.418
R3740 VSS.n376 VSS.t479 77.0434
R3741 VSS.n412 VSS.t2373 77.0434
R3742 VSS.n469 VSS.t1494 77.0434
R3743 VSS.n493 VSS.t1700 77.0434
R3744 VSS.n501 VSS.t1755 77.0434
R3745 VSS.n508 VSS.t186 77.0434
R3746 VSS.n2020 VSS.t1098 77.0434
R3747 VSS.n1182 VSS.t3443 77.0434
R3748 VSS.n1169 VSS.t207 77.0434
R3749 VSS.t2303 VSS.t2301 76.7706
R3750 VSS.t2301 VSS.t2305 76.7706
R3751 VSS.t2305 VSS.t2299 76.7706
R3752 VSS.t1501 VSS.t1499 76.7706
R3753 VSS.t1499 VSS.t1495 76.7706
R3754 VSS.t1495 VSS.t1497 76.7706
R3755 VSS.t3596 VSS.t1147 75.8626
R3756 VSS.t1208 VSS.t1366 75.8626
R3757 VSS.t2003 VSS.t169 75.8626
R3758 VSS.t924 VSS.t2271 75.8626
R3759 VSS.t2123 VSS.t805 75.8626
R3760 VSS.t2829 VSS.t2253 75.8626
R3761 VSS.t2828 VSS.t334 75.8626
R3762 VSS.t694 VSS.t3422 75.8626
R3763 VSS.t2711 VSS.t1200 75.8626
R3764 VSS.t991 VSS.t2964 75.8626
R3765 VSS.t1778 VSS.t2726 74.9853
R3766 VSS.t104 VSS.t106 74.9853
R3767 VSS.t106 VSS.t110 74.9853
R3768 VSS.t110 VSS.t108 74.9853
R3769 VSS.t3553 VSS.t1821 74.9853
R3770 VSS.n3874 VSS.n3813 74.8536
R3771 VSS.n91 VSS.t1702 74.2862
R3772 VSS.n119 VSS.t1695 74.2862
R3773 VSS.n125 VSS.t2365 74.2862
R3774 VSS.n140 VSS.t1767 74.2862
R3775 VSS.n332 VSS.t1818 74.2862
R3776 VSS.n382 VSS.t477 74.2862
R3777 VSS.n418 VSS.t2375 74.2862
R3778 VSS.n446 VSS.t2453 74.2862
R3779 VSS.n463 VSS.t1492 74.2862
R3780 VSS.n483 VSS.t946 74.2862
R3781 VSS.n496 VSS.t1769 74.2862
R3782 VSS.n497 VSS.t1689 74.2862
R3783 VSS.n513 VSS.t188 74.2862
R3784 VSS.n10 VSS.t1217 74.2862
R3785 VSS.n2257 VSS.t1100 74.2862
R3786 VSS.n1949 VSS.t3581 74.2862
R3787 VSS.n2788 VSS.t3466 74.2862
R3788 VSS.n1179 VSS.t3445 74.2862
R3789 VSS.n1173 VSS.t198 74.2862
R3790 VSS.n1450 VSS.t2082 74.2862
R3791 VSS.n1593 VSS.t1088 74.2862
R3792 VSS.n4240 VSS.n4212 73.4123
R3793 VSS.n4246 VSS.n4211 73.4123
R3794 VSS.n4263 VSS.n4262 73.1255
R3795 VSS.n4262 VSS.n4261 73.1255
R3796 VSS.n4283 VSS.n4282 73.1255
R3797 VSS.n4282 VSS.n4281 73.1255
R3798 VSS.n4257 VSS.n4248 73.1255
R3799 VSS.n4257 VSS.n4256 73.1255
R3800 VSS.n4251 VSS.n4247 73.1255
R3801 VSS.n4252 VSS.n4251 73.1255
R3802 VSS.n4275 VSS.n4274 73.1255
R3803 VSS.n4276 VSS.n4275 73.1255
R3804 VSS.n4296 VSS.n3877 73.1255
R3805 VSS.n3878 VSS.n3875 73.1255
R3806 VSS.n4170 VSS.n3931 73.1255
R3807 VSS.n4171 VSS.n4170 73.1255
R3808 VSS.n4200 VSS.n4199 73.1255
R3809 VSS.n4201 VSS.n4200 73.1255
R3810 VSS.n5199 VSS.t1567 72.8576
R3811 VSS.n5162 VSS.t1561 72.8576
R3812 VSS.n189 VSS.t1565 72.8576
R3813 VSS.n232 VSS.t3302 72.8576
R3814 VSS.n328 VSS.t1601 72.8576
R3815 VSS.n343 VSS.t3371 72.8576
R3816 VSS.n413 VSS.t1609 72.8576
R3817 VSS.n422 VSS.t2864 72.8576
R3818 VSS.n437 VSS.t1603 72.8576
R3819 VSS.n454 VSS.t1613 72.8576
R3820 VSS.n480 VSS.t2756 72.8576
R3821 VSS.n510 VSS.t3316 72.8576
R3822 VSS.n526 VSS.t1559 72.8576
R3823 VSS.n534 VSS.t3342 72.8576
R3824 VSS.n561 VSS.t3340 72.8576
R3825 VSS.n5378 VSS.t1563 72.8576
R3826 VSS.n5386 VSS.t3338 72.8576
R3827 VSS.n2049 VSS.t3369 72.8576
R3828 VSS.n2137 VSS.t2721 72.8576
R3829 VSS.n2149 VSS.t3300 72.8576
R3830 VSS.n1941 VSS.t1046 72.8576
R3831 VSS.n2642 VSS.t3310 72.8576
R3832 VSS.n2645 VSS.t3334 72.8576
R3833 VSS.n2838 VSS.t3326 72.8576
R3834 VSS.n2845 VSS.t3328 72.8576
R3835 VSS.n2914 VSS.t3344 72.8576
R3836 VSS.n2930 VSS.t3332 72.8576
R3837 VSS.n3326 VSS.t1623 72.8576
R3838 VSS.n3128 VSS.t3362 72.8576
R3839 VSS.n3170 VSS.t3350 72.8576
R3840 VSS.n3236 VSS.t1615 72.8576
R3841 VSS.n1175 VSS.t1569 72.8576
R3842 VSS.n1382 VSS.t1556 72.8576
R3843 VSS.n1394 VSS.t1571 72.8576
R3844 VSS.n1397 VSS.t2750 72.8576
R3845 VSS.n1065 VSS.t3366 72.8576
R3846 VSS.n1014 VSS.t3356 72.8576
R3847 VSS.n995 VSS.t3360 72.8576
R3848 VSS.n3680 VSS.t1621 72.8576
R3849 VSS.n3769 VSS.t1323 72.8576
R3850 VSS.n3733 VSS.t3447 72.8576
R3851 VSS.n3996 VSS.t3153 72.5303
R3852 VSS.t1646 VSS.t2520 72.437
R3853 VSS.n4168 VSS.t2430 72.3506
R3854 VSS.t3477 VSS.n3956 70.7543
R3855 VSS.n4044 VSS.t3568 70.7543
R3856 VSS.n4044 VSS.t3560 70.7543
R3857 VSS.n4051 VSS.t3481 70.7543
R3858 VSS.t3479 VSS.n4051 70.7543
R3859 VSS.n3718 VSS.t1037 70.3474
R3860 VSS.n235 VSS.t711 70.0005
R3861 VSS.n325 VSS.t1300 70.0005
R3862 VSS.n338 VSS.t589 70.0005
R3863 VSS.n403 VSS.t618 70.0005
R3864 VSS.n430 VSS.t2547 70.0005
R3865 VSS.n461 VSS.t2268 70.0005
R3866 VSS.n475 VSS.t723 70.0005
R3867 VSS.n504 VSS.t1287 70.0005
R3868 VSS.n529 VSS.t870 70.0005
R3869 VSS.n557 VSS.t1268 70.0005
R3870 VSS.n5381 VSS.t2203 70.0005
R3871 VSS.n2121 VSS.t2423 70.0005
R3872 VSS.n2154 VSS.t803 70.0005
R3873 VSS.n2638 VSS.t361 70.0005
R3874 VSS.n2641 VSS.t985 70.0005
R3875 VSS.n2795 VSS.t2481 70.0005
R3876 VSS.n2854 VSS.t631 70.0005
R3877 VSS.n2917 VSS.t678 70.0005
R3878 VSS.n2934 VSS.t1257 70.0005
R3879 VSS.n2951 VSS.t734 70.0005
R3880 VSS.n3004 VSS.t1874 70.0005
R3881 VSS.n3161 VSS.t123 70.0005
R3882 VSS.n3231 VSS.t2356 70.0005
R3883 VSS.n1391 VSS.t748 70.0005
R3884 VSS.n1048 VSS.t2092 70.0005
R3885 VSS.n1009 VSS.t2135 70.0005
R3886 VSS.n1701 VSS.t1526 70.0005
R3887 VSS.n3675 VSS.t1422 70.0005
R3888 VSS.n2278 VSS.t65 69.0554
R3889 VSS.n2278 VSS.t1435 68.7993
R3890 VSS.n1868 VSS.t3714 68.6994
R3891 VSS.n3830 VSS.n1722 68.5181
R3892 VSS.n3836 VSS.n3835 68.5181
R3893 VSS.n3835 VSS.n3829 68.5181
R3894 VSS.n4895 VSS.n1722 68.5181
R3895 VSS.t3347 VSS.t2715 68.4179
R3896 VSS.n1499 VSS.t2416 68.3082
R3897 VSS.n1514 VSS.t2382 68.3082
R3898 VSS.n3694 VSS.t3666 68.3082
R3899 VSS.n4033 VSS.n3956 67.8062
R3900 VSS.t2132 VSS.t687 67.4335
R3901 VSS.t1976 VSS.t459 67.4335
R3902 VSS.t302 VSS.t696 67.4335
R3903 VSS.t543 VSS.t1841 67.4335
R3904 VSS.t1252 VSS.n2942 67.4335
R3905 VSS.t677 VSS.t1648 67.4335
R3906 VSS.t1652 VSS.t1680 67.4335
R3907 VSS.t1350 VSS.t3403 67.4335
R3908 VSS.t2383 VSS.t502 67.4335
R3909 VSS.t3006 VSS.t2562 67.4335
R3910 VSS.t2194 VSS.t3471 67.4335
R3911 VSS.t1293 VSS.t2021 67.4335
R3912 VSS.t3485 VSS.t1115 67.4335
R3913 VSS.t3412 VSS.t3457 67.4335
R3914 VSS.t1476 VSS.t3089 67.4335
R3915 VSS.n4883 VSS.n4882 67.2005
R3916 VSS.n4882 VSS.n1731 67.2005
R3917 VSS.n4871 VSS.n4870 67.2005
R3918 VSS.n4870 VSS.n4869 67.2005
R3919 VSS.n4869 VSS.n1742 67.2005
R3920 VSS.n4029 VSS.n4028 67.2005
R3921 VSS.n4028 VSS.n4027 67.2005
R3922 VSS.n4027 VSS.n3946 67.2005
R3923 VSS.n4148 VSS.n4147 67.2005
R3924 VSS.n4147 VSS.n3948 67.2005
R3925 VSS.n2281 VSS.t2984 67.1434
R3926 VSS.n4261 VSS.t250 67.0365
R3927 VSS.n1740 VSS.n1731 66.8805
R3928 VSS.n4149 VSS.n4148 66.8805
R3929 VSS.n2554 VSS.n2553 66.462
R3930 VSS.n2459 VSS.n2458 66.462
R3931 VSS.n2312 VSS.n2311 66.462
R3932 VSS.t255 VSS.t3375 65.6822
R3933 VSS.t2639 VSS.t2636 65.0051
R3934 VSS.t2634 VSS.t2635 65.0051
R3935 VSS.t2632 VSS.t2633 65.0051
R3936 VSS.n4019 VSS.n4018 65.0005
R3937 VSS.n4018 VSS.n4017 65.0005
R3938 VSS.n4015 VSS.n4014 65.0005
R3939 VSS.n4016 VSS.n4015 65.0005
R3940 VSS.n4857 VSS.n4856 65.0005
R3941 VSS.n4858 VSS.n4857 65.0005
R3942 VSS.n4860 VSS.n4859 65.0005
R3943 VSS.n4859 VSS.n4858 65.0005
R3944 VSS.t1819 VSS.t2067 64.8806
R3945 VSS.t2723 VSS.t2655 64.2732
R3946 VSS.t3687 VSS.t3635 64.2732
R3947 VSS.t1169 VSS.t138 64.1585
R3948 VSS.t1175 VSS.t140 64.1585
R3949 VSS.n1869 VSS.n1849 62.9556
R3950 VSS.n406 VSS.n405 62.7697
R3951 VSS.n348 VSS.n347 62.7697
R3952 VSS.n2491 VSS.n2490 62.7697
R3953 VSS.n2423 VSS.n2422 62.7697
R3954 VSS.n3524 VSS.n3523 62.7697
R3955 VSS.n2882 VSS.n2881 62.7697
R3956 VSS.n3185 VSS.n3184 62.7697
R3957 VSS.n3084 VSS.n3083 62.7697
R3958 VSS.n1161 VSS.n1160 62.7697
R3959 VSS.t3392 VSS.t1237 62.2966
R3960 VSS.n4238 VSS.n4237 61.7917
R3961 VSS.n5255 VSS.t1893 61.4291
R3962 VSS.n5286 VSS.t2262 61.4291
R3963 VSS.n5303 VSS.t1304 61.4291
R3964 VSS.n5361 VSS.t2289 61.4291
R3965 VSS.n565 VSS.t1221 61.4291
R3966 VSS.n702 VSS.t948 61.4291
R3967 VSS.n754 VSS.t2457 61.4291
R3968 VSS.n923 VSS.t1538 61.4291
R3969 VSS.n2718 VSS.t2479 61.4291
R3970 VSS.n3472 VSS.t497 61.4291
R3971 VSS.n1459 VSS.t2575 61.4291
R3972 VSS.n1602 VSS.t2463 61.4291
R3973 VSS.t1395 VSS.t1039 60.9277
R3974 VSS.n232 VSS.t1514 60.5809
R3975 VSS.n328 VSS.t2597 60.5809
R3976 VSS.n343 VSS.t1860 60.5809
R3977 VSS.n413 VSS.t811 60.5809
R3978 VSS.n437 VSS.t1226 60.5809
R3979 VSS.n454 VSS.t382 60.5809
R3980 VSS.n480 VSS.t235 60.5809
R3981 VSS.n510 VSS.t996 60.5809
R3982 VSS.n534 VSS.t2525 60.5809
R3983 VSS.n561 VSS.t2000 60.5809
R3984 VSS.n5386 VSS.t3292 60.5809
R3985 VSS.n2049 VSS.t989 60.5809
R3986 VSS.n2149 VSS.t2530 60.5809
R3987 VSS.n2642 VSS.t262 60.5809
R3988 VSS.n2645 VSS.t157 60.5809
R3989 VSS.n2838 VSS.t2170 60.5809
R3990 VSS.n2845 VSS.t1062 60.5809
R3991 VSS.n2914 VSS.t1393 60.5809
R3992 VSS.n2930 VSS.t1993 60.5809
R3993 VSS.n3326 VSS.t2621 60.5809
R3994 VSS.n3128 VSS.t2296 60.5809
R3995 VSS.n3170 VSS.t807 60.5809
R3996 VSS.n3236 VSS.t1316 60.5809
R3997 VSS.n1397 VSS.t289 60.5809
R3998 VSS.n1065 VSS.t352 60.5809
R3999 VSS.n1014 VSS.t3269 60.5809
R4000 VSS.n995 VSS.t2227 60.5809
R4001 VSS.n3680 VSS.t2557 60.5809
R4002 VSS.n4191 VSS.n3912 59.4829
R4003 VSS.n4191 VSS.n4190 59.4829
R4004 VSS.n4190 VSS.n3918 59.4829
R4005 VSS.n4181 VSS.n3918 59.4829
R4006 VSS.n4181 VSS.n4180 59.4829
R4007 VSS.n4180 VSS.n3930 59.4829
R4008 VSS.n4233 VSS.n4221 59.4829
R4009 VSS.n4234 VSS.n4233 59.4829
R4010 VSS.n3102 VSS.t1321 59.0774
R4011 VSS.t3594 VSS.t395 59.0043
R4012 VSS.t148 VSS.t2443 59.0043
R4013 VSS.t1469 VSS.t2669 59.0043
R4014 VSS.t3679 VSS.t2566 59.0043
R4015 VSS.t3492 VSS.t573 59.0043
R4016 VSS.t10 VSS.n2634 59.0043
R4017 VSS.t3677 VSS.t1960 59.0043
R4018 VSS.t1225 VSS.t3434 59.0043
R4019 VSS.t154 VSS.t2638 58.9109
R4020 VSS.n320 VSS.n318 58.8805
R4021 VSS.n260 VSS.t1332 58.5719
R4022 VSS.n352 VSS.t2891 58.5719
R4023 VSS.n545 VSS.t758 58.5719
R4024 VSS.n2105 VSS.t2713 58.5719
R4025 VSS.n2344 VSS.t3093 58.5719
R4026 VSS.n2410 VSS.t1579 58.5719
R4027 VSS.n1259 VSS.t3381 58.5719
R4028 VSS.n1198 VSS.t3643 58.5719
R4029 VSS.n1152 VSS.t1691 58.5719
R4030 VSS.n1375 VSS.t1765 58.5719
R4031 VSS.n1508 VSS.t3056 58.5719
R4032 VSS.n1518 VSS.t3547 58.5719
R4033 VSS.n1027 VSS.t71 58.5719
R4034 VSS.n1038 VSS.t2897 58.5719
R4035 VSS.n3702 VSS.t1751 58.5719
R4036 VSS.n2955 VSS.t329 57.875
R4037 VSS.n3150 VSS.t81 57.875
R4038 VSS.n3223 VSS.t3543 57.875
R4039 VSS.n3593 VSS.t1753 57.875
R4040 VSS.n3625 VSS.t1577 57.875
R4041 VSS.n3653 VSS.t3065 57.875
R4042 VSS.n4584 VSS.t3376 57.875
R4043 VSS.t741 VSS.t255 56.8795
R4044 VSS.n4880 VSS.t3697 56.7747
R4045 VSS.n4880 VSS.t3699 56.7747
R4046 VSS.n4873 VSS.t2927 56.7747
R4047 VSS.n4873 VSS.t2922 56.7747
R4048 VSS.n4867 VSS.t3701 56.7747
R4049 VSS.n4867 VSS.t3703 56.7747
R4050 VSS.n3102 VSS.t229 56.3082
R4051 VSS.n38 VSS.t240 55.7148
R4052 VSS.n98 VSS.t2060 55.7148
R4053 VSS.n111 VSS.t1858 55.7148
R4054 VSS.n132 VSS.t2143 55.7148
R4055 VSS.n149 VSS.t1146 55.7148
R4056 VSS.n158 VSS.t552 55.7148
R4057 VSS.n173 VSS.t1012 55.7148
R4058 VSS.n192 VSS.t281 55.7148
R4059 VSS.n246 VSS.t1863 55.7148
R4060 VSS.n250 VSS.t1910 55.7148
R4061 VSS.n531 VSS.t1969 55.7148
R4062 VSS.n2517 VSS.t3607 55.7148
R4063 VSS.n1961 VSS.t489 55.7148
R4064 VSS.n2568 VSS.t1107 55.7148
R4065 VSS.n2605 VSS.t3609 55.7148
R4066 VSS.n3790 VSS.t1040 55.7148
R4067 VSS.t2836 VSS.n4143 54.5685
R4068 VSS.n4840 VSS.t2852 54.5685
R4069 VSS.n3894 VSS.t63 53.7941
R4070 VSS.n364 VSS.t1922 52.8576
R4071 VSS.n395 VSS.t992 52.8576
R4072 VSS.n426 VSS.t655 52.8576
R4073 VSS.n458 VSS.t769 52.8576
R4074 VSS.n2399 VSS.t782 52.8576
R4075 VSS.n2404 VSS.t912 52.8576
R4076 VSS.n1973 VSS.t1118 52.8576
R4077 VSS.n2763 VSS.t3461 52.8576
R4078 VSS.n2779 VSS.t514 52.8576
R4079 VSS.n1205 VSS.t501 52.8576
R4080 VSS.n1098 VSS.t2234 52.8576
R4081 VSS.n1019 VSS.t3597 52.8576
R4082 VSS.n4671 VSS.t2248 52.8576
R4083 VSS.n4884 VSS.n4883 52.0324
R4084 VSS.n4128 VSS.n3948 52.0324
R4085 VSS.n4176 VSS.n4175 51.7539
R4086 VSS.n1040 VSS.t44 51.6928
R4087 VSS.n35 VSS.t3579 51.4291
R4088 VSS.n32 VSS.t1848 51.4291
R4089 VSS.n222 VSS.t2748 51.4291
R4090 VSS.n254 VSS.t1197 51.4291
R4091 VSS.n283 VSS.t1081 51.4291
R4092 VSS.n4920 VSS.t3634 51.4291
R4093 VSS.n303 VSS.t2577 51.4291
R4094 VSS.n287 VSS.t1726 51.4291
R4095 VSS.n288 VSS.t3571 51.4291
R4096 VSS.n312 VSS.t1824 51.4291
R4097 VSS.n315 VSS.t1749 51.4291
R4098 VSS.n516 VSS.t1633 51.4291
R4099 VSS.n5394 VSS.t1739 51.4291
R4100 VSS.n5397 VSS.t2617 51.4291
R4101 VSS.n5398 VSS.t2615 51.4291
R4102 VSS.n5401 VSS.t1792 51.4291
R4103 VSS.n5402 VSS.t2502 51.4291
R4104 VSS.n2059 VSS.t1718 51.4291
R4105 VSS.n2063 VSS.t1840 51.4291
R4106 VSS.n2064 VSS.t975 51.4291
R4107 VSS.n2056 VSS.t3585 51.4291
R4108 VSS.n2409 VSS.t775 51.4291
R4109 VSS.n2653 VSS.t2833 51.4291
R4110 VSS.n2656 VSS.t3640 51.4291
R4111 VSS.n2657 VSS.t1543 51.4291
R4112 VSS.n3031 VSS.t1574 51.4291
R4113 VSS.n3035 VSS.t2725 51.4291
R4114 VSS.n3036 VSS.t1785 51.4291
R4115 VSS.n2814 VSS.t2821 51.4291
R4116 VSS.n2815 VSS.t1733 51.4291
R4117 VSS.n2804 VSS.t1737 51.4291
R4118 VSS.n2865 VSS.t2485 51.4291
R4119 VSS.n2756 VSS.t503 51.4291
R4120 VSS.n2937 VSS.t1631 51.4291
R4121 VSS.n3027 VSS.t1781 51.4291
R4122 VSS.n3028 VSS.t1232 51.4291
R4123 VSS.n3024 VSS.t1794 51.4291
R4124 VSS.n3067 VSS.t2316 51.4291
R4125 VSS.n3021 VSS.t1783 51.4291
R4126 VSS.n3073 VSS.t2605 51.4291
R4127 VSS.n3110 VSS.t2428 51.4291
R4128 VSS.n1185 VSS.t205 51.4291
R4129 VSS.n1357 VSS.t260 51.4291
R4130 VSS.n1148 VSS.t3654 51.4291
R4131 VSS.n1034 VSS.t1166 51.4291
R4132 VSS.n1045 VSS.t1712 51.4291
R4133 VSS.n1643 VSS.t3593 51.4291
R4134 VSS.n998 VSS.t1334 51.4291
R4135 VSS.n1710 VSS.t3040 51.4291
R4136 VSS.n1711 VSS.t174 51.4291
R4137 VSS.n977 VSS.t1797 51.4291
R4138 VSS.n961 VSS.t2877 51.4291
R4139 VSS.n962 VSS.t1666 51.4291
R4140 VSS.n1273 VSS.t1773 51.4291
R4141 VSS.n1274 VSS.t3421 51.4291
R4142 VSS.n1276 VSS.t3624 51.4291
R4143 VSS.n1277 VSS.t973 51.4291
R4144 VSS.n3596 VSS.t1508 51.4291
R4145 VSS.n3607 VSS.t2501 51.4291
R4146 VSS.n3621 VSS.t2338 51.4291
R4147 VSS.n3635 VSS.t2517 51.4291
R4148 VSS.n3648 VSS.t265 51.4291
R4149 VSS.n3664 VSS.t2507 51.4291
R4150 VSS.n3688 VSS.t367 51.4291
R4151 VSS.n3704 VSS.t1914 51.4291
R4152 VSS.n3707 VSS.t3489 51.4291
R4153 VSS.n3744 VSS.t3660 51.4291
R4154 VSS.n3756 VSS.t1831 51.4291
R4155 VSS.n4592 VSS.t1154 51.4291
R4156 VSS.n3565 VSS.t97 51.4291
R4157 VSS.n3562 VSS.t505 51.4291
R4158 VSS.n4632 VSS.t3473 51.4291
R4159 VSS.n4649 VSS.t1949 51.4291
R4160 VSS.n4668 VSS.t2308 51.4291
R4161 VSS.n4674 VSS.t46 51.4291
R4162 VSS.n4677 VSS.t2835 51.4291
R4163 VSS.n4680 VSS.t2521 51.4291
R4164 VSS.n4683 VSS.t3577 51.4291
R4165 VSS.t3477 VSS.n4034 51.3
R4166 VSS.n4041 VSS.t3568 51.3
R4167 VSS.t3560 VSS.n4041 51.3
R4168 VSS.n4145 VSS.t3481 51.3
R4169 VSS.n4145 VSS.t3479 51.3
R4170 VSS.n4281 VSS.t741 50.7854
R4171 VSS.t1515 VSS.t3175 50.5752
R4172 VSS.t425 VSS.t815 50.5752
R4173 VSS.t1641 VSS.t330 50.5752
R4174 VSS.t2332 VSS.t617 50.5752
R4175 VSS.t1894 VSS.t596 50.5752
R4176 VSS.t1770 VSS.t1286 50.5752
R4177 VSS.t210 VSS.t2542 50.5752
R4178 VSS.n4157 VSS.t1808 50.3389
R4179 VSS.n4017 VSS.n3969 50.1178
R4180 VSS.n4159 VSS.t1806 49.813
R4181 VSS.n4732 VSS.n1919 49.7947
R4182 VSS.n4283 VSS.n3907 49.6897
R4183 VSS.n3891 VSS.t60 49.2941
R4184 VSS.n4034 VSS.n4033 49.1625
R4185 VSS.n4185 VSS.n4184 48.7505
R4186 VSS.n4184 VSS.n4183 48.7505
R4187 VSS.n3915 VSS.n3914 48.7505
R4188 VSS.n4183 VSS.n3915 48.7505
R4189 VSS.t2065 VSS.t2061 48.5195
R4190 VSS.t2063 VSS.t2065 48.5195
R4191 VSS.t2067 VSS.t2063 48.5195
R4192 VSS.n1116 VSS.t42 48.2862
R4193 VSS.n1108 VSS.t460 48.2862
R4194 VSS.n3885 VSS.t1931 47.2331
R4195 VSS.n3884 VSS.t1929 47.2331
R4196 VSS.n3883 VSS.t1936 47.2331
R4197 VSS.t1237 VSS.t2634 46.7226
R4198 VSS.n4197 VSS.n3914 46.6799
R4199 VSS.n3103 VSS.n3102 46.2505
R4200 VSS.n4286 VSS.n3904 46.1526
R4201 VSS.n4198 VSS.n3913 45.7304
R4202 VSS.n275 VSS.t1629 45.7148
R4203 VSS.n4960 VSS.t1741 45.7148
R4204 VSS.n4968 VSS.t2411 45.7148
R4205 VSS.n543 VSS.t258 45.7148
R4206 VSS.n597 VSS.t211 45.7148
R4207 VSS.n604 VSS.t2571 45.7148
R4208 VSS.n2389 VSS.t1722 45.7148
R4209 VSS.n2382 VSS.t1090 45.7148
R4210 VSS.n2374 VSS.t93 45.7148
R4211 VSS.n2128 VSS.t2418 45.7148
R4212 VSS.n2151 VSS.t1130 45.7148
R4213 VSS.n2996 VSS.t2272 45.7148
R4214 VSS.n994 VSS.t2177 45.7148
R4215 VSS.n4294 VSS.n3880 43.6225
R4216 VSS.n210 VSS.t2976 43.3851
R4217 VSS.n3893 VSS.n3892 43.373
R4218 VSS.n3881 VSS.t1927 42.9573
R4219 VSS.n3882 VSS.t1934 42.8802
R4220 VSS.n3882 VSS.t1933 42.7331
R4221 VSS.n3881 VSS.t1926 42.6862
R4222 VSS.t250 VSS.t2632 42.6598
R4223 VSS.t2432 VSS.n3995 42.2975
R4224 VSS.t2716 VSS.t1087 42.1461
R4225 VSS.t1187 VSS.t247 42.1461
R4226 VSS.t1793 VSS.t2550 42.1461
R4227 VSS.t2315 VSS.t764 42.1461
R4228 VSS.t2531 VSS.t2806 42.1461
R4229 VSS.t2766 VSS.t1487 42.1461
R4230 VSS.t2251 VSS.t1878 42.1461
R4231 VSS.t3050 VSS.t3638 42.1461
R4232 VSS.t102 VSS.t2894 42.1461
R4233 VSS.t1093 VSS.t1432 42.1461
R4234 VSS.t2998 VSS.t3487 42.1461
R4235 VSS.t1558 VSS.t3313 42.1461
R4236 VSS.n4286 VSS.n4285 42.0061
R4237 VSS.n4038 VSS.n3955 41.7862
R4238 VSS.n4038 VSS.n4037 41.7862
R4239 VSS.n4042 VSS.n3947 41.7862
R4240 VSS.n4048 VSS.n3950 41.7862
R4241 VSS.n4144 VSS.n3950 41.7862
R4242 VSS.n4026 VSS.n4025 41.7862
R4243 VSS.n4025 VSS.n3957 41.7862
R4244 VSS.n4878 VSS.n4877 41.7862
R4245 VSS.n4879 VSS.n4878 41.7862
R4246 VSS.n1744 VSS.n1741 41.7862
R4247 VSS.n1745 VSS.n1744 41.7862
R4248 VSS.n1746 VSS.n1743 41.7862
R4249 VSS.n4866 VSS.n1743 41.7862
R4250 VSS.n1732 VSS.n1730 41.7862
R4251 VSS.n4838 VSS.n1732 41.7862
R4252 VSS.n405 VSS.t1595 41.539
R4253 VSS.n406 VSS.t2333 41.539
R4254 VSS.n347 VSS.t691 41.539
R4255 VSS.n348 VSS.t1211 41.539
R4256 VSS.n2491 VSS.t1306 41.539
R4257 VSS.n2490 VSS.t53 41.539
R4258 VSS.n2423 VSS.t1587 41.539
R4259 VSS.n2422 VSS.t559 41.539
R4260 VSS.n3524 VSS.t3439 41.539
R4261 VSS.n3523 VSS.t7 41.539
R4262 VSS.n2882 VSS.t2394 41.539
R4263 VSS.n2881 VSS.t2396 41.539
R4264 VSS.n3184 VSS.t1242 41.539
R4265 VSS.n3185 VSS.t386 41.539
R4266 VSS.n3083 VSS.t2314 41.539
R4267 VSS.n3084 VSS.t531 41.539
R4268 VSS.n1160 VSS.t1589 41.539
R4269 VSS.n1161 VSS.t3420 41.539
R4270 VSS.t1171 VSS.t2834 41.3928
R4271 VSS.n4893 VSS.n4892 40.9835
R4272 VSS.t1842 VSS.t1819 40.6211
R4273 VSS.n2553 VSS.t151 40.6159
R4274 VSS.n2554 VSS.t2120 40.6159
R4275 VSS.n2459 VSS.t574 40.6159
R4276 VSS.n2458 VSS.t3423 40.6159
R4277 VSS.n2312 VSS.t465 40.6159
R4278 VSS.n2311 VSS.t1102 40.6159
R4279 VSS.n52 VSS.t242 40.0005
R4280 VSS.n52 VSS.t244 40.0005
R4281 VSS.n38 VSS.t2392 40.0005
R4282 VSS.n98 VSS.t3433 40.0005
R4283 VSS.n100 VSS.t2054 40.0005
R4284 VSS.n100 VSS.t2058 40.0005
R4285 VSS.n111 VSS.t2104 40.0005
R4286 VSS.n114 VSS.t1856 40.0005
R4287 VSS.n114 VSS.t1854 40.0005
R4288 VSS.n132 VSS.t1410 40.0005
R4289 VSS.n135 VSS.t2147 40.0005
R4290 VSS.n135 VSS.t2145 40.0005
R4291 VSS.n148 VSS.t1142 40.0005
R4292 VSS.n148 VSS.t1144 40.0005
R4293 VSS.n149 VSS.t2752 40.0005
R4294 VSS.n158 VSS.t1987 40.0005
R4295 VSS.n161 VSS.t556 40.0005
R4296 VSS.n161 VSS.t550 40.0005
R4297 VSS.n173 VSS.t1939 40.0005
R4298 VSS.n175 VSS.t1014 40.0005
R4299 VSS.n175 VSS.t1018 40.0005
R4300 VSS.n192 VSS.t2270 40.0005
R4301 VSS.n193 VSS.t279 40.0005
R4302 VSS.n193 VSS.t285 40.0005
R4303 VSS.n243 VSS.t1867 40.0005
R4304 VSS.n243 VSS.t1869 40.0005
R4305 VSS.n246 VSS.t1619 40.0005
R4306 VSS.n249 VSS.t1912 40.0005
R4307 VSS.n249 VSS.t1906 40.0005
R4308 VSS.n250 VSS.t1383 40.0005
R4309 VSS.n364 VSS.t2015 40.0005
R4310 VSS.n372 VSS.t884 40.0005
R4311 VSS.n372 VSS.t872 40.0005
R4312 VSS.n373 VSS.t882 40.0005
R4313 VSS.n373 VSS.t890 40.0005
R4314 VSS.n377 VSS.t898 40.0005
R4315 VSS.n377 VSS.t888 40.0005
R4316 VSS.n378 VSS.t886 40.0005
R4317 VSS.n381 VSS.t874 40.0005
R4318 VSS.n381 VSS.t902 40.0005
R4319 VSS.n385 VSS.t896 40.0005
R4320 VSS.n385 VSS.t892 40.0005
R4321 VSS.n390 VSS.t900 40.0005
R4322 VSS.n390 VSS.t3015 40.0005
R4323 VSS.n387 VSS.t876 40.0005
R4324 VSS.n387 VSS.t880 40.0005
R4325 VSS.n394 VSS.t3021 40.0005
R4326 VSS.n394 VSS.t2997 40.0005
R4327 VSS.n395 VSS.t1745 40.0005
R4328 VSS.n426 VSS.t1743 40.0005
R4329 VSS.n458 VSS.t1635 40.0005
R4330 VSS.n531 VSS.t3090 40.0005
R4331 VSS.n535 VSS.t1971 40.0005
R4332 VSS.n535 VSS.t1973 40.0005
R4333 VSS.n2037 VSS.t432 40.0005
R4334 VSS.n2037 VSS.t426 40.0005
R4335 VSS.n2214 VSS.t422 40.0005
R4336 VSS.n2214 VSS.t434 40.0005
R4337 VSS.n2034 VSS.t440 40.0005
R4338 VSS.n2034 VSS.t424 40.0005
R4339 VSS.n2221 VSS.t416 40.0005
R4340 VSS.n2031 VSS.t436 40.0005
R4341 VSS.n2031 VSS.t438 40.0005
R4342 VSS.n2228 VSS.t420 40.0005
R4343 VSS.n2228 VSS.t444 40.0005
R4344 VSS.n2027 VSS.t418 40.0005
R4345 VSS.n2027 VSS.t414 40.0005
R4346 VSS.n2024 VSS.t428 40.0005
R4347 VSS.n2024 VSS.t3009 40.0005
R4348 VSS.n2023 VSS.t3019 40.0005
R4349 VSS.n2023 VSS.t3011 40.0005
R4350 VSS.n2413 VSS.t825 40.0005
R4351 VSS.n2413 VSS.t843 40.0005
R4352 VSS.n2416 VSS.t839 40.0005
R4353 VSS.n2416 VSS.t849 40.0005
R4354 VSS.n2417 VSS.t821 40.0005
R4355 VSS.n2417 VSS.t831 40.0005
R4356 VSS.n1993 VSS.t823 40.0005
R4357 VSS.n1990 VSS.t835 40.0005
R4358 VSS.n1990 VSS.t851 40.0005
R4359 VSS.n1989 VSS.t845 40.0005
R4360 VSS.n1989 VSS.t841 40.0005
R4361 VSS.n2485 VSS.t837 40.0005
R4362 VSS.n2485 VSS.t827 40.0005
R4363 VSS.n2488 VSS.t833 40.0005
R4364 VSS.n2488 VSS.t3013 40.0005
R4365 VSS.n2497 VSS.t3003 40.0005
R4366 VSS.n2497 VSS.t3001 40.0005
R4367 VSS.n1973 VSS.t2487 40.0005
R4368 VSS.n1961 VSS.t1724 40.0005
R4369 VSS.n2570 VSS.t491 40.0005
R4370 VSS.n2570 VSS.t493 40.0005
R4371 VSS.n1954 VSS.t2996 40.0005
R4372 VSS.n1954 VSS.t2994 40.0005
R4373 VSS.n2584 VSS.t2999 40.0005
R4374 VSS.n2584 VSS.t21 40.0005
R4375 VSS.n2587 VSS.t15 40.0005
R4376 VSS.n2587 VSS.t39 40.0005
R4377 VSS.n1951 VSS.t11 40.0005
R4378 VSS.n1951 VSS.t17 40.0005
R4379 VSS.n2593 VSS.t19 40.0005
R4380 VSS.n2593 VSS.t33 40.0005
R4381 VSS.n2597 VSS.t9 40.0005
R4382 VSS.n2598 VSS.t13 40.0005
R4383 VSS.n2598 VSS.t25 40.0005
R4384 VSS.n2600 VSS.t29 40.0005
R4385 VSS.n2600 VSS.t31 40.0005
R4386 VSS.n2604 VSS.t37 40.0005
R4387 VSS.n2604 VSS.t23 40.0005
R4388 VSS.n1125 VSS.t324 40.0005
R4389 VSS.n1125 VSS.t312 40.0005
R4390 VSS.n1205 VSS.t248 40.0005
R4391 VSS.n1483 VSS.t305 40.0005
R4392 VSS.n1483 VSS.t301 40.0005
R4393 VSS.n1490 VSS.t316 40.0005
R4394 VSS.n1490 VSS.t303 40.0005
R4395 VSS.n1119 VSS.t320 40.0005
R4396 VSS.n1098 VSS.t2873 40.0005
R4397 VSS.n1496 VSS.t299 40.0005
R4398 VSS.n1496 VSS.t307 40.0005
R4399 VSS.n1558 VSS.t318 40.0005
R4400 VSS.n1558 VSS.t295 40.0005
R4401 VSS.n1500 VSS.t314 40.0005
R4402 VSS.n1500 VSS.t311 40.0005
R4403 VSS.n1501 VSS.t3629 40.0005
R4404 VSS.n1501 VSS.t322 40.0005
R4405 VSS.n1504 VSS.t3631 40.0005
R4406 VSS.n1504 VSS.t3627 40.0005
R4407 VSS.n3790 VSS.t2327 40.0005
R4408 VSS.n3791 VSS.t1034 40.0005
R4409 VSS.n3791 VSS.t1036 40.0005
R4410 VSS.n4671 VSS.t1707 40.0005
R4411 VSS.n1040 VSS.t57 39.6928
R4412 VSS.n1856 VSS.t2068 39.6928
R4413 VSS.n4740 VSS.t1345 39.6928
R4414 VSS.n4741 VSS.t2109 39.6928
R4415 VSS.n4753 VSS.t2273 39.6928
R4416 VSS.n4754 VSS.t1182 39.6928
R4417 VSS.n4089 VSS.t2300 39.6928
R4418 VSS.n4093 VSS.t1498 39.6928
R4419 VSS.n4774 VSS.t164 39.6928
R4420 VSS.n4775 VSS.t599 39.6928
R4421 VSS.n4769 VSS.t1362 39.6928
R4422 VSS.n4770 VSS.t192 39.6928
R4423 VSS.n4238 VSS.t564 39.2687
R4424 VSS.n3967 VSS.n3964 39.0005
R4425 VSS.n4022 VSS.n3962 39.0005
R4426 VSS.n3962 VSS.n3960 39.0005
R4427 VSS.n4864 VSS.n4863 39.0005
R4428 VSS.n4865 VSS.n4864 39.0005
R4429 VSS.n1757 VSS.n1752 39.0005
R4430 VSS.n1757 VSS.n1756 39.0005
R4431 VSS.n1755 VSS.n1753 39.0005
R4432 VSS.n4298 VSS.n4297 39.0005
R4433 VSS.t1928 VSS.n4298 39.0005
R4434 VSS.n3879 VSS.n3876 39.0005
R4435 VSS.t1928 VSS.n3876 39.0005
R4436 VSS.n3966 VSS.n3965 39.0005
R4437 VSS.n3995 VSS.n3966 39.0005
R4438 VSS.n359 VSS.t3453 38.7697
R4439 VSS.n556 VSS.t2221 38.7697
R4440 VSS.n2028 VSS.t1190 38.7697
R4441 VSS.n1995 VSS.t121 38.7697
R4442 VSS.n2606 VSS.t789 38.7697
R4443 VSS.n2894 VSS.t1223 38.7697
R4444 VSS.n2929 VSS.t2496 38.7697
R4445 VSS.n3099 VSS.t1109 38.7697
R4446 VSS.n3099 VSS.t3662 38.7697
R4447 VSS.n3207 VSS.t641 38.7697
R4448 VSS.n3227 VSS.t2323 38.7697
R4449 VSS.n1188 VSS.t3441 38.7697
R4450 VSS.n1166 VSS.t512 38.7697
R4451 VSS.n1163 VSS.t378 38.7697
R4452 VSS.n1378 VSS.t170 38.7697
R4453 VSS.n1133 VSS.t773 38.7697
R4454 VSS.n1131 VSS.t2348 38.7697
R4455 VSS.n1128 VSS.t343 38.7697
R4456 VSS.n1511 VSS.t1367 38.7697
R4457 VSS.n1605 VSS.t2042 38.7697
R4458 VSS.n1611 VSS.t2589 38.7697
R4459 VSS.n1856 VSS.t1820 38.7697
R4460 VSS.n4740 VSS.t2680 38.7697
R4461 VSS.n4741 VSS.t2874 38.7697
R4462 VSS.n4753 VSS.t3023 38.7697
R4463 VSS.n4754 VSS.t3696 38.7697
R4464 VSS.n4089 VSS.t2724 38.7697
R4465 VSS.n4093 VSS.t3688 38.7697
R4466 VSS.n4774 VSS.t2858 38.7697
R4467 VSS.n4775 VSS.t1720 38.7697
R4468 VSS.n4769 VSS.t3529 38.7697
R4469 VSS.n4770 VSS.t3522 38.7697
R4470 VSS.n5254 VSS.t1763 38.5719
R4471 VSS.n5285 VSS.t2363 38.5719
R4472 VSS.n5302 VSS.t1687 38.5719
R4473 VSS.n5360 VSS.t1698 38.5719
R4474 VSS.n227 VSS.t1510 38.5719
R4475 VSS.n227 VSS.t2951 38.5719
R4476 VSS.n18 VSS.t1954 38.5719
R4477 VSS.n18 VSS.t3674 38.5719
R4478 VSS.n566 VSS.t1219 38.5719
R4479 VSS.n701 VSS.t944 38.5719
R4480 VSS.n753 VSS.t2455 38.5719
R4481 VSS.n922 VSS.t1810 38.5719
R4482 VSS.n335 VSS.t1002 38.5719
R4483 VSS.n335 VSS.t2963 38.5719
R4484 VSS.n353 VSS.t2211 38.5719
R4485 VSS.n353 VSS.t2947 38.5719
R4486 VSS.n378 VSS.t894 38.5719
R4487 VSS.n423 VSS.t1414 38.5719
R4488 VSS.n423 VSS.t2953 38.5719
R4489 VSS.n443 VSS.t457 38.5719
R4490 VSS.n443 VSS.t2961 38.5719
R4491 VSS.n447 VSS.t2959 38.5719
R4492 VSS.n447 VSS.t527 38.5719
R4493 VSS.n487 VSS.t904 38.5719
R4494 VSS.n487 VSS.t2911 38.5719
R4495 VSS.n517 VSS.t2217 38.5719
R4496 VSS.n517 VSS.t2876 38.5719
R4497 VSS.n540 VSS.t2543 38.5719
R4498 VSS.n540 VSS.t3668 38.5719
R4499 VSS.n5395 VSS.t1376 38.5719
R4500 VSS.n5395 VSS.t3672 38.5719
R4501 VSS.n2717 VSS.t3583 38.5719
R4502 VSS.n2195 VSS.t2498 38.5719
R4503 VSS.n2196 VSS.t3039 38.5719
R4504 VSS.n2097 VSS.t2941 38.5719
R4505 VSS.n2097 VSS.t1440 38.5719
R4506 VSS.n2118 VSS.t1326 38.5719
R4507 VSS.n2118 VSS.t1924 38.5719
R4508 VSS.n2140 VSS.t2929 38.5719
R4509 VSS.n2140 VSS.t2407 38.5719
R4510 VSS.n2157 VSS.t2129 38.5719
R4511 VSS.n2157 VSS.t2017 38.5719
R4512 VSS.n2221 VSS.t430 38.5719
R4513 VSS.n2401 VSS.t1759 38.5719
R4514 VSS.n2401 VSS.t1714 38.5719
R4515 VSS.n2405 VSS.t2659 38.5719
R4516 VSS.n2405 VSS.t1058 38.5719
R4517 VSS.n2408 VSS.t3 38.5719
R4518 VSS.n2408 VSS.t2668 38.5719
R4519 VSS.n1993 VSS.t829 38.5719
R4520 VSS.n2597 VSS.t35 38.5719
R4521 VSS.n2649 VSS.t1389 38.5719
R4522 VSS.n2649 VSS.t3676 38.5719
R4523 VSS.n2652 VSS.t1120 38.5719
R4524 VSS.n2652 VSS.t3678 38.5719
R4525 VSS.n3473 VSS.t3468 38.5719
R4526 VSS.n2803 VSS.t2438 38.5719
R4527 VSS.n2803 VSS.t3680 38.5719
R4528 VSS.n2829 VSS.t1124 38.5719
R4529 VSS.n2829 VSS.t3670 38.5719
R4530 VSS.n2754 VSS.t2764 38.5719
R4531 VSS.n2754 VSS.t406 38.5719
R4532 VSS.n2764 VSS.t3617 38.5719
R4533 VSS.n2764 VSS.t791 38.5719
R4534 VSS.n2776 VSS.t793 38.5719
R4535 VSS.n2776 VSS.t2252 38.5719
R4536 VSS.n2905 VSS.t2185 38.5719
R4537 VSS.n2905 VSS.t2907 38.5719
R4538 VSS.n2924 VSS.t1466 38.5719
R4539 VSS.n2924 VSS.t2913 38.5719
R4540 VSS.n2965 VSS.t2945 38.5719
R4541 VSS.n2965 VSS.t2448 38.5719
R4542 VSS.n3243 VSS.t1459 38.5719
R4543 VSS.n3243 VSS.t2939 38.5719
R4544 VSS.n3130 VSS.t648 38.5719
R4545 VSS.n3130 VSS.t756 38.5719
R4546 VSS.n2993 VSS.t923 38.5719
R4547 VSS.n2993 VSS.t2933 38.5719
R4548 VSS.n2980 VSS.t1488 38.5719
R4549 VSS.n2980 VSS.t2935 38.5719
R4550 VSS.n1460 VSS.t2080 38.5719
R4551 VSS.n1184 VSS.t3645 38.5719
R4552 VSS.n1184 VSS.t2519 38.5719
R4553 VSS.n1153 VSS.t580 38.5719
R4554 VSS.n1153 VSS.t3383 38.5719
R4555 VSS.n1139 VSS.t2909 38.5719
R4556 VSS.n1139 VSS.t2492 38.5719
R4557 VSS.n1119 VSS.t309 38.5719
R4558 VSS.n1603 VSS.t1086 38.5719
R4559 VSS.n1116 VSS.t3545 38.5719
R4560 VSS.n1108 VSS.t79 38.5719
R4561 VSS.n1031 VSS.t3538 38.5719
R4562 VSS.n1031 VSS.t394 38.5719
R4563 VSS.n1037 VSS.t349 38.5719
R4564 VSS.n1037 VSS.t2949 38.5719
R4565 VSS.n1049 VSS.t2256 38.5719
R4566 VSS.n1049 VSS.t2593 38.5719
R4567 VSS.n1634 VSS.t666 38.5719
R4568 VSS.n1634 VSS.t2595 38.5719
R4569 VSS.n1641 VSS.t2087 38.5719
R4570 VSS.n1641 VSS.t2955 38.5719
R4571 VSS.n1648 VSS.t2116 38.5719
R4572 VSS.n1648 VSS.t67 38.5719
R4573 VSS.n1677 VSS.t2223 38.5719
R4574 VSS.n1677 VSS.t2957 38.5719
R4575 VSS.n1702 VSS.t3290 38.5719
R4576 VSS.n1702 VSS.t2175 38.5719
R4577 VSS.n3685 VSS.t2931 38.5719
R4578 VSS.n3685 VSS.t2258 38.5719
R4579 VSS.n4624 VSS.t2505 38.5719
R4580 VSS.n4624 VSS.t602 38.5719
R4581 VSS.n4855 VSS.n1760 38.4005
R4582 VSS.n4013 VSS.n3963 38.4005
R4583 VSS.t2196 VSS.t3138 37.2536
R4584 VSS.n2783 VSS.t2773 36.9236
R4585 VSS.n2777 VSS.t3044 36.9236
R4586 VSS.n3995 VSS.n3994 36.7321
R4587 VSS.t1423 VSS.n4300 36.7011
R4588 VSS.n3722 VSS.n3721 36.4703
R4589 VSS.n2350 VSS.t2889 36.0005
R4590 VSS.n2003 VSS.t952 36.0005
R4591 VSS.n2003 VSS.t1585 36.0005
R4592 VSS.n2396 VSS.t3493 36.0005
R4593 VSS.n2510 VSS.t2537 36.0005
R4594 VSS.n1957 VSS.t1996 36.0005
R4595 VSS.n2594 VSS.t475 36.0005
R4596 VSS.n1379 VSS.t2004 36.0005
R4597 VSS.n1122 VSS.t168 36.0005
R4598 VSS.n2783 VSS.t469 35.0774
R4599 VSS.n2777 VSS.t1876 35.0774
R4600 VSS.n806 VSS.n805 34.6358
R4601 VSS.n679 VSS.n494 34.6358
R4602 VSS.n2609 VSS.n2608 34.6358
R4603 VSS.n3287 VSS.n3286 34.6358
R4604 VSS.n1335 VSS.n1334 34.6358
R4605 VSS.n1339 VSS.n1338 34.6358
R4606 VSS.n1474 VSS.n1473 34.6358
R4607 VSS.n1478 VSS.n1477 34.6358
R4608 VSS.n1560 VSS.n1557 34.6358
R4609 VSS.n71 VSS.n70 34.6358
R4610 VSS.n5367 VSS.n94 34.6358
R4611 VSS.n5368 VSS.n5367 34.6358
R4612 VSS.n5369 VSS.n5368 34.6358
R4613 VSS.n5357 VSS.n96 34.6358
R4614 VSS.n5358 VSS.n5357 34.6358
R4615 VSS.n5306 VSS.n5305 34.6358
R4616 VSS.n5306 VSS.n120 34.6358
R4617 VSS.n5310 VSS.n120 34.6358
R4618 VSS.n5295 VSS.n123 34.6358
R4619 VSS.n5300 VSS.n123 34.6358
R4620 VSS.n5289 VSS.n5288 34.6358
R4621 VSS.n5289 VSS.n126 34.6358
R4622 VSS.n5293 VSS.n126 34.6358
R4623 VSS.n5283 VSS.n129 34.6358
R4624 VSS.n5258 VSS.n5257 34.6358
R4625 VSS.n5258 VSS.n141 34.6358
R4626 VSS.n5262 VSS.n141 34.6358
R4627 VSS.n5252 VSS.n144 34.6358
R4628 VSS.n5231 VSS.n5230 34.6358
R4629 VSS.n5232 VSS.n5231 34.6358
R4630 VSS.n5205 VSS.n164 34.6358
R4631 VSS.n5206 VSS.n5205 34.6358
R4632 VSS.n5207 VSS.n5206 34.6358
R4633 VSS.n5201 VSS.n5198 34.6358
R4634 VSS.n5168 VSS.n179 34.6358
R4635 VSS.n5161 VSS.n5160 34.6358
R4636 VSS.n5164 VSS.n5161 34.6358
R4637 VSS.n5139 VSS.n5138 34.6358
R4638 VSS.n5139 VSS.n187 34.6358
R4639 VSS.n5132 VSS.n190 34.6358
R4640 VSS.n5136 VSS.n190 34.6358
R4641 VSS.n5086 VSS.n5085 34.6358
R4642 VSS.n5092 VSS.n5091 34.6358
R4643 VSS.n5063 VSS.n225 34.6358
R4644 VSS.n5067 VSS.n225 34.6358
R4645 VSS.n5051 VSS.n5050 34.6358
R4646 VSS.n5051 VSS.n230 34.6358
R4647 VSS.n5055 VSS.n230 34.6358
R4648 VSS.n5056 VSS.n5055 34.6358
R4649 VSS.n5057 VSS.n5056 34.6358
R4650 VSS.n5043 VSS.n5042 34.6358
R4651 VSS.n5044 VSS.n5043 34.6358
R4652 VSS.n5044 VSS.n233 34.6358
R4653 VSS.n5048 VSS.n233 34.6358
R4654 VSS.n5038 VSS.n5037 34.6358
R4655 VSS.n5039 VSS.n5038 34.6358
R4656 VSS.n5013 VSS.n5012 34.6358
R4657 VSS.n5000 VSS.n4999 34.6358
R4658 VSS.n5000 VSS.n257 34.6358
R4659 VSS.n5004 VSS.n257 34.6358
R4660 VSS.n5005 VSS.n5004 34.6358
R4661 VSS.n5006 VSS.n5005 34.6358
R4662 VSS.n4997 VSS.n261 34.6358
R4663 VSS.n4967 VSS.n4966 34.6358
R4664 VSS.n4959 VSS.n4958 34.6358
R4665 VSS.n4962 VSS.n4959 34.6358
R4666 VSS.n4954 VSS.n4953 34.6358
R4667 VSS.n4955 VSS.n4954 34.6358
R4668 VSS.n4947 VSS.n281 34.6358
R4669 VSS.n4948 VSS.n4947 34.6358
R4670 VSS.n4949 VSS.n4948 34.6358
R4671 VSS.n4935 VSS.n4918 34.6358
R4672 VSS.n929 VSS.n928 34.6358
R4673 VSS.n921 VSS.n920 34.6358
R4674 VSS.n917 VSS.n916 34.6358
R4675 VSS.n914 VSS.n333 34.6358
R4676 VSS.n902 VSS.n341 34.6358
R4677 VSS.n898 VSS.n341 34.6358
R4678 VSS.n895 VSS.n894 34.6358
R4679 VSS.n889 VSS.n888 34.6358
R4680 VSS.n869 VSS.n360 34.6358
R4681 VSS.n841 VSS.n379 34.6358
R4682 VSS.n839 VSS.n838 34.6358
R4683 VSS.n818 VSS.n817 34.6358
R4684 VSS.n810 VSS.n410 34.6358
R4685 VSS.n805 VSS.n804 34.6358
R4686 VSS.n804 VSS.n416 34.6358
R4687 VSS.n800 VSS.n416 34.6358
R4688 VSS.n797 VSS.n420 34.6358
R4689 VSS.n793 VSS.n792 34.6358
R4690 VSS.n792 VSS.n791 34.6358
R4691 VSS.n777 VSS.n435 34.6358
R4692 VSS.n773 VSS.n772 34.6358
R4693 VSS.n772 VSS.n771 34.6358
R4694 VSS.n767 VSS.n766 34.6358
R4695 VSS.n751 VSS.n451 34.6358
R4696 VSS.n747 VSS.n451 34.6358
R4697 VSS.n709 VSS.n708 34.6358
R4698 VSS.n708 VSS.n707 34.6358
R4699 VSS.n698 VSS.n481 34.6358
R4700 VSS.n694 VSS.n481 34.6358
R4701 VSS.n692 VSS.n484 34.6358
R4702 VSS.n675 VSS.n494 34.6358
R4703 VSS.n669 VSS.n668 34.6358
R4704 VSS.n666 VSS.n502 34.6358
R4705 VSS.n658 VSS.n506 34.6358
R4706 VSS.n652 VSS.n651 34.6358
R4707 VSS.n651 VSS.n511 34.6358
R4708 VSS.n647 VSS.n511 34.6358
R4709 VSS.n626 VSS.n625 34.6358
R4710 VSS.n625 VSS.n624 34.6358
R4711 VSS.n621 VSS.n620 34.6358
R4712 VSS.n620 VSS.n619 34.6358
R4713 VSS.n612 VSS.n611 34.6358
R4714 VSS.n595 VSS.n541 34.6358
R4715 VSS.n591 VSS.n590 34.6358
R4716 VSS.n584 VSS.n583 34.6358
R4717 VSS.n580 VSS.n552 34.6358
R4718 VSS.n576 VSS.n575 34.6358
R4719 VSS.n572 VSS.n558 34.6358
R4720 VSS.n568 VSS.n558 34.6358
R4721 VSS.n5477 VSS.n9 34.6358
R4722 VSS.n5477 VSS.n5476 34.6358
R4723 VSS.n5448 VSS.n5447 34.6358
R4724 VSS.n5444 VSS.n5443 34.6358
R4725 VSS.n5443 VSS.n5442 34.6358
R4726 VSS.n2110 VSS.n2050 34.6358
R4727 VSS.n2111 VSS.n2110 34.6358
R4728 VSS.n2114 VSS.n2047 34.6358
R4729 VSS.n2123 VSS.n2120 34.6358
R4730 VSS.n2127 VSS.n2045 34.6358
R4731 VSS.n2202 VSS.n2135 34.6358
R4732 VSS.n2187 VSS.n2144 34.6358
R4733 VSS.n2182 VSS.n2181 34.6358
R4734 VSS.n2181 VSS.n2147 34.6358
R4735 VSS.n2169 VSS.n2168 34.6358
R4736 VSS.n2168 VSS.n2155 34.6358
R4737 VSS.n2162 VSS.n2161 34.6358
R4738 VSS.n2161 VSS.n2040 34.6358
R4739 VSS.n2227 VSS.n2226 34.6358
R4740 VSS.n2237 VSS.n2235 34.6358
R4741 VSS.n2255 VSS.n2018 34.6358
R4742 VSS.n2256 VSS.n2255 34.6358
R4743 VSS.n2260 VSS.n2256 34.6358
R4744 VSS.n2334 VSS.n2264 34.6358
R4745 VSS.n2308 VSS.n2272 34.6358
R4746 VSS.n2286 VSS.n2283 34.6358
R4747 VSS.n2283 VSS.n2015 34.6358
R4748 VSS.n2349 VSS.n2011 34.6358
R4749 VSS.n2352 VSS.n2009 34.6358
R4750 VSS.n2356 VSS.n2009 34.6358
R4751 VSS.n2357 VSS.n2356 34.6358
R4752 VSS.n2366 VSS.n2365 34.6358
R4753 VSS.n2380 VSS.n2001 34.6358
R4754 VSS.n2392 VSS.n2391 34.6358
R4755 VSS.n2471 VSS.n1997 34.6358
R4756 VSS.n2467 VSS.n1997 34.6358
R4757 VSS.n2479 VSS.n2478 34.6358
R4758 VSS.n2512 VSS.n1977 34.6358
R4759 VSS.n2516 VSS.n1977 34.6358
R4760 VSS.n2633 VSS.n1950 34.6358
R4761 VSS.n2630 VSS.n2629 34.6358
R4762 VSS.n2730 VSS.n2729 34.6358
R4763 VSS.n2729 VSS.n1939 34.6358
R4764 VSS.n2725 VSS.n2724 34.6358
R4765 VSS.n2724 VSS.n2723 34.6358
R4766 VSS.n2714 VSS.n1945 34.6358
R4767 VSS.n2701 VSS.n2700 34.6358
R4768 VSS.n2700 VSS.n2639 34.6358
R4769 VSS.n2696 VSS.n2639 34.6358
R4770 VSS.n2692 VSS.n2643 34.6358
R4771 VSS.n2688 VSS.n2643 34.6358
R4772 VSS.n2688 VSS.n2687 34.6358
R4773 VSS.n2685 VSS.n2646 34.6358
R4774 VSS.n2674 VSS.n2673 34.6358
R4775 VSS.n3050 VSS.n3049 34.6358
R4776 VSS.n2825 VSS.n2824 34.6358
R4777 VSS.n2837 VSS.n2836 34.6358
R4778 VSS.n2836 VSS.n2799 34.6358
R4779 VSS.n2844 VSS.n2797 34.6358
R4780 VSS.n2840 VSS.n2797 34.6358
R4781 VSS.n2848 VSS.n2847 34.6358
R4782 VSS.n2853 VSS.n2852 34.6358
R4783 VSS.n2852 VSS.n2793 34.6358
R4784 VSS.n2868 VSS.n2749 34.6358
R4785 VSS.n3514 VSS.n3513 34.6358
R4786 VSS.n3504 VSS.n3503 34.6358
R4787 VSS.n3492 VSS.n3491 34.6358
R4788 VSS.n3493 VSS.n3492 34.6358
R4789 VSS.n3493 VSS.n2771 34.6358
R4790 VSS.n3497 VSS.n2771 34.6358
R4791 VSS.n3498 VSS.n3497 34.6358
R4792 VSS.n3481 VSS.n2780 34.6358
R4793 VSS.n3485 VSS.n2780 34.6358
R4794 VSS.n3479 VSS.n2784 34.6358
R4795 VSS.n3465 VSS.n2786 34.6358
R4796 VSS.n3469 VSS.n2786 34.6358
R4797 VSS.n3470 VSS.n3469 34.6358
R4798 VSS.n3457 VSS.n2789 34.6358
R4799 VSS.n3461 VSS.n2789 34.6358
R4800 VSS.n3395 VSS.n2918 34.6358
R4801 VSS.n3399 VSS.n2918 34.6358
R4802 VSS.n3378 VSS.n2927 34.6358
R4803 VSS.n3379 VSS.n3378 34.6358
R4804 VSS.n3380 VSS.n3379 34.6358
R4805 VSS.n3367 VSS.n2931 34.6358
R4806 VSS.n3371 VSS.n2931 34.6358
R4807 VSS.n3348 VSS.n3346 34.6358
R4808 VSS.n3352 VSS.n2944 34.6358
R4809 VSS.n3339 VSS.n3338 34.6358
R4810 VSS.n3340 VSS.n3339 34.6358
R4811 VSS.n3333 VSS.n3332 34.6358
R4812 VSS.n3329 VSS.n3328 34.6358
R4813 VSS.n3088 VSS.n3016 34.6358
R4814 VSS.n3122 VSS.n3121 34.6358
R4815 VSS.n3123 VSS.n3122 34.6358
R4816 VSS.n3127 VSS.n3126 34.6358
R4817 VSS.n3135 VSS.n2999 34.6358
R4818 VSS.n3136 VSS.n3135 34.6358
R4819 VSS.n3137 VSS.n3136 34.6358
R4820 VSS.n3153 VSS.n3149 34.6358
R4821 VSS.n3157 VSS.n2990 34.6358
R4822 VSS.n3176 VSS.n2986 34.6358
R4823 VSS.n3177 VSS.n3176 34.6358
R4824 VSS.n3201 VSS.n2975 34.6358
R4825 VSS.n3213 VSS.n3212 34.6358
R4826 VSS.n3214 VSS.n3213 34.6358
R4827 VSS.n3281 VSS.n3280 34.6358
R4828 VSS.n3274 VSS.n3273 34.6358
R4829 VSS.n3273 VSS.n3272 34.6358
R4830 VSS.n3269 VSS.n3268 34.6358
R4831 VSS.n1319 VSS.n1318 34.6358
R4832 VSS.n1326 VSS.n1177 34.6358
R4833 VSS.n1322 VSS.n1177 34.6358
R4834 VSS.n1250 VSS.n1249 34.6358
R4835 VSS.n1334 VSS.n1333 34.6358
R4836 VSS.n1333 VSS.n1171 34.6358
R4837 VSS.n1352 VSS.n1351 34.6358
R4838 VSS.n1363 VSS.n1150 34.6358
R4839 VSS.n1364 VSS.n1363 34.6358
R4840 VSS.n1438 VSS.n1437 34.6358
R4841 VSS.n1434 VSS.n1380 34.6358
R4842 VSS.n1430 VSS.n1429 34.6358
R4843 VSS.n1430 VSS.n1380 34.6358
R4844 VSS.n1423 VSS.n1422 34.6358
R4845 VSS.n1409 VSS.n1408 34.6358
R4846 VSS.n1410 VSS.n1409 34.6358
R4847 VSS.n1405 VSS.n1404 34.6358
R4848 VSS.n1399 VSS.n1144 34.6358
R4849 VSS.n1467 VSS.n1466 34.6358
R4850 VSS.n1466 VSS.n1136 34.6358
R4851 VSS.n1462 VSS.n1136 34.6358
R4852 VSS.n1473 VSS.n1472 34.6358
R4853 VSS.n1486 VSS.n1485 34.6358
R4854 VSS.n1564 VSS.n1497 34.6358
R4855 VSS.n1545 VSS.n1543 34.6358
R4856 VSS.n1537 VSS.n1509 34.6358
R4857 VSS.n1541 VSS.n1509 34.6358
R4858 VSS.n1531 VSS.n1530 34.6358
R4859 VSS.n1528 VSS.n1516 34.6358
R4860 VSS.n1523 VSS.n1522 34.6358
R4861 VSS.n1587 VSS.n1586 34.6358
R4862 VSS.n1596 VSS.n1595 34.6358
R4863 VSS.n1610 VSS.n1101 34.6358
R4864 VSS.n1618 VSS.n1617 34.6358
R4865 VSS.n1617 VSS.n1099 34.6358
R4866 VSS.n1095 VSS.n1093 34.6358
R4867 VSS.n1093 VSS.n1092 34.6358
R4868 VSS.n1084 VSS.n1035 34.6358
R4869 VSS.n1071 VSS.n1043 34.6358
R4870 VSS.n1072 VSS.n1071 34.6358
R4871 VSS.n1073 VSS.n1072 34.6358
R4872 VSS.n1056 VSS.n1050 34.6358
R4873 VSS.n1651 VSS.n1650 34.6358
R4874 VSS.n1665 VSS.n1664 34.6358
R4875 VSS.n1664 VSS.n1663 34.6358
R4876 VSS.n1663 VSS.n1012 34.6358
R4877 VSS.n1659 VSS.n1012 34.6358
R4878 VSS.n1684 VSS.n1683 34.6358
R4879 VSS.n1700 VSS.n992 34.6358
R4880 VSS.n1696 VSS.n992 34.6358
R4881 VSS.n1696 VSS.n1695 34.6358
R4882 VSS.n4005 VSS.n4001 34.6358
R4883 VSS.n4009 VSS.n4001 34.6358
R4884 VSS.n1827 VSS.n1826 34.6358
R4885 VSS.n4752 VSS.n4738 34.6358
R4886 VSS.n1901 VSS.n1900 34.6358
R4887 VSS.n1911 VSS.n1889 34.6358
R4888 VSS.n1914 VSS.n1913 34.6358
R4889 VSS.n4064 VSS.n4063 34.6358
R4890 VSS.n4074 VSS.n4055 34.6358
R4891 VSS.n4079 VSS.n4076 34.6358
R4892 VSS.n4101 VSS.n4090 34.6358
R4893 VSS.n1805 VSS.n1804 34.6358
R4894 VSS.n1809 VSS.n1808 34.6358
R4895 VSS.n1796 VSS.n1795 34.6358
R4896 VSS.n4785 VSS.n4784 34.6358
R4897 VSS.n4559 VSS.n3585 34.6358
R4898 VSS.n4552 VSS.n4551 34.6358
R4899 VSS.n4553 VSS.n4552 34.6358
R4900 VSS.n4548 VSS.n4547 34.6358
R4901 VSS.n4541 VSS.n3594 34.6358
R4902 VSS.n4545 VSS.n3594 34.6358
R4903 VSS.n4522 VSS.n4521 34.6358
R4904 VSS.n4493 VSS.n3619 34.6358
R4905 VSS.n4486 VSS.n3623 34.6358
R4906 VSS.n4482 VSS.n4479 34.6358
R4907 VSS.n4477 VSS.n3626 34.6358
R4908 VSS.n4467 VSS.n4466 34.6358
R4909 VSS.n4467 VSS.n3629 34.6358
R4910 VSS.n4471 VSS.n3629 34.6358
R4911 VSS.n4448 VSS.n3638 34.6358
R4912 VSS.n4452 VSS.n3638 34.6358
R4913 VSS.n4440 VSS.n3643 34.6358
R4914 VSS.n4441 VSS.n4440 34.6358
R4915 VSS.n4442 VSS.n4441 34.6358
R4916 VSS.n4435 VSS.n4434 34.6358
R4917 VSS.n4429 VSS.n4428 34.6358
R4918 VSS.n4430 VSS.n4429 34.6358
R4919 VSS.n4418 VSS.n3651 34.6358
R4920 VSS.n4422 VSS.n3651 34.6358
R4921 VSS.n4416 VSS.n4415 34.6358
R4922 VSS.n4412 VSS.n4411 34.6358
R4923 VSS.n4405 VSS.n4404 34.6358
R4924 VSS.n4405 VSS.n3658 34.6358
R4925 VSS.n4409 VSS.n3658 34.6358
R4926 VSS.n4398 VSS.n3662 34.6358
R4927 VSS.n4402 VSS.n3662 34.6358
R4928 VSS.n4392 VSS.n4391 34.6358
R4929 VSS.n4377 VSS.n4376 34.6358
R4930 VSS.n4379 VSS.n4377 34.6358
R4931 VSS.n4383 VSS.n3673 34.6358
R4932 VSS.n4386 VSS.n4385 34.6358
R4933 VSS.n4367 VSS.n3678 34.6358
R4934 VSS.n4371 VSS.n3678 34.6358
R4935 VSS.n4372 VSS.n4371 34.6358
R4936 VSS.n4373 VSS.n4372 34.6358
R4937 VSS.n4359 VSS.n4358 34.6358
R4938 VSS.n4360 VSS.n4359 34.6358
R4939 VSS.n4360 VSS.n3681 34.6358
R4940 VSS.n4364 VSS.n3681 34.6358
R4941 VSS.n4365 VSS.n4364 34.6358
R4942 VSS.n4336 VSS.n4335 34.6358
R4943 VSS.n4336 VSS.n3692 34.6358
R4944 VSS.n4340 VSS.n3692 34.6358
R4945 VSS.n4328 VSS.n4327 34.6358
R4946 VSS.n4329 VSS.n4328 34.6358
R4947 VSS.n4329 VSS.n3696 34.6358
R4948 VSS.n4333 VSS.n3696 34.6358
R4949 VSS.n4321 VSS.n3700 34.6358
R4950 VSS.n4322 VSS.n4321 34.6358
R4951 VSS.n4310 VSS.n4309 34.6358
R4952 VSS.n3751 VSS.n3750 34.6358
R4953 VSS.n3768 VSS.n3737 34.6358
R4954 VSS.n3764 VSS.n3737 34.6358
R4955 VSS.n3778 VSS.n3777 34.6358
R4956 VSS.n3777 VSS.n3776 34.6358
R4957 VSS.n3776 VSS.n3735 34.6358
R4958 VSS.n3772 VSS.n3735 34.6358
R4959 VSS.n3772 VSS.n3771 34.6358
R4960 VSS.n3782 VSS.n3731 34.6358
R4961 VSS.n3723 VSS.n3722 34.6358
R4962 VSS.n4906 VSS.n4901 34.6358
R4963 VSS.n3810 VSS.n3788 34.6358
R4964 VSS.n4565 VSS.n4564 34.6358
R4965 VSS.n4570 VSS.n4569 34.6358
R4966 VSS.n4571 VSS.n4570 34.6358
R4967 VSS.n4571 VSS.n3580 34.6358
R4968 VSS.n4579 VSS.n4576 34.6358
R4969 VSS.n4583 VSS.n3578 34.6358
R4970 VSS.n4587 VSS.n4586 34.6358
R4971 VSS.n4605 VSS.n4604 34.6358
R4972 VSS.n4613 VSS.n4612 34.6358
R4973 VSS.n4626 VSS.n3560 34.6358
R4974 VSS.n4656 VSS.n1922 34.6358
R4975 VSS.n4660 VSS.n1922 34.6358
R4976 VSS.n4661 VSS.n4660 34.6358
R4977 VSS.n4718 VSS.n4717 34.6358
R4978 VSS.n4717 VSS.n4716 34.6358
R4979 VSS.n275 VSS.t2151 34.506
R4980 VSS.n4960 VSS.t1193 34.506
R4981 VSS.n4968 VSS.t2413 34.506
R4982 VSS.n543 VSS.t1178 34.506
R4983 VSS.n597 VSS.t2569 34.506
R4984 VSS.n604 VSS.t3282 34.506
R4985 VSS.n2389 VSS.t1443 34.506
R4986 VSS.n2382 VSS.t1951 34.506
R4987 VSS.n2374 VSS.t95 34.506
R4988 VSS.n2128 VSS.t3284 34.506
R4989 VSS.n2151 VSS.t570 34.506
R4990 VSS.n2996 VSS.t1479 34.506
R4991 VSS.n994 VSS.t1050 34.506
R4992 VSS.n5153 VSS.t3734 34.2973
R4993 VSS.n5191 VSS.t3712 34.2973
R4994 VSS.n4984 VSS.t3746 34.2973
R4995 VSS.n5391 VSS.t3726 34.2973
R4996 VSS.n937 VSS.t3732 34.2973
R4997 VSS.n3319 VSS.t3763 34.2973
R4998 VSS.n3417 VSS.t3730 34.2973
R4999 VSS.n1267 VSS.t3750 34.2973
R5000 VSS.n1830 VSS.n1821 34.2593
R5001 VSS.n1904 VSS.n1893 34.2593
R5002 VSS.n1917 VSS.n1885 34.2593
R5003 VSS.n4067 VSS.n4058 34.2593
R5004 VSS.n4078 VSS.n4052 34.2593
R5005 VSS.n1811 VSS.n1810 34.2593
R5006 VSS.n1798 VSS.n1797 34.2593
R5007 VSS.n2244 VSS.n2021 34.2593
R5008 VSS.n2499 VSS.n1983 34.2593
R5009 VSS.t2700 VSS.n3872 34.0246
R5010 VSS.n3975 VSS.t2698 34.0246
R5011 VSS.n2076 VSS.n2075 33.8829
R5012 VSS.n2366 VSS.n2004 33.8829
R5013 VSS.n2579 VSS.n2578 33.8829
R5014 VSS.n2627 VSS.n2595 33.8829
R5015 VSS.n3048 VSS.n3047 33.8829
R5016 VSS.n3499 VSS.n3498 33.8829
R5017 VSS.n3506 VSS.n3505 33.8829
R5018 VSS.n3465 VSS.n3464 33.8829
R5019 VSS.n3462 VSS.n3461 33.8829
R5020 VSS.n3392 VSS.n3391 33.8829
R5021 VSS.n3388 VSS.n3387 33.8829
R5022 VSS.n3117 VSS.n3116 33.8829
R5023 VSS.n3126 VSS.n3002 33.8829
R5024 VSS.n3147 VSS.n2994 33.8829
R5025 VSS.n3194 VSS.n3193 33.8829
R5026 VSS.n1399 VSS.n1398 33.8829
R5027 VSS.n1531 VSS.n1512 33.8829
R5028 VSS.n1588 VSS.n1587 33.8829
R5029 VSS.n1656 VSS.n1655 33.8829
R5030 VSS.t2222 VSS.t1111 33.717
R5031 VSS.t2956 VSS.t3663 33.717
R5032 VSS.t1228 VSS.t2948 33.717
R5033 VSS.t1974 VSS.t3102 33.717
R5034 VSS.t3653 VSS.t374 33.717
R5035 VSS.t498 VSS.t199 33.717
R5036 VSS.t1782 VSS.t2604 33.717
R5037 VSS.t2790 VSS.t2722 33.717
R5038 VSS.t3448 VSS.t2704 33.717
R5039 VSS.t1826 VSS.t2184 33.717
R5040 VSS.t3438 VSS.t3636 33.717
R5041 VSS.t1736 VSS.t2437 33.717
R5042 VSS.t2707 VSS.t2940 33.717
R5043 VSS.t2499 VSS.t2406 33.717
R5044 VSS.t2886 VSS.t421 33.717
R5045 VSS.t3092 VSS.t3527 33.717
R5046 VSS.t30 VSS.t2776 33.717
R5047 VSS.t2832 VSS.t1119 33.717
R5048 VSS.t654 VSS.t2548 33.717
R5049 VSS.t1003 VSS.t2960 33.717
R5050 VSS.n871 VSS.n870 33.5064
R5051 VSS.n2303 VSS.n2302 33.5064
R5052 VSS.n2450 VSS.n2449 33.5064
R5053 VSS.n72 VSS.t2215 33.462
R5054 VSS.n72 VSS.t1704 33.462
R5055 VSS.n217 VSS.t233 33.462
R5056 VSS.n217 VSS.t1545 33.462
R5057 VSS.n263 VSS.t2611 33.462
R5058 VSS.n263 VSS.t2539 33.462
R5059 VSS.n278 VSS.t2613 33.462
R5060 VSS.n278 VSS.t865 33.462
R5061 VSS.n4917 VSS.t3504 33.462
R5062 VSS.n4917 VSS.t495 33.462
R5063 VSS.n311 VSS.t2609 33.462
R5064 VSS.n311 VSS.t1319 33.462
R5065 VSS.n2085 VSS.t1989 33.462
R5066 VSS.n2085 VSS.t3506 33.462
R5067 VSS.n3222 VSS.t3028 33.462
R5068 VSS.n3222 VSS.t2329 33.462
R5069 VSS.n2895 VSS.t3373 33.462
R5070 VSS.n2895 VSS.t1023 33.462
R5071 VSS.n3076 VSS.t2807 33.462
R5072 VSS.n3076 VSS.t942 33.462
R5073 VSS.n2972 VSS.t2626 33.462
R5074 VSS.n2972 VSS.t546 33.462
R5075 VSS.n1268 VSS.t2870 33.462
R5076 VSS.n1268 VSS.t2388 33.462
R5077 VSS.n3599 VSS.t1804 33.462
R5078 VSS.n3599 VSS.t2039 33.462
R5079 VSS.n3614 VSS.t1056 33.462
R5080 VSS.n3614 VSS.t3029 33.462
R5081 VSS.n3618 VSS.t1979 33.462
R5082 VSS.n3618 VSS.t3611 33.462
R5083 VSS.n3640 VSS.t1846 33.462
R5084 VSS.n3640 VSS.t2291 33.462
R5085 VSS.n3691 VSS.t2122 33.462
R5086 VSS.n3691 VSS.t2693 33.462
R5087 VSS.n3571 VSS.t1486 33.462
R5088 VSS.n3571 VSS.t1730 33.462
R5089 VSS.n4606 VSS.t3532 33.462
R5090 VSS.n4606 VSS.t2591 33.462
R5091 VSS.n1982 VSS.t2563 33.2313
R5092 VSS.n2586 VSS.t971 33.2313
R5093 VSS.n2603 VSS.t2244 33.2313
R5094 VSS.n2606 VSS.t1044 33.2313
R5095 VSS.n1166 VSS.t153 33.2313
R5096 VSS.n1378 VSS.t3049 33.2313
R5097 VSS.n1383 VSS.t1887 33.2313
R5098 VSS.n1133 VSS.t576 33.2313
R5099 VSS.n1128 VSS.t3496 33.2313
R5100 VSS.n1511 VSS.t1637 33.2313
R5101 VSS.n1820 VSS.t2687 33.2313
R5102 VSS.n1892 VSS.t3024 33.2313
R5103 VSS.n1891 VSS.t1788 33.2313
R5104 VSS.n1884 VSS.t2630 33.2313
R5105 VSS.n1883 VSS.t1777 33.2313
R5106 VSS.n4057 VSS.t1779 33.2313
R5107 VSS.n4077 VSS.t3554 33.2313
R5108 VSS.n1780 VSS.t2800 33.2313
R5109 VSS.n1779 VSS.t2642 33.2313
R5110 VSS.n1788 VSS.t2860 33.2313
R5111 VSS.n1787 VSS.t2847 33.2313
R5112 VSS.n818 VSS.n399 33.1299
R5113 VSS.n2484 VSS.n1987 33.1299
R5114 VSS.n1006 VSS.n1003 33.1299
R5115 VSS.n2079 VSS.n2078 33.1299
R5116 VSS.n2241 VSS.n2240 33.1299
R5117 VSS.n2163 VSS.n2162 32.7534
R5118 VSS.n1085 VSS.n1084 32.7534
R5119 VSS.n4267 VSS.t2635 32.5028
R5120 VSS.n4260 VSS.t2637 32.5028
R5121 VSS.n5090 VSS.n5089 32.377
R5122 VSS.n780 VSS.n779 32.377
R5123 VSS.n1548 VSS.n1505 32.377
R5124 VSS.n2244 VSS.n2243 32.377
R5125 VSS.n2146 VSS.t2789 32.3082
R5126 VSS.n2041 VSS.t3081 32.3082
R5127 VSS.n2250 VSS.t3076 32.3082
R5128 VSS.n2269 VSS.t3086 32.3082
R5129 VSS.n2864 VSS.t1833 32.3082
R5130 VSS.n2902 VSS.t3404 32.3082
R5131 VSS.n2908 VSS.t1827 32.3082
R5132 VSS.n2920 VSS.t1835 32.3082
R5133 VSS.n2947 VSS.t3395 32.3082
R5134 VSS.n3168 VSS.t1829 32.3082
R5135 VSS.n1387 VSS.t1279 32.3082
R5136 VSS.n1820 VSS.t1176 32.3082
R5137 VSS.n1892 VSS.t525 32.3082
R5138 VSS.n1891 VSS.t2399 32.3082
R5139 VSS.n1884 VSS.t1404 32.3082
R5140 VSS.n1883 VSS.t698 32.3082
R5141 VSS.n4057 VSS.t964 32.3082
R5142 VSS.n4077 VSS.t109 32.3082
R5143 VSS.n1780 VSS.t1898 32.3082
R5144 VSS.n1779 VSS.t541 32.3082
R5145 VSS.n1788 VSS.t223 32.3082
R5146 VSS.n1787 VSS.t863 32.3082
R5147 VSS.n3631 VSS.t2796 32.3082
R5148 VSS.n3645 VSS.t2792 32.3082
R5149 VSS.n3660 VSS.t2799 32.3082
R5150 VSS.n3582 VSS.t3393 32.3082
R5151 VSS.n4662 VSS.t1837 32.3082
R5152 VSS.n4284 VSS.n4283 32.1808
R5153 VSS.n1751 VSS.n1742 32.0005
R5154 VSS.n2119 VSS.n2047 32.0005
R5155 VSS.n2671 VSS.n2670 32.0005
R5156 VSS.n2822 VSS.n2821 32.0005
R5157 VSS.n1704 VSS.n1703 32.0005
R5158 VSS.n4030 VSS.n4029 32.0005
R5159 VSS.n1554 VSS.n1502 31.624
R5160 VSS.n1869 VSS.n1868 31.4781
R5161 VSS.n1868 VSS.n1867 31.4781
R5162 VSS.n2441 VSS.n2440 31.2476
R5163 VSS.n1826 VSS.n1825 31.2476
R5164 VSS.n1900 VSS.n1899 31.2476
R5165 VSS.n1913 VSS.n1912 31.2476
R5166 VSS.n4063 VSS.n4062 31.2476
R5167 VSS.n4076 VSS.n4075 31.2476
R5168 VSS.n1808 VSS.n1783 31.2476
R5169 VSS.n1795 VSS.n1791 31.2476
R5170 VSS.n5089 VSS.n214 30.8711
R5171 VSS.n2175 VSS.n2152 30.8711
R5172 VSS.n2504 VSS.n2503 30.8711
R5173 VSS.n1489 VSS.n1123 30.8711
R5174 VSS.n1088 VSS.n1087 30.8711
R5175 VSS.n890 VSS.n889 30.7665
R5176 VSS.n813 VSS.n812 30.7665
R5177 VSS.n2888 VSS.n2860 30.7665
R5178 VSS.n3530 VSS.n2757 30.7665
R5179 VSS.n3081 VSS.n3019 30.7665
R5180 VSS.n3182 VSS.n2984 30.7665
R5181 VSS.n1346 VSS.n1345 30.7665
R5182 VSS.n5376 VSS.t3147 30.5899
R5183 VSS.n2388 VSS.n1999 30.4946
R5184 VSS.n2447 VSS.n2446 30.4946
R5185 VSS.n2436 VSS.n2435 30.4946
R5186 VSS.n3511 VSS.n3510 30.4946
R5187 VSS.n1479 VSS.n1478 30.4946
R5188 VSS.n1980 VSS.t1294 30.462
R5189 VSS.n2750 VSS.t2783 30.462
R5190 VSS.n1023 VSS.t1583 30.462
R5191 VSS.n2309 VSS.n2308 30.2506
R5192 VSS.n2557 VSS.n2556 30.2506
R5193 VSS.n2194 VSS.n2193 29.8804
R5194 VSS.t1760 VSS.n4255 29.7943
R5195 VSS.n5061 VSS.n228 29.7417
R5196 VSS.n909 VSS.n908 29.7417
R5197 VSS.n798 VSS.n797 29.7417
R5198 VSS.n757 VSS.n756 29.7417
R5199 VSS.n2189 VSS.n2188 29.7417
R5200 VSS.n2622 VSS.n2621 29.7417
R5201 VSS.n2681 VSS.n2680 29.7417
R5202 VSS.n2674 VSS.n2650 29.7417
R5203 VSS.n2825 VSS.n2801 29.7417
R5204 VSS.n2832 VSS.n2831 29.7417
R5205 VSS.n3384 VSS.n2925 29.7417
R5206 VSS.n3142 VSS.n3141 29.7417
R5207 VSS.n1453 VSS.n1452 29.7417
R5208 VSS.n1492 VSS.n1491 29.7417
R5209 VSS.n4354 VSS.n3683 29.7417
R5210 VSS.n1980 VSS.t673 29.539
R5211 VSS.n2750 VSS.t853 29.539
R5212 VSS.n1023 VSS.t1314 29.539
R5213 VSS.t2154 VSS.t961 29.4244
R5214 VSS.t2152 VSS.t959 29.4244
R5215 VSS.t2158 VSS.t957 29.4244
R5216 VSS.n4732 VSS.t718 29.3883
R5217 VSS.n509 VSS.n506 29.3652
R5218 VSS.n872 VSS.n871 29.3652
R5219 VSS.n681 VSS.n680 29.3652
R5220 VSS.n2230 VSS.n2029 29.3652
R5221 VSS.n2248 VSS.n2247 29.3652
R5222 VSS.n2392 VSS.n1996 29.3652
R5223 VSS.n3456 VSS.n3455 29.3652
R5224 VSS.n3198 VSS.n2977 29.3652
R5225 VSS.n1437 VSS.n1436 29.3652
R5226 VSS.n1109 VSS.n1106 29.3652
R5227 VSS.n4285 VSS.n4284 29.2561
R5228 VSS.n876 VSS.n357 28.9887
R5229 VSS.n2209 VSS.n2038 28.9887
R5230 VSS.n2434 VSS.n2414 28.9887
R5231 VSS.n2509 VSS.n1979 28.9887
R5232 VSS.n2615 VSS.n2614 28.9887
R5233 VSS.n3367 VSS.n3366 28.9887
R5234 VSS.n4165 VSS.n4164 28.9887
R5235 VSS.n4163 VSS.n3938 28.9887
R5236 VSS.n35 VSS.t662 28.7917
R5237 VSS.n32 VSS.t979 28.7917
R5238 VSS.n222 VSS.t627 28.7917
R5239 VSS.n254 VSS.t271 28.7917
R5240 VSS.n283 VSS.t2013 28.7917
R5241 VSS.n4920 VSS.t2320 28.7917
R5242 VSS.n303 VSS.t1472 28.7917
R5243 VSS.n287 VSS.t763 28.7917
R5244 VSS.n288 VSS.t1956 28.7917
R5245 VSS.n312 VSS.t1134 28.7917
R5246 VSS.n315 VSS.t1066 28.7917
R5247 VSS.n516 VSS.t1138 28.7917
R5248 VSS.n5394 VSS.t3274 28.7917
R5249 VSS.n5397 VSS.t388 28.7917
R5250 VSS.n5398 VSS.t1520 28.7917
R5251 VSS.n5401 VSS.t938 28.7917
R5252 VSS.n5402 VSS.t1206 28.7917
R5253 VSS.n2059 VSS.t410 28.7917
R5254 VSS.n2063 VSS.t217 28.7917
R5255 VSS.n2064 VSS.t976 28.7917
R5256 VSS.n2056 VSS.t1076 28.7917
R5257 VSS.n2653 VSS.t1961 28.7917
R5258 VSS.n2656 VSS.t1904 28.7917
R5259 VSS.n2657 VSS.t275 28.7917
R5260 VSS.n3031 VSS.t2285 28.7917
R5261 VSS.n3035 VSS.t2179 28.7917
R5262 VSS.n3036 VSS.t3277 28.7917
R5263 VSS.n2814 VSS.t115 28.7917
R5264 VSS.n2815 VSS.t1155 28.7917
R5265 VSS.n2804 VSS.t2567 28.7917
R5266 VSS.n2865 VSS.t928 28.7917
R5267 VSS.n2937 VSS.t713 28.7917
R5268 VSS.n3027 VSS.t1355 28.7917
R5269 VSS.n3028 VSS.t1236 28.7917
R5270 VSS.n3024 VSS.t1881 28.7917
R5271 VSS.n3067 VSS.t2553 28.7917
R5272 VSS.n3021 VSS.t767 28.7917
R5273 VSS.n3073 VSS.t2534 28.7917
R5274 VSS.n3110 VSS.t563 28.7917
R5275 VSS.n1148 VSS.t2444 28.7917
R5276 VSS.n998 VSS.t1889 28.7917
R5277 VSS.n1710 VSS.t1230 28.7917
R5278 VSS.n1711 VSS.t1028 28.7917
R5279 VSS.n977 VSS.t2029 28.7917
R5280 VSS.n961 VSS.t293 28.7917
R5281 VSS.n962 VSS.t391 28.7917
R5282 VSS.n1273 VSS.t2277 28.7917
R5283 VSS.n1274 VSS.t967 28.7917
R5284 VSS.n1276 VSS.t2325 28.7917
R5285 VSS.n1277 VSS.t83 28.7917
R5286 VSS.n3596 VSS.t2599 28.7917
R5287 VSS.n3607 VSS.t729 28.7917
R5288 VSS.n3621 VSS.t1203 28.7917
R5289 VSS.n3635 VSS.t2161 28.7917
R5290 VSS.n3648 VSS.t267 28.7917
R5291 VSS.n3664 VSS.t2511 28.7917
R5292 VSS.n3688 VSS.t369 28.7917
R5293 VSS.n3704 VSS.t1918 28.7917
R5294 VSS.n3707 VSS.t91 28.7917
R5295 VSS.n3744 VSS.t1965 28.7917
R5296 VSS.n3756 VSS.t1519 28.7917
R5297 VSS.n4592 VSS.t48 28.7917
R5298 VSS.n3565 VSS.t99 28.7917
R5299 VSS.n4632 VSS.t799 28.7917
R5300 VSS.n4649 VSS.t593 28.7917
R5301 VSS.n4668 VSS.t2312 28.7917
R5302 VSS.n4674 VSS.t719 28.7917
R5303 VSS.n4677 VSS.t139 28.7917
R5304 VSS.n4680 VSS.t2199 28.7917
R5305 VSS.n4683 VSS.t746 28.7917
R5306 VSS.n2319 VSS.t1096 28.6159
R5307 VSS.n2319 VSS.t3605 28.6159
R5308 VSS.n2275 VSS.t1094 28.6159
R5309 VSS.n2275 VSS.t3619 28.6159
R5310 VSS.n2395 VSS.t1092 28.6159
R5311 VSS.n2395 VSS.t3615 28.6159
R5312 VSS.n2545 VSS.t3470 28.6159
R5313 VSS.n2545 VSS.t3623 28.6159
R5314 VSS.n2281 VSS.t3069 28.6159
R5315 VSS.n2409 VSS.t1 28.3801
R5316 VSS.n2756 VSS.t408 28.3801
R5317 VSS.n1185 VSS.t2450 28.3801
R5318 VSS.n1357 VSS.t582 28.3801
R5319 VSS.n1034 VSS.t396 28.3801
R5320 VSS.n1045 VSS.t568 28.3801
R5321 VSS.n1643 VSS.t2118 28.3801
R5322 VSS.n3562 VSS.t603 28.3801
R5323 VSS.n2763 VSS.t1902 28.3166
R5324 VSS.n86 VSS.n85 28.2358
R5325 VSS.n5278 VSS.n129 28.2358
R5326 VSS.n5230 VSS.n152 28.2358
R5327 VSS.n5219 VSS.n155 28.2358
R5328 VSS.n5207 VSS.n162 28.2358
R5329 VSS.n5170 VSS.n176 28.2358
R5330 VSS.n5106 VSS.n203 28.2358
R5331 VSS.n5098 VSS.n5097 28.2358
R5332 VSS.n5023 VSS.n247 28.2358
R5333 VSS.n877 VSS.n876 28.2358
R5334 VSS.n725 VSS.n470 28.2358
R5335 VSS.n659 VSS.n658 28.2358
R5336 VSS.n607 VSS.n536 28.2358
R5337 VSS.n2091 VSS.n2090 28.2358
R5338 VSS.n2365 VSS.n2364 28.2358
R5339 VSS.n2534 VSS.n2533 28.2358
R5340 VSS.n1345 VSS.n1344 28.2358
R5341 VSS.n2274 VSS.n2272 28.2358
R5342 VSS.n1671 VSS.n1670 28.2358
R5343 VSS.t96 VSS.t504 28.2056
R5344 VSS.n576 VSS.n554 27.8593
R5345 VSS.n2240 VSS.n2025 27.8593
R5346 VSS.n2525 VSS.n2524 27.8593
R5347 VSS.n3514 VSS.n2760 27.8593
R5348 VSS.n3503 VSS.n2769 27.8593
R5349 VSS.n3395 VSS.n3394 27.8593
R5350 VSS.n3340 VSS.n2949 27.8593
R5351 VSS.n3274 VSS.n3229 27.8593
R5352 VSS.n4748 VSS.n4738 27.8593
R5353 VSS.n4097 VSS.n4090 27.8593
R5354 VSS.n4784 VSS.n4783 27.8593
R5355 VSS.n4379 VSS.n4378 27.8593
R5356 VSS.n4016 VSS.n4012 27.7877
R5357 VSS.n4256 VSS.t1760 27.7629
R5358 VSS.n894 VSS.n344 27.6711
R5359 VSS.n817 VSS.n816 27.6711
R5360 VSS.n2493 VSS.n2487 27.6711
R5361 VSS.n2884 VSS.n2877 27.6711
R5362 VSS.n3188 VSS.n3187 27.6711
R5363 VSS.n3932 VSS.n3914 27.6576
R5364 VSS.n2399 VSS.t695 27.5691
R5365 VSS.n2404 VSS.t2020 27.5691
R5366 VSS.n2779 VSS.t2254 27.5691
R5367 VSS.n1019 VSS.t669 27.5691
R5368 VSS.n363 VSS.n360 27.4829
R5369 VSS.n2259 VSS.n2258 27.4829
R5370 VSS.n2505 VSS.n2504 27.4829
R5371 VSS.n3374 VSS.n3373 27.4829
R5372 VSS.n1243 VSS.n1242 27.4829
R5373 VSS.n1472 VSS.n1134 27.4829
R5374 VSS.n1530 VSS.n1529 27.4829
R5375 VSS.n1612 VSS.n1610 27.4829
R5376 VSS.n1077 VSS.n1041 27.4829
R5377 VSS.n4335 VSS.n4334 27.4829
R5378 VSS.n2576 VSS.n2575 27.4829
R5379 VSS.n3521 VSS.n3520 27.434
R5380 VSS.n4966 VSS.n273 27.2385
R5381 VSS.n2381 VSS.n2380 27.2385
R5382 VSS.n2158 VSS.n2155 27.1064
R5383 VSS.n2583 VSS.n1955 27.1064
R5384 VSS.n1550 VSS.n1549 27.1064
R5385 VSS.n4822 VSS.n4821 26.9005
R5386 VSS.n3858 VSS.n3822 26.9005
R5387 VSS.n2517 VSS.t956 26.8576
R5388 VSS.n2568 VSS.t1068 26.8576
R5389 VSS.n2605 VSS.t857 26.8576
R5390 VSS.n210 VSS.t611 26.7697
R5391 VSS.n1499 VSS.t934 26.7697
R5392 VSS.n1514 VSS.t2360 26.7697
R5393 VSS.n3694 VSS.t1114 26.7697
R5394 VSS.n5324 VSS.n5323 26.7299
R5395 VSS.n5276 VSS.n5275 26.7299
R5396 VSS.n882 VSS.n354 26.7299
R5397 VSS.n747 VSS.n746 26.7299
R5398 VSS.n662 VSS.n502 26.7299
R5399 VSS.n2104 VSS.n2103 26.7299
R5400 VSS.n3519 VSS.n3518 26.7299
R5401 VSS.n1340 VSS.n1339 26.7299
R5402 VSS.n3268 VSS.n3267 26.6009
R5403 VSS.t1705 VSS.t2326 26.4906
R5404 VSS.n4998 VSS.n4997 26.3534
R5405 VSS.n864 VSS.n863 26.3534
R5406 VSS.n1438 VSS.n1376 26.3534
R5407 VSS.n1620 VSS.n1619 26.3534
R5408 VSS.n1695 VSS.n1694 26.3534
R5409 VSS.n5102 VSS.n207 25.977
R5410 VSS.n5103 VSS.n5102 25.977
R5411 VSS.n5096 VSS.n211 25.977
R5412 VSS.n2351 VSS.n2349 25.977
R5413 VSS.n2562 VSS.n2561 25.977
R5414 VSS.n3547 VSS.n3546 25.977
R5415 VSS.n3205 VSS.n2975 25.977
R5416 VSS.n1250 VSS.n1180 25.977
R5417 VSS.n1365 VSS.n1364 25.977
R5418 VSS.n1423 VSS.n1384 25.977
R5419 VSS.n1629 VSS.n1022 25.977
R5420 VSS.n1651 VSS.n1015 25.977
R5421 VSS.n1831 VSS.n1830 25.977
R5422 VSS.n1905 VSS.n1904 25.977
R5423 VSS.n1918 VSS.n1917 25.977
R5424 VSS.n4068 VSS.n4067 25.977
R5425 VSS.n4083 VSS.n4052 25.977
R5426 VSS.n1811 VSS.n1776 25.977
R5427 VSS.n1798 VSS.n1785 25.977
R5428 VSS.n4557 VSS.n3588 25.977
R5429 VSS.n4529 VSS.n3600 25.977
R5430 VSS.n4526 VSS.n3603 25.977
R5431 VSS.n4499 VSS.n3616 25.977
R5432 VSS.n4460 VSS.n4459 25.977
R5433 VSS.n3763 VSS.n3762 25.977
R5434 VSS.n3784 VSS.n3783 25.977
R5435 VSS.n4598 VSS.n3574 25.977
R5436 VSS.n4630 VSS.n3560 25.977
R5437 VSS.n2141 VSS.t2500 25.9346
R5438 VSS.n2933 VSS.t2189 25.9346
R5439 VSS.n4111 VSS.t1778 25.8881
R5440 VSS.n433 VSS.t1163 25.8467
R5441 VSS.n433 VSS.t1430 25.8467
R5442 VSS.n2773 VSS.t1879 25.8467
R5443 VSS.n2773 VSS.t3047 25.8467
R5444 VSS.n2782 VSS.t471 25.8467
R5445 VSS.n2782 VSS.t2775 25.8467
R5446 VSS.n3018 VSS.t452 25.8467
R5447 VSS.n3018 VSS.t450 25.8467
R5448 VSS.n3013 VSS.t1812 25.8467
R5449 VSS.n3013 VSS.t2898 25.8467
R5450 VSS.n1854 VSS.t2066 25.8467
R5451 VSS.n1854 VSS.t2064 25.8467
R5452 VSS.n4744 VSS.t1347 25.8467
R5453 VSS.n4744 VSS.t1341 25.8467
R5454 VSS.n4745 VSS.t2111 25.8467
R5455 VSS.n4745 VSS.t2110 25.8467
R5456 VSS.n4734 VSS.t2275 25.8467
R5457 VSS.n4734 VSS.t2276 25.8467
R5458 VSS.n4735 VSS.t1186 25.8467
R5459 VSS.n4735 VSS.t1180 25.8467
R5460 VSS.n4086 VSS.t2302 25.8467
R5461 VSS.n4086 VSS.t2306 25.8467
R5462 VSS.n4092 VSS.t1500 25.8467
R5463 VSS.n4092 VSS.t1496 25.8467
R5464 VSS.n4777 VSS.t166 25.8467
R5465 VSS.n4777 VSS.t162 25.8467
R5466 VSS.n4778 VSS.t601 25.8467
R5467 VSS.n4778 VSS.t600 25.8467
R5468 VSS.n4790 VSS.t1364 25.8467
R5469 VSS.n4790 VSS.t1363 25.8467
R5470 VSS.n4791 VSS.t196 25.8467
R5471 VSS.n4791 VSS.t190 25.8467
R5472 VSS.n5247 VSS.n144 25.7355
R5473 VSS.n5083 VSS.n218 25.7355
R5474 VSS.n631 VSS.n630 25.7355
R5475 VSS.n2328 VSS.n2266 25.7355
R5476 VSS.n3453 VSS.n2897 25.7355
R5477 VSS.n77 VSS.n30 25.6926
R5478 VSS.n85 VSS.n27 25.6926
R5479 VSS.n5181 VSS.n171 25.6926
R5480 VSS.n5143 VSS.n187 25.6926
R5481 VSS.n5110 VSS.n203 25.6926
R5482 VSS.n4974 VSS.n271 25.6926
R5483 VSS.n950 VSS.n313 25.6926
R5484 VSS.n835 VSS.n834 25.6926
R5485 VSS.n5472 VSS.n5471 25.6926
R5486 VSS.n5442 VSS.n5383 25.6926
R5487 VSS.n2302 VSS.n2301 25.6926
R5488 VSS.n1219 VSS.n1218 25.6926
R5489 VSS.n4506 VSS.n3612 25.6926
R5490 VSS.n53 VSS.n51 25.6005
R5491 VSS.n60 VSS.n59 25.6005
R5492 VSS.n66 VSS.n65 25.6005
R5493 VSS.n5351 VSS.n5350 25.6005
R5494 VSS.n5318 VSS.n5317 25.6005
R5495 VSS.n5270 VSS.n5269 25.6005
R5496 VSS.n5238 VSS.n5237 25.6005
R5497 VSS.n5212 VSS.n5211 25.6005
R5498 VSS.n5175 VSS.n5174 25.6005
R5499 VSS.n5126 VSS.n194 25.6005
R5500 VSS.n5069 VSS.n5068 25.6005
R5501 VSS.n5029 VSS.n244 25.6005
R5502 VSS.n5019 VSS.n5018 25.6005
R5503 VSS.n5011 VSS.n5010 25.6005
R5504 VSS.n4942 VSS.n4941 25.6005
R5505 VSS.n4930 VSS.n4929 25.6005
R5506 VSS.n295 VSS.n294 25.6005
R5507 VSS.n5415 VSS.n5414 25.6005
R5508 VSS.n5409 VSS.n5408 25.6005
R5509 VSS.n2071 VSS.n2070 25.6005
R5510 VSS.n2571 VSS.n1958 25.6005
R5511 VSS.n2670 VSS.n2654 25.6005
R5512 VSS.n2664 VSS.n2658 25.6005
R5513 VSS.n3043 VSS.n3042 25.6005
R5514 VSS.n2813 VSS.n2807 25.6005
R5515 VSS.n2821 VSS.n2805 25.6005
R5516 VSS.n3361 VSS.n3360 25.6005
R5517 VSS.n3056 VSS.n3055 25.6005
R5518 VSS.n3062 VSS.n3061 25.6005
R5519 VSS.n1371 VSS.n1370 25.6005
R5520 VSS.n1689 VSS.n1688 25.6005
R5521 VSS.n1713 VSS.n958 25.6005
R5522 VSS.n969 VSS.n968 25.6005
R5523 VSS.n1290 VSS.n1289 25.6005
R5524 VSS.n1284 VSS.n1283 25.6005
R5525 VSS.n4539 VSS.n3597 25.6005
R5526 VSS.n4515 VSS.n4514 25.6005
R5527 VSS.n4488 VSS.n4487 25.6005
R5528 VSS.n4454 VSS.n4453 25.6005
R5529 VSS.n4424 VSS.n4423 25.6005
R5530 VSS.n4397 VSS.n4396 25.6005
R5531 VSS.n4348 VSS.n3686 25.6005
R5532 VSS.n4315 VSS.n4314 25.6005
R5533 VSS.n4307 VSS.n3709 25.6005
R5534 VSS.n3749 VSS.n3743 25.6005
R5535 VSS.n3755 VSS.n3741 25.6005
R5536 VSS.n3804 VSS.n3803 25.6005
R5537 VSS.n4591 VSS.n3576 25.6005
R5538 VSS.n4618 VSS.n4617 25.6005
R5539 VSS.n4647 VSS.n1926 25.6005
R5540 VSS.n4654 VSS.n1924 25.6005
R5541 VSS.n4729 VSS.n4728 25.6005
R5542 VSS.n4712 VSS.n4711 25.6005
R5543 VSS.n4706 VSS.n4705 25.6005
R5544 VSS.n4700 VSS.n4699 25.6005
R5545 VSS.n4694 VSS.n4693 25.6005
R5546 VSS.n300 VSS.n299 25.5964
R5547 VSS.n974 VSS.n973 25.5964
R5548 VSS.n4273 VSS.n4246 25.4945
R5549 VSS.n91 VSS.t1337 25.4291
R5550 VSS.n119 VSS.t1504 25.4291
R5551 VSS.n125 VSS.t485 25.4291
R5552 VSS.n140 VSS.t1381 25.4291
R5553 VSS.n332 VSS.t2238 25.4291
R5554 VSS.n382 VSS.t1373 25.4291
R5555 VSS.n418 VSS.t1412 25.4291
R5556 VSS.n446 VSS.t1004 25.4291
R5557 VSS.n463 VSS.t587 25.4291
R5558 VSS.n483 VSS.t660 25.4291
R5559 VSS.n496 VSS.t2131 25.4291
R5560 VSS.n497 VSS.t2587 25.4291
R5561 VSS.n513 VSS.t404 25.4291
R5562 VSS.n10 VSS.t176 25.4291
R5563 VSS.n2105 VSS.t2168 25.4291
R5564 VSS.n2257 VSS.t346 25.4291
R5565 VSS.n1949 VSS.t1030 25.4291
R5566 VSS.n2788 VSS.t2052 25.4291
R5567 VSS.n1179 VSS.t2555 25.4291
R5568 VSS.n1173 VSS.t1188 25.4291
R5569 VSS.n1450 VSS.t3427 25.4291
R5570 VSS.n1508 VSS.t2173 25.4291
R5571 VSS.n1518 VSS.t2370 25.4291
R5572 VSS.n1593 VSS.t1975 25.4291
R5573 VSS.n1038 VSS.t1901 25.4291
R5574 VSS.n3702 VSS.t1531 25.4291
R5575 VSS.n4970 VSS.n271 25.3891
R5576 VSS.n607 VSS.n606 25.3891
R5577 VSS.n2376 VSS.n2371 25.3891
R5578 VSS.t2759 VSS.n4035 25.3345
R5579 VSS.t2515 VSS.t931 25.2879
R5580 VSS.t1746 VSS.t2286 25.2879
R5581 VSS.t649 VSS.t2284 25.2879
R5582 VSS.t530 VSS.t449 25.2879
R5583 VSS.t2793 VSS.t1813 25.2879
R5584 VSS.t1871 VSS.t562 25.2879
R5585 VSS.t1674 VSS.t2934 25.2879
R5586 VSS.t792 VSS.t1875 25.2879
R5587 VSS.t1075 VSS.t3505 25.2879
R5588 VSS.t3062 VSS.t2022 25.2879
R5589 VSS.t1884 VSS.t838 25.2879
R5590 VSS.t557 VSS.t848 25.2879
R5591 VSS.t3004 VSS.t1995 25.2879
R5592 VSS.t2243 VSS.t36 25.2879
R5593 VSS.t1318 VSS.t1133 25.2879
R5594 VSS.t1436 VSS.t455 25.2879
R5595 VSS.n87 VSS.n25 25.224
R5596 VSS.n87 VSS.n86 25.224
R5597 VSS.n5325 VSS.n5324 25.224
R5598 VSS.n5325 VSS.n109 25.224
R5599 VSS.n5277 VSS.n5276 25.224
R5600 VSS.n5278 VSS.n5277 25.224
R5601 VSS.n5226 VSS.n5225 25.224
R5602 VSS.n5226 VSS.n152 25.224
R5603 VSS.n5223 VSS.n155 25.224
R5604 VSS.n5224 VSS.n5223 25.224
R5605 VSS.n5105 VSS.n5104 25.224
R5606 VSS.n5106 VSS.n5105 25.224
R5607 VSS.n878 VSS.n354 25.224
R5608 VSS.n878 VSS.n877 25.224
R5609 VSS.n851 VSS.n374 25.224
R5610 VSS.n847 VSS.n374 25.224
R5611 VSS.n746 VSS.n745 25.224
R5612 VSS.n721 VSS.n470 25.224
R5613 VSS.n660 VSS.n659 25.224
R5614 VSS.n2092 VSS.n2091 25.224
R5615 VSS.n2364 VSS.n2006 25.224
R5616 VSS.n2429 VSS.n2428 25.224
R5617 VSS.n2547 VSS.n1966 25.224
R5618 VSS.n2563 VSS.n2562 25.224
R5619 VSS.n2623 VSS.n2622 25.224
R5620 VSS.n2620 VSS.n2601 25.224
R5621 VSS.n3520 VSS.n3519 25.224
R5622 VSS.n3441 VSS.n2900 25.224
R5623 VSS.n3442 VSS.n3441 25.224
R5624 VSS.n3193 VSS.n3192 25.224
R5625 VSS.n3291 VSS.n3290 25.224
R5626 VSS.n1213 VSS.n1212 25.224
R5627 VSS.n1356 VSS.n1156 25.224
R5628 VSS.n1670 VSS.n1669 25.224
R5629 VSS.n1669 VSS.n1007 25.224
R5630 VSS.n1907 VSS.n1905 25.224
R5631 VSS.n1906 VSS.n1889 25.224
R5632 VSS.n4070 VSS.n4068 25.224
R5633 VSS.n4069 VSS.n4055 25.224
R5634 VSS.n1802 VSS.n1785 25.224
R5635 VSS.n1804 VSS.n1803 25.224
R5636 VSS.n4553 VSS.n3588 25.224
R5637 VSS.n4533 VSS.n3600 25.224
R5638 VSS.n4522 VSS.n3603 25.224
R5639 VSS.n4495 VSS.n3616 25.224
R5640 VSS.n4459 VSS.n4458 25.224
R5641 VSS.n3764 VSS.n3763 25.224
R5642 VSS.n3783 VSS.n3782 25.224
R5643 VSS.n4594 VSS.n3574 25.224
R5644 VSS.n5198 VSS.n5197 24.9894
R5645 VSS.n5160 VSS.n181 24.9894
R5646 VSS.n1295 VSS.n1270 24.9894
R5647 VSS.n1762 VSS.t1451 24.9236
R5648 VSS.n1762 VSS.t1455 24.9236
R5649 VSS.n4835 VSS.t2839 24.9236
R5650 VSS.n4835 VSS.t2853 24.9236
R5651 VSS.n209 VSS.t2629 24.9236
R5652 VSS.n209 VSS.t1850 24.9236
R5653 VSS.n213 VSS.t609 24.9236
R5654 VSS.n213 VSS.t607 24.9236
R5655 VSS.n22 VSS.t2209 24.9236
R5656 VSS.n22 VSS.t2205 24.9236
R5657 VSS.n356 VSS.t2969 24.9236
R5658 VSS.n356 VSS.t2972 24.9236
R5659 VSS.n359 VSS.t2127 24.9236
R5660 VSS.n362 VSS.t2982 24.9236
R5661 VSS.n362 VSS.t2703 24.9236
R5662 VSS.n551 VSS.t1272 24.9236
R5663 VSS.n551 VSS.t1264 24.9236
R5664 VSS.n556 VSS.t55 24.9236
R5665 VSS.n2146 VSS.t2183 24.9236
R5666 VSS.n2041 VSS.t1428 24.9236
R5667 VSS.n2028 VSS.t3656 24.9236
R5668 VSS.n2250 VSS.t1523 24.9236
R5669 VSS.n2269 VSS.t103 24.9236
R5670 VSS.n2350 VSS.t2824 24.9236
R5671 VSS.n2008 VSS.t950 24.9236
R5672 VSS.n2008 VSS.t1052 24.9236
R5673 VSS.n2372 VSS.t1651 24.9236
R5674 VSS.n2372 VSS.t2467 24.9236
R5675 VSS.n1995 VSS.t3084 24.9236
R5676 VSS.n2396 VSS.t2023 24.9236
R5677 VSS.n1982 VSS.t3491 24.9236
R5678 VSS.n2510 VSS.t3425 24.9236
R5679 VSS.n2520 VSS.t1060 24.9236
R5680 VSS.n2520 VSS.t2657 24.9236
R5681 VSS.n1963 VSS.t3397 24.9236
R5682 VSS.n1963 VSS.t3413 24.9236
R5683 VSS.n1957 VSS.t2545 24.9236
R5684 VSS.n2586 VSS.t3042 24.9236
R5685 VSS.n2594 VSS.t2242 24.9236
R5686 VSS.n2603 VSS.t2777 24.9236
R5687 VSS.n1947 VSS.t359 24.9236
R5688 VSS.n1947 VSS.t357 24.9236
R5689 VSS.n2878 VSS.t635 24.9236
R5690 VSS.n2878 VSS.t633 24.9236
R5691 VSS.n2864 VSS.t400 24.9236
R5692 VSS.n2762 VSS.t2250 24.9236
R5693 VSS.n2762 VSS.t787 24.9236
R5694 VSS.n2767 VSS.t3402 24.9236
R5695 VSS.n2767 VSS.t3415 24.9236
R5696 VSS.n2768 VSS.t3411 24.9236
R5697 VSS.n2768 VSS.t3406 24.9236
R5698 VSS.n2894 VSS.t3408 24.9236
R5699 VSS.n2902 VSS.t1353 24.9236
R5700 VSS.n2908 VSS.t1215 24.9236
R5701 VSS.n2920 VSS.t1308 24.9236
R5702 VSS.n2921 VSS.t676 24.9236
R5703 VSS.n2921 VSS.t682 24.9236
R5704 VSS.n2940 VSS.t1253 24.9236
R5705 VSS.n2940 VSS.t1259 24.9236
R5706 VSS.n2946 VSS.t732 24.9236
R5707 VSS.n2946 VSS.t736 24.9236
R5708 VSS.n2947 VSS.t1339 24.9236
R5709 VSS.n2954 VSS.t1054 24.9236
R5710 VSS.n2954 VSS.t133 24.9236
R5711 VSS.n3001 VSS.t2900 24.9236
R5712 VSS.n3001 VSS.t1483 24.9236
R5713 VSS.n2992 VSS.t129 24.9236
R5714 VSS.n2992 VSS.t131 24.9236
R5715 VSS.n3158 VSS.t814 24.9236
R5716 VSS.n3158 VSS.t2025 24.9236
R5717 VSS.n3168 VSS.t2124 24.9236
R5718 VSS.n3199 VSS.t3589 24.9236
R5719 VSS.n3199 VSS.t3603 24.9236
R5720 VSS.n3219 VSS.t620 24.9236
R5721 VSS.n3219 VSS.t548 24.9236
R5722 VSS.n3226 VSS.t2354 24.9236
R5723 VSS.n3226 VSS.t2352 24.9236
R5724 VSS.n1188 VSS.t544 24.9236
R5725 VSS.n1163 VSS.t3399 24.9236
R5726 VSS.n1379 VSS.t1597 24.9236
R5727 VSS.n1383 VSS.t2677 24.9236
R5728 VSS.n1387 VSS.t920 24.9236
R5729 VSS.n1131 VSS.t3088 24.9236
R5730 VSS.n1122 VSS.t3502 24.9236
R5731 VSS.n1011 VSS.t1330 24.9236
R5732 VSS.n1011 VSS.t1328 24.9236
R5733 VSS.n1605 VSS.t3079 24.9236
R5734 VSS.n1611 VSS.t3658 24.9236
R5735 VSS.n4000 VSS.t1008 24.9236
R5736 VSS.n4000 VSS.t1007 24.9236
R5737 VSS.n3999 VSS.t178 24.9236
R5738 VSS.n3999 VSS.t184 24.9236
R5739 VSS.n1823 VSS.t1172 24.9236
R5740 VSS.n1823 VSS.t1170 24.9236
R5741 VSS.n1896 VSS.t519 24.9236
R5742 VSS.n1896 VSS.t523 24.9236
R5743 VSS.n1895 VSS.t2401 24.9236
R5744 VSS.n1895 VSS.t2402 24.9236
R5745 VSS.n1888 VSS.t1402 24.9236
R5746 VSS.n1888 VSS.t1401 24.9236
R5747 VSS.n1887 VSS.t700 24.9236
R5748 VSS.n1887 VSS.t702 24.9236
R5749 VSS.n4060 VSS.t960 24.9236
R5750 VSS.n4060 VSS.t958 24.9236
R5751 VSS.n4054 VSS.t107 24.9236
R5752 VSS.n4054 VSS.t111 24.9236
R5753 VSS.n1782 VSS.t1897 24.9236
R5754 VSS.n1782 VSS.t1899 24.9236
R5755 VSS.n1781 VSS.t537 24.9236
R5756 VSS.n1781 VSS.t539 24.9236
R5757 VSS.n1790 VSS.t227 24.9236
R5758 VSS.n1790 VSS.t221 24.9236
R5759 VSS.n1789 VSS.t862 24.9236
R5760 VSS.n1789 VSS.t861 24.9236
R5761 VSS.n3590 VSS.t2040 24.9236
R5762 VSS.n3590 VSS.t2535 24.9236
R5763 VSS.n4480 VSS.t1981 24.9236
R5764 VSS.n4480 VSS.t3280 24.9236
R5765 VSS.n3631 VSS.t2340 24.9236
R5766 VSS.n3645 VSS.t686 24.9236
R5767 VSS.n3654 VSS.t1070 24.9236
R5768 VSS.n3654 VSS.t2085 24.9236
R5769 VSS.n3660 VSS.t1445 24.9236
R5770 VSS.n3672 VSS.t1424 24.9236
R5771 VSS.n3672 VSS.t1426 24.9236
R5772 VSS.n3582 VSS.t1238 24.9236
R5773 VSS.n4577 VSS.t2345 24.9236
R5774 VSS.n4577 VSS.t742 24.9236
R5775 VSS.n4662 VSS.t1249 24.9236
R5776 VSS.n4113 VSS.t2837 24.9236
R5777 VSS.n4113 VSS.t2857 24.9236
R5778 VSS.n4115 VSS.t2155 24.9236
R5779 VSS.n4115 VSS.t2153 24.9236
R5780 VSS.n3936 VSS.t2436 24.9236
R5781 VSS.n3936 VSS.t2433 24.9236
R5782 VSS.n3937 VSS.t2434 24.9236
R5783 VSS.n3937 VSS.t2390 24.9236
R5784 VSS.n3104 VSS.n3101 24.8682
R5785 VSS.n64 VSS.n36 24.8476
R5786 VSS.n70 VSS.n33 24.8476
R5787 VSS.n5073 VSS.n223 24.8476
R5788 VSS.n5037 VSS.n238 24.8476
R5789 VSS.n5006 VSS.n255 24.8476
R5790 VSS.n4943 VSS.n281 24.8476
R5791 VSS.n4931 VSS.n4918 24.8476
R5792 VSS.n299 VSS.n289 24.8476
R5793 VSS.n951 VSS.n950 24.8476
R5794 VSS.n784 VSS.n431 24.8476
R5795 VSS.n732 VSS.n464 24.8476
R5796 VSS.n714 VSS.n473 24.8476
R5797 VSS.n626 VSS.n524 24.8476
R5798 VSS.n5419 VSS.n5399 24.8476
R5799 VSS.n5413 VSS.n5403 24.8476
R5800 VSS.n2075 VSS.n2065 24.8476
R5801 VSS.n2090 VSS.n2057 24.8476
R5802 VSS.n2704 VSS.n2703 24.8476
R5803 VSS.n2666 VSS.n2665 24.8476
R5804 VSS.n3047 VSS.n3037 24.8476
R5805 VSS.n2817 VSS.n2816 24.8476
R5806 VSS.n2869 VSS.n2868 24.8476
R5807 VSS.n3356 VSS.n2938 24.8476
R5808 VSS.n3060 VSS.n3029 24.8476
R5809 VSS.n3066 VSS.n3025 24.8476
R5810 VSS.n3069 VSS.n3068 24.8476
R5811 VSS.n1415 VSS.n1389 24.8476
R5812 VSS.n1052 VSS.n1050 24.8476
R5813 VSS.n1684 VSS.n999 24.8476
R5814 VSS.n1712 VSS.n1709 24.8476
R5815 VSS.n973 VSS.n963 24.8476
R5816 VSS.n1291 VSS.n1270 24.8476
R5817 VSS.n1288 VSS.n1278 24.8476
R5818 VSS.n4541 VSS.n4540 24.8476
R5819 VSS.n4519 VSS.n3608 24.8476
R5820 VSS.n4489 VSS.n3619 24.8476
R5821 VSS.n4458 VSS.n3636 24.8476
R5822 VSS.n4428 VSS.n3649 24.8476
R5823 VSS.n4392 VSS.n3665 24.8476
R5824 VSS.n4347 VSS.n4346 24.8476
R5825 VSS.n4309 VSS.n4308 24.8476
R5826 VSS.n4310 VSS.n3705 24.8476
R5827 VSS.n3745 VSS.n3711 24.8476
R5828 VSS.n3758 VSS.n3757 24.8476
R5829 VSS.n4594 VSS.n4593 24.8476
R5830 VSS.n4613 VSS.n3566 24.8476
R5831 VSS.n4633 VSS.n4631 24.8476
R5832 VSS.n4650 VSS.n4648 24.8476
R5833 VSS.n4724 VSS.n4669 24.8476
R5834 VSS.n4716 VSS.n4675 24.8476
R5835 VSS.n4710 VSS.n4678 24.8476
R5836 VSS.n4704 VSS.n4681 24.8476
R5837 VSS.n4698 VSS.n4684 24.8476
R5838 VSS.n2955 VSS.t3097 24.6931
R5839 VSS.n3150 VSS.t3591 24.6931
R5840 VSS.n3223 VSS.t1161 24.6931
R5841 VSS.n3593 VSS.t918 24.6931
R5842 VSS.n3625 VSS.t780 24.6931
R5843 VSS.n3653 VSS.t3101 24.6931
R5844 VSS.n4584 VSS.t256 24.6931
R5845 VSS.n54 VSS.n53 24.4711
R5846 VSS.n58 VSS.n39 24.4711
R5847 VSS.n5353 VSS.n96 24.4711
R5848 VSS.n5352 VSS.n5351 24.4711
R5849 VSS.n5323 VSS.n112 24.4711
R5850 VSS.n5319 VSS.n5318 24.4711
R5851 VSS.n5275 VSS.n133 24.4711
R5852 VSS.n5271 VSS.n5270 24.4711
R5853 VSS.n5237 VSS.n5236 24.4711
R5854 VSS.n5232 VSS.n150 24.4711
R5855 VSS.n5217 VSS.n159 24.4711
R5856 VSS.n5213 VSS.n5212 24.4711
R5857 VSS.n5177 VSS.n171 24.4711
R5858 VSS.n5176 VSS.n5175 24.4711
R5859 VSS.n5132 VSS.n5131 24.4711
R5860 VSS.n5130 VSS.n194 24.4711
R5861 VSS.n5098 VSS.n207 24.4711
R5862 VSS.n5025 VSS.n244 24.4711
R5863 VSS.n5024 VSS.n5023 24.4711
R5864 VSS.n5018 VSS.n5017 24.4711
R5865 VSS.n5013 VSS.n251 24.4711
R5866 VSS.n861 VSS.n365 24.4711
R5867 VSS.n791 VSS.n427 24.4711
R5868 VSS.n778 VSS.n777 24.4711
R5869 VSS.n736 VSS.n459 24.4711
R5870 VSS.n619 VSS.n532 24.4711
R5871 VSS.n2092 VSS.n2054 24.4711
R5872 VSS.n2096 VSS.n2054 24.4711
R5873 VSS.n2533 VSS.n2532 24.4711
R5874 VSS.n2557 VSS.n1964 24.4711
R5875 VSS.n2561 VSS.n1964 24.4711
R5876 VSS.n3486 VSS.n3485 24.4711
R5877 VSS.n3214 VSS.n2970 24.4711
R5878 VSS.n1314 VSS.n1260 24.4711
R5879 VSS.n1318 VSS.n1260 24.4711
R5880 VSS.n4756 VSS.n4755 24.4711
R5881 VSS.n4103 VSS.n4102 24.4711
R5882 VSS.n4789 VSS.n4771 24.4711
R5883 VSS.n4559 VSS.n4558 24.4711
R5884 VSS.n4558 VSS.n4557 24.4711
R5885 VSS.n4529 VSS.n4528 24.4711
R5886 VSS.n4527 VSS.n4526 24.4711
R5887 VSS.n4501 VSS.n4500 24.4711
R5888 VSS.n4500 VSS.n4499 24.4711
R5889 VSS.n4464 VSS.n3633 24.4711
R5890 VSS.n4460 VSS.n3633 24.4711
R5891 VSS.n3758 VSS.n3739 24.4711
R5892 VSS.n3762 VSS.n3739 24.4711
R5893 VSS.n3784 VSS.n3729 24.4711
R5894 VSS.n3806 VSS.n3788 24.4711
R5895 VSS.n3805 VSS.n3804 24.4711
R5896 VSS.n4599 VSS.n4598 24.4711
R5897 VSS.n4600 VSS.n4599 24.4711
R5898 VSS.n4718 VSS.n4672 24.4711
R5899 VSS.n54 VSS.n39 24.0946
R5900 VSS.n59 VSS.n58 24.0946
R5901 VSS.n65 VSS.n64 24.0946
R5902 VSS.n5353 VSS.n5352 24.0946
R5903 VSS.n5319 VSS.n112 24.0946
R5904 VSS.n5271 VSS.n133 24.0946
R5905 VSS.n5236 VSS.n150 24.0946
R5906 VSS.n5213 VSS.n159 24.0946
R5907 VSS.n5177 VSS.n5176 24.0946
R5908 VSS.n5131 VSS.n5130 24.0946
R5909 VSS.n5068 VSS.n5067 24.0946
R5910 VSS.n5025 VSS.n5024 24.0946
R5911 VSS.n5017 VSS.n251 24.0946
R5912 VSS.n5012 VSS.n5011 24.0946
R5913 VSS.n863 VSS.n862 24.0946
R5914 VSS.n857 VSS.n365 24.0946
R5915 VSS.n742 VSS.n741 24.0946
R5916 VSS.n740 VSS.n459 24.0946
R5917 VSS.n615 VSS.n532 24.0946
R5918 VSS.n5420 VSS.n5419 24.0946
R5919 VSS.n5414 VSS.n5413 24.0946
R5920 VSS.n2176 VSS.n2175 24.0946
R5921 VSS.n2216 VSS.n2215 24.0946
R5922 VSS.n2528 VSS.n2527 24.0946
R5923 VSS.n2567 VSS.n2566 24.0946
R5924 VSS.n2666 VSS.n2654 24.0946
R5925 VSS.n2817 VSS.n2805 24.0946
R5926 VSS.n3531 VSS.n3530 24.0946
R5927 VSS.n3435 VSS.n2903 24.0946
R5928 VSS.n3362 VSS.n3361 24.0946
R5929 VSS.n3354 VSS.n3353 24.0946
R5930 VSS.n3061 VSS.n3060 24.0946
R5931 VSS.n3116 VSS.n3115 24.0946
R5932 VSS.n3178 VSS.n2984 24.0946
R5933 VSS.n1243 VSS.n1186 24.0946
R5934 VSS.n1207 VSS.n1206 24.0946
R5935 VSS.n1170 VSS.n1167 24.0946
R5936 VSS.n1358 VSS.n1356 24.0946
R5937 VSS.n1371 VSS.n1145 24.0946
R5938 VSS.n1414 VSS.n1413 24.0946
R5939 VSS.n1132 VSS.n1129 24.0946
R5940 VSS.n1624 VSS.n1029 24.0946
R5941 VSS.n1063 VSS.n1046 24.0946
R5942 VSS.n1640 VSS.n1020 24.0946
R5943 VSS.n1690 VSS.n1689 24.0946
R5944 VSS.n1289 VSS.n1288 24.0946
R5945 VSS.n4535 VSS.n3597 24.0946
R5946 VSS.n4487 VSS.n4486 24.0946
R5947 VSS.n4453 VSS.n4452 24.0946
R5948 VSS.n4446 VSS.n3641 24.0946
R5949 VSS.n4423 VSS.n4422 24.0946
R5950 VSS.n4411 VSS.n4410 24.0946
R5951 VSS.n4398 VSS.n4397 24.0946
R5952 VSS.n4352 VSS.n3686 24.0946
R5953 VSS.n4316 VSS.n4315 24.0946
R5954 VSS.n3751 VSS.n3741 24.0946
R5955 VSS.n3750 VSS.n3749 24.0946
R5956 VSS.n3806 VSS.n3805 24.0946
R5957 VSS.n4576 VSS.n4575 24.0946
R5958 VSS.n4587 VSS.n3576 24.0946
R5959 VSS.n4619 VSS.n4618 24.0946
R5960 VSS.n4619 VSS.n3563 24.0946
R5961 VSS.n4648 VSS.n4647 24.0946
R5962 VSS.n4724 VSS.n4723 24.0946
R5963 VSS.n4722 VSS.n4672 24.0946
R5964 VSS.n4711 VSS.n4710 24.0946
R5965 VSS.n4705 VSS.n4704 24.0946
R5966 VSS.n4699 VSS.n4698 24.0946
R5967 VSS.n260 VSS.t1387 24.0005
R5968 VSS.n352 VSS.t3601 24.0005
R5969 VSS.n545 VSS.t2820 24.0005
R5970 VSS.n2344 VSS.t335 24.0005
R5971 VSS.n2410 VSS.t917 24.0005
R5972 VSS.n1259 VSS.t510 24.0005
R5973 VSS.n1198 VSS.t203 24.0005
R5974 VSS.n1152 VSS.t252 24.0005
R5975 VSS.n1375 VSS.t2672 24.0005
R5976 VSS.n1027 VSS.t1159 24.0005
R5977 VSS.n682 VSS.n681 23.7181
R5978 VSS.n2335 VSS.n2016 23.7181
R5979 VSS.n5374 VSS.n5373 23.7181
R5980 VSS.n5313 VSS.n5312 23.7181
R5981 VSS.n5265 VSS.n5264 23.7181
R5982 VSS.n5219 VSS.n5218 23.7181
R5983 VSS.n5218 VSS.n5217 23.7181
R5984 VSS.n5170 VSS.n5169 23.7181
R5985 VSS.n5169 VSS.n5168 23.7181
R5986 VSS.n5074 VSS.n5073 23.7181
R5987 VSS.n4992 VSS.n4991 23.7181
R5988 VSS.n4937 VSS.n4915 23.7181
R5989 VSS.n904 VSS.n903 23.7181
R5990 VSS.n903 VSS.n902 23.7181
R5991 VSS.n812 VSS.n811 23.7181
R5992 VSS.n811 VSS.n810 23.7181
R5993 VSS.n771 VSS.n439 23.7181
R5994 VSS.n767 VSS.n439 23.7181
R5995 VSS.n721 VSS.n720 23.7181
R5996 VSS.n714 VSS.n713 23.7181
R5997 VSS.n588 VSS.n587 23.7181
R5998 VSS.n5449 VSS.n5448 23.7181
R5999 VSS.n2204 VSS.n2043 23.7181
R6000 VSS.n2330 VSS.n2264 23.7181
R6001 VSS.n2329 VSS.n2328 23.7181
R6002 VSS.n2288 VSS.n2287 23.7181
R6003 VSS.n2338 VSS.n2015 23.7181
R6004 VSS.n2338 VSS.n2013 23.7181
R6005 VSS.n2475 VSS.n1994 23.7181
R6006 VSS.n2708 VSS.n2636 23.7181
R6007 VSS.n2704 VSS.n2636 23.7181
R6008 VSS.n2890 VSS.n2791 23.7181
R6009 VSS.n3480 VSS.n3479 23.7181
R6010 VSS.n3430 VSS.n3429 23.7181
R6011 VSS.n3163 VSS.n2988 23.7181
R6012 VSS.n3167 VSS.n2988 23.7181
R6013 VSS.n1314 VSS.n1313 23.7181
R6014 VSS.n1254 VSS.n1180 23.7181
R6015 VSS.n1212 VSS.n1202 23.7181
R6016 VSS.n1329 VSS.n1171 23.7181
R6017 VSS.n1443 VSS.n1145 23.7181
R6018 VSS.n1443 VSS.n1442 23.7181
R6019 VSS.n1446 VSS.n1144 23.7181
R6020 VSS.n1446 VSS.n1142 23.7181
R6021 VSS.n1566 VSS.n1120 23.7181
R6022 VSS.n1064 VSS.n1063 23.7181
R6023 VSS.n1627 VSS.n1025 23.7181
R6024 VSS.n1655 VSS.n1015 23.7181
R6025 VSS.n1675 VSS.n1003 23.7181
R6026 VSS.n1704 VSS.n990 23.7181
R6027 VSS.n1709 VSS.n986 23.7181
R6028 VSS.n4563 VSS.n3585 23.7181
R6029 VSS.n4521 VSS.n4520 23.7181
R6030 VSS.n4520 VSS.n4519 23.7181
R6031 VSS.n4473 VSS.n3626 23.7181
R6032 VSS.n4434 VSS.n3646 23.7181
R6033 VSS.n4430 VSS.n3646 23.7181
R6034 VSS.n4391 VSS.n4390 23.7181
R6035 VSS.n4390 VSS.n4389 23.7181
R6036 VSS.n4346 VSS.n3689 23.7181
R6037 VSS.n4342 VSS.n3689 23.7181
R6038 VSS.n4303 VSS.n3711 23.7181
R6039 VSS.n4907 VSS.n4906 23.7181
R6040 VSS.n3811 VSS.n3810 23.7181
R6041 VSS.n4564 VSS.n4563 23.7181
R6042 VSS.n4611 VSS.n3568 23.7181
R6043 VSS.n4612 VSS.n4611 23.7181
R6044 VSS.n4631 VSS.n4630 23.7181
R6045 VSS.n4730 VSS.n1920 23.7181
R6046 VSS.n4821 VSS.n4820 23.7005
R6047 VSS.n3823 VSS.n3822 23.7005
R6048 VSS.n3819 VSS.n3817 23.4005
R6049 VSS.n3817 VSS.n3816 23.4005
R6050 VSS.n3864 VSS.n3815 23.4005
R6051 VSS.n3815 VSS.n3813 23.4005
R6052 VSS.n3989 VSS.n3988 23.4005
R6053 VSS.n3990 VSS.n3989 23.4005
R6054 VSS.n3978 VSS.n3977 23.4005
R6055 VSS.n3977 VSS.n3976 23.4005
R6056 VSS.n2235 VSS.n2234 23.3417
R6057 VSS.n2467 VSS.n2466 23.3417
R6058 VSS.n3546 VSS.n2751 23.3417
R6059 VSS.n1555 VSS.n1554 23.3417
R6060 VSS.n1859 VSS.n1855 23.3417
R6061 VSS.n4747 VSS.n4746 23.3417
R6062 VSS.n4760 VSS.n4736 23.3417
R6063 VSS.n4107 VSS.n4087 23.3417
R6064 VSS.n4096 VSS.n4095 23.3417
R6065 VSS.n4779 VSS.n4773 23.3417
R6066 VSS.n4793 VSS.n4792 23.3417
R6067 VSS.n2498 VSS.n2496 23.2371
R6068 VSS.n3873 VSS.t2652 23.1369
R6069 VSS.n3991 VSS.t2684 23.1369
R6070 VSS.n4969 VSS.n4967 23.0907
R6071 VSS.n605 VSS.n603 23.0907
R6072 VSS.n5369 VSS.n92 22.9652
R6073 VSS.n5311 VSS.n5310 22.9652
R6074 VSS.n5294 VSS.n5293 22.9652
R6075 VSS.n5263 VSS.n5262 22.9652
R6076 VSS.n5062 VSS.n5061 22.9652
R6077 VSS.n5033 VSS.n5032 22.9652
R6078 VSS.n916 VSS.n915 22.9652
R6079 VSS.n908 VSS.n336 22.9652
R6080 VSS.n800 VSS.n799 22.9652
R6081 VSS.n762 VSS.n761 22.9652
R6082 VSS.n757 VSS.n448 22.9652
R6083 VSS.n733 VSS.n732 22.9652
R6084 VSS.n728 VSS.n727 22.9652
R6085 VSS.n719 VSS.n718 22.9652
R6086 VSS.n694 VSS.n693 22.9652
R6087 VSS.n674 VSS.n673 22.9652
R6088 VSS.n673 VSS.n498 22.9652
R6089 VSS.n647 VSS.n646 22.9652
R6090 VSS.n5476 VSS.n11 22.9652
R6091 VSS.n2183 VSS.n2182 22.9652
R6092 VSS.n2251 VSS.n2018 22.9652
R6093 VSS.n2360 VSS.n2358 22.9652
R6094 VSS.n2360 VSS.n2359 22.9652
R6095 VSS.n2505 VSS.n1979 22.9652
R6096 VSS.n2710 VSS.n2709 22.9652
R6097 VSS.n2680 VSS.n2679 22.9652
R6098 VSS.n2831 VSS.n2830 22.9652
R6099 VSS.n2871 VSS.n2870 22.9652
R6100 VSS.n3172 VSS.n3169 22.9652
R6101 VSS.n3188 VSS.n2981 22.9652
R6102 VSS.n3201 VSS.n3200 22.9652
R6103 VSS.n1255 VSS.n1254 22.9652
R6104 VSS.n1420 VSS.n1419 22.9652
R6105 VSS.n1453 VSS.n1140 22.9652
R6106 VSS.n1596 VSS.n1104 22.9652
R6107 VSS.n1595 VSS.n1594 22.9652
R6108 VSS.n1092 VSS.n1032 22.9652
R6109 VSS.n1057 VSS.n1056 22.9652
R6110 VSS.n1650 VSS.n1649 22.9652
R6111 VSS.n4466 VSS.n4465 22.9652
R6112 VSS.n4436 VSS.n3643 22.9652
R6113 VSS.n4404 VSS.n4403 22.9652
R6114 VSS.n4354 VSS.n4353 22.9652
R6115 VSS.n4569 VSS.n3583 22.9652
R6116 VSS.n4626 VSS.n4625 22.9652
R6117 VSS.n4663 VSS.n4661 22.9652
R6118 VSS.n2320 VSS.n2318 22.9145
R6119 VSS.n2428 VSS.n2418 22.6609
R6120 VSS.n4849 VSS.t3698 22.6141
R6121 VSS.n4833 VSS.t3700 22.6141
R6122 VSS.n4832 VSS.t3702 22.6141
R6123 VSS.n4831 VSS.t3704 22.6141
R6124 VSS.n4131 VSS.t3480 22.6141
R6125 VSS.n3943 VSS.t3476 22.6141
R6126 VSS.n3944 VSS.t3478 22.6141
R6127 VSS.n4132 VSS.t3482 22.6141
R6128 VSS.n823 VSS.n822 22.5887
R6129 VSS.n2499 VSS.n2498 22.5887
R6130 VSS.n2579 VSS.n1955 22.5887
R6131 VSS.n1549 VSS.n1548 22.5887
R6132 VSS.n4280 VSS.n3904 22.5005
R6133 VSS.n4281 VSS.n4280 22.5005
R6134 VSS.n4220 VSS.n4215 22.5005
R6135 VSS.n4237 VSS.n4215 22.5005
R6136 VSS.n4226 VSS.n4225 22.5005
R6137 VSS.n4229 VSS.n4226 22.5005
R6138 VSS.n4206 VSS.n4205 22.5005
R6139 VSS.t564 VSS.n4206 22.5005
R6140 VSS.n599 VSS.n538 22.3444
R6141 VSS.n5199 VSS.t2294 22.3257
R6142 VSS.n5162 VSS.t1032 22.3257
R6143 VSS.n189 VSS.t2298 22.3257
R6144 VSS.n422 VSS.t2280 22.3257
R6145 VSS.n526 VSS.t2470 22.3257
R6146 VSS.n5378 VSS.t454 22.3257
R6147 VSS.n2137 VSS.t2425 22.3257
R6148 VSS.n1941 VSS.t3451 22.3257
R6149 VSS.n1175 VSS.t2006 22.3257
R6150 VSS.n1382 VSS.t940 22.3257
R6151 VSS.n1394 VSS.t1072 22.3257
R6152 VSS.n3769 VSS.t2035 22.3257
R6153 VSS.n3733 VSS.t954 22.3257
R6154 VSS.n5362 VSS.n94 22.2496
R6155 VSS.n5305 VSS.n5304 22.2496
R6156 VSS.n5288 VSS.n5287 22.2496
R6157 VSS.n5257 VSS.n5256 22.2496
R6158 VSS.n924 VSS.n921 22.2496
R6159 VSS.n703 VSS.n700 22.2496
R6160 VSS.n564 VSS.n563 22.2496
R6161 VSS.n2719 VSS.n2716 22.2496
R6162 VSS.n3471 VSS.n3470 22.2496
R6163 VSS.n1458 VSS.n1457 22.2496
R6164 VSS.n1601 VSS.n1600 22.2496
R6165 VSS.n73 VSS.n71 22.2123
R6166 VSS.n73 VSS.n30 22.2123
R6167 VSS.n5085 VSS.n5084 22.2123
R6168 VSS.n5084 VSS.n5083 22.2123
R6169 VSS.n4993 VSS.n261 22.2123
R6170 VSS.n4993 VSS.n4992 22.2123
R6171 VSS.n4953 VSS.n279 22.2123
R6172 VSS.n4949 VSS.n279 22.2123
R6173 VSS.n4937 VSS.n4936 22.2123
R6174 VSS.n4936 VSS.n4935 22.2123
R6175 VSS.n713 VSS.n712 22.2123
R6176 VSS.n2335 VSS.n2334 22.2123
R6177 VSS.n2287 VSS.n2286 22.2123
R6178 VSS.n2342 VSS.n2013 22.2123
R6179 VSS.n2454 VSS.n2402 22.2123
R6180 VSS.n2450 VSS.n2402 22.2123
R6181 VSS.n2446 VSS.n2406 22.2123
R6182 VSS.n2875 VSS.n2862 22.2123
R6183 VSS.n3510 VSS.n2765 22.2123
R6184 VSS.n3506 VSS.n2765 22.2123
R6185 VSS.n3488 VSS.n3487 22.2123
R6186 VSS.n3481 VSS.n3480 22.2123
R6187 VSS.n3455 VSS.n3454 22.2123
R6188 VSS.n3454 VSS.n3453 22.2123
R6189 VSS.n3431 VSS.n3430 22.2123
R6190 VSS.n3077 VSS.n3075 22.2123
R6191 VSS.n3077 VSS.n3019 22.2123
R6192 VSS.n3092 VSS.n3016 22.2123
R6193 VSS.n3212 VSS.n2973 22.2123
R6194 VSS.n1241 VSS.n1189 22.2123
R6195 VSS.n1215 VSS.n1214 22.2123
R6196 VSS.n1352 VSS.n1156 22.2123
R6197 VSS.n1468 VSS.n1467 22.2123
R6198 VSS.n4005 VSS.n4004 22.2123
R6199 VSS.n4010 VSS.n4009 22.2123
R6200 VSS.n4535 VSS.n4534 22.2123
R6201 VSS.n4534 VSS.n4533 22.2123
R6202 VSS.n4502 VSS.n3612 22.2123
R6203 VSS.n4502 VSS.n4501 22.2123
R6204 VSS.n4495 VSS.n4494 22.2123
R6205 VSS.n4494 VSS.n4493 22.2123
R6206 VSS.n4448 VSS.n4447 22.2123
R6207 VSS.n4447 VSS.n4446 22.2123
R6208 VSS.n4342 VSS.n4341 22.2123
R6209 VSS.n4341 VSS.n4340 22.2123
R6210 VSS.n3723 VSS.n3719 22.2123
R6211 VSS.n4600 VSS.n3572 22.2123
R6212 VSS.n4604 VSS.n3572 22.2123
R6213 VSS.n4607 VSS.n4605 22.2123
R6214 VSS.n4607 VSS.n3568 22.2123
R6215 VSS.n2710 VSS.n1948 21.8358
R6216 VSS.n3391 VSS.n2922 21.8358
R6217 VSS.n3356 VSS.n3355 21.8358
R6218 VSS.n3149 VSS.n3148 21.8358
R6219 VSS.n4384 VSS.n4383 21.8358
R6220 VSS.n2979 VSS.t5 21.795
R6221 VSS.n5373 VSS.n92 21.4593
R6222 VSS.n5312 VSS.n5311 21.4593
R6223 VSS.n5295 VSS.n5294 21.4593
R6224 VSS.n5264 VSS.n5263 21.4593
R6225 VSS.n5063 VSS.n5062 21.4593
R6226 VSS.n5033 VSS.n238 21.4593
R6227 VSS.n915 VSS.n914 21.4593
R6228 VSS.n910 VSS.n333 21.4593
R6229 VSS.n884 VSS.n350 21.4593
R6230 VSS.n883 VSS.n882 21.4593
R6231 VSS.n761 VSS.n448 21.4593
R6232 VSS.n734 VSS.n733 21.4593
R6233 VSS.n728 VSS.n464 21.4593
R6234 VSS.n718 VSS.n473 21.4593
R6235 VSS.n693 VSS.n692 21.4593
R6236 VSS.n675 VSS.n674 21.4593
R6237 VSS.n669 VSS.n498 21.4593
R6238 VSS.n646 VSS.n645 21.4593
R6239 VSS.n630 VSS.n524 21.4593
R6240 VSS.n596 VSS.n595 21.4593
R6241 VSS.n5472 VSS.n11 21.4593
R6242 VSS.n5463 VSS.n5462 21.4593
R6243 VSS.n2098 VSS.n2096 21.4593
R6244 VSS.n2106 VSS.n2104 21.4593
R6245 VSS.n2130 VSS.n2043 21.4593
R6246 VSS.n2189 VSS.n2142 21.4593
R6247 VSS.n2183 VSS.n2144 21.4593
R6248 VSS.n2207 VSS.n2040 21.4593
R6249 VSS.n2251 VSS.n2249 21.4593
R6250 VSS.n2318 VSS.n2270 21.4593
R6251 VSS.n2442 VSS.n2441 21.4593
R6252 VSS.n2512 VSS.n2511 21.4593
R6253 VSS.n2521 VSS.n2519 21.4593
R6254 VSS.n2709 VSS.n2708 21.4593
R6255 VSS.n2679 VSS.n2678 21.4593
R6256 VSS.n2856 VSS.n2791 21.4593
R6257 VSS.n3488 VSS.n2774 21.4593
R6258 VSS.n3436 VSS.n3435 21.4593
R6259 VSS.n3429 VSS.n2906 21.4593
R6260 VSS.n3374 VSS.n2927 21.4593
R6261 VSS.n3366 VSS.n3365 21.4593
R6262 VSS.n3344 VSS.n3343 21.4593
R6263 VSS.n3169 VSS.n3167 21.4593
R6264 VSS.n3200 VSS.n3198 21.4593
R6265 VSS.n3278 VSS.n3277 21.4593
R6266 VSS.n1256 VSS.n1255 21.4593
R6267 VSS.n1422 VSS.n1421 21.4593
R6268 VSS.n1419 VSS.n1389 21.4593
R6269 VSS.n1451 VSS.n1142 21.4593
R6270 VSS.n1457 VSS.n1140 21.4593
R6271 VSS.n1543 VSS.n1542 21.4593
R6272 VSS.n1524 VSS.n1516 21.4593
R6273 VSS.n1586 VSS.n1110 21.4593
R6274 VSS.n1594 VSS.n1106 21.4593
R6275 VSS.n1600 VSS.n1104 21.4593
R6276 VSS.n1088 VSS.n1032 21.4593
R6277 VSS.n1080 VSS.n1035 21.4593
R6278 VSS.n1052 VSS.n1025 21.4593
R6279 VSS.n1642 VSS.n1640 21.4593
R6280 VSS.n4465 VSS.n4464 21.4593
R6281 VSS.n4436 VSS.n4435 21.4593
R6282 VSS.n4403 VSS.n4402 21.4593
R6283 VSS.n4353 VSS.n4352 21.4593
R6284 VSS.n4317 VSS.n4316 21.4593
R6285 VSS.n4565 VSS.n3583 21.4593
R6286 VSS.n4625 VSS.n4623 21.4593
R6287 VSS.n4663 VSS.n1920 21.4593
R6288 VSS.n4898 VSS.n4896 21.3456
R6289 VSS.n853 VSS.n852 21.0829
R6290 VSS.n2130 VSS.n2129 21.0829
R6291 VSS.n2466 VSS.n2465 21.0829
R6292 VSS.n2547 VSS.n2546 21.0829
R6293 VSS.n4756 VSS.n4736 21.0829
R6294 VSS.n4103 VSS.n4087 21.0829
R6295 VSS.n4792 VSS.n4789 21.0829
R6296 VSS.n852 VSS.n851 20.7064
R6297 VSS.n846 VSS.n845 20.7064
R6298 VSS.n668 VSS.n667 20.7064
R6299 VSS.n2213 VSS.n2038 20.7064
R6300 VSS.n2216 VSS.n2035 20.7064
R6301 VSS.n2436 VSS.n2411 20.7064
R6302 VSS.n2621 VSS.n2620 20.7064
R6303 VSS.n3094 VSS.n3014 20.7064
R6304 VSS.n1249 VSS.n1248 20.7064
R6305 VSS.n1359 VSS.n1155 20.7064
R6306 VSS.n1485 VSS.n1484 20.7064
R6307 VSS.n1491 VSS.n1489 20.7064
R6308 VSS.t728 VSS.n3605 20.6942
R6309 VSS.n4962 VSS.n4961 20.4554
R6310 VSS.n2384 VSS.n2383 20.4554
R6311 VSS.n896 VSS.n895 20.3299
R6312 VSS.n745 VSS.n455 20.3299
R6313 VSS.n653 VSS.n652 20.3299
R6314 VSS.n2099 VSS.n2052 20.3299
R6315 VSS.n2112 VSS.n2111 20.3299
R6316 VSS.n2539 VSS.n2538 20.3299
R6317 VSS.n1321 VSS.n1320 20.3299
R6318 VSS.n1403 VSS.n1402 20.3299
R6319 VSS.n1658 VSS.n1657 20.3299
R6320 VSS.n1682 VSS.n1001 20.3299
R6321 VSS.n1690 VSS.n996 20.3299
R6322 VSS.n1764 VSS.n1763 20.3039
R6323 VSS.n4890 VSS.n4889 20.3039
R6324 VSS.n4124 VSS.n4121 20.3039
R6325 VSS.n4119 VSS.n4116 20.3039
R6326 VSS.n2456 VSS.n2455 20.0859
R6327 VSS.n51 VSS.n41 19.9534
R6328 VSS.n5350 VSS.n101 19.9534
R6329 VSS.n5317 VSS.n115 19.9534
R6330 VSS.n5269 VSS.n136 19.9534
R6331 VSS.n5238 VSS.n146 19.9534
R6332 VSS.n5211 VSS.n162 19.9534
R6333 VSS.n5174 VSS.n176 19.9534
R6334 VSS.n5126 VSS.n5125 19.9534
R6335 VSS.n5030 VSS.n5029 19.9534
R6336 VSS.n5019 VSS.n247 19.9534
R6337 VSS.n857 VSS.n856 19.9534
R6338 VSS.n779 VSS.n778 19.9534
R6339 VSS.n741 VSS.n740 19.9534
R6340 VSS.n641 VSS.n514 19.9534
R6341 VSS.n614 VSS.n613 19.9534
R6342 VSS.n611 VSS.n536 19.9534
R6343 VSS.n5422 VSS.n5392 19.9534
R6344 VSS.n2575 VSS.n1958 19.9534
R6345 VSS.n1208 VSS.n1207 19.9534
R6346 VSS.n1537 VSS.n1536 19.9534
R6347 VSS.n1522 VSS.n1519 19.9534
R6348 VSS.n1620 VSS.n1029 19.9534
R6349 VSS.n1067 VSS.n1064 19.9534
R6350 VSS.n1629 VSS.n1628 19.9534
R6351 VSS.n4755 VSS.n4752 19.9534
R6352 VSS.n4102 VSS.n4101 19.9534
R6353 VSS.n4785 VSS.n4771 19.9534
R6354 VSS.n4327 VSS.n3698 19.9534
R6355 VSS.n4323 VSS.n4322 19.9534
R6356 VSS.n3803 VSS.n3793 19.9534
R6357 VSS.n4723 VSS.n4722 19.9534
R6358 VSS.n4886 VSS.n4885 19.8626
R6359 VSS.n4127 VSS.n4126 19.8626
R6360 VSS.t2636 VSS.n3586 19.6373
R6361 VSS.t2633 VSS.t376 19.6373
R6362 VSS.n60 VSS.n36 19.577
R6363 VSS.n66 VSS.n33 19.577
R6364 VSS.n5069 VSS.n223 19.577
R6365 VSS.n5010 VSS.n255 19.577
R6366 VSS.n4943 VSS.n4942 19.577
R6367 VSS.n4931 VSS.n4930 19.577
R6368 VSS.n295 VSS.n289 19.577
R6369 VSS.n855 VSS.n854 19.577
R6370 VSS.n5415 VSS.n5399 19.577
R6371 VSS.n5409 VSS.n5403 19.577
R6372 VSS.n2079 VSS.n2060 19.577
R6373 VSS.n2071 VSS.n2065 19.577
R6374 VSS.n2289 VSS.n2279 19.577
R6375 VSS.n2370 VSS.n2369 19.577
R6376 VSS.n2665 VSS.n2664 19.577
R6377 VSS.n3050 VSS.n3032 19.577
R6378 VSS.n3043 VSS.n3037 19.577
R6379 VSS.n2816 VSS.n2813 19.577
R6380 VSS.n2870 VSS.n2869 19.577
R6381 VSS.n3360 VSS.n2938 19.577
R6382 VSS.n3056 VSS.n3029 19.577
R6383 VSS.n3062 VSS.n3025 19.577
R6384 VSS.n3068 VSS.n3066 19.577
R6385 VSS.n3069 VSS.n3022 19.577
R6386 VSS.n3075 VSS.n3074 19.577
R6387 VSS.n1370 VSS.n1369 19.577
R6388 VSS.n1094 VSS.n1028 19.577
R6389 VSS.n1688 VSS.n999 19.577
R6390 VSS.n1713 VSS.n1712 19.577
R6391 VSS.n969 VSS.n963 19.577
R6392 VSS.n1291 VSS.n1290 19.577
R6393 VSS.n1284 VSS.n1278 19.577
R6394 VSS.n4540 VSS.n4539 19.577
R6395 VSS.n4515 VSS.n3608 19.577
R6396 VSS.n4489 VSS.n4488 19.577
R6397 VSS.n4454 VSS.n3636 19.577
R6398 VSS.n4424 VSS.n3649 19.577
R6399 VSS.n4396 VSS.n3665 19.577
R6400 VSS.n4348 VSS.n4347 19.577
R6401 VSS.n4314 VSS.n3705 19.577
R6402 VSS.n4308 VSS.n4307 19.577
R6403 VSS.n3745 VSS.n3743 19.577
R6404 VSS.n3757 VSS.n3755 19.577
R6405 VSS.n4593 VSS.n4591 19.577
R6406 VSS.n4617 VSS.n3566 19.577
R6407 VSS.n4633 VSS.n1926 19.577
R6408 VSS.n4650 VSS.n1924 19.577
R6409 VSS.n4728 VSS.n4669 19.577
R6410 VSS.n4712 VSS.n4675 19.577
R6411 VSS.n4706 VSS.n4678 19.577
R6412 VSS.n4700 VSS.n4681 19.577
R6413 VSS.n4694 VSS.n4684 19.577
R6414 VSS.n4174 VSS.n3932 19.5165
R6415 VSS.n4886 VSS.n1728 19.4212
R6416 VSS.n4126 VSS.n4125 19.4212
R6417 VSS.n47 VSS.n41 19.3355
R6418 VSS.n5334 VSS.n101 19.3355
R6419 VSS.n5329 VSS.n109 19.3355
R6420 VSS.n5242 VSS.n146 19.3355
R6421 VSS.n5125 VSS.n5124 19.3355
R6422 VSS.n3799 VSS.n3793 19.3355
R6423 VSS.n3094 VSS.n3093 19.2005
R6424 VSS.n1764 VSS.n1726 18.9798
R6425 VSS.n3088 VSS.n3087 18.9221
R6426 VSS.n5225 VSS.n5224 18.824
R6427 VSS.n835 VSS.n386 18.824
R6428 VSS.n587 VSS.n549 18.824
R6429 VSS.n5447 VSS.n5379 18.824
R6430 VSS.n2208 VSS.n2207 18.824
R6431 VSS.n2481 VSS.n2480 18.824
R6432 VSS.n2633 VSS.n1952 18.824
R6433 VSS.n2607 VSS.n1938 18.824
R6434 VSS.n2716 VSS.n2715 18.824
R6435 VSS.n2876 VSS.n2875 18.824
R6436 VSS.n3385 VSS.n3384 18.824
R6437 VSS.n3347 VSS.n2944 18.824
R6438 VSS.n3143 VSS.n3142 18.824
R6439 VSS.n3290 VSS.n3220 18.824
R6440 VSS.n3284 VSS.n3224 18.824
R6441 VSS.n1256 VSS.n1176 18.824
R6442 VSS.n1536 VSS.n1535 18.824
R6443 VSS.n4389 VSS.n3670 18.824
R6444 VSS.n4120 VSS.n4119 18.7591
R6445 VSS.n5462 VSS.n5461 18.7296
R6446 VSS.n786 VSS.n785 18.4476
R6447 VSS.n2352 VSS.n2351 18.4476
R6448 VSS.n2465 VSS.n2397 18.4476
R6449 VSS.n1427 VSS.n1384 18.4476
R6450 VSS.n1861 VSS.n1860 18.2129
R6451 VSS.n827 VSS.n826 18.1632
R6452 VSS.n3997 VSS.n3996 18.0884
R6453 VSS.n4999 VSS.n4998 18.0711
R6454 VSS.n425 VSS.n424 18.0711
R6455 VSS.n590 VSS.n589 18.0711
R6456 VSS.n2106 VSS.n2050 18.0711
R6457 VSS.n2345 VSS.n2011 18.0711
R6458 VSS.n2544 VSS.n1968 18.0711
R6459 VSS.n2585 VSS.n2583 18.0711
R6460 VSS.n1340 VSS.n1164 18.0711
R6461 VSS.n1442 VSS.n1376 18.0711
R6462 VSS.n1550 VSS.n1502 18.0711
R6463 VSS.n1542 VSS.n1541 18.0711
R6464 VSS.n1524 VSS.n1523 18.0711
R6465 VSS.n1573 VSS.n1115 18.0711
R6466 VSS.n4317 VSS.n3700 18.0711
R6467 VSS.n4036 VSS.t1836 17.9597
R6468 VSS.n4843 VSS.n4842 17.9205
R6469 VSS.n4137 VSS.n4112 17.9205
R6470 VSS.n2551 VSS.n1966 17.9177
R6471 VSS.n1575 VSS.n1574 17.7867
R6472 VSS.n5039 VSS.n236 17.6946
R6473 VSS.n735 VSS.n734 17.6946
R6474 VSS.n712 VSS.n476 17.6946
R6475 VSS.n2122 VSS.n2045 17.6946
R6476 VSS.n2170 VSS.n2169 17.6946
R6477 VSS.n2696 VSS.n2695 17.6946
R6478 VSS.n2796 VSS.n2793 17.6946
R6479 VSS.n3400 VSS.n3399 17.6946
R6480 VSS.n3362 VSS.n2935 17.6946
R6481 VSS.n3338 VSS.n2952 17.6946
R6482 VSS.n3118 VSS.n3005 17.6946
R6483 VSS.n3162 VSS.n3160 17.6946
R6484 VSS.n3272 VSS.n3232 17.6946
R6485 VSS.n1413 VSS.n1392 17.6946
R6486 VSS.n4376 VSS.n3676 17.6946
R6487 VSS.n5313 VSS.n115 17.3181
R6488 VSS.n5265 VSS.n136 17.3181
R6489 VSS.n5031 VSS.n5030 17.3181
R6490 VSS.n765 VSS.n764 17.3181
R6491 VSS.n2220 VSS.n2035 17.3181
R6492 VSS.n3533 VSS.n2751 17.3181
R6493 VSS.n1569 VSS.n1115 17.3181
R6494 VSS.n4011 VSS.n4010 17.3181
R6495 VSS.n3887 VSS.n3879 17.1349
R6496 VSS.n4295 VSS.n3879 17.119
R6497 VSS.n1840 VSS.n1838 17.1007
R6498 VSS.n4842 VSS.n4841 17.0672
R6499 VSS.n4142 VSS.n4112 17.0672
R6500 VSS.n575 VSS.n574 16.9417
R6501 VSS.n2120 VSS.n2119 16.9417
R6502 VSS.n2890 VSS.n2889 16.9417
R6503 VSS.n3131 VSS.n2999 16.9417
R6504 VSS.n1247 VSS.n1186 16.9417
R6505 VSS.n1242 VSS.n1241 16.9417
R6506 VSS.n1359 VSS.n1358 16.9417
R6507 VSS.n1529 VSS.n1528 16.9417
R6508 VSS.n1606 VSS.n1101 16.9417
R6509 VSS.n1073 VSS.n1041 16.9417
R6510 VSS.n1059 VSS.n1046 16.9417
R6511 VSS.n1635 VSS.n1633 16.9417
R6512 VSS.n4762 VSS.n4761 16.9417
R6513 VSS.n4109 VSS.n4108 16.9417
R6514 VSS.n4797 VSS.n1777 16.9417
R6515 VSS.n4334 VSS.n4333 16.9417
R6516 VSS.n4623 VSS.n3563 16.9417
R6517 VSS.t1327 VSS.t2089 16.8587
R6518 VSS.t348 VSS.t2896 16.8587
R6519 VSS.t41 VSS.t3533 16.8587
R6520 VSS.t1586 VSS.t820 16.8587
R6521 VSS.t156 VSS.t353 16.8587
R6522 VSS.t1301 VSS.t3141 16.8587
R6523 VSS.t3216 VSS.t2910 16.8587
R6524 VSS.t1699 VSS.n492 16.8587
R6525 VSS.t997 VSS.t1656 16.8587
R6526 VSS.n4172 VSS.t1805 16.7248
R6527 VSS.n5032 VSS.n5031 16.5652
R6528 VSS.n2099 VSS.n2098 16.5652
R6529 VSS.n3425 VSS.n3424 16.5652
R6530 VSS.n3208 VSS.n3206 16.5652
R6531 VSS.n1079 VSS.n1078 16.5652
R6532 VSS.n1860 VSS.n1859 16.5652
R6533 VSS.n4748 VSS.n4747 16.5652
R6534 VSS.n4761 VSS.n4760 16.5652
R6535 VSS.n4108 VSS.n4107 16.5652
R6536 VSS.n4097 VSS.n4096 16.5652
R6537 VSS.n4783 VSS.n4773 16.5652
R6538 VSS.n4793 VSS.n1777 16.5652
R6539 VSS.n1832 VSS.n1831 16.3238
R6540 VSS.n5097 VSS.n5096 16.1887
R6541 VSS.n845 VSS.n379 16.1887
R6542 VSS.n2209 VSS.n2208 16.1887
R6543 VSS.n2455 VSS.n2454 16.1887
R6544 VSS.n2435 VSS.n2434 16.1887
R6545 VSS.n2518 VSS.n2516 16.1887
R6546 VSS.n2614 VSS.n2611 16.1887
R6547 VSS.n3487 VSS.n3486 16.1887
R6548 VSS.n1492 VSS.n1120 16.1887
R6549 VSS.n4273 VSS.n4272 16.1856
R6550 VSS.n4269 VSS.n4249 16.1856
R6551 VSS.n4249 VSS.n3907 16.1856
R6552 VSS.n4270 VSS.n4269 16.1529
R6553 VSS.n4175 VSS.n4174 16.126
R6554 VSS.n4272 VSS.n4271 16.0673
R6555 VSS.n3098 VSS.n3014 16.0566
R6556 VSS.t2140 VSS.n3812 15.8945
R6557 VSS.n5374 VSS.n25 15.8123
R6558 VSS.n5104 VSS.n5103 15.8123
R6559 VSS.n793 VSS.n425 15.8123
R6560 VSS.n624 VSS.n527 15.8123
R6561 VSS.n584 VSS.n549 15.8123
R6562 VSS.n2204 VSS.n2203 15.8123
R6563 VSS.n2480 VSS.n2479 15.8123
R6564 VSS.n2630 VSS.n1952 15.8123
R6565 VSS.n2715 VSS.n2714 15.8123
R6566 VSS.n2877 VSS.n2876 15.8123
R6567 VSS.n3437 VSS.n2900 15.8123
R6568 VSS.n3386 VSS.n3385 15.8123
R6569 VSS.n3348 VSS.n3347 15.8123
R6570 VSS.n3093 VSS.n3092 15.8123
R6571 VSS.n3115 VSS.n3007 15.8123
R6572 VSS.n3144 VSS.n3143 15.8123
R6573 VSS.n3287 VSS.n3220 15.8123
R6574 VSS.n3281 VSS.n3224 15.8123
R6575 VSS.n1326 VSS.n1176 15.8123
R6576 VSS.n1214 VSS.n1213 15.8123
R6577 VSS.n1421 VSS.n1420 15.8123
R6578 VSS.n4386 VSS.n3670 15.8123
R6579 VSS.n486 VSS.n484 15.6771
R6580 VSS.n2461 VSS.n2397 15.6589
R6581 VSS.n3299 VSS.n2967 15.5708
R6582 VSS.n785 VSS.n784 15.4358
R6583 VSS.n589 VSS.n588 15.4358
R6584 VSS.n2193 VSS.n2142 15.4358
R6585 VSS.n2589 VSS.n2585 15.4358
R6586 VSS.n4164 VSS.n4163 15.4358
R6587 VSS.n1351 VSS.n1350 15.3347
R6588 VSS.n4198 VSS.n4197 15.2301
R6589 VSS.n4929 VSS.n4928 15.1944
R6590 VSS.n4693 VSS.n4692 15.1944
R6591 VSS.n4514 VSS.n4513 15.1514
R6592 VSS.n386 VSS.n383 15.0593
R6593 VSS.n415 VSS.n414 15.0593
R6594 VSS.n720 VSS.n719 15.0593
R6595 VSS.n2371 VSS.n2370 15.0593
R6596 VSS.n2540 VSS.n2539 15.0593
R6597 VSS.n2540 VSS.n1968 15.0593
R6598 VSS.n3074 VSS.n3022 15.0593
R6599 VSS.n3152 VSS.n3151 15.0593
R6600 VSS.n3292 VSS.n3291 15.0593
R6601 VSS.n3295 VSS.n2969 15.0593
R6602 VSS.n5118 VSS.n5117 14.8179
R6603 VSS.n5075 VSS.n5074 14.8179
R6604 VSS.n956 VSS.n284 14.8179
R6605 VSS.n638 VSS.n637 14.8179
R6606 VSS.n1717 VSS.n959 14.8179
R6607 VSS.n2293 VSS.n2279 14.775
R6608 VSS.n3406 VSS.n2915 14.775
R6609 VSS.n1231 VSS.n1189 14.775
R6610 VSS.n4245 VSS.n4212 14.7155
R6611 VSS.n4246 VSS.n4245 14.7155
R6612 VSS.n5092 VSS.n211 14.6829
R6613 VSS.n5057 VSS.n228 14.6829
R6614 VSS.n888 VSS.n350 14.6829
R6615 VSS.n766 VSS.n765 14.6829
R6616 VSS.n645 VSS.n514 14.6829
R6617 VSS.n603 VSS.n538 14.6829
R6618 VSS.n2188 VSS.n2187 14.6829
R6619 VSS.n2681 VSS.n2646 14.6829
R6620 VSS.n2678 VSS.n2650 14.6829
R6621 VSS.n2832 VSS.n2799 14.6829
R6622 VSS.n3380 VSS.n2925 14.6829
R6623 VSS.n3279 VSS.n3278 14.6829
R6624 VSS.n1078 VSS.n1077 14.6829
R6625 VSS.n1683 VSS.n1682 14.6829
R6626 VSS.n4358 VSS.n3683 14.6829
R6627 VSS.n3994 VSS.t2435 14.4705
R6628 VSS.n654 VSS.n653 14.3064
R6629 VSS.n2534 VSS.n1970 14.3064
R6630 VSS.n2538 VSS.n1970 14.3064
R6631 VSS.n1678 VSS.n1001 14.3064
R6632 VSS.n1693 VSS.n996 14.3064
R6633 VSS.n4762 VSS.n1918 14.3064
R6634 VSS.n4109 VSS.n4083 14.3064
R6635 VSS.n4797 VSS.n1776 14.3064
R6636 VSS.n4528 VSS.n4527 14.3064
R6637 VSS.n414 VSS.n410 14.3064
R6638 VSS.n615 VSS.n614 14.3064
R6639 VSS.n1404 VSS.n1403 14.3064
R6640 VSS.n1659 VSS.n1658 14.3064
R6641 VSS.n4903 VSS.n4902 14.2403
R6642 VSS.n3108 VSS.n3009 14.2278
R6643 VSS.n4991 VSS.n4990 14.0717
R6644 VSS.n3308 VSS.n2963 14.022
R6645 VSS.n2083 VSS.n2060 13.9299
R6646 VSS.n2129 VSS.n2127 13.9299
R6647 VSS.n2171 VSS.n2152 13.9299
R6648 VSS.n2223 VSS.n2222 13.9299
R6649 VSS.n2345 VSS.n2343 13.9299
R6650 VSS.n2384 VSS.n1999 13.9299
R6651 VSS.n2439 VSS.n2411 13.9299
R6652 VSS.n2532 VSS.n1972 13.9299
R6653 VSS.n2546 VSS.n2544 13.9299
R6654 VSS.n3054 VSS.n3032 13.9299
R6655 VSS.n3111 VSS.n3109 13.9299
R6656 VSS.n3137 VSS.n2997 13.9299
R6657 VSS.n1322 VSS.n1321 13.9299
R6658 VSS.n1613 VSS.n1099 13.9299
R6659 VSS.n1624 VSS.n1028 13.9299
R6660 VSS.n4323 VSS.n3698 13.9299
R6661 VSS.n4194 VSS.t86 13.684
R6662 VSS.n727 VSS.n726 13.5534
R6663 VSS.n582 VSS.n581 13.5534
R6664 VSS.n2487 VSS.n2486 13.5534
R6665 VSS.n3292 VSS.n2970 13.5534
R6666 VSS.n3295 VSS.n2967 13.5534
R6667 VSS.n1676 VSS.n1675 13.5534
R6668 VSS.n3811 VSS.n3729 13.5534
R6669 VSS.n4655 VSS.n4654 13.5534
R6670 VSS.n5449 VSS.n23 13.417
R6671 VSS.n4941 VSS.n4915 13.177
R6672 VSS.n956 VSS.n285 13.177
R6673 VSS.n952 VSS.n285 13.177
R6674 VSS.n856 VSS.n855 13.177
R6675 VSS.n639 VSS.n638 13.177
R6676 VSS.n2084 VSS.n2083 13.177
R6677 VSS.n2086 VSS.n2084 13.177
R6678 VSS.n3548 VSS.n3547 13.177
R6679 VSS.n3402 VSS.n2915 13.177
R6680 VSS.n3055 VSS.n3054 13.177
R6681 VSS.n1155 VSS.n1154 13.177
R6682 VSS.n1569 VSS.n1118 13.177
R6683 VSS.n1717 VSS.n958 13.177
R6684 VSS.n4473 VSS.n4472 13.177
R6685 VSS.n4303 VSS.n3709 13.177
R6686 VSS.n4730 VSS.n4729 13.177
R6687 VSS.t3187 VSS.t728 12.9341
R6688 VSS.t1507 VSS.t1055 12.9341
R6689 VSS.n4267 VSS.n3586 12.866
R6690 VSS.t376 VSS.n4260 12.866
R6691 VSS.n4819 VSS.n1773 12.8005
R6692 VSS.n3843 VSS.n3824 12.8005
R6693 VSS.n5117 VSS.n5116 12.8005
R6694 VSS.n897 VSS.n896 12.8005
R6695 VSS.n457 VSS.n455 12.8005
R6696 VSS.n583 VSS.n582 12.8005
R6697 VSS.n2343 VSS.n2342 12.8005
R6698 VSS.n2430 VSS.n2429 12.8005
R6699 VSS.n1948 VSS.n1945 12.8005
R6700 VSS.n3388 VSS.n2922 12.8005
R6701 VSS.n3355 VSS.n3354 12.8005
R6702 VSS.n3346 VSS.n3345 12.8005
R6703 VSS.n3148 VSS.n3147 12.8005
R6704 VSS.n3151 VSS.n2990 12.8005
R6705 VSS.n3206 VSS.n3205 12.8005
R6706 VSS.n3280 VSS.n3279 12.8005
R6707 VSS.n1365 VSS.n1147 12.8005
R6708 VSS.n1613 VSS.n1612 12.8005
R6709 VSS.n1628 VSS.n1627 12.8005
R6710 VSS.n4385 VSS.n4384 12.8005
R6711 VSS.n3727 VSS.n3719 12.8005
R6712 VSS.n3716 VSS.n3715 12.8005
R6713 VSS.n2314 VSS.n2270 12.6471
R6714 VSS.n4818 VSS.n1775 12.561
R6715 VSS.n3845 VSS.n3844 12.56
R6716 VSS.n826 VSS.n825 12.424
R6717 VSS.n640 VSS.n639 12.424
R6718 VSS.n5421 VSS.n5420 12.424
R6719 VSS.n2113 VSS.n2112 12.424
R6720 VSS.n2203 VSS.n2202 12.424
R6721 VSS.n2289 VSS.n2288 12.424
R6722 VSS.n3109 VSS.n3108 12.424
R6723 VSS.n1369 VSS.n1147 12.424
R6724 VSS.n1644 VSS.n1642 12.424
R6725 VSS.n2420 VSS.n1994 12.3195
R6726 VSS.n4253 VSS.n4203 12.1744
R6727 VSS.n4183 VSS.n3926 12.1636
R6728 VSS.n825 VSS.n824 12.0476
R6729 VSS.n764 VSS.n763 12.0476
R6730 VSS.n2373 VSS.n2001 12.0476
R6731 VSS.n2616 VSS.n2615 12.0476
R6732 VSS.n2611 VSS.n2610 12.0476
R6733 VSS.n2871 VSS.n2862 12.0476
R6734 VSS.n3245 VSS.n2969 12.0476
R6735 VSS.n1329 VSS.n1174 12.0476
R6736 VSS.n1479 VSS.n1126 12.0476
R6737 VSS.n1644 VSS.n1017 12.0476
R6738 VSS.n4255 VSS.n4253 11.9432
R6739 VSS.n5359 VSS.n5358 11.7085
R6740 VSS.n5301 VSS.n5300 11.7085
R6741 VSS.n5284 VSS.n5283 11.7085
R6742 VSS.n5253 VSS.n5252 11.7085
R6743 VSS.n928 VSS.n326 11.7085
R6744 VSS.n752 VSS.n751 11.7085
R6745 VSS.n707 VSS.n478 11.7085
R6746 VSS.n568 VSS.n567 11.7085
R6747 VSS.n2723 VSS.n1943 11.7085
R6748 VSS.n3474 VSS.n2784 11.7085
R6749 VSS.n1462 VSS.n1461 11.7085
R6750 VSS.n841 VSS.n840 11.6711
R6751 VSS.n2511 VSS.n2509 11.6711
R6752 VSS.n2628 VSS.n2627 11.6711
R6753 VSS.n1208 VSS.n1202 11.6711
R6754 VSS.n939 VSS.n320 11.5456
R6755 VSS.n1898 VSS.n1897 11.4713
R6756 VSS.n1793 VSS.n1792 11.4713
R6757 VSS.n2234 VSS.n2233 11.2946
R6758 VSS.n2430 VSS.n2414 11.2946
R6759 VSS.n3425 VSS.n2906 11.2946
R6760 VSS.n1206 VSS.n1174 11.2946
R6761 VSS.n1678 VSS.n1676 11.2946
R6762 VSS.n2375 VSS.n2373 11.0436
R6763 VSS.n4844 VSS.n4843 11.0072
R6764 VSS.n4138 VSS.n4137 11.0072
R6765 VSS.n787 VSS.n427 10.9181
R6766 VSS.n2177 VSS.n2176 10.9181
R6767 VSS.n2215 VSS.n2213 10.9181
R6768 VSS.n3548 VSS.n2749 10.9181
R6769 VSS.n3431 VSS.n2903 10.9181
R6770 VSS.n3402 VSS.n3401 10.9181
R6771 VSS.n3353 VSS.n3352 10.9181
R6772 VSS.n3141 VSS.n2997 10.9181
R6773 VSS.n3178 VSS.n3177 10.9181
R6774 VSS.n1415 VSS.n1414 10.9181
R6775 VSS.n4472 VSS.n4471 10.9181
R6776 VSS.n4442 VSS.n3641 10.9181
R6777 VSS.n4410 VSS.n4409 10.9181
R6778 VSS.n4575 VSS.n3580 10.9181
R6779 VSS.n4656 VSS.n4655 10.9181
R6780 VSS.t87 VSS.n3927 10.6432
R6781 VSS.n4900 VSS.n4899 10.5934
R6782 VSS.n862 VSS.n861 10.5417
R6783 VSS.n574 VSS.n573 10.5417
R6784 VSS.n2442 VSS.n2406 10.5417
R6785 VSS.n3437 VSS.n3436 10.5417
R6786 VSS.n4902 VSS.n4901 10.5417
R6787 VSS.n2730 VSS.n1938 10.5417
R6788 VSS.n3712 VSS.n1720 10.4684
R6789 VSS.n3892 VSS.t2106 10.4216
R6790 VSS.n3892 VSS.t2108 10.4216
R6791 VSS.n1825 VSS.n1824 10.4058
R6792 VSS.n1899 VSS.n1898 10.4058
R6793 VSS.n4062 VSS.n4061 10.4058
R6794 VSS.n1793 VSS.n1791 10.4058
R6795 VSS.n3890 VSS.t1547 10.219
R6796 VSS.n847 VSS.n846 10.1652
R6797 VSS.n787 VSS.n786 10.1652
R6798 VSS.n726 VSS.n725 10.1652
R6799 VSS.n667 VSS.n666 10.1652
R6800 VSS.n3345 VSS.n3344 10.1652
R6801 VSS.n1248 VSS.n1247 10.1652
R6802 VSS.n1636 VSS.n1635 10.1652
R6803 VSS.n4958 VSS.n276 10.0265
R6804 VSS.n544 VSS.n541 10.0265
R6805 VSS.n2390 VSS.n2388 10.0265
R6806 VSS.n43 VSS.n42 9.83768
R6807 VSS.n4926 VSS.n4923 9.83768
R6808 VSS.n3795 VSS.n3794 9.83768
R6809 VSS.n4690 VSS.n4687 9.83768
R6810 VSS.n781 VSS.n431 9.78874
R6811 VSS.n621 VSS.n530 9.78874
R6812 VSS.n5444 VSS.n5382 9.78874
R6813 VSS.n2330 VSS.n2329 9.78874
R6814 VSS.n2528 VSS.n1972 9.78874
R6815 VSS.n3533 VSS.n3532 9.78874
R6816 VSS.n3532 VSS.n3531 9.78874
R6817 VSS.n1519 VSS.n1118 9.78874
R6818 VSS.n1010 VSS.n1007 9.78874
R6819 VSS.n3101 VSS.n3100 9.61041
R6820 VSS.n4899 VSS.n4898 9.48661
R6821 VSS.n4907 VSS.n4900 9.41378
R6822 VSS.n5201 VSS.n5200 9.41227
R6823 VSS.n5163 VSS.n179 9.41227
R6824 VSS.n5137 VSS.n5136 9.41227
R6825 VSS.n2624 VSS.n2623 9.41227
R6826 VSS.n1942 VSS.n1939 9.41227
R6827 VSS.n3329 VSS.n2956 9.41227
R6828 VSS.n3285 VSS.n3284 9.41227
R6829 VSS.n1429 VSS.n1428 9.41227
R6830 VSS.n1405 VSS.n1395 9.41227
R6831 VSS.n1636 VSS.n1020 9.41227
R6832 VSS.n1907 VSS.n1906 9.41227
R6833 VSS.n4070 VSS.n4069 9.41227
R6834 VSS.n1803 VSS.n1802 9.41227
R6835 VSS.n4546 VSS.n4545 9.41227
R6836 VSS.n4478 VSS.n4477 9.41227
R6837 VSS.n4418 VSS.n4417 9.41227
R6838 VSS.n3771 VSS.n3770 9.41227
R6839 VSS.n3734 VSS.n3731 9.41227
R6840 VSS.n4586 VSS.n4585 9.41227
R6841 VSS.n4165 VSS.n3934 9.41227
R6842 VSS.n3716 VSS.n3712 9.32264
R6843 VSS.n4842 VSS.n4834 9.3005
R6844 VSS.n1765 VSS.n1764 9.3005
R6845 VSS.n4890 VSS.n1727 9.3005
R6846 VSS.n4889 VSS.n4888 9.3005
R6847 VSS.n4887 VSS.n4886 9.3005
R6848 VSS.n4884 VSS.n1729 9.3005
R6849 VSS.n4926 VSS.n4925 9.3005
R6850 VSS.n4928 VSS.n4927 9.3005
R6851 VSS.n4929 VSS.n4921 9.3005
R6852 VSS.n4930 VSS.n4919 9.3005
R6853 VSS.n4932 VSS.n4931 9.3005
R6854 VSS.n4933 VSS.n4918 9.3005
R6855 VSS.n4935 VSS.n4934 9.3005
R6856 VSS.n4936 VSS.n4916 9.3005
R6857 VSS.n4938 VSS.n4937 9.3005
R6858 VSS.n4941 VSS.n4940 9.3005
R6859 VSS.n4942 VSS.n282 9.3005
R6860 VSS.n4944 VSS.n4943 9.3005
R6861 VSS.n4945 VSS.n281 9.3005
R6862 VSS.n4947 VSS.n4946 9.3005
R6863 VSS.n4948 VSS.n280 9.3005
R6864 VSS.n4950 VSS.n4949 9.3005
R6865 VSS.n4951 VSS.n279 9.3005
R6866 VSS.n4953 VSS.n4952 9.3005
R6867 VSS.n4954 VSS.n277 9.3005
R6868 VSS.n4956 VSS.n4955 9.3005
R6869 VSS.n4958 VSS.n4957 9.3005
R6870 VSS.n4959 VSS.n274 9.3005
R6871 VSS.n4963 VSS.n4962 9.3005
R6872 VSS.n4964 VSS.n273 9.3005
R6873 VSS.n4966 VSS.n4965 9.3005
R6874 VSS.n4967 VSS.n272 9.3005
R6875 VSS.n4971 VSS.n4970 9.3005
R6876 VSS.n4972 VSS.n271 9.3005
R6877 VSS.n4974 VSS.n4973 9.3005
R6878 VSS.n4976 VSS.n270 9.3005
R6879 VSS.n4978 VSS.n4977 9.3005
R6880 VSS.n4979 VSS.n269 9.3005
R6881 VSS.n4981 VSS.n4980 9.3005
R6882 VSS.n4982 VSS.n267 9.3005
R6883 VSS.n4988 VSS.n4987 9.3005
R6884 VSS.n4990 VSS.n4989 9.3005
R6885 VSS.n4991 VSS.n264 9.3005
R6886 VSS.n4992 VSS.n262 9.3005
R6887 VSS.n4994 VSS.n4993 9.3005
R6888 VSS.n4995 VSS.n261 9.3005
R6889 VSS.n4997 VSS.n4996 9.3005
R6890 VSS.n4998 VSS.n259 9.3005
R6891 VSS.n4999 VSS.n258 9.3005
R6892 VSS.n5001 VSS.n5000 9.3005
R6893 VSS.n5002 VSS.n257 9.3005
R6894 VSS.n5004 VSS.n5003 9.3005
R6895 VSS.n5005 VSS.n256 9.3005
R6896 VSS.n5007 VSS.n5006 9.3005
R6897 VSS.n5008 VSS.n255 9.3005
R6898 VSS.n5010 VSS.n5009 9.3005
R6899 VSS.n5011 VSS.n253 9.3005
R6900 VSS.n5012 VSS.n252 9.3005
R6901 VSS.n5014 VSS.n5013 9.3005
R6902 VSS.n5015 VSS.n251 9.3005
R6903 VSS.n5017 VSS.n5016 9.3005
R6904 VSS.n5018 VSS.n248 9.3005
R6905 VSS.n5020 VSS.n5019 9.3005
R6906 VSS.n5021 VSS.n247 9.3005
R6907 VSS.n5023 VSS.n5022 9.3005
R6908 VSS.n5024 VSS.n245 9.3005
R6909 VSS.n5026 VSS.n5025 9.3005
R6910 VSS.n5027 VSS.n244 9.3005
R6911 VSS.n5029 VSS.n5028 9.3005
R6912 VSS.n5030 VSS.n242 9.3005
R6913 VSS.n5031 VSS.n240 9.3005
R6914 VSS.n5032 VSS.n239 9.3005
R6915 VSS.n5034 VSS.n5033 9.3005
R6916 VSS.n5035 VSS.n238 9.3005
R6917 VSS.n5037 VSS.n5036 9.3005
R6918 VSS.n5038 VSS.n237 9.3005
R6919 VSS.n5040 VSS.n5039 9.3005
R6920 VSS.n5042 VSS.n5041 9.3005
R6921 VSS.n5043 VSS.n234 9.3005
R6922 VSS.n5045 VSS.n5044 9.3005
R6923 VSS.n5046 VSS.n233 9.3005
R6924 VSS.n5048 VSS.n5047 9.3005
R6925 VSS.n5050 VSS.n231 9.3005
R6926 VSS.n5052 VSS.n5051 9.3005
R6927 VSS.n5053 VSS.n230 9.3005
R6928 VSS.n5055 VSS.n5054 9.3005
R6929 VSS.n5056 VSS.n229 9.3005
R6930 VSS.n5058 VSS.n5057 9.3005
R6931 VSS.n5059 VSS.n228 9.3005
R6932 VSS.n5061 VSS.n5060 9.3005
R6933 VSS.n5062 VSS.n226 9.3005
R6934 VSS.n5064 VSS.n5063 9.3005
R6935 VSS.n5065 VSS.n225 9.3005
R6936 VSS.n5067 VSS.n5066 9.3005
R6937 VSS.n5068 VSS.n224 9.3005
R6938 VSS.n5070 VSS.n5069 9.3005
R6939 VSS.n5071 VSS.n223 9.3005
R6940 VSS.n5073 VSS.n5072 9.3005
R6941 VSS.n5074 VSS.n220 9.3005
R6942 VSS.n5075 VSS.n219 9.3005
R6943 VSS.n5080 VSS.n5079 9.3005
R6944 VSS.n5081 VSS.n218 9.3005
R6945 VSS.n5083 VSS.n5082 9.3005
R6946 VSS.n5084 VSS.n216 9.3005
R6947 VSS.n5085 VSS.n215 9.3005
R6948 VSS.n5087 VSS.n5086 9.3005
R6949 VSS.n5089 VSS.n5088 9.3005
R6950 VSS.n5091 VSS.n212 9.3005
R6951 VSS.n5093 VSS.n5092 9.3005
R6952 VSS.n5094 VSS.n211 9.3005
R6953 VSS.n5096 VSS.n5095 9.3005
R6954 VSS.n5097 VSS.n208 9.3005
R6955 VSS.n5099 VSS.n5098 9.3005
R6956 VSS.n5100 VSS.n207 9.3005
R6957 VSS.n5102 VSS.n5101 9.3005
R6958 VSS.n5103 VSS.n206 9.3005
R6959 VSS.n5104 VSS.n205 9.3005
R6960 VSS.n5105 VSS.n204 9.3005
R6961 VSS.n5107 VSS.n5106 9.3005
R6962 VSS.n5108 VSS.n203 9.3005
R6963 VSS.n5110 VSS.n5109 9.3005
R6964 VSS.n5112 VSS.n202 9.3005
R6965 VSS.n5114 VSS.n5113 9.3005
R6966 VSS.n5117 VSS.n198 9.3005
R6967 VSS.n5118 VSS.n197 9.3005
R6968 VSS.n5122 VSS.n5121 9.3005
R6969 VSS.n5124 VSS.n5123 9.3005
R6970 VSS.n5125 VSS.n195 9.3005
R6971 VSS.n5127 VSS.n5126 9.3005
R6972 VSS.n5128 VSS.n194 9.3005
R6973 VSS.n5130 VSS.n5129 9.3005
R6974 VSS.n5131 VSS.n191 9.3005
R6975 VSS.n5133 VSS.n5132 9.3005
R6976 VSS.n5134 VSS.n190 9.3005
R6977 VSS.n5136 VSS.n5135 9.3005
R6978 VSS.n5138 VSS.n188 9.3005
R6979 VSS.n5140 VSS.n5139 9.3005
R6980 VSS.n5141 VSS.n187 9.3005
R6981 VSS.n5143 VSS.n5142 9.3005
R6982 VSS.n5145 VSS.n186 9.3005
R6983 VSS.n5147 VSS.n5146 9.3005
R6984 VSS.n5148 VSS.n185 9.3005
R6985 VSS.n5150 VSS.n5149 9.3005
R6986 VSS.n5151 VSS.n182 9.3005
R6987 VSS.n5157 VSS.n5156 9.3005
R6988 VSS.n5158 VSS.n181 9.3005
R6989 VSS.n5160 VSS.n5159 9.3005
R6990 VSS.n5161 VSS.n180 9.3005
R6991 VSS.n5165 VSS.n5164 9.3005
R6992 VSS.n5166 VSS.n179 9.3005
R6993 VSS.n5168 VSS.n5167 9.3005
R6994 VSS.n5169 VSS.n177 9.3005
R6995 VSS.n5171 VSS.n5170 9.3005
R6996 VSS.n5172 VSS.n176 9.3005
R6997 VSS.n5174 VSS.n5173 9.3005
R6998 VSS.n5175 VSS.n174 9.3005
R6999 VSS.n5176 VSS.n172 9.3005
R7000 VSS.n5178 VSS.n5177 9.3005
R7001 VSS.n5179 VSS.n171 9.3005
R7002 VSS.n5181 VSS.n5180 9.3005
R7003 VSS.n5183 VSS.n170 9.3005
R7004 VSS.n5185 VSS.n5184 9.3005
R7005 VSS.n5186 VSS.n169 9.3005
R7006 VSS.n5188 VSS.n5187 9.3005
R7007 VSS.n5189 VSS.n167 9.3005
R7008 VSS.n5195 VSS.n5194 9.3005
R7009 VSS.n5197 VSS.n5196 9.3005
R7010 VSS.n5198 VSS.n165 9.3005
R7011 VSS.n5202 VSS.n5201 9.3005
R7012 VSS.n5203 VSS.n164 9.3005
R7013 VSS.n5205 VSS.n5204 9.3005
R7014 VSS.n5206 VSS.n163 9.3005
R7015 VSS.n5208 VSS.n5207 9.3005
R7016 VSS.n5209 VSS.n162 9.3005
R7017 VSS.n5211 VSS.n5210 9.3005
R7018 VSS.n5212 VSS.n160 9.3005
R7019 VSS.n5214 VSS.n5213 9.3005
R7020 VSS.n5215 VSS.n159 9.3005
R7021 VSS.n5217 VSS.n5216 9.3005
R7022 VSS.n5218 VSS.n156 9.3005
R7023 VSS.n5220 VSS.n5219 9.3005
R7024 VSS.n5221 VSS.n155 9.3005
R7025 VSS.n5223 VSS.n5222 9.3005
R7026 VSS.n5224 VSS.n154 9.3005
R7027 VSS.n5225 VSS.n153 9.3005
R7028 VSS.n5227 VSS.n5226 9.3005
R7029 VSS.n5228 VSS.n152 9.3005
R7030 VSS.n5230 VSS.n5229 9.3005
R7031 VSS.n5231 VSS.n151 9.3005
R7032 VSS.n5233 VSS.n5232 9.3005
R7033 VSS.n5234 VSS.n150 9.3005
R7034 VSS.n5236 VSS.n5235 9.3005
R7035 VSS.n5237 VSS.n147 9.3005
R7036 VSS.n5239 VSS.n5238 9.3005
R7037 VSS.n5240 VSS.n146 9.3005
R7038 VSS.n5242 VSS.n5241 9.3005
R7039 VSS.n5244 VSS.n145 9.3005
R7040 VSS.n5248 VSS.n5247 9.3005
R7041 VSS.n5249 VSS.n144 9.3005
R7042 VSS.n5252 VSS.n5251 9.3005
R7043 VSS.n5250 VSS.n143 9.3005
R7044 VSS.n5257 VSS.n142 9.3005
R7045 VSS.n5259 VSS.n5258 9.3005
R7046 VSS.n5260 VSS.n141 9.3005
R7047 VSS.n5262 VSS.n5261 9.3005
R7048 VSS.n5263 VSS.n139 9.3005
R7049 VSS.n5264 VSS.n137 9.3005
R7050 VSS.n5266 VSS.n5265 9.3005
R7051 VSS.n5267 VSS.n136 9.3005
R7052 VSS.n5269 VSS.n5268 9.3005
R7053 VSS.n5270 VSS.n134 9.3005
R7054 VSS.n5272 VSS.n5271 9.3005
R7055 VSS.n5273 VSS.n133 9.3005
R7056 VSS.n5275 VSS.n5274 9.3005
R7057 VSS.n5276 VSS.n131 9.3005
R7058 VSS.n5277 VSS.n130 9.3005
R7059 VSS.n5279 VSS.n5278 9.3005
R7060 VSS.n5280 VSS.n129 9.3005
R7061 VSS.n5283 VSS.n5282 9.3005
R7062 VSS.n5281 VSS.n128 9.3005
R7063 VSS.n5288 VSS.n127 9.3005
R7064 VSS.n5290 VSS.n5289 9.3005
R7065 VSS.n5291 VSS.n126 9.3005
R7066 VSS.n5293 VSS.n5292 9.3005
R7067 VSS.n5294 VSS.n124 9.3005
R7068 VSS.n5296 VSS.n5295 9.3005
R7069 VSS.n5297 VSS.n123 9.3005
R7070 VSS.n5300 VSS.n5299 9.3005
R7071 VSS.n5298 VSS.n122 9.3005
R7072 VSS.n5305 VSS.n121 9.3005
R7073 VSS.n5307 VSS.n5306 9.3005
R7074 VSS.n5308 VSS.n120 9.3005
R7075 VSS.n5310 VSS.n5309 9.3005
R7076 VSS.n5311 VSS.n118 9.3005
R7077 VSS.n5312 VSS.n116 9.3005
R7078 VSS.n5314 VSS.n5313 9.3005
R7079 VSS.n5315 VSS.n115 9.3005
R7080 VSS.n5317 VSS.n5316 9.3005
R7081 VSS.n5318 VSS.n113 9.3005
R7082 VSS.n5320 VSS.n5319 9.3005
R7083 VSS.n5321 VSS.n112 9.3005
R7084 VSS.n5323 VSS.n5322 9.3005
R7085 VSS.n5324 VSS.n110 9.3005
R7086 VSS.n5326 VSS.n5325 9.3005
R7087 VSS.n5327 VSS.n109 9.3005
R7088 VSS.n5329 VSS.n5328 9.3005
R7089 VSS.n5331 VSS.n108 9.3005
R7090 VSS.n5335 VSS.n5334 9.3005
R7091 VSS.n5339 VSS.n101 9.3005
R7092 VSS.n5350 VSS.n5349 9.3005
R7093 VSS.n5351 VSS.n99 9.3005
R7094 VSS.n5352 VSS.n97 9.3005
R7095 VSS.n5354 VSS.n5353 9.3005
R7096 VSS.n5355 VSS.n96 9.3005
R7097 VSS.n5357 VSS.n5356 9.3005
R7098 VSS.n5358 VSS.n95 9.3005
R7099 VSS.n5364 VSS.n5363 9.3005
R7100 VSS.n5365 VSS.n94 9.3005
R7101 VSS.n5367 VSS.n5366 9.3005
R7102 VSS.n5368 VSS.n93 9.3005
R7103 VSS.n5370 VSS.n5369 9.3005
R7104 VSS.n5371 VSS.n92 9.3005
R7105 VSS.n5373 VSS.n5372 9.3005
R7106 VSS.n5374 VSS.n90 9.3005
R7107 VSS.n89 VSS.n25 9.3005
R7108 VSS.n88 VSS.n87 9.3005
R7109 VSS.n86 VSS.n26 9.3005
R7110 VSS.n85 VSS.n84 9.3005
R7111 VSS.n83 VSS.n27 9.3005
R7112 VSS.n82 VSS.n81 9.3005
R7113 VSS.n80 VSS.n28 9.3005
R7114 VSS.n77 VSS.n76 9.3005
R7115 VSS.n75 VSS.n30 9.3005
R7116 VSS.n74 VSS.n73 9.3005
R7117 VSS.n71 VSS.n31 9.3005
R7118 VSS.n70 VSS.n69 9.3005
R7119 VSS.n68 VSS.n33 9.3005
R7120 VSS.n67 VSS.n66 9.3005
R7121 VSS.n65 VSS.n34 9.3005
R7122 VSS.n64 VSS.n63 9.3005
R7123 VSS.n62 VSS.n36 9.3005
R7124 VSS.n61 VSS.n60 9.3005
R7125 VSS.n59 VSS.n37 9.3005
R7126 VSS.n58 VSS.n57 9.3005
R7127 VSS.n56 VSS.n39 9.3005
R7128 VSS.n55 VSS.n54 9.3005
R7129 VSS.n53 VSS.n40 9.3005
R7130 VSS.n51 VSS.n50 9.3005
R7131 VSS.n49 VSS.n41 9.3005
R7132 VSS.n48 VSS.n47 9.3005
R7133 VSS.n45 VSS.n42 9.3005
R7134 VSS.n4939 VSS.n4915 9.3005
R7135 VSS.n296 VSS.n295 9.3005
R7136 VSS.n297 VSS.n289 9.3005
R7137 VSS.n299 VSS.n298 9.3005
R7138 VSS.n301 VSS.n286 9.3005
R7139 VSS.n308 VSS.n307 9.3005
R7140 VSS.n309 VSS.n284 9.3005
R7141 VSS.n954 VSS.n285 9.3005
R7142 VSS.n953 VSS.n952 9.3005
R7143 VSS.n951 VSS.n310 9.3005
R7144 VSS.n950 VSS.n949 9.3005
R7145 VSS.n948 VSS.n313 9.3005
R7146 VSS.n947 VSS.n946 9.3005
R7147 VSS.n945 VSS.n314 9.3005
R7148 VSS.n943 VSS.n942 9.3005
R7149 VSS.n941 VSS.n940 9.3005
R7150 VSS.n321 VSS.n319 9.3005
R7151 VSS.n934 VSS.n933 9.3005
R7152 VSS.n932 VSS.n931 9.3005
R7153 VSS.n929 VSS.n323 9.3005
R7154 VSS.n928 VSS.n927 9.3005
R7155 VSS.n926 VSS.n925 9.3005
R7156 VSS.n921 VSS.n327 9.3005
R7157 VSS.n920 VSS.n919 9.3005
R7158 VSS.n918 VSS.n917 9.3005
R7159 VSS.n916 VSS.n330 9.3005
R7160 VSS.n915 VSS.n331 9.3005
R7161 VSS.n914 VSS.n913 9.3005
R7162 VSS.n912 VSS.n333 9.3005
R7163 VSS.n911 VSS.n910 9.3005
R7164 VSS.n909 VSS.n334 9.3005
R7165 VSS.n908 VSS.n907 9.3005
R7166 VSS.n906 VSS.n336 9.3005
R7167 VSS.n905 VSS.n904 9.3005
R7168 VSS.n903 VSS.n337 9.3005
R7169 VSS.n902 VSS.n901 9.3005
R7170 VSS.n900 VSS.n341 9.3005
R7171 VSS.n899 VSS.n898 9.3005
R7172 VSS.n895 VSS.n342 9.3005
R7173 VSS.n894 VSS.n893 9.3005
R7174 VSS.n892 VSS.n344 9.3005
R7175 VSS.n891 VSS.n890 9.3005
R7176 VSS.n889 VSS.n345 9.3005
R7177 VSS.n888 VSS.n887 9.3005
R7178 VSS.n886 VSS.n350 9.3005
R7179 VSS.n885 VSS.n884 9.3005
R7180 VSS.n883 VSS.n351 9.3005
R7181 VSS.n882 VSS.n881 9.3005
R7182 VSS.n880 VSS.n354 9.3005
R7183 VSS.n879 VSS.n878 9.3005
R7184 VSS.n877 VSS.n355 9.3005
R7185 VSS.n876 VSS.n875 9.3005
R7186 VSS.n874 VSS.n873 9.3005
R7187 VSS.n871 VSS.n358 9.3005
R7188 VSS.n869 VSS.n868 9.3005
R7189 VSS.n867 VSS.n360 9.3005
R7190 VSS.n866 VSS.n865 9.3005
R7191 VSS.n863 VSS.n361 9.3005
R7192 VSS.n861 VSS.n860 9.3005
R7193 VSS.n859 VSS.n365 9.3005
R7194 VSS.n858 VSS.n857 9.3005
R7195 VSS.n856 VSS.n366 9.3005
R7196 VSS.n855 VSS.n367 9.3005
R7197 VSS.n854 VSS.n369 9.3005
R7198 VSS.n853 VSS.n370 9.3005
R7199 VSS.n852 VSS.n371 9.3005
R7200 VSS.n851 VSS.n850 9.3005
R7201 VSS.n849 VSS.n374 9.3005
R7202 VSS.n848 VSS.n847 9.3005
R7203 VSS.n846 VSS.n375 9.3005
R7204 VSS.n845 VSS.n844 9.3005
R7205 VSS.n843 VSS.n379 9.3005
R7206 VSS.n842 VSS.n841 9.3005
R7207 VSS.n839 VSS.n380 9.3005
R7208 VSS.n838 VSS.n837 9.3005
R7209 VSS.n836 VSS.n835 9.3005
R7210 VSS.n834 VSS.n384 9.3005
R7211 VSS.n831 VSS.n830 9.3005
R7212 VSS.n829 VSS.n388 9.3005
R7213 VSS.n828 VSS.n827 9.3005
R7214 VSS.n826 VSS.n389 9.3005
R7215 VSS.n825 VSS.n396 9.3005
R7216 VSS.n824 VSS.n397 9.3005
R7217 VSS.n823 VSS.n398 9.3005
R7218 VSS.n821 VSS.n820 9.3005
R7219 VSS.n819 VSS.n818 9.3005
R7220 VSS.n817 VSS.n400 9.3005
R7221 VSS.n816 VSS.n815 9.3005
R7222 VSS.n814 VSS.n813 9.3005
R7223 VSS.n812 VSS.n402 9.3005
R7224 VSS.n811 VSS.n409 9.3005
R7225 VSS.n810 VSS.n809 9.3005
R7226 VSS.n808 VSS.n410 9.3005
R7227 VSS.n807 VSS.n806 9.3005
R7228 VSS.n805 VSS.n411 9.3005
R7229 VSS.n804 VSS.n803 9.3005
R7230 VSS.n802 VSS.n416 9.3005
R7231 VSS.n801 VSS.n800 9.3005
R7232 VSS.n799 VSS.n417 9.3005
R7233 VSS.n798 VSS.n419 9.3005
R7234 VSS.n797 VSS.n796 9.3005
R7235 VSS.n795 VSS.n420 9.3005
R7236 VSS.n794 VSS.n793 9.3005
R7237 VSS.n792 VSS.n421 9.3005
R7238 VSS.n791 VSS.n790 9.3005
R7239 VSS.n789 VSS.n427 9.3005
R7240 VSS.n788 VSS.n787 9.3005
R7241 VSS.n786 VSS.n428 9.3005
R7242 VSS.n785 VSS.n429 9.3005
R7243 VSS.n784 VSS.n783 9.3005
R7244 VSS.n782 VSS.n781 9.3005
R7245 VSS.n779 VSS.n432 9.3005
R7246 VSS.n778 VSS.n434 9.3005
R7247 VSS.n777 VSS.n776 9.3005
R7248 VSS.n775 VSS.n435 9.3005
R7249 VSS.n774 VSS.n773 9.3005
R7250 VSS.n772 VSS.n436 9.3005
R7251 VSS.n771 VSS.n770 9.3005
R7252 VSS.n769 VSS.n439 9.3005
R7253 VSS.n768 VSS.n767 9.3005
R7254 VSS.n766 VSS.n440 9.3005
R7255 VSS.n765 VSS.n441 9.3005
R7256 VSS.n764 VSS.n442 9.3005
R7257 VSS.n763 VSS.n444 9.3005
R7258 VSS.n762 VSS.n445 9.3005
R7259 VSS.n761 VSS.n760 9.3005
R7260 VSS.n759 VSS.n448 9.3005
R7261 VSS.n758 VSS.n757 9.3005
R7262 VSS.n756 VSS.n449 9.3005
R7263 VSS.n452 VSS.n450 9.3005
R7264 VSS.n751 VSS.n750 9.3005
R7265 VSS.n749 VSS.n451 9.3005
R7266 VSS.n748 VSS.n747 9.3005
R7267 VSS.n746 VSS.n453 9.3005
R7268 VSS.n745 VSS.n744 9.3005
R7269 VSS.n743 VSS.n742 9.3005
R7270 VSS.n741 VSS.n456 9.3005
R7271 VSS.n740 VSS.n739 9.3005
R7272 VSS.n738 VSS.n459 9.3005
R7273 VSS.n737 VSS.n736 9.3005
R7274 VSS.n734 VSS.n460 9.3005
R7275 VSS.n733 VSS.n462 9.3005
R7276 VSS.n732 VSS.n731 9.3005
R7277 VSS.n730 VSS.n464 9.3005
R7278 VSS.n729 VSS.n728 9.3005
R7279 VSS.n727 VSS.n465 9.3005
R7280 VSS.n726 VSS.n468 9.3005
R7281 VSS.n725 VSS.n724 9.3005
R7282 VSS.n723 VSS.n470 9.3005
R7283 VSS.n722 VSS.n721 9.3005
R7284 VSS.n720 VSS.n471 9.3005
R7285 VSS.n719 VSS.n472 9.3005
R7286 VSS.n718 VSS.n717 9.3005
R7287 VSS.n716 VSS.n473 9.3005
R7288 VSS.n715 VSS.n714 9.3005
R7289 VSS.n713 VSS.n474 9.3005
R7290 VSS.n712 VSS.n711 9.3005
R7291 VSS.n710 VSS.n709 9.3005
R7292 VSS.n708 VSS.n477 9.3005
R7293 VSS.n707 VSS.n706 9.3005
R7294 VSS.n705 VSS.n704 9.3005
R7295 VSS.n700 VSS.n479 9.3005
R7296 VSS.n698 VSS.n697 9.3005
R7297 VSS.n696 VSS.n481 9.3005
R7298 VSS.n695 VSS.n694 9.3005
R7299 VSS.n693 VSS.n482 9.3005
R7300 VSS.n692 VSS.n691 9.3005
R7301 VSS.n690 VSS.n484 9.3005
R7302 VSS.n689 VSS.n688 9.3005
R7303 VSS.n686 VSS.n485 9.3005
R7304 VSS.n685 VSS.n684 9.3005
R7305 VSS.n681 VSS.n489 9.3005
R7306 VSS.n679 VSS.n678 9.3005
R7307 VSS.n677 VSS.n494 9.3005
R7308 VSS.n676 VSS.n675 9.3005
R7309 VSS.n674 VSS.n495 9.3005
R7310 VSS.n673 VSS.n672 9.3005
R7311 VSS.n671 VSS.n498 9.3005
R7312 VSS.n670 VSS.n669 9.3005
R7313 VSS.n668 VSS.n499 9.3005
R7314 VSS.n667 VSS.n500 9.3005
R7315 VSS.n666 VSS.n665 9.3005
R7316 VSS.n664 VSS.n502 9.3005
R7317 VSS.n663 VSS.n662 9.3005
R7318 VSS.n660 VSS.n503 9.3005
R7319 VSS.n659 VSS.n505 9.3005
R7320 VSS.n658 VSS.n657 9.3005
R7321 VSS.n656 VSS.n506 9.3005
R7322 VSS.n655 VSS.n654 9.3005
R7323 VSS.n652 VSS.n507 9.3005
R7324 VSS.n651 VSS.n650 9.3005
R7325 VSS.n649 VSS.n511 9.3005
R7326 VSS.n648 VSS.n647 9.3005
R7327 VSS.n646 VSS.n512 9.3005
R7328 VSS.n645 VSS.n644 9.3005
R7329 VSS.n643 VSS.n514 9.3005
R7330 VSS.n642 VSS.n641 9.3005
R7331 VSS.n640 VSS.n515 9.3005
R7332 VSS.n639 VSS.n518 9.3005
R7333 VSS.n638 VSS.n520 9.3005
R7334 VSS.n637 VSS.n636 9.3005
R7335 VSS.n635 VSS.n634 9.3005
R7336 VSS.n631 VSS.n522 9.3005
R7337 VSS.n630 VSS.n629 9.3005
R7338 VSS.n628 VSS.n524 9.3005
R7339 VSS.n627 VSS.n626 9.3005
R7340 VSS.n625 VSS.n525 9.3005
R7341 VSS.n624 VSS.n623 9.3005
R7342 VSS.n622 VSS.n621 9.3005
R7343 VSS.n620 VSS.n528 9.3005
R7344 VSS.n619 VSS.n618 9.3005
R7345 VSS.n617 VSS.n532 9.3005
R7346 VSS.n616 VSS.n615 9.3005
R7347 VSS.n612 VSS.n533 9.3005
R7348 VSS.n611 VSS.n610 9.3005
R7349 VSS.n609 VSS.n536 9.3005
R7350 VSS.n608 VSS.n607 9.3005
R7351 VSS.n606 VSS.n537 9.3005
R7352 VSS.n603 VSS.n602 9.3005
R7353 VSS.n601 VSS.n538 9.3005
R7354 VSS.n600 VSS.n599 9.3005
R7355 VSS.n596 VSS.n539 9.3005
R7356 VSS.n595 VSS.n594 9.3005
R7357 VSS.n593 VSS.n541 9.3005
R7358 VSS.n592 VSS.n591 9.3005
R7359 VSS.n590 VSS.n542 9.3005
R7360 VSS.n589 VSS.n546 9.3005
R7361 VSS.n588 VSS.n547 9.3005
R7362 VSS.n587 VSS.n586 9.3005
R7363 VSS.n585 VSS.n584 9.3005
R7364 VSS.n583 VSS.n550 9.3005
R7365 VSS.n580 VSS.n579 9.3005
R7366 VSS.n578 VSS.n552 9.3005
R7367 VSS.n577 VSS.n576 9.3005
R7368 VSS.n575 VSS.n553 9.3005
R7369 VSS.n574 VSS.n555 9.3005
R7370 VSS.n572 VSS.n571 9.3005
R7371 VSS.n570 VSS.n558 9.3005
R7372 VSS.n569 VSS.n568 9.3005
R7373 VSS.n560 VSS.n559 9.3005
R7374 VSS.n563 VSS.n5 9.3005
R7375 VSS.n9 VSS.n6 9.3005
R7376 VSS.n5478 VSS.n5477 9.3005
R7377 VSS.n5476 VSS.n5475 9.3005
R7378 VSS.n5474 VSS.n11 9.3005
R7379 VSS.n5473 VSS.n5472 9.3005
R7380 VSS.n5471 VSS.n12 9.3005
R7381 VSS.n5468 VSS.n5467 9.3005
R7382 VSS.n5466 VSS.n13 9.3005
R7383 VSS.n5465 VSS.n5464 9.3005
R7384 VSS.n5462 VSS.n14 9.3005
R7385 VSS.n5460 VSS.n5459 9.3005
R7386 VSS.n5458 VSS.n5457 9.3005
R7387 VSS.n5455 VSS.n21 9.3005
R7388 VSS.n5452 VSS.n5451 9.3005
R7389 VSS.n5450 VSS.n5449 9.3005
R7390 VSS.n5448 VSS.n24 9.3005
R7391 VSS.n5447 VSS.n5446 9.3005
R7392 VSS.n5445 VSS.n5444 9.3005
R7393 VSS.n5443 VSS.n5380 9.3005
R7394 VSS.n5442 VSS.n5441 9.3005
R7395 VSS.n5440 VSS.n5383 9.3005
R7396 VSS.n5439 VSS.n5438 9.3005
R7397 VSS.n5436 VSS.n5384 9.3005
R7398 VSS.n5435 VSS.n5434 9.3005
R7399 VSS.n5433 VSS.n5387 9.3005
R7400 VSS.n5432 VSS.n5431 9.3005
R7401 VSS.n5390 VSS.n5388 9.3005
R7402 VSS.n5426 VSS.n5425 9.3005
R7403 VSS.n5424 VSS.n5392 9.3005
R7404 VSS.n5423 VSS.n5422 9.3005
R7405 VSS.n5421 VSS.n5393 9.3005
R7406 VSS.n5420 VSS.n5396 9.3005
R7407 VSS.n5419 VSS.n5418 9.3005
R7408 VSS.n5417 VSS.n5399 9.3005
R7409 VSS.n5416 VSS.n5415 9.3005
R7410 VSS.n5414 VSS.n5400 9.3005
R7411 VSS.n5413 VSS.n5412 9.3005
R7412 VSS.n5411 VSS.n5403 9.3005
R7413 VSS.n5410 VSS.n5409 9.3005
R7414 VSS.n956 VSS.n955 9.3005
R7415 VSS.n2072 VSS.n2071 9.3005
R7416 VSS.n2073 VSS.n2065 9.3005
R7417 VSS.n2075 VSS.n2074 9.3005
R7418 VSS.n2077 VSS.n2062 9.3005
R7419 VSS.n2080 VSS.n2079 9.3005
R7420 VSS.n2081 VSS.n2060 9.3005
R7421 VSS.n2084 VSS.n2058 9.3005
R7422 VSS.n2087 VSS.n2086 9.3005
R7423 VSS.n2088 VSS.n2057 9.3005
R7424 VSS.n2090 VSS.n2089 9.3005
R7425 VSS.n2091 VSS.n2055 9.3005
R7426 VSS.n2093 VSS.n2092 9.3005
R7427 VSS.n2094 VSS.n2054 9.3005
R7428 VSS.n2096 VSS.n2095 9.3005
R7429 VSS.n2098 VSS.n2053 9.3005
R7430 VSS.n2100 VSS.n2099 9.3005
R7431 VSS.n2101 VSS.n2052 9.3005
R7432 VSS.n2103 VSS.n2102 9.3005
R7433 VSS.n2104 VSS.n2051 9.3005
R7434 VSS.n2107 VSS.n2106 9.3005
R7435 VSS.n2108 VSS.n2050 9.3005
R7436 VSS.n2110 VSS.n2109 9.3005
R7437 VSS.n2111 VSS.n2048 9.3005
R7438 VSS.n2115 VSS.n2114 9.3005
R7439 VSS.n2116 VSS.n2047 9.3005
R7440 VSS.n2119 VSS.n2117 9.3005
R7441 VSS.n2120 VSS.n2046 9.3005
R7442 VSS.n2124 VSS.n2123 9.3005
R7443 VSS.n2125 VSS.n2045 9.3005
R7444 VSS.n2127 VSS.n2126 9.3005
R7445 VSS.n2129 VSS.n2044 9.3005
R7446 VSS.n2131 VSS.n2130 9.3005
R7447 VSS.n2132 VSS.n2043 9.3005
R7448 VSS.n2204 VSS.n2133 9.3005
R7449 VSS.n2203 VSS.n2134 9.3005
R7450 VSS.n2202 VSS.n2201 9.3005
R7451 VSS.n2200 VSS.n2135 9.3005
R7452 VSS.n2199 VSS.n2198 9.3005
R7453 VSS.n2194 VSS.n2136 9.3005
R7454 VSS.n2193 VSS.n2192 9.3005
R7455 VSS.n2191 VSS.n2142 9.3005
R7456 VSS.n2190 VSS.n2189 9.3005
R7457 VSS.n2188 VSS.n2143 9.3005
R7458 VSS.n2187 VSS.n2186 9.3005
R7459 VSS.n2185 VSS.n2144 9.3005
R7460 VSS.n2184 VSS.n2183 9.3005
R7461 VSS.n2182 VSS.n2145 9.3005
R7462 VSS.n2181 VSS.n2180 9.3005
R7463 VSS.n2179 VSS.n2147 9.3005
R7464 VSS.n2178 VSS.n2177 9.3005
R7465 VSS.n2176 VSS.n2148 9.3005
R7466 VSS.n2175 VSS.n2174 9.3005
R7467 VSS.n2173 VSS.n2152 9.3005
R7468 VSS.n2172 VSS.n2171 9.3005
R7469 VSS.n2169 VSS.n2153 9.3005
R7470 VSS.n2168 VSS.n2167 9.3005
R7471 VSS.n2166 VSS.n2155 9.3005
R7472 VSS.n2165 VSS.n2164 9.3005
R7473 VSS.n2162 VSS.n2156 9.3005
R7474 VSS.n2161 VSS.n2160 9.3005
R7475 VSS.n2159 VSS.n2040 9.3005
R7476 VSS.n2207 VSS.n2042 9.3005
R7477 VSS.n2208 VSS.n2039 9.3005
R7478 VSS.n2210 VSS.n2209 9.3005
R7479 VSS.n2211 VSS.n2038 9.3005
R7480 VSS.n2213 VSS.n2212 9.3005
R7481 VSS.n2215 VSS.n2036 9.3005
R7482 VSS.n2217 VSS.n2216 9.3005
R7483 VSS.n2218 VSS.n2035 9.3005
R7484 VSS.n2220 VSS.n2219 9.3005
R7485 VSS.n2222 VSS.n2033 9.3005
R7486 VSS.n2224 VSS.n2223 9.3005
R7487 VSS.n2226 VSS.n2225 9.3005
R7488 VSS.n2227 VSS.n2030 9.3005
R7489 VSS.n2231 VSS.n2230 9.3005
R7490 VSS.n2233 VSS.n2232 9.3005
R7491 VSS.n2235 VSS.n2026 9.3005
R7492 VSS.n2238 VSS.n2237 9.3005
R7493 VSS.n2240 VSS.n2239 9.3005
R7494 VSS.n2242 VSS.n2022 9.3005
R7495 VSS.n2245 VSS.n2244 9.3005
R7496 VSS.n2247 VSS.n2246 9.3005
R7497 VSS.n2249 VSS.n2019 9.3005
R7498 VSS.n2252 VSS.n2251 9.3005
R7499 VSS.n2253 VSS.n2018 9.3005
R7500 VSS.n2255 VSS.n2254 9.3005
R7501 VSS.n2256 VSS.n2017 9.3005
R7502 VSS.n2261 VSS.n2260 9.3005
R7503 VSS.n2262 VSS.n2016 9.3005
R7504 VSS.n2335 VSS.n2263 9.3005
R7505 VSS.n2334 VSS.n2333 9.3005
R7506 VSS.n2332 VSS.n2264 9.3005
R7507 VSS.n2331 VSS.n2330 9.3005
R7508 VSS.n2329 VSS.n2265 9.3005
R7509 VSS.n2328 VSS.n2327 9.3005
R7510 VSS.n2326 VSS.n2266 9.3005
R7511 VSS.n2325 VSS.n2324 9.3005
R7512 VSS.n2321 VSS.n2267 9.3005
R7513 VSS.n2318 VSS.n2317 9.3005
R7514 VSS.n2316 VSS.n2270 9.3005
R7515 VSS.n2315 VSS.n2314 9.3005
R7516 VSS.n2309 VSS.n2271 9.3005
R7517 VSS.n2308 VSS.n2307 9.3005
R7518 VSS.n2306 VSS.n2272 9.3005
R7519 VSS.n2305 VSS.n2304 9.3005
R7520 VSS.n2302 VSS.n2273 9.3005
R7521 VSS.n2301 VSS.n2300 9.3005
R7522 VSS.n2299 VSS.n2298 9.3005
R7523 VSS.n2296 VSS.n2277 9.3005
R7524 VSS.n2293 VSS.n2292 9.3005
R7525 VSS.n2291 VSS.n2279 9.3005
R7526 VSS.n2290 VSS.n2289 9.3005
R7527 VSS.n2288 VSS.n2280 9.3005
R7528 VSS.n2287 VSS.n2282 9.3005
R7529 VSS.n2286 VSS.n2285 9.3005
R7530 VSS.n2284 VSS.n2283 9.3005
R7531 VSS.n2015 VSS.n2014 9.3005
R7532 VSS.n2339 VSS.n2338 9.3005
R7533 VSS.n2340 VSS.n2013 9.3005
R7534 VSS.n2342 VSS.n2341 9.3005
R7535 VSS.n2343 VSS.n2012 9.3005
R7536 VSS.n2346 VSS.n2345 9.3005
R7537 VSS.n2347 VSS.n2011 9.3005
R7538 VSS.n2349 VSS.n2348 9.3005
R7539 VSS.n2351 VSS.n2010 9.3005
R7540 VSS.n2353 VSS.n2352 9.3005
R7541 VSS.n2354 VSS.n2009 9.3005
R7542 VSS.n2356 VSS.n2355 9.3005
R7543 VSS.n2357 VSS.n2007 9.3005
R7544 VSS.n2361 VSS.n2360 9.3005
R7545 VSS.n2362 VSS.n2006 9.3005
R7546 VSS.n2364 VSS.n2363 9.3005
R7547 VSS.n2365 VSS.n2005 9.3005
R7548 VSS.n2367 VSS.n2366 9.3005
R7549 VSS.n2369 VSS.n2368 9.3005
R7550 VSS.n2371 VSS.n2002 9.3005
R7551 VSS.n2377 VSS.n2376 9.3005
R7552 VSS.n2378 VSS.n2001 9.3005
R7553 VSS.n2380 VSS.n2379 9.3005
R7554 VSS.n2381 VSS.n2000 9.3005
R7555 VSS.n2385 VSS.n2384 9.3005
R7556 VSS.n2386 VSS.n1999 9.3005
R7557 VSS.n2388 VSS.n2387 9.3005
R7558 VSS.n2391 VSS.n1998 9.3005
R7559 VSS.n2393 VSS.n2392 9.3005
R7560 VSS.n2471 VSS.n2470 9.3005
R7561 VSS.n2469 VSS.n1997 9.3005
R7562 VSS.n2468 VSS.n2467 9.3005
R7563 VSS.n2466 VSS.n2394 9.3005
R7564 VSS.n2465 VSS.n2464 9.3005
R7565 VSS.n2463 VSS.n2397 9.3005
R7566 VSS.n2462 VSS.n2461 9.3005
R7567 VSS.n2456 VSS.n2398 9.3005
R7568 VSS.n2455 VSS.n2400 9.3005
R7569 VSS.n2454 VSS.n2453 9.3005
R7570 VSS.n2452 VSS.n2402 9.3005
R7571 VSS.n2451 VSS.n2450 9.3005
R7572 VSS.n2448 VSS.n2403 9.3005
R7573 VSS.n2446 VSS.n2445 9.3005
R7574 VSS.n2444 VSS.n2406 9.3005
R7575 VSS.n2443 VSS.n2442 9.3005
R7576 VSS.n2441 VSS.n2407 9.3005
R7577 VSS.n2439 VSS.n2438 9.3005
R7578 VSS.n2437 VSS.n2436 9.3005
R7579 VSS.n2435 VSS.n2412 9.3005
R7580 VSS.n2434 VSS.n2433 9.3005
R7581 VSS.n2432 VSS.n2414 9.3005
R7582 VSS.n2431 VSS.n2430 9.3005
R7583 VSS.n2429 VSS.n2415 9.3005
R7584 VSS.n2428 VSS.n2427 9.3005
R7585 VSS.n2426 VSS.n2425 9.3005
R7586 VSS.n2420 VSS.n2419 9.3005
R7587 VSS.n1994 VSS.n1992 9.3005
R7588 VSS.n2476 VSS.n2475 9.3005
R7589 VSS.n2478 VSS.n2477 9.3005
R7590 VSS.n2479 VSS.n1988 9.3005
R7591 VSS.n2482 VSS.n2481 9.3005
R7592 VSS.n2484 VSS.n2483 9.3005
R7593 VSS.n2487 VSS.n1986 9.3005
R7594 VSS.n2494 VSS.n2493 9.3005
R7595 VSS.n2496 VSS.n2495 9.3005
R7596 VSS.n2498 VSS.n1984 9.3005
R7597 VSS.n2500 VSS.n2499 9.3005
R7598 VSS.n2502 VSS.n2501 9.3005
R7599 VSS.n2504 VSS.n1981 9.3005
R7600 VSS.n2506 VSS.n2505 9.3005
R7601 VSS.n2507 VSS.n1979 9.3005
R7602 VSS.n2509 VSS.n2508 9.3005
R7603 VSS.n2511 VSS.n1978 9.3005
R7604 VSS.n2513 VSS.n2512 9.3005
R7605 VSS.n2514 VSS.n1977 9.3005
R7606 VSS.n2516 VSS.n2515 9.3005
R7607 VSS.n2519 VSS.n1976 9.3005
R7608 VSS.n2522 VSS.n2521 9.3005
R7609 VSS.n2524 VSS.n2523 9.3005
R7610 VSS.n2527 VSS.n1974 9.3005
R7611 VSS.n2529 VSS.n2528 9.3005
R7612 VSS.n2530 VSS.n1972 9.3005
R7613 VSS.n2532 VSS.n2531 9.3005
R7614 VSS.n2533 VSS.n1971 9.3005
R7615 VSS.n2535 VSS.n2534 9.3005
R7616 VSS.n2536 VSS.n1970 9.3005
R7617 VSS.n2538 VSS.n2537 9.3005
R7618 VSS.n2539 VSS.n1969 9.3005
R7619 VSS.n2541 VSS.n2540 9.3005
R7620 VSS.n2542 VSS.n1968 9.3005
R7621 VSS.n2544 VSS.n2543 9.3005
R7622 VSS.n2546 VSS.n1967 9.3005
R7623 VSS.n2548 VSS.n2547 9.3005
R7624 VSS.n2549 VSS.n1966 9.3005
R7625 VSS.n2551 VSS.n2550 9.3005
R7626 VSS.n2556 VSS.n1965 9.3005
R7627 VSS.n2558 VSS.n2557 9.3005
R7628 VSS.n2559 VSS.n1964 9.3005
R7629 VSS.n2561 VSS.n2560 9.3005
R7630 VSS.n2562 VSS.n1962 9.3005
R7631 VSS.n2564 VSS.n2563 9.3005
R7632 VSS.n2566 VSS.n2565 9.3005
R7633 VSS.n2567 VSS.n1959 9.3005
R7634 VSS.n2572 VSS.n2571 9.3005
R7635 VSS.n2573 VSS.n1958 9.3005
R7636 VSS.n2575 VSS.n2574 9.3005
R7637 VSS.n2577 VSS.n1956 9.3005
R7638 VSS.n2580 VSS.n2579 9.3005
R7639 VSS.n2581 VSS.n1955 9.3005
R7640 VSS.n2583 VSS.n2582 9.3005
R7641 VSS.n2585 VSS.n1953 9.3005
R7642 VSS.n2590 VSS.n2589 9.3005
R7643 VSS.n2591 VSS.n1950 9.3005
R7644 VSS.n2633 VSS.n2632 9.3005
R7645 VSS.n2631 VSS.n2630 9.3005
R7646 VSS.n2629 VSS.n2592 9.3005
R7647 VSS.n2627 VSS.n2626 9.3005
R7648 VSS.n2625 VSS.n2624 9.3005
R7649 VSS.n2622 VSS.n2596 9.3005
R7650 VSS.n2621 VSS.n2599 9.3005
R7651 VSS.n2620 VSS.n2619 9.3005
R7652 VSS.n2618 VSS.n2601 9.3005
R7653 VSS.n2617 VSS.n2616 9.3005
R7654 VSS.n2615 VSS.n2602 9.3005
R7655 VSS.n2614 VSS.n2613 9.3005
R7656 VSS.n2612 VSS.n2611 9.3005
R7657 VSS.n2609 VSS.n1934 9.3005
R7658 VSS.n2608 VSS.n1935 9.3005
R7659 VSS.n2731 VSS.n2730 9.3005
R7660 VSS.n2729 VSS.n2728 9.3005
R7661 VSS.n2727 VSS.n1939 9.3005
R7662 VSS.n2726 VSS.n2725 9.3005
R7663 VSS.n2724 VSS.n1940 9.3005
R7664 VSS.n2723 VSS.n2722 9.3005
R7665 VSS.n2721 VSS.n2720 9.3005
R7666 VSS.n2716 VSS.n1944 9.3005
R7667 VSS.n2714 VSS.n2713 9.3005
R7668 VSS.n2712 VSS.n1945 9.3005
R7669 VSS.n2711 VSS.n2710 9.3005
R7670 VSS.n2709 VSS.n1946 9.3005
R7671 VSS.n2708 VSS.n2707 9.3005
R7672 VSS.n2706 VSS.n2636 9.3005
R7673 VSS.n2705 VSS.n2704 9.3005
R7674 VSS.n2701 VSS.n2637 9.3005
R7675 VSS.n2700 VSS.n2699 9.3005
R7676 VSS.n2698 VSS.n2639 9.3005
R7677 VSS.n2697 VSS.n2696 9.3005
R7678 VSS.n2694 VSS.n2640 9.3005
R7679 VSS.n2692 VSS.n2691 9.3005
R7680 VSS.n2690 VSS.n2643 9.3005
R7681 VSS.n2689 VSS.n2688 9.3005
R7682 VSS.n2687 VSS.n2644 9.3005
R7683 VSS.n2685 VSS.n2684 9.3005
R7684 VSS.n2683 VSS.n2646 9.3005
R7685 VSS.n2682 VSS.n2681 9.3005
R7686 VSS.n2680 VSS.n2647 9.3005
R7687 VSS.n2679 VSS.n2648 9.3005
R7688 VSS.n2678 VSS.n2677 9.3005
R7689 VSS.n2676 VSS.n2650 9.3005
R7690 VSS.n2675 VSS.n2674 9.3005
R7691 VSS.n2673 VSS.n2651 9.3005
R7692 VSS.n2670 VSS.n2669 9.3005
R7693 VSS.n2668 VSS.n2654 9.3005
R7694 VSS.n2667 VSS.n2666 9.3005
R7695 VSS.n2665 VSS.n2655 9.3005
R7696 VSS.n2664 VSS.n2663 9.3005
R7697 VSS.n2083 VSS.n2082 9.3005
R7698 VSS.n3296 VSS.n3295 9.3005
R7699 VSS.n3306 VSS.n3305 9.3005
R7700 VSS.n3386 VSS.n2923 9.3005
R7701 VSS.n3393 VSS.n2919 9.3005
R7702 VSS.n3403 VSS.n3402 9.3005
R7703 VSS.n3404 VSS.n2915 9.3005
R7704 VSS.n3406 VSS.n3405 9.3005
R7705 VSS.n3408 VSS.n2913 9.3005
R7706 VSS.n3411 VSS.n3410 9.3005
R7707 VSS.n3412 VSS.n2912 9.3005
R7708 VSS.n3414 VSS.n3413 9.3005
R7709 VSS.n3415 VSS.n2910 9.3005
R7710 VSS.n3421 VSS.n3420 9.3005
R7711 VSS.n3423 VSS.n3422 9.3005
R7712 VSS.n3426 VSS.n3425 9.3005
R7713 VSS.n3433 VSS.n2903 9.3005
R7714 VSS.n3436 VSS.n2901 9.3005
R7715 VSS.n3444 VSS.n2898 9.3005
R7716 VSS.n3458 VSS.n3457 9.3005
R7717 VSS.n3463 VSS.n2787 9.3005
R7718 VSS.n3476 VSS.n3475 9.3005
R7719 VSS.n3480 VSS.n2781 9.3005
R7720 VSS.n3486 VSS.n2778 9.3005
R7721 VSS.n3489 VSS.n3488 9.3005
R7722 VSS.n3508 VSS.n2765 9.3005
R7723 VSS.n3513 VSS.n2761 9.3005
R7724 VSS.n3527 VSS.n3526 9.3005
R7725 VSS.n3531 VSS.n2755 9.3005
R7726 VSS.n3534 VSS.n3533 9.3005
R7727 VSS.n3547 VSS.n2747 9.3005
R7728 VSS.n3549 VSS.n3548 9.3005
R7729 VSS.n2872 VSS.n2871 9.3005
R7730 VSS.n2830 VSS.n2828 9.3005
R7731 VSS.n2824 VSS.n2802 9.3005
R7732 VSS.n2819 VSS.n2805 9.3005
R7733 VSS.n2816 VSS.n2806 9.3005
R7734 VSS.n2813 VSS.n2812 9.3005
R7735 VSS.n2818 VSS.n2817 9.3005
R7736 VSS.n2821 VSS.n2820 9.3005
R7737 VSS.n2826 VSS.n2825 9.3005
R7738 VSS.n2827 VSS.n2801 9.3005
R7739 VSS.n2831 VSS.n2800 9.3005
R7740 VSS.n2833 VSS.n2832 9.3005
R7741 VSS.n2834 VSS.n2799 9.3005
R7742 VSS.n2836 VSS.n2835 9.3005
R7743 VSS.n2837 VSS.n2798 9.3005
R7744 VSS.n2841 VSS.n2840 9.3005
R7745 VSS.n2842 VSS.n2797 9.3005
R7746 VSS.n2844 VSS.n2843 9.3005
R7747 VSS.n2847 VSS.n2794 9.3005
R7748 VSS.n2849 VSS.n2848 9.3005
R7749 VSS.n2850 VSS.n2793 9.3005
R7750 VSS.n2852 VSS.n2851 9.3005
R7751 VSS.n2853 VSS.n2792 9.3005
R7752 VSS.n2857 VSS.n2856 9.3005
R7753 VSS.n2858 VSS.n2791 9.3005
R7754 VSS.n2890 VSS.n2859 9.3005
R7755 VSS.n2888 VSS.n2887 9.3005
R7756 VSS.n2886 VSS.n2860 9.3005
R7757 VSS.n2885 VSS.n2884 9.3005
R7758 VSS.n2877 VSS.n2861 9.3005
R7759 VSS.n2875 VSS.n2874 9.3005
R7760 VSS.n2873 VSS.n2862 9.3005
R7761 VSS.n2870 VSS.n2863 9.3005
R7762 VSS.n2869 VSS.n2866 9.3005
R7763 VSS.n2868 VSS.n2867 9.3005
R7764 VSS.n2749 VSS.n2748 9.3005
R7765 VSS.n3546 VSS.n3545 9.3005
R7766 VSS.n3535 VSS.n2751 9.3005
R7767 VSS.n3532 VSS.n2753 9.3005
R7768 VSS.n3530 VSS.n3529 9.3005
R7769 VSS.n3528 VSS.n2757 9.3005
R7770 VSS.n3520 VSS.n2758 9.3005
R7771 VSS.n3519 VSS.n2759 9.3005
R7772 VSS.n3517 VSS.n3516 9.3005
R7773 VSS.n3515 VSS.n3514 9.3005
R7774 VSS.n3510 VSS.n3509 9.3005
R7775 VSS.n3507 VSS.n3506 9.3005
R7776 VSS.n3504 VSS.n2766 9.3005
R7777 VSS.n3503 VSS.n3502 9.3005
R7778 VSS.n3501 VSS.n3500 9.3005
R7779 VSS.n3498 VSS.n2770 9.3005
R7780 VSS.n3497 VSS.n3496 9.3005
R7781 VSS.n3495 VSS.n2771 9.3005
R7782 VSS.n3494 VSS.n3493 9.3005
R7783 VSS.n3492 VSS.n2772 9.3005
R7784 VSS.n3491 VSS.n3490 9.3005
R7785 VSS.n3487 VSS.n2775 9.3005
R7786 VSS.n3485 VSS.n3484 9.3005
R7787 VSS.n3483 VSS.n2780 9.3005
R7788 VSS.n3482 VSS.n3481 9.3005
R7789 VSS.n3479 VSS.n3478 9.3005
R7790 VSS.n3477 VSS.n2784 9.3005
R7791 VSS.n3470 VSS.n2785 9.3005
R7792 VSS.n3469 VSS.n3468 9.3005
R7793 VSS.n3467 VSS.n2786 9.3005
R7794 VSS.n3466 VSS.n3465 9.3005
R7795 VSS.n3461 VSS.n3460 9.3005
R7796 VSS.n3459 VSS.n2789 9.3005
R7797 VSS.n3455 VSS.n2790 9.3005
R7798 VSS.n3454 VSS.n2896 9.3005
R7799 VSS.n3453 VSS.n3452 9.3005
R7800 VSS.n3451 VSS.n2897 9.3005
R7801 VSS.n3450 VSS.n3449 9.3005
R7802 VSS.n3442 VSS.n2899 9.3005
R7803 VSS.n3441 VSS.n3440 9.3005
R7804 VSS.n3439 VSS.n2900 9.3005
R7805 VSS.n3438 VSS.n3437 9.3005
R7806 VSS.n3435 VSS.n3434 9.3005
R7807 VSS.n3432 VSS.n3431 9.3005
R7808 VSS.n3430 VSS.n2904 9.3005
R7809 VSS.n3429 VSS.n3428 9.3005
R7810 VSS.n3427 VSS.n2906 9.3005
R7811 VSS.n3424 VSS.n2907 9.3005
R7812 VSS.n3401 VSS.n2916 9.3005
R7813 VSS.n3399 VSS.n3398 9.3005
R7814 VSS.n3397 VSS.n2918 9.3005
R7815 VSS.n3396 VSS.n3395 9.3005
R7816 VSS.n3391 VSS.n3390 9.3005
R7817 VSS.n3389 VSS.n3388 9.3005
R7818 VSS.n3384 VSS.n3383 9.3005
R7819 VSS.n3382 VSS.n2925 9.3005
R7820 VSS.n3381 VSS.n3380 9.3005
R7821 VSS.n3379 VSS.n2926 9.3005
R7822 VSS.n3378 VSS.n3377 9.3005
R7823 VSS.n3376 VSS.n2927 9.3005
R7824 VSS.n3375 VSS.n3374 9.3005
R7825 VSS.n3373 VSS.n2928 9.3005
R7826 VSS.n3371 VSS.n3370 9.3005
R7827 VSS.n3369 VSS.n2931 9.3005
R7828 VSS.n3368 VSS.n3367 9.3005
R7829 VSS.n3366 VSS.n2932 9.3005
R7830 VSS.n3365 VSS.n3364 9.3005
R7831 VSS.n3363 VSS.n3362 9.3005
R7832 VSS.n3361 VSS.n2936 9.3005
R7833 VSS.n3360 VSS.n3359 9.3005
R7834 VSS.n3358 VSS.n2938 9.3005
R7835 VSS.n3357 VSS.n3356 9.3005
R7836 VSS.n3354 VSS.n2939 9.3005
R7837 VSS.n3353 VSS.n2943 9.3005
R7838 VSS.n3352 VSS.n3351 9.3005
R7839 VSS.n3350 VSS.n2944 9.3005
R7840 VSS.n3349 VSS.n3348 9.3005
R7841 VSS.n3346 VSS.n2945 9.3005
R7842 VSS.n3344 VSS.n2948 9.3005
R7843 VSS.n3343 VSS.n3342 9.3005
R7844 VSS.n3341 VSS.n3340 9.3005
R7845 VSS.n3339 VSS.n2950 9.3005
R7846 VSS.n3338 VSS.n3337 9.3005
R7847 VSS.n3336 VSS.n3335 9.3005
R7848 VSS.n3333 VSS.n2953 9.3005
R7849 VSS.n3332 VSS.n3331 9.3005
R7850 VSS.n3330 VSS.n3329 9.3005
R7851 VSS.n3328 VSS.n2957 9.3005
R7852 VSS.n3325 VSS.n3324 9.3005
R7853 VSS.n3323 VSS.n3322 9.3005
R7854 VSS.n3317 VSS.n2959 9.3005
R7855 VSS.n3316 VSS.n3315 9.3005
R7856 VSS.n3314 VSS.n2961 9.3005
R7857 VSS.n3313 VSS.n3312 9.3005
R7858 VSS.n3310 VSS.n2962 9.3005
R7859 VSS.n3308 VSS.n3307 9.3005
R7860 VSS.n3301 VSS.n2964 9.3005
R7861 VSS.n3299 VSS.n3298 9.3005
R7862 VSS.n3297 VSS.n2967 9.3005
R7863 VSS.n2969 VSS.n2968 9.3005
R7864 VSS.n3247 VSS.n3246 9.3005
R7865 VSS.n3249 VSS.n3248 9.3005
R7866 VSS.n3250 VSS.n3240 9.3005
R7867 VSS.n3253 VSS.n3252 9.3005
R7868 VSS.n3255 VSS.n3254 9.3005
R7869 VSS.n3256 VSS.n3238 9.3005
R7870 VSS.n3258 VSS.n3257 9.3005
R7871 VSS.n3259 VSS.n3237 9.3005
R7872 VSS.n3261 VSS.n3260 9.3005
R7873 VSS.n3263 VSS.n3235 9.3005
R7874 VSS.n3265 VSS.n3264 9.3005
R7875 VSS.n3267 VSS.n3266 9.3005
R7876 VSS.n3044 VSS.n3043 9.3005
R7877 VSS.n3045 VSS.n3037 9.3005
R7878 VSS.n3047 VSS.n3046 9.3005
R7879 VSS.n3049 VSS.n3034 9.3005
R7880 VSS.n3051 VSS.n3050 9.3005
R7881 VSS.n3052 VSS.n3032 9.3005
R7882 VSS.n3055 VSS.n3030 9.3005
R7883 VSS.n3057 VSS.n3056 9.3005
R7884 VSS.n3058 VSS.n3029 9.3005
R7885 VSS.n3060 VSS.n3059 9.3005
R7886 VSS.n3061 VSS.n3026 9.3005
R7887 VSS.n3063 VSS.n3062 9.3005
R7888 VSS.n3064 VSS.n3025 9.3005
R7889 VSS.n3066 VSS.n3065 9.3005
R7890 VSS.n3068 VSS.n3023 9.3005
R7891 VSS.n3070 VSS.n3069 9.3005
R7892 VSS.n3071 VSS.n3022 9.3005
R7893 VSS.n3074 VSS.n3072 9.3005
R7894 VSS.n3075 VSS.n3020 9.3005
R7895 VSS.n3078 VSS.n3077 9.3005
R7896 VSS.n3079 VSS.n3019 9.3005
R7897 VSS.n3081 VSS.n3080 9.3005
R7898 VSS.n3086 VSS.n3017 9.3005
R7899 VSS.n3089 VSS.n3088 9.3005
R7900 VSS.n3090 VSS.n3016 9.3005
R7901 VSS.n3092 VSS.n3091 9.3005
R7902 VSS.n3093 VSS.n3015 9.3005
R7903 VSS.n3095 VSS.n3094 9.3005
R7904 VSS.n3096 VSS.n3014 9.3005
R7905 VSS.n3098 VSS.n3097 9.3005
R7906 VSS.n3101 VSS.n3012 9.3005
R7907 VSS.n3105 VSS.n3104 9.3005
R7908 VSS.n3106 VSS.n3009 9.3005
R7909 VSS.n3108 VSS.n3107 9.3005
R7910 VSS.n3109 VSS.n3008 9.3005
R7911 VSS.n3112 VSS.n3111 9.3005
R7912 VSS.n3113 VSS.n3007 9.3005
R7913 VSS.n3115 VSS.n3114 9.3005
R7914 VSS.n3116 VSS.n3006 9.3005
R7915 VSS.n3119 VSS.n3118 9.3005
R7916 VSS.n3121 VSS.n3120 9.3005
R7917 VSS.n3122 VSS.n3003 9.3005
R7918 VSS.n3124 VSS.n3123 9.3005
R7919 VSS.n3126 VSS.n3125 9.3005
R7920 VSS.n3127 VSS.n3000 9.3005
R7921 VSS.n3132 VSS.n3131 9.3005
R7922 VSS.n3133 VSS.n2999 9.3005
R7923 VSS.n3135 VSS.n3134 9.3005
R7924 VSS.n3136 VSS.n2998 9.3005
R7925 VSS.n3138 VSS.n3137 9.3005
R7926 VSS.n3139 VSS.n2997 9.3005
R7927 VSS.n3141 VSS.n3140 9.3005
R7928 VSS.n3142 VSS.n2995 9.3005
R7929 VSS.n3145 VSS.n3144 9.3005
R7930 VSS.n3147 VSS.n3146 9.3005
R7931 VSS.n3149 VSS.n2991 9.3005
R7932 VSS.n3154 VSS.n3153 9.3005
R7933 VSS.n3155 VSS.n2990 9.3005
R7934 VSS.n3157 VSS.n3156 9.3005
R7935 VSS.n3160 VSS.n2989 9.3005
R7936 VSS.n3164 VSS.n3163 9.3005
R7937 VSS.n3165 VSS.n2988 9.3005
R7938 VSS.n3167 VSS.n3166 9.3005
R7939 VSS.n3169 VSS.n2987 9.3005
R7940 VSS.n3173 VSS.n3172 9.3005
R7941 VSS.n3174 VSS.n2986 9.3005
R7942 VSS.n3176 VSS.n3175 9.3005
R7943 VSS.n3177 VSS.n2985 9.3005
R7944 VSS.n3179 VSS.n3178 9.3005
R7945 VSS.n3180 VSS.n2984 9.3005
R7946 VSS.n3182 VSS.n3181 9.3005
R7947 VSS.n3187 VSS.n2982 9.3005
R7948 VSS.n3189 VSS.n3188 9.3005
R7949 VSS.n3190 VSS.n2981 9.3005
R7950 VSS.n3192 VSS.n3191 9.3005
R7951 VSS.n3193 VSS.n2978 9.3005
R7952 VSS.n3196 VSS.n3195 9.3005
R7953 VSS.n3198 VSS.n3197 9.3005
R7954 VSS.n3200 VSS.n2976 9.3005
R7955 VSS.n3202 VSS.n3201 9.3005
R7956 VSS.n3203 VSS.n2975 9.3005
R7957 VSS.n3205 VSS.n3204 9.3005
R7958 VSS.n3206 VSS.n2974 9.3005
R7959 VSS.n3209 VSS.n3208 9.3005
R7960 VSS.n3210 VSS.n2973 9.3005
R7961 VSS.n3212 VSS.n3211 9.3005
R7962 VSS.n3213 VSS.n2971 9.3005
R7963 VSS.n3215 VSS.n3214 9.3005
R7964 VSS.n3216 VSS.n2970 9.3005
R7965 VSS.n3292 VSS.n3217 9.3005
R7966 VSS.n3291 VSS.n3218 9.3005
R7967 VSS.n3290 VSS.n3289 9.3005
R7968 VSS.n3288 VSS.n3287 9.3005
R7969 VSS.n3286 VSS.n3221 9.3005
R7970 VSS.n3284 VSS.n3283 9.3005
R7971 VSS.n3282 VSS.n3281 9.3005
R7972 VSS.n3280 VSS.n3225 9.3005
R7973 VSS.n3278 VSS.n3228 9.3005
R7974 VSS.n3277 VSS.n3276 9.3005
R7975 VSS.n3275 VSS.n3274 9.3005
R7976 VSS.n3273 VSS.n3230 9.3005
R7977 VSS.n3272 VSS.n3271 9.3005
R7978 VSS.n3270 VSS.n3269 9.3005
R7979 VSS.n3268 VSS.n3233 9.3005
R7980 VSS.n3054 VSS.n3053 9.3005
R7981 VSS.n970 VSS.n969 9.3005
R7982 VSS.n971 VSS.n963 9.3005
R7983 VSS.n973 VSS.n972 9.3005
R7984 VSS.n975 VSS.n960 9.3005
R7985 VSS.n982 VSS.n981 9.3005
R7986 VSS.n983 VSS.n959 9.3005
R7987 VSS.n1715 VSS.n958 9.3005
R7988 VSS.n1714 VSS.n1713 9.3005
R7989 VSS.n1712 VSS.n984 9.3005
R7990 VSS.n1709 VSS.n1708 9.3005
R7991 VSS.n1705 VSS.n1704 9.3005
R7992 VSS.n1703 VSS.n991 9.3005
R7993 VSS.n1700 VSS.n1699 9.3005
R7994 VSS.n1698 VSS.n992 9.3005
R7995 VSS.n1697 VSS.n1696 9.3005
R7996 VSS.n1695 VSS.n993 9.3005
R7997 VSS.n1693 VSS.n1692 9.3005
R7998 VSS.n1691 VSS.n1690 9.3005
R7999 VSS.n1689 VSS.n997 9.3005
R8000 VSS.n1688 VSS.n1687 9.3005
R8001 VSS.n1686 VSS.n999 9.3005
R8002 VSS.n1685 VSS.n1684 9.3005
R8003 VSS.n1683 VSS.n1000 9.3005
R8004 VSS.n1682 VSS.n1681 9.3005
R8005 VSS.n1680 VSS.n1001 9.3005
R8006 VSS.n1679 VSS.n1678 9.3005
R8007 VSS.n1676 VSS.n1002 9.3005
R8008 VSS.n1675 VSS.n1674 9.3005
R8009 VSS.n1673 VSS.n1003 9.3005
R8010 VSS.n1672 VSS.n1671 9.3005
R8011 VSS.n1670 VSS.n1005 9.3005
R8012 VSS.n1669 VSS.n1668 9.3005
R8013 VSS.n1667 VSS.n1007 9.3005
R8014 VSS.n1666 VSS.n1665 9.3005
R8015 VSS.n1664 VSS.n1008 9.3005
R8016 VSS.n1663 VSS.n1662 9.3005
R8017 VSS.n1661 VSS.n1012 9.3005
R8018 VSS.n1660 VSS.n1659 9.3005
R8019 VSS.n1657 VSS.n1013 9.3005
R8020 VSS.n1655 VSS.n1654 9.3005
R8021 VSS.n1653 VSS.n1015 9.3005
R8022 VSS.n1652 VSS.n1651 9.3005
R8023 VSS.n1650 VSS.n1016 9.3005
R8024 VSS.n1649 VSS.n1647 9.3005
R8025 VSS.n1646 VSS.n1017 9.3005
R8026 VSS.n1645 VSS.n1644 9.3005
R8027 VSS.n1642 VSS.n1018 9.3005
R8028 VSS.n1640 VSS.n1639 9.3005
R8029 VSS.n1638 VSS.n1020 9.3005
R8030 VSS.n1637 VSS.n1636 9.3005
R8031 VSS.n1635 VSS.n1021 9.3005
R8032 VSS.n1633 VSS.n1632 9.3005
R8033 VSS.n1631 VSS.n1022 9.3005
R8034 VSS.n1630 VSS.n1629 9.3005
R8035 VSS.n1628 VSS.n1024 9.3005
R8036 VSS.n1627 VSS.n1026 9.3005
R8037 VSS.n1051 VSS.n1025 9.3005
R8038 VSS.n1053 VSS.n1052 9.3005
R8039 VSS.n1054 VSS.n1050 9.3005
R8040 VSS.n1056 VSS.n1055 9.3005
R8041 VSS.n1057 VSS.n1047 9.3005
R8042 VSS.n1060 VSS.n1059 9.3005
R8043 VSS.n1061 VSS.n1046 9.3005
R8044 VSS.n1063 VSS.n1062 9.3005
R8045 VSS.n1064 VSS.n1044 9.3005
R8046 VSS.n1068 VSS.n1067 9.3005
R8047 VSS.n1069 VSS.n1043 9.3005
R8048 VSS.n1071 VSS.n1070 9.3005
R8049 VSS.n1072 VSS.n1042 9.3005
R8050 VSS.n1074 VSS.n1073 9.3005
R8051 VSS.n1075 VSS.n1041 9.3005
R8052 VSS.n1077 VSS.n1076 9.3005
R8053 VSS.n1078 VSS.n1039 9.3005
R8054 VSS.n1079 VSS.n1036 9.3005
R8055 VSS.n1081 VSS.n1080 9.3005
R8056 VSS.n1082 VSS.n1035 9.3005
R8057 VSS.n1084 VSS.n1083 9.3005
R8058 VSS.n1086 VSS.n1033 9.3005
R8059 VSS.n1089 VSS.n1088 9.3005
R8060 VSS.n1090 VSS.n1032 9.3005
R8061 VSS.n1092 VSS.n1091 9.3005
R8062 VSS.n1093 VSS.n1030 9.3005
R8063 VSS.n1096 VSS.n1095 9.3005
R8064 VSS.n1624 VSS.n1623 9.3005
R8065 VSS.n1622 VSS.n1029 9.3005
R8066 VSS.n1621 VSS.n1620 9.3005
R8067 VSS.n1618 VSS.n1097 9.3005
R8068 VSS.n1617 VSS.n1616 9.3005
R8069 VSS.n1615 VSS.n1099 9.3005
R8070 VSS.n1614 VSS.n1613 9.3005
R8071 VSS.n1612 VSS.n1100 9.3005
R8072 VSS.n1610 VSS.n1609 9.3005
R8073 VSS.n1608 VSS.n1101 9.3005
R8074 VSS.n1607 VSS.n1606 9.3005
R8075 VSS.n1103 VSS.n1102 9.3005
R8076 VSS.n1600 VSS.n1599 9.3005
R8077 VSS.n1598 VSS.n1104 9.3005
R8078 VSS.n1597 VSS.n1596 9.3005
R8079 VSS.n1595 VSS.n1105 9.3005
R8080 VSS.n1594 VSS.n1592 9.3005
R8081 VSS.n1591 VSS.n1106 9.3005
R8082 VSS.n1590 VSS.n1589 9.3005
R8083 VSS.n1587 VSS.n1107 9.3005
R8084 VSS.n1586 VSS.n1585 9.3005
R8085 VSS.n1584 VSS.n1583 9.3005
R8086 VSS.n1579 VSS.n1111 9.3005
R8087 VSS.n1578 VSS.n1577 9.3005
R8088 VSS.n1576 VSS.n1575 9.3005
R8089 VSS.n1574 VSS.n1113 9.3005
R8090 VSS.n1573 VSS.n1572 9.3005
R8091 VSS.n1571 VSS.n1115 9.3005
R8092 VSS.n1570 VSS.n1569 9.3005
R8093 VSS.n1118 VSS.n1117 9.3005
R8094 VSS.n1520 VSS.n1519 9.3005
R8095 VSS.n1522 VSS.n1521 9.3005
R8096 VSS.n1523 VSS.n1517 9.3005
R8097 VSS.n1525 VSS.n1524 9.3005
R8098 VSS.n1526 VSS.n1516 9.3005
R8099 VSS.n1528 VSS.n1527 9.3005
R8100 VSS.n1529 VSS.n1515 9.3005
R8101 VSS.n1530 VSS.n1513 9.3005
R8102 VSS.n1532 VSS.n1531 9.3005
R8103 VSS.n1534 VSS.n1533 9.3005
R8104 VSS.n1536 VSS.n1510 9.3005
R8105 VSS.n1538 VSS.n1537 9.3005
R8106 VSS.n1539 VSS.n1509 9.3005
R8107 VSS.n1541 VSS.n1540 9.3005
R8108 VSS.n1542 VSS.n1507 9.3005
R8109 VSS.n1543 VSS.n1506 9.3005
R8110 VSS.n1546 VSS.n1545 9.3005
R8111 VSS.n1548 VSS.n1547 9.3005
R8112 VSS.n1549 VSS.n1503 9.3005
R8113 VSS.n1551 VSS.n1550 9.3005
R8114 VSS.n1552 VSS.n1502 9.3005
R8115 VSS.n1554 VSS.n1553 9.3005
R8116 VSS.n1557 VSS.n1498 9.3005
R8117 VSS.n1561 VSS.n1560 9.3005
R8118 VSS.n1562 VSS.n1497 9.3005
R8119 VSS.n1564 VSS.n1563 9.3005
R8120 VSS.n1566 VSS.n1495 9.3005
R8121 VSS.n1494 VSS.n1120 9.3005
R8122 VSS.n1493 VSS.n1492 9.3005
R8123 VSS.n1491 VSS.n1121 9.3005
R8124 VSS.n1489 VSS.n1488 9.3005
R8125 VSS.n1487 VSS.n1486 9.3005
R8126 VSS.n1485 VSS.n1124 9.3005
R8127 VSS.n1484 VSS.n1482 9.3005
R8128 VSS.n1481 VSS.n1126 9.3005
R8129 VSS.n1480 VSS.n1479 9.3005
R8130 VSS.n1478 VSS.n1127 9.3005
R8131 VSS.n1477 VSS.n1476 9.3005
R8132 VSS.n1475 VSS.n1474 9.3005
R8133 VSS.n1473 VSS.n1130 9.3005
R8134 VSS.n1472 VSS.n1471 9.3005
R8135 VSS.n1470 VSS.n1134 9.3005
R8136 VSS.n1469 VSS.n1468 9.3005
R8137 VSS.n1467 VSS.n1135 9.3005
R8138 VSS.n1466 VSS.n1465 9.3005
R8139 VSS.n1464 VSS.n1136 9.3005
R8140 VSS.n1463 VSS.n1462 9.3005
R8141 VSS.n1138 VSS.n1137 9.3005
R8142 VSS.n1457 VSS.n1456 9.3005
R8143 VSS.n1455 VSS.n1140 9.3005
R8144 VSS.n1454 VSS.n1453 9.3005
R8145 VSS.n1452 VSS.n1141 9.3005
R8146 VSS.n1451 VSS.n1449 9.3005
R8147 VSS.n1448 VSS.n1142 9.3005
R8148 VSS.n1447 VSS.n1446 9.3005
R8149 VSS.n1144 VSS.n1143 9.3005
R8150 VSS.n1400 VSS.n1399 9.3005
R8151 VSS.n1402 VSS.n1401 9.3005
R8152 VSS.n1404 VSS.n1396 9.3005
R8153 VSS.n1406 VSS.n1405 9.3005
R8154 VSS.n1408 VSS.n1407 9.3005
R8155 VSS.n1409 VSS.n1393 9.3005
R8156 VSS.n1411 VSS.n1410 9.3005
R8157 VSS.n1413 VSS.n1412 9.3005
R8158 VSS.n1414 VSS.n1390 9.3005
R8159 VSS.n1416 VSS.n1415 9.3005
R8160 VSS.n1417 VSS.n1389 9.3005
R8161 VSS.n1419 VSS.n1418 9.3005
R8162 VSS.n1420 VSS.n1388 9.3005
R8163 VSS.n1421 VSS.n1386 9.3005
R8164 VSS.n1422 VSS.n1385 9.3005
R8165 VSS.n1424 VSS.n1423 9.3005
R8166 VSS.n1425 VSS.n1384 9.3005
R8167 VSS.n1427 VSS.n1426 9.3005
R8168 VSS.n1429 VSS.n1381 9.3005
R8169 VSS.n1431 VSS.n1430 9.3005
R8170 VSS.n1432 VSS.n1380 9.3005
R8171 VSS.n1434 VSS.n1433 9.3005
R8172 VSS.n1437 VSS.n1377 9.3005
R8173 VSS.n1439 VSS.n1438 9.3005
R8174 VSS.n1440 VSS.n1376 9.3005
R8175 VSS.n1442 VSS.n1441 9.3005
R8176 VSS.n1443 VSS.n1374 9.3005
R8177 VSS.n1373 VSS.n1145 9.3005
R8178 VSS.n1372 VSS.n1371 9.3005
R8179 VSS.n1370 VSS.n1146 9.3005
R8180 VSS.n1369 VSS.n1368 9.3005
R8181 VSS.n1367 VSS.n1147 9.3005
R8182 VSS.n1366 VSS.n1365 9.3005
R8183 VSS.n1364 VSS.n1149 9.3005
R8184 VSS.n1363 VSS.n1362 9.3005
R8185 VSS.n1361 VSS.n1150 9.3005
R8186 VSS.n1360 VSS.n1359 9.3005
R8187 VSS.n1358 VSS.n1151 9.3005
R8188 VSS.n1356 VSS.n1355 9.3005
R8189 VSS.n1354 VSS.n1156 9.3005
R8190 VSS.n1353 VSS.n1352 9.3005
R8191 VSS.n1351 VSS.n1157 9.3005
R8192 VSS.n1349 VSS.n1348 9.3005
R8193 VSS.n1347 VSS.n1346 9.3005
R8194 VSS.n1345 VSS.n1159 9.3005
R8195 VSS.n1344 VSS.n1343 9.3005
R8196 VSS.n1342 VSS.n1164 9.3005
R8197 VSS.n1341 VSS.n1340 9.3005
R8198 VSS.n1339 VSS.n1165 9.3005
R8199 VSS.n1338 VSS.n1337 9.3005
R8200 VSS.n1336 VSS.n1335 9.3005
R8201 VSS.n1334 VSS.n1168 9.3005
R8202 VSS.n1333 VSS.n1332 9.3005
R8203 VSS.n1331 VSS.n1171 9.3005
R8204 VSS.n1330 VSS.n1329 9.3005
R8205 VSS.n1174 VSS.n1172 9.3005
R8206 VSS.n1206 VSS.n1204 9.3005
R8207 VSS.n1207 VSS.n1203 9.3005
R8208 VSS.n1209 VSS.n1208 9.3005
R8209 VSS.n1210 VSS.n1202 9.3005
R8210 VSS.n1212 VSS.n1211 9.3005
R8211 VSS.n1213 VSS.n1201 9.3005
R8212 VSS.n1214 VSS.n1200 9.3005
R8213 VSS.n1216 VSS.n1215 9.3005
R8214 VSS.n1218 VSS.n1217 9.3005
R8215 VSS.n1219 VSS.n1197 9.3005
R8216 VSS.n1222 VSS.n1221 9.3005
R8217 VSS.n1228 VSS.n1227 9.3005
R8218 VSS.n1232 VSS.n1231 9.3005
R8219 VSS.n1190 VSS.n1189 9.3005
R8220 VSS.n1241 VSS.n1240 9.3005
R8221 VSS.n1242 VSS.n1187 9.3005
R8222 VSS.n1244 VSS.n1243 9.3005
R8223 VSS.n1245 VSS.n1186 9.3005
R8224 VSS.n1247 VSS.n1246 9.3005
R8225 VSS.n1248 VSS.n1183 9.3005
R8226 VSS.n1249 VSS.n1181 9.3005
R8227 VSS.n1251 VSS.n1250 9.3005
R8228 VSS.n1252 VSS.n1180 9.3005
R8229 VSS.n1254 VSS.n1253 9.3005
R8230 VSS.n1255 VSS.n1178 9.3005
R8231 VSS.n1257 VSS.n1256 9.3005
R8232 VSS.n1326 VSS.n1325 9.3005
R8233 VSS.n1324 VSS.n1177 9.3005
R8234 VSS.n1323 VSS.n1322 9.3005
R8235 VSS.n1319 VSS.n1258 9.3005
R8236 VSS.n1318 VSS.n1317 9.3005
R8237 VSS.n1316 VSS.n1260 9.3005
R8238 VSS.n1315 VSS.n1314 9.3005
R8239 VSS.n1311 VSS.n1310 9.3005
R8240 VSS.n1309 VSS.n1308 9.3005
R8241 VSS.n1307 VSS.n1264 9.3005
R8242 VSS.n1305 VSS.n1304 9.3005
R8243 VSS.n1303 VSS.n1302 9.3005
R8244 VSS.n1300 VSS.n1266 9.3005
R8245 VSS.n1271 VSS.n1269 9.3005
R8246 VSS.n1295 VSS.n1294 9.3005
R8247 VSS.n1293 VSS.n1270 9.3005
R8248 VSS.n1292 VSS.n1291 9.3005
R8249 VSS.n1290 VSS.n1272 9.3005
R8250 VSS.n1289 VSS.n1275 9.3005
R8251 VSS.n1288 VSS.n1287 9.3005
R8252 VSS.n1286 VSS.n1278 9.3005
R8253 VSS.n1285 VSS.n1284 9.3005
R8254 VSS.n1717 VSS.n1716 9.3005
R8255 VSS.n4009 VSS.n4008 9.3005
R8256 VSS.n4007 VSS.n4001 9.3005
R8257 VSS.n4006 VSS.n4005 9.3005
R8258 VSS.n4010 VSS.n3998 9.3005
R8259 VSS.n4011 VSS.n3939 9.3005
R8260 VSS.n1826 VSS.n1822 9.3005
R8261 VSS.n1828 VSS.n1827 9.3005
R8262 VSS.n1830 VSS.n1829 9.3005
R8263 VSS.n1831 VSS.n1819 9.3005
R8264 VSS.n1833 VSS.n1832 9.3005
R8265 VSS.n1835 VSS.n1834 9.3005
R8266 VSS.n1838 VSS.n1817 9.3005
R8267 VSS.n1841 VSS.n1840 9.3005
R8268 VSS.n1842 VSS.n1816 9.3005
R8269 VSS.n1844 VSS.n1843 9.3005
R8270 VSS.n1845 VSS.n1814 9.3005
R8271 VSS.n1877 VSS.n1876 9.3005
R8272 VSS.n1875 VSS.n1815 9.3005
R8273 VSS.n1874 VSS.n1873 9.3005
R8274 VSS.n1872 VSS.n1871 9.3005
R8275 VSS.n1848 VSS.n1847 9.3005
R8276 VSS.n1865 VSS.n1864 9.3005
R8277 VSS.n1863 VSS.n1851 9.3005
R8278 VSS.n1862 VSS.n1861 9.3005
R8279 VSS.n1860 VSS.n1852 9.3005
R8280 VSS.n1859 VSS.n1858 9.3005
R8281 VSS.n4761 VSS.n1882 9.3005
R8282 VSS.n4758 VSS.n4736 9.3005
R8283 VSS.n4755 VSS.n4737 9.3005
R8284 VSS.n4749 VSS.n4748 9.3005
R8285 VSS.n4747 VSS.n4739 9.3005
R8286 VSS.n4750 VSS.n4738 9.3005
R8287 VSS.n4752 VSS.n4751 9.3005
R8288 VSS.n4757 VSS.n4756 9.3005
R8289 VSS.n4760 VSS.n4759 9.3005
R8290 VSS.n4763 VSS.n4762 9.3005
R8291 VSS.n1900 VSS.n1894 9.3005
R8292 VSS.n1902 VSS.n1901 9.3005
R8293 VSS.n1904 VSS.n1903 9.3005
R8294 VSS.n1905 VSS.n1890 9.3005
R8295 VSS.n1908 VSS.n1907 9.3005
R8296 VSS.n1909 VSS.n1889 9.3005
R8297 VSS.n1911 VSS.n1910 9.3005
R8298 VSS.n1913 VSS.n1886 9.3005
R8299 VSS.n1915 VSS.n1914 9.3005
R8300 VSS.n1917 VSS.n1916 9.3005
R8301 VSS.n1918 VSS.n1881 9.3005
R8302 VSS.n4096 VSS.n4091 9.3005
R8303 VSS.n4098 VSS.n4097 9.3005
R8304 VSS.n4099 VSS.n4090 9.3005
R8305 VSS.n4101 VSS.n4100 9.3005
R8306 VSS.n4102 VSS.n4088 9.3005
R8307 VSS.n4104 VSS.n4103 9.3005
R8308 VSS.n4105 VSS.n4087 9.3005
R8309 VSS.n4107 VSS.n4106 9.3005
R8310 VSS.n4108 VSS.n4085 9.3005
R8311 VSS.n4109 VSS.n4084 9.3005
R8312 VSS.n4063 VSS.n4059 9.3005
R8313 VSS.n4065 VSS.n4064 9.3005
R8314 VSS.n4067 VSS.n4066 9.3005
R8315 VSS.n4068 VSS.n4056 9.3005
R8316 VSS.n4071 VSS.n4070 9.3005
R8317 VSS.n4072 VSS.n4055 9.3005
R8318 VSS.n4074 VSS.n4073 9.3005
R8319 VSS.n4076 VSS.n4053 9.3005
R8320 VSS.n4080 VSS.n4079 9.3005
R8321 VSS.n4081 VSS.n4052 9.3005
R8322 VSS.n4083 VSS.n4082 9.3005
R8323 VSS.n4795 VSS.n1777 9.3005
R8324 VSS.n4792 VSS.n4768 9.3005
R8325 VSS.n4787 VSS.n4771 9.3005
R8326 VSS.n4783 VSS.n4782 9.3005
R8327 VSS.n4781 VSS.n4773 9.3005
R8328 VSS.n4784 VSS.n4772 9.3005
R8329 VSS.n4786 VSS.n4785 9.3005
R8330 VSS.n4789 VSS.n4788 9.3005
R8331 VSS.n4794 VSS.n4793 9.3005
R8332 VSS.n1795 VSS.n1794 9.3005
R8333 VSS.n1796 VSS.n1786 9.3005
R8334 VSS.n1799 VSS.n1798 9.3005
R8335 VSS.n1800 VSS.n1785 9.3005
R8336 VSS.n1802 VSS.n1801 9.3005
R8337 VSS.n1804 VSS.n1784 9.3005
R8338 VSS.n1806 VSS.n1805 9.3005
R8339 VSS.n1808 VSS.n1807 9.3005
R8340 VSS.n1809 VSS.n1778 9.3005
R8341 VSS.n1812 VSS.n1811 9.3005
R8342 VSS.n1813 VSS.n1776 9.3005
R8343 VSS.n4797 VSS.n4796 9.3005
R8344 VSS.n4906 VSS.n4905 9.3005
R8345 VSS.n4904 VSS.n4901 9.3005
R8346 VSS.n3725 VSS.n3719 9.3005
R8347 VSS.n3724 VSS.n3723 9.3005
R8348 VSS.n3722 VSS.n3720 9.3005
R8349 VSS.n3727 VSS.n3726 9.3005
R8350 VSS.n4690 VSS.n4689 9.3005
R8351 VSS.n4692 VSS.n4691 9.3005
R8352 VSS.n3797 VSS.n3794 9.3005
R8353 VSS.n3800 VSS.n3799 9.3005
R8354 VSS.n3801 VSS.n3793 9.3005
R8355 VSS.n3803 VSS.n3802 9.3005
R8356 VSS.n3804 VSS.n3792 9.3005
R8357 VSS.n3805 VSS.n3789 9.3005
R8358 VSS.n3807 VSS.n3806 9.3005
R8359 VSS.n3808 VSS.n3788 9.3005
R8360 VSS.n3810 VSS.n3809 9.3005
R8361 VSS.n3811 VSS.n3787 9.3005
R8362 VSS.n3786 VSS.n3729 9.3005
R8363 VSS.n3785 VSS.n3784 9.3005
R8364 VSS.n3783 VSS.n3730 9.3005
R8365 VSS.n3782 VSS.n3781 9.3005
R8366 VSS.n3780 VSS.n3731 9.3005
R8367 VSS.n3779 VSS.n3778 9.3005
R8368 VSS.n3777 VSS.n3732 9.3005
R8369 VSS.n3776 VSS.n3775 9.3005
R8370 VSS.n3774 VSS.n3735 9.3005
R8371 VSS.n3773 VSS.n3772 9.3005
R8372 VSS.n3771 VSS.n3736 9.3005
R8373 VSS.n3768 VSS.n3767 9.3005
R8374 VSS.n3766 VSS.n3737 9.3005
R8375 VSS.n3765 VSS.n3764 9.3005
R8376 VSS.n3763 VSS.n3738 9.3005
R8377 VSS.n3762 VSS.n3761 9.3005
R8378 VSS.n3760 VSS.n3739 9.3005
R8379 VSS.n3759 VSS.n3758 9.3005
R8380 VSS.n3757 VSS.n3740 9.3005
R8381 VSS.n3755 VSS.n3754 9.3005
R8382 VSS.n3753 VSS.n3741 9.3005
R8383 VSS.n3752 VSS.n3751 9.3005
R8384 VSS.n3750 VSS.n3742 9.3005
R8385 VSS.n3749 VSS.n3748 9.3005
R8386 VSS.n3747 VSS.n3743 9.3005
R8387 VSS.n3746 VSS.n3745 9.3005
R8388 VSS.n3711 VSS.n3710 9.3005
R8389 VSS.n4304 VSS.n4303 9.3005
R8390 VSS.n4305 VSS.n3709 9.3005
R8391 VSS.n4307 VSS.n4306 9.3005
R8392 VSS.n4308 VSS.n3708 9.3005
R8393 VSS.n4309 VSS.n3706 9.3005
R8394 VSS.n4311 VSS.n4310 9.3005
R8395 VSS.n4312 VSS.n3705 9.3005
R8396 VSS.n4314 VSS.n4313 9.3005
R8397 VSS.n4315 VSS.n3703 9.3005
R8398 VSS.n4316 VSS.n3701 9.3005
R8399 VSS.n4318 VSS.n4317 9.3005
R8400 VSS.n4319 VSS.n3700 9.3005
R8401 VSS.n4321 VSS.n4320 9.3005
R8402 VSS.n4322 VSS.n3699 9.3005
R8403 VSS.n4324 VSS.n4323 9.3005
R8404 VSS.n4325 VSS.n3698 9.3005
R8405 VSS.n4327 VSS.n4326 9.3005
R8406 VSS.n4328 VSS.n3697 9.3005
R8407 VSS.n4330 VSS.n4329 9.3005
R8408 VSS.n4331 VSS.n3696 9.3005
R8409 VSS.n4333 VSS.n4332 9.3005
R8410 VSS.n4334 VSS.n3695 9.3005
R8411 VSS.n4335 VSS.n3693 9.3005
R8412 VSS.n4337 VSS.n4336 9.3005
R8413 VSS.n4338 VSS.n3692 9.3005
R8414 VSS.n4340 VSS.n4339 9.3005
R8415 VSS.n4341 VSS.n3690 9.3005
R8416 VSS.n4343 VSS.n4342 9.3005
R8417 VSS.n4344 VSS.n3689 9.3005
R8418 VSS.n4346 VSS.n4345 9.3005
R8419 VSS.n4347 VSS.n3687 9.3005
R8420 VSS.n4349 VSS.n4348 9.3005
R8421 VSS.n4350 VSS.n3686 9.3005
R8422 VSS.n4352 VSS.n4351 9.3005
R8423 VSS.n4353 VSS.n3684 9.3005
R8424 VSS.n4355 VSS.n4354 9.3005
R8425 VSS.n4356 VSS.n3683 9.3005
R8426 VSS.n4358 VSS.n4357 9.3005
R8427 VSS.n4359 VSS.n3682 9.3005
R8428 VSS.n4361 VSS.n4360 9.3005
R8429 VSS.n4362 VSS.n3681 9.3005
R8430 VSS.n4364 VSS.n4363 9.3005
R8431 VSS.n4365 VSS.n3679 9.3005
R8432 VSS.n4368 VSS.n4367 9.3005
R8433 VSS.n4369 VSS.n3678 9.3005
R8434 VSS.n4371 VSS.n4370 9.3005
R8435 VSS.n4372 VSS.n3677 9.3005
R8436 VSS.n4374 VSS.n4373 9.3005
R8437 VSS.n4376 VSS.n4375 9.3005
R8438 VSS.n4377 VSS.n3674 9.3005
R8439 VSS.n4380 VSS.n4379 9.3005
R8440 VSS.n4381 VSS.n3673 9.3005
R8441 VSS.n4383 VSS.n4382 9.3005
R8442 VSS.n4385 VSS.n3671 9.3005
R8443 VSS.n4387 VSS.n4386 9.3005
R8444 VSS.n4389 VSS.n4388 9.3005
R8445 VSS.n4390 VSS.n3669 9.3005
R8446 VSS.n4391 VSS.n3666 9.3005
R8447 VSS.n4393 VSS.n4392 9.3005
R8448 VSS.n4394 VSS.n3665 9.3005
R8449 VSS.n4396 VSS.n4395 9.3005
R8450 VSS.n4397 VSS.n3663 9.3005
R8451 VSS.n4399 VSS.n4398 9.3005
R8452 VSS.n4400 VSS.n3662 9.3005
R8453 VSS.n4402 VSS.n4401 9.3005
R8454 VSS.n4403 VSS.n3661 9.3005
R8455 VSS.n4404 VSS.n3659 9.3005
R8456 VSS.n4406 VSS.n4405 9.3005
R8457 VSS.n4407 VSS.n3658 9.3005
R8458 VSS.n4409 VSS.n4408 9.3005
R8459 VSS.n4410 VSS.n3657 9.3005
R8460 VSS.n4411 VSS.n3656 9.3005
R8461 VSS.n4413 VSS.n4412 9.3005
R8462 VSS.n4415 VSS.n4414 9.3005
R8463 VSS.n4416 VSS.n3652 9.3005
R8464 VSS.n4419 VSS.n4418 9.3005
R8465 VSS.n4420 VSS.n3651 9.3005
R8466 VSS.n4422 VSS.n4421 9.3005
R8467 VSS.n4423 VSS.n3650 9.3005
R8468 VSS.n4425 VSS.n4424 9.3005
R8469 VSS.n4426 VSS.n3649 9.3005
R8470 VSS.n4428 VSS.n4427 9.3005
R8471 VSS.n4429 VSS.n3647 9.3005
R8472 VSS.n4431 VSS.n4430 9.3005
R8473 VSS.n4432 VSS.n3646 9.3005
R8474 VSS.n4434 VSS.n4433 9.3005
R8475 VSS.n4435 VSS.n3644 9.3005
R8476 VSS.n4437 VSS.n4436 9.3005
R8477 VSS.n4438 VSS.n3643 9.3005
R8478 VSS.n4440 VSS.n4439 9.3005
R8479 VSS.n4441 VSS.n3642 9.3005
R8480 VSS.n4443 VSS.n4442 9.3005
R8481 VSS.n4444 VSS.n3641 9.3005
R8482 VSS.n4446 VSS.n4445 9.3005
R8483 VSS.n4447 VSS.n3639 9.3005
R8484 VSS.n4449 VSS.n4448 9.3005
R8485 VSS.n4450 VSS.n3638 9.3005
R8486 VSS.n4452 VSS.n4451 9.3005
R8487 VSS.n4453 VSS.n3637 9.3005
R8488 VSS.n4455 VSS.n4454 9.3005
R8489 VSS.n4456 VSS.n3636 9.3005
R8490 VSS.n4458 VSS.n4457 9.3005
R8491 VSS.n4459 VSS.n3634 9.3005
R8492 VSS.n4461 VSS.n4460 9.3005
R8493 VSS.n4462 VSS.n3633 9.3005
R8494 VSS.n4464 VSS.n4463 9.3005
R8495 VSS.n4465 VSS.n3632 9.3005
R8496 VSS.n4466 VSS.n3630 9.3005
R8497 VSS.n4468 VSS.n4467 9.3005
R8498 VSS.n4469 VSS.n3629 9.3005
R8499 VSS.n4471 VSS.n4470 9.3005
R8500 VSS.n4472 VSS.n3627 9.3005
R8501 VSS.n4474 VSS.n4473 9.3005
R8502 VSS.n4475 VSS.n3626 9.3005
R8503 VSS.n4477 VSS.n4476 9.3005
R8504 VSS.n4479 VSS.n3624 9.3005
R8505 VSS.n4483 VSS.n4482 9.3005
R8506 VSS.n4484 VSS.n3623 9.3005
R8507 VSS.n4486 VSS.n4485 9.3005
R8508 VSS.n4487 VSS.n3622 9.3005
R8509 VSS.n4488 VSS.n3620 9.3005
R8510 VSS.n4490 VSS.n4489 9.3005
R8511 VSS.n4491 VSS.n3619 9.3005
R8512 VSS.n4493 VSS.n4492 9.3005
R8513 VSS.n4494 VSS.n3617 9.3005
R8514 VSS.n4496 VSS.n4495 9.3005
R8515 VSS.n4497 VSS.n3616 9.3005
R8516 VSS.n4499 VSS.n4498 9.3005
R8517 VSS.n4500 VSS.n3615 9.3005
R8518 VSS.n4501 VSS.n3613 9.3005
R8519 VSS.n4503 VSS.n4502 9.3005
R8520 VSS.n4504 VSS.n3612 9.3005
R8521 VSS.n4506 VSS.n4505 9.3005
R8522 VSS.n4508 VSS.n3611 9.3005
R8523 VSS.n4511 VSS.n4510 9.3005
R8524 VSS.n4513 VSS.n4512 9.3005
R8525 VSS.n4514 VSS.n3609 9.3005
R8526 VSS.n4516 VSS.n4515 9.3005
R8527 VSS.n4517 VSS.n3608 9.3005
R8528 VSS.n4519 VSS.n4518 9.3005
R8529 VSS.n4520 VSS.n3606 9.3005
R8530 VSS.n4521 VSS.n3604 9.3005
R8531 VSS.n4523 VSS.n4522 9.3005
R8532 VSS.n4524 VSS.n3603 9.3005
R8533 VSS.n4526 VSS.n4525 9.3005
R8534 VSS.n4527 VSS.n3602 9.3005
R8535 VSS.n4528 VSS.n3601 9.3005
R8536 VSS.n4530 VSS.n4529 9.3005
R8537 VSS.n4531 VSS.n3600 9.3005
R8538 VSS.n4533 VSS.n4532 9.3005
R8539 VSS.n4534 VSS.n3598 9.3005
R8540 VSS.n4536 VSS.n4535 9.3005
R8541 VSS.n4537 VSS.n3597 9.3005
R8542 VSS.n4539 VSS.n4538 9.3005
R8543 VSS.n4540 VSS.n3595 9.3005
R8544 VSS.n4542 VSS.n4541 9.3005
R8545 VSS.n4543 VSS.n3594 9.3005
R8546 VSS.n4545 VSS.n4544 9.3005
R8547 VSS.n4547 VSS.n3592 9.3005
R8548 VSS.n4549 VSS.n4548 9.3005
R8549 VSS.n4551 VSS.n4550 9.3005
R8550 VSS.n4552 VSS.n3589 9.3005
R8551 VSS.n4554 VSS.n4553 9.3005
R8552 VSS.n4555 VSS.n3588 9.3005
R8553 VSS.n4557 VSS.n4556 9.3005
R8554 VSS.n4558 VSS.n3587 9.3005
R8555 VSS.n4560 VSS.n4559 9.3005
R8556 VSS.n4561 VSS.n3585 9.3005
R8557 VSS.n4564 VSS.n3584 9.3005
R8558 VSS.n4566 VSS.n4565 9.3005
R8559 VSS.n4567 VSS.n3583 9.3005
R8560 VSS.n4569 VSS.n4568 9.3005
R8561 VSS.n4570 VSS.n3581 9.3005
R8562 VSS.n4572 VSS.n4571 9.3005
R8563 VSS.n4573 VSS.n3580 9.3005
R8564 VSS.n4575 VSS.n4574 9.3005
R8565 VSS.n4576 VSS.n3579 9.3005
R8566 VSS.n4580 VSS.n4579 9.3005
R8567 VSS.n4581 VSS.n3578 9.3005
R8568 VSS.n4583 VSS.n4582 9.3005
R8569 VSS.n4586 VSS.n3577 9.3005
R8570 VSS.n4588 VSS.n4587 9.3005
R8571 VSS.n4589 VSS.n3576 9.3005
R8572 VSS.n4591 VSS.n4590 9.3005
R8573 VSS.n4593 VSS.n3575 9.3005
R8574 VSS.n4595 VSS.n4594 9.3005
R8575 VSS.n4596 VSS.n3574 9.3005
R8576 VSS.n4598 VSS.n4597 9.3005
R8577 VSS.n4599 VSS.n3573 9.3005
R8578 VSS.n4601 VSS.n4600 9.3005
R8579 VSS.n4602 VSS.n3572 9.3005
R8580 VSS.n4604 VSS.n4603 9.3005
R8581 VSS.n4605 VSS.n3570 9.3005
R8582 VSS.n4608 VSS.n4607 9.3005
R8583 VSS.n4609 VSS.n3568 9.3005
R8584 VSS.n4611 VSS.n4610 9.3005
R8585 VSS.n4612 VSS.n3567 9.3005
R8586 VSS.n4614 VSS.n4613 9.3005
R8587 VSS.n4615 VSS.n3566 9.3005
R8588 VSS.n4617 VSS.n4616 9.3005
R8589 VSS.n4618 VSS.n3564 9.3005
R8590 VSS.n4620 VSS.n4619 9.3005
R8591 VSS.n4621 VSS.n3563 9.3005
R8592 VSS.n4623 VSS.n4622 9.3005
R8593 VSS.n4625 VSS.n3561 9.3005
R8594 VSS.n4627 VSS.n4626 9.3005
R8595 VSS.n4628 VSS.n3560 9.3005
R8596 VSS.n4630 VSS.n4629 9.3005
R8597 VSS.n4631 VSS.n3558 9.3005
R8598 VSS.n4634 VSS.n4633 9.3005
R8599 VSS.n1927 VSS.n1926 9.3005
R8600 VSS.n4647 VSS.n4646 9.3005
R8601 VSS.n4648 VSS.n1925 9.3005
R8602 VSS.n4651 VSS.n4650 9.3005
R8603 VSS.n4652 VSS.n1924 9.3005
R8604 VSS.n4654 VSS.n4653 9.3005
R8605 VSS.n4655 VSS.n1923 9.3005
R8606 VSS.n4657 VSS.n4656 9.3005
R8607 VSS.n4658 VSS.n1922 9.3005
R8608 VSS.n4660 VSS.n4659 9.3005
R8609 VSS.n4661 VSS.n1921 9.3005
R8610 VSS.n4664 VSS.n4663 9.3005
R8611 VSS.n4665 VSS.n1920 9.3005
R8612 VSS.n4730 VSS.n4666 9.3005
R8613 VSS.n4729 VSS.n4667 9.3005
R8614 VSS.n4728 VSS.n4727 9.3005
R8615 VSS.n4726 VSS.n4669 9.3005
R8616 VSS.n4725 VSS.n4724 9.3005
R8617 VSS.n4723 VSS.n4670 9.3005
R8618 VSS.n4722 VSS.n4721 9.3005
R8619 VSS.n4720 VSS.n4672 9.3005
R8620 VSS.n4719 VSS.n4718 9.3005
R8621 VSS.n4717 VSS.n4673 9.3005
R8622 VSS.n4716 VSS.n4715 9.3005
R8623 VSS.n4714 VSS.n4675 9.3005
R8624 VSS.n4713 VSS.n4712 9.3005
R8625 VSS.n4711 VSS.n4676 9.3005
R8626 VSS.n4710 VSS.n4709 9.3005
R8627 VSS.n4708 VSS.n4678 9.3005
R8628 VSS.n4707 VSS.n4706 9.3005
R8629 VSS.n4705 VSS.n4679 9.3005
R8630 VSS.n4704 VSS.n4703 9.3005
R8631 VSS.n4702 VSS.n4681 9.3005
R8632 VSS.n4701 VSS.n4700 9.3005
R8633 VSS.n4699 VSS.n4682 9.3005
R8634 VSS.n4698 VSS.n4697 9.3005
R8635 VSS.n4696 VSS.n4684 9.3005
R8636 VSS.n4695 VSS.n4694 9.3005
R8637 VSS.n4693 VSS.n4685 9.3005
R8638 VSS.n4563 VSS.n4562 9.3005
R8639 VSS.n4129 VSS.n4128 9.3005
R8640 VSS.n4126 VSS.n4114 9.3005
R8641 VSS.n4124 VSS.n4123 9.3005
R8642 VSS.n4122 VSS.n4121 9.3005
R8643 VSS.n4119 VSS.n4118 9.3005
R8644 VSS.n4139 VSS.n4112 9.3005
R8645 VSS.n4163 VSS.n4162 9.3005
R8646 VSS.n4164 VSS.n3935 9.3005
R8647 VSS.n4166 VSS.n4165 9.3005
R8648 VSS.n3605 VSS.t1752 9.054
R8649 VSS.n824 VSS.n823 9.03579
R8650 VSS.n530 VSS.n527 9.03579
R8651 VSS.n2230 VSS.n2229 9.03579
R8652 VSS.n2616 VSS.n2601 9.03579
R8653 VSS.n3192 VSS.n2981 9.03579
R8654 VSS.n3208 VSS.n2973 9.03579
R8655 VSS.n1560 VSS.n1559 9.03579
R8656 VSS.n3982 VSS.n3974 8.88145
R8657 VSS.n3868 VSS.n3820 8.88145
R8658 VSS.n4279 VSS.n3905 8.86414
R8659 VSS.n4279 VSS.n4278 8.86414
R8660 VSS.n4204 VSS.n4203 8.86414
R8661 VSS.n3986 VSS.n3974 8.8249
R8662 VSS.n3868 VSS.n3867 8.8249
R8663 VSS.n598 VSS.n596 8.78481
R8664 VSS.n2198 VSS.n2197 8.64611
R8665 VSS.n4187 VSS.n3913 8.64324
R8666 VSS.n4187 VSS.n4186 8.64324
R8667 VSS.n4176 VSS.n3922 8.64324
R8668 VSS.n4003 VSS.n4002 8.58762
R8669 VSS.n4012 VSS.n3997 8.55042
R8670 VSS.n3983 VSS.n3982 8.54514
R8671 VSS.n3862 VSS.n3820 8.54514
R8672 VSS.n2313 VSS.n2310 8.53383
R8673 VSS.n2460 VSS.n2457 8.53383
R8674 VSS.n2555 VSS.n2552 8.53383
R8675 VSS.t3357 VSS.t3289 8.42962
R8676 VSS.t350 VSS.t567 8.42962
R8677 VSS.t377 VSS.t3620 8.42962
R8678 VSS.t3602 VSS.t51 8.42962
R8679 VSS.t929 VSS.t1832 8.42962
R8680 VSS.t447 VSS.t411 8.42962
R8681 VSS.t445 VSS.t409 8.42962
R8682 VSS.t1988 VSS.t1073 8.42962
R8683 VSS.t3614 VSS.t2826 8.42962
R8684 VSS.t3622 VSS.t142 8.42962
R8685 VSS.t144 VSS.t2670 8.42962
R8686 VSS.t1131 VSS.t2608 8.42962
R8687 VSS.t3600 VSS.t2210 8.42962
R8688 VSS.t2125 VSS.t2946 8.42962
R8689 VSS.t2216 VSS.t1137 8.42962
R8690 VSS.t2875 VSS.t1135 8.42962
R8691 VSS.t3273 VSS.t1375 8.42962
R8692 VSS.t3275 VSS.t3671 8.42962
R8693 VSS.n3714 VSS.n3713 8.32651
R8694 VSS.n865 VSS.n864 8.28285
R8695 VSS.n763 VSS.n762 8.28285
R8696 VSS.n662 VSS.n661 8.28285
R8697 VSS.n581 VSS.n580 8.28285
R8698 VSS.n2703 VSS.n2702 8.28285
R8699 VSS.n1215 VSS.n1199 8.28285
R8700 VSS.n1484 VSS.n1126 8.28285
R8701 VSS.n1619 VSS.n1618 8.28285
R8702 VSS.n1694 VSS.n1693 8.28285
R8703 VSS.n3264 VSS.n3263 8.23546
R8704 VSS.n3261 VSS.n3237 8.23546
R8705 VSS.n3257 VSS.n3237 8.23546
R8706 VSS.n3257 VSS.n3256 8.23546
R8707 VSS.n3256 VSS.n3255 8.23546
R8708 VSS.n3250 VSS.n3249 8.23546
R8709 VSS.n4185 VSS.n3922 8.20563
R8710 VSS.n19 VSS.n17 8.10717
R8711 VSS.n3244 VSS.n3242 8.10717
R8712 VSS.n1582 VSS.n1581 8.10717
R8713 VSS.n349 VSS.n346 8.05976
R8714 VSS.n2424 VSS.n2421 8.05976
R8715 VSS.n3525 VSS.n3522 8.05976
R8716 VSS.n3085 VSS.n3082 8.05976
R8717 VSS.n1162 VSS.n1158 8.05976
R8718 VSS.n931 VSS.n930 8.0482
R8719 VSS.n5050 VSS.n5049 7.90638
R8720 VSS.n917 VSS.n329 7.90638
R8721 VSS.n773 VSS.n438 7.90638
R8722 VSS.n699 VSS.n698 7.90638
R8723 VSS.n641 VSS.n640 7.90638
R8724 VSS.n562 VSS.n9 7.90638
R8725 VSS.n5422 VSS.n5421 7.90638
R8726 VSS.n2150 VSS.n2147 7.90638
R8727 VSS.n2693 VSS.n2692 7.90638
R8728 VSS.n2686 VSS.n2685 7.90638
R8729 VSS.n2839 VSS.n2837 7.90638
R8730 VSS.n2846 VSS.n2844 7.90638
R8731 VSS.n2856 VSS.n2855 7.90638
R8732 VSS.n3373 VSS.n3372 7.90638
R8733 VSS.n3171 VSS.n2986 7.90638
R8734 VSS.n1066 VSS.n1043 7.90638
R8735 VSS.n4366 VSS.n4365 7.90638
R8736 VSS.n3264 VSS.n3234 7.6984
R8737 VSS.n3249 VSS.n3241 7.6984
R8738 VSS.n4195 VSS.t1807 7.60243
R8739 VSS.n3304 VSS.n2966 7.6005
R8740 VSS.n2164 VSS.n2158 7.52991
R8741 VSS.n2223 VSS.n2032 7.52991
R8742 VSS.n1344 VSS.n1164 7.52991
R8743 VSS.n1574 VSS.n1573 7.52991
R8744 VSS.n4219 VSS.n3880 7.26779
R8745 VSS.n4161 VSS.n3938 7.16275
R8746 VSS.n952 VSS.n951 7.15344
R8747 VSS.n865 VSS.n363 7.15344
R8748 VSS.n2086 VSS.n2057 7.15344
R8749 VSS.n1633 VSS.n1022 7.15344
R8750 VSS.n4004 VSS.n4003 7.15034
R8751 VSS.n404 VSS.n401 7.11161
R8752 VSS.n3715 VSS.n3714 7.02466
R8753 VSS.n854 VSS.n853 6.77697
R8754 VSS.n554 VSS.n552 6.77697
R8755 VSS.n2889 VSS.n2888 6.77697
R8756 VSS.n3517 VSS.n2760 6.77697
R8757 VSS.n3500 VSS.n2769 6.77697
R8758 VSS.n3394 VSS.n3393 6.77697
R8759 VSS.n3343 VSS.n2949 6.77697
R8760 VSS.n3153 VSS.n3152 6.77697
R8761 VSS.n3277 VSS.n3229 6.77697
R8762 VSS.n4378 VSS.n3673 6.77697
R8763 VSS.n5461 VSS.n5460 6.7747
R8764 VSS.n2489 VSS.n1985 6.63754
R8765 VSS.n4095 VSS.n4094 6.5783
R8766 VSS.n4746 VSS.n4743 6.57826
R8767 VSS.n4780 VSS.n4779 6.57826
R8768 VSS.n1857 VSS.n1855 6.57825
R8769 VSS.n4817 VSS.n4816 6.57154
R8770 VSS.n3850 VSS.n3840 6.57154
R8771 VSS.n2138 VSS.n2135 6.52992
R8772 VSS.n3252 VSS.n3251 6.44526
R8773 VSS.n5200 VSS.n164 6.4005
R8774 VSS.n5164 VSS.n5163 6.4005
R8775 VSS.n5138 VSS.n5137 6.4005
R8776 VSS.n884 VSS.n883 6.4005
R8777 VSS.n2258 VSS.n2016 6.4005
R8778 VSS.n2304 VSS.n2274 6.4005
R8779 VSS.n2526 VSS.n2525 6.4005
R8780 VSS.n2725 VSS.n1942 6.4005
R8781 VSS.n3335 VSS.n3334 6.4005
R8782 VSS.n3111 VSS.n3007 6.4005
R8783 VSS.n3160 VSS.n3159 6.4005
R8784 VSS.n3183 VSS.n2983 6.4005
R8785 VSS.n1428 VSS.n1427 6.4005
R8786 VSS.n1408 VSS.n1395 6.4005
R8787 VSS.n1080 VSS.n1079 6.4005
R8788 VSS.n4551 VSS.n3591 6.4005
R8789 VSS.n4481 VSS.n3623 6.4005
R8790 VSS.n4412 VSS.n3655 6.4005
R8791 VSS.n3770 VSS.n3768 6.4005
R8792 VSS.n3778 VSS.n3734 6.4005
R8793 VSS.n4579 VSS.n4578 6.4005
R8794 VSS.n81 VSS.n80 6.26433
R8795 VSS.n5184 VSS.n5183 6.26433
R8796 VSS.n5184 VSS.n169 6.26433
R8797 VSS.n5146 VSS.n5145 6.26433
R8798 VSS.n5146 VSS.n185 6.26433
R8799 VSS.n5113 VSS.n5112 6.26433
R8800 VSS.n4977 VSS.n4976 6.26433
R8801 VSS.n4977 VSS.n269 6.26433
R8802 VSS.n946 VSS.n945 6.26433
R8803 VSS.n831 VSS.n388 6.26433
R8804 VSS.n686 VSS.n685 6.26433
R8805 VSS.n5468 VSS.n13 6.26433
R8806 VSS.n5436 VSS.n5435 6.26433
R8807 VSS.n3410 VSS.n2912 6.26433
R8808 VSS.n3312 VSS.n2961 6.26433
R8809 VSS.n1579 VSS.n1578 6.26433
R8810 VSS.n1844 VSS.n1816 6.26433
R8811 VSS.n1845 VSS.n1844 6.26433
R8812 VSS.n1876 VSS.n1845 6.26433
R8813 VSS.n1876 VSS.n1875 6.26433
R8814 VSS.n4510 VSS.n4508 6.26433
R8815 VSS.n4141 VSS.n4140 6.21883
R8816 VSS.n4117 VSS.n4116 6.21725
R8817 VSS.n1763 VSS.n1761 6.21725
R8818 VSS.n4837 VSS.n4836 6.20545
R8819 VSS.n944 VSS.n943 6.12816
R8820 VSS.t2637 VSS.t154 6.09468
R8821 VSS.n4281 VSS.t2344 6.09468
R8822 VSS.n5382 VSS.n5379 6.02403
R8823 VSS.n2229 VSS.n2227 6.02403
R8824 VSS.n2236 VSS.n2025 6.02403
R8825 VSS.n2571 VSS.n2569 6.02403
R8826 VSS.n1468 VSS.n1134 6.02403
R8827 VSS.n1559 VSS.n1497 6.02403
R8828 VSS.n1556 VSS.n1555 6.02403
R8829 VSS.n3844 VSS.n3843 6.0005
R8830 VSS.n4819 VSS.n4818 6.0005
R8831 VSS.n4816 VSS.n4815 5.99811
R8832 VSS.n3850 VSS.n3849 5.99811
R8833 VSS.n46 VSS.n45 5.98311
R8834 VSS.n5331 VSS.n5330 5.98311
R8835 VSS.n5244 VSS.n5243 5.98311
R8836 VSS.n5121 VSS.n5119 5.98311
R8837 VSS.n5079 VSS.n5076 5.98311
R8838 VSS.n4925 VSS.n4922 5.98311
R8839 VSS.n307 VSS.n302 5.98311
R8840 VSS.n634 VSS.n523 5.98311
R8841 VSS.n2324 VSS.n2268 5.98311
R8842 VSS.n3449 VSS.n3445 5.98311
R8843 VSS.n3301 VSS.n3300 5.98311
R8844 VSS.n981 VSS.n976 5.98311
R8845 VSS.n1835 VSS.n1818 5.98311
R8846 VSS.n3798 VSS.n3797 5.98311
R8847 VSS.n4689 VSS.n4686 5.98311
R8848 VSS.n4816 VSS.n4809 5.92155
R8849 VSS.n3851 VSS.n3850 5.92155
R8850 VSS.n3443 VSS.n3442 5.88425
R8851 VSS.n81 VSS.n29 5.85582
R8852 VSS.n5183 VSS.n5182 5.85582
R8853 VSS.n5145 VSS.n5144 5.85582
R8854 VSS.n5112 VSS.n5111 5.85582
R8855 VSS.n4976 VSS.n4975 5.85582
R8856 VSS.n687 VSS.n686 5.85582
R8857 VSS.n5457 VSS.n20 5.85582
R8858 VSS.n5438 VSS.n5385 5.85582
R8859 VSS.n2298 VSS.n2276 5.85582
R8860 VSS.n3408 VSS.n3407 5.85582
R8861 VSS.n3310 VSS.n3309 5.85582
R8862 VSS.n1221 VSS.n1220 5.85582
R8863 VSS.n1580 VSS.n1579 5.85582
R8864 VSS.n1839 VSS.n1816 5.85582
R8865 VSS.n4508 VSS.n4507 5.85582
R8866 VSS.n946 VSS.n317 5.78773
R8867 VSS.n5188 VSS.n169 5.65809
R8868 VSS.n5150 VSS.n185 5.65809
R8869 VSS.n4981 VSS.n269 5.65809
R8870 VSS.n5435 VSS.n5387 5.65809
R8871 VSS.n3414 VSS.n2912 5.65809
R8872 VSS.n3316 VSS.n2961 5.65809
R8873 VSS.n873 VSS.n357 5.64756
R8874 VSS.n1875 VSS.n1874 5.60959
R8875 VSS.n4167 VSS.n3934 5.5751
R8876 VSS.n3981 VSS.n3980 5.48621
R8877 VSS.n3870 VSS.n3818 5.48621
R8878 VSS.n4743 VSS.n4742 5.47169
R8879 VSS.n4780 VSS.n4776 5.47169
R8880 VSS.n4898 VSS.n4897 5.438
R8881 VSS.n873 VSS.n872 5.27109
R8882 VSS.n806 VSS.n415 5.27109
R8883 VSS.n680 VSS.n679 5.27109
R8884 VSS.n654 VSS.n509 5.27109
R8885 VSS.n2103 VSS.n2052 5.27109
R8886 VSS.n2222 VSS.n2220 5.27109
R8887 VSS.n2233 VSS.n2029 5.27109
R8888 VSS.n2249 VSS.n2248 5.27109
R8889 VSS.n2471 VSS.n1996 5.27109
R8890 VSS.n2608 VSS.n2607 5.27109
R8891 VSS.n3457 VSS.n3456 5.27109
R8892 VSS.n3131 VSS.n3129 5.27109
R8893 VSS.n3195 VSS.n2977 5.27109
R8894 VSS.n1338 VSS.n1167 5.27109
R8895 VSS.n1335 VSS.n1170 5.27109
R8896 VSS.n1477 VSS.n1129 5.27109
R8897 VSS.n1474 VSS.n1132 5.27109
R8898 VSS.n1557 VSS.n1556 5.27109
R8899 VSS.n1535 VSS.n1534 5.27109
R8900 VSS.n1589 VSS.n1109 5.27109
R8901 VSS.n3895 VSS.n3894 5.22706
R8902 VSS.n3865 VSS.n3814 5.22371
R8903 VSS.n3872 VSS.n3814 5.22371
R8904 VSS.n3871 VSS.n3870 5.22371
R8905 VSS.n3872 VSS.n3871 5.22371
R8906 VSS.n3973 VSS.n3971 5.22371
R8907 VSS.n3975 VSS.n3971 5.22371
R8908 VSS.n3980 VSS.n3970 5.22371
R8909 VSS.n3975 VSS.n3970 5.22371
R8910 VSS.n292 VSS.n290 5.13108
R8911 VSS.n292 VSS.n291 5.13108
R8912 VSS.n5406 VSS.n5404 5.13108
R8913 VSS.n5406 VSS.n5405 5.13108
R8914 VSS.n2068 VSS.n2066 5.13108
R8915 VSS.n2068 VSS.n2067 5.13108
R8916 VSS.n2661 VSS.n2659 5.13108
R8917 VSS.n2661 VSS.n2660 5.13108
R8918 VSS.n3040 VSS.n3038 5.13108
R8919 VSS.n3040 VSS.n3039 5.13108
R8920 VSS.n2810 VSS.n2808 5.13108
R8921 VSS.n2810 VSS.n2809 5.13108
R8922 VSS.n986 VSS.n985 5.13108
R8923 VSS.n966 VSS.n964 5.13108
R8924 VSS.n966 VSS.n965 5.13108
R8925 VSS.n1313 VSS.n1262 5.13108
R8926 VSS.n1281 VSS.n1279 5.13108
R8927 VSS.n1281 VSS.n1280 5.13108
R8928 VSS.n3883 VSS.n3882 5.063
R8929 VSS.n3886 VSS.n3885 5.063
R8930 VSS.n5426 VSS.n5392 5.03644
R8931 VSS.n3424 VSS.n3423 5.03644
R8932 VSS.n3721 VSS.n1767 4.99908
R8933 VSS.n3312 VSS.n3311 4.90263
R8934 VSS.n910 VSS.n909 4.89462
R8935 VSS.n2566 VSS.n1960 4.89462
R8936 VSS.n2589 VSS.n2588 4.89462
R8937 VSS.n3985 VSS.n3984 4.8755
R8938 VSS.n5154 VSS.n5153 4.85762
R8939 VSS.n5192 VSS.n5191 4.85762
R8940 VSS.n4985 VSS.n4984 4.85762
R8941 VSS.n5429 VSS.n5391 4.85762
R8942 VSS.n937 VSS.n936 4.85762
R8943 VSS.n3320 VSS.n3319 4.85762
R8944 VSS.n3418 VSS.n3417 4.85762
R8945 VSS.n1298 VSS.n1267 4.85762
R8946 VSS.n3262 VSS.n3261 4.83407
R8947 VSS.n45 VSS.n44 4.8005
R8948 VSS.n5332 VSS.n5331 4.8005
R8949 VSS.n5245 VSS.n5244 4.8005
R8950 VSS.n5121 VSS.n5120 4.8005
R8951 VSS.n5079 VSS.n5078 4.8005
R8952 VSS.n4925 VSS.n4924 4.8005
R8953 VSS.n307 VSS.n306 4.8005
R8954 VSS.n634 VSS.n633 4.8005
R8955 VSS.n2324 VSS.n2323 4.8005
R8956 VSS.n3449 VSS.n3448 4.8005
R8957 VSS.n3302 VSS.n3301 4.8005
R8958 VSS.n981 VSS.n980 4.8005
R8959 VSS.n1836 VSS.n1835 4.8005
R8960 VSS.n3797 VSS.n3796 4.8005
R8961 VSS.n4689 VSS.n4688 4.8005
R8962 VSS.n3893 VSS.n3891 4.79738
R8963 VSS.n1221 VSS.n1196 4.76646
R8964 VSS.n294 VSS.n293 4.75748
R8965 VSS.n5408 VSS.n5407 4.75748
R8966 VSS.n2070 VSS.n2069 4.75748
R8967 VSS.n2662 VSS.n2658 4.75748
R8968 VSS.n3042 VSS.n3041 4.75748
R8969 VSS.n968 VSS.n967 4.75748
R8970 VSS.n1283 VSS.n1282 4.75748
R8971 VSS.n2811 VSS.n2807 4.75739
R8972 VSS.n4811 VSS.n4810 4.7489
R8973 VSS.n3842 VSS.n3841 4.7489
R8974 VSS.n2880 VSS.n2879 4.74124
R8975 VSS.n4807 VSS.n4802 4.6799
R8976 VSS.n3853 VSS.n3825 4.6799
R8977 VSS.n4803 VSS.n4802 4.58401
R8978 VSS.n3826 VSS.n3825 4.58401
R8979 VSS.n4813 VSS.n4810 4.57445
R8980 VSS.n3847 VSS.n3841 4.57445
R8981 VSS.n1606 VSS.n1604 4.55553
R8982 VSS.n339 VSS.n336 4.51815
R8983 VSS.n840 VSS.n839 4.51815
R8984 VSS.n2226 VSS.n2032 4.51815
R8985 VSS.n2478 VSS.n1991 4.51815
R8986 VSS.n2629 VSS.n2628 4.51815
R8987 VSS.n1436 VSS.n1435 4.51815
R8988 VSS.n1565 VSS.n1564 4.51815
R8989 VSS.n1058 VSS.n1057 4.51815
R8990 VSS.n5342 VSS.n5336 4.51401
R8991 VSS.n5346 VSS.n104 4.51401
R8992 VSS.n5487 VSS.n3 4.51401
R8993 VSS.n8 VSS.n7 4.51401
R8994 VSS.n2740 VSS.n1932 4.51401
R8995 VSS.n1937 VSS.n1936 4.51401
R8996 VSS.n3537 VSS.n3536 4.51401
R8997 VSS.n3551 VSS.n3550 4.51401
R8998 VSS.n1226 VSS.n1225 4.51401
R8999 VSS.n1239 VSS.n1238 4.51401
R9000 VSS.n4640 VSS.n3556 4.51401
R9001 VSS.n4645 VSS.n4644 4.51401
R9002 VSS.n4823 VSS.n4822 4.5005
R9003 VSS.n4820 VSS.n1770 4.5005
R9004 VSS.n4806 VSS.n4805 4.5005
R9005 VSS.n4809 VSS.n4808 4.5005
R9006 VSS.n4815 VSS.n4814 4.5005
R9007 VSS.n4812 VSS.n1775 4.5005
R9008 VSS.n3823 VSS.n3821 4.5005
R9009 VSS.n3859 VSS.n3858 4.5005
R9010 VSS.n3855 VSS.n3854 4.5005
R9011 VSS.n3852 VSS.n3851 4.5005
R9012 VSS.n3849 VSS.n3848 4.5005
R9013 VSS.n3846 VSS.n3845 4.5005
R9014 VSS.n5341 VSS.n5340 4.5005
R9015 VSS.n5337 VSS.n102 4.5005
R9016 VSS.n5348 VSS.n5347 4.5005
R9017 VSS.n5486 VSS.n5485 4.5005
R9018 VSS.n5484 VSS.n5483 4.5005
R9019 VSS.n5480 VSS.n5479 4.5005
R9020 VSS.n2739 VSS.n2738 4.5005
R9021 VSS.n2737 VSS.n2736 4.5005
R9022 VSS.n2733 VSS.n2732 4.5005
R9023 VSS.n3543 VSS.n3542 4.5005
R9024 VSS.n3544 VSS.n2746 4.5005
R9025 VSS.n3538 VSS.n2752 4.5005
R9026 VSS.n1223 VSS.n1194 4.5005
R9027 VSS.n1234 VSS.n1233 4.5005
R9028 VSS.n1195 VSS.n1191 4.5005
R9029 VSS.n4639 VSS.n4638 4.5005
R9030 VSS.n4637 VSS.n4636 4.5005
R9031 VSS.n3559 VSS.n1928 4.5005
R9032 VSS.n5470 VSS.n5469 4.49412
R9033 VSS.n3889 VSS.n3888 4.43994
R9034 VSS.n5363 VSS.n5359 4.35795
R9035 VSS.n5301 VSS.n122 4.35795
R9036 VSS.n5284 VSS.n128 4.35795
R9037 VSS.n5253 VSS.n143 4.35795
R9038 VSS.n925 VSS.n326 4.35795
R9039 VSS.n752 VSS.n450 4.35795
R9040 VSS.n704 VSS.n478 4.35795
R9041 VSS.n567 VSS.n560 4.35795
R9042 VSS.n2720 VSS.n1943 4.35795
R9043 VSS.n3475 VSS.n3474 4.35795
R9044 VSS.n1461 VSS.n1138 4.35795
R9045 VSS.n1604 VSS.n1103 4.35795
R9046 VSS.n5113 VSS.n201 4.28986
R9047 VSS.n4955 VSS.n276 4.26717
R9048 VSS.n591 VSS.n544 4.26717
R9049 VSS.n2391 VSS.n2390 4.26717
R9050 VSS.n4765 VSS.n1880 4.25685
R9051 VSS.n943 VSS.n318 4.22178
R9052 VSS.n832 VSS.n831 4.22178
R9053 VSS.n491 VSS.n488 4.15369
R9054 VSS.n2448 VSS.n2447 4.14168
R9055 VSS.n3255 VSS.n3239 4.11798
R9056 VSS.n3252 VSS.n3239 4.11798
R9057 VSS.n5116 VSS.n201 4.07323
R9058 VSS.n682 VSS.n491 4.07323
R9059 VSS.n990 VSS.n989 4.07323
R9060 VSS.n988 VSS.n986 4.07323
R9061 VSS.n1313 VSS.n1312 4.07323
R9062 VSS.n1865 VSS.n1851 4.03338
R9063 VSS.n1879 VSS.n1878 3.9555
R9064 VSS.n4765 VSS.n4764 3.9555
R9065 VSS.n4767 VSS.n4766 3.9555
R9066 VSS.n5456 VSS.n5455 3.94944
R9067 VSS.n3104 VSS.n3103 3.93896
R9068 VSS.n4219 VSS.n4212 3.91766
R9069 VSS.n2297 VSS.n2296 3.88135
R9070 VSS.t1055 VSS.t3187 3.88057
R9071 VSS.n5086 VSS.n214 3.76521
R9072 VSS.n2358 VSS.n2357 3.76521
R9073 VSS.n2503 VSS.n2502 3.76521
R9074 VSS.n1486 VSS.n1123 3.76521
R9075 VSS.n1087 VSS.n1086 3.76521
R9076 VSS.n5437 VSS.n5436 3.6771
R9077 VSS.n3410 VSS.n3409 3.6771
R9078 VSS.n3857 VSS.n3856 3.60014
R9079 VSS.n4804 VSS.n1772 3.59914
R9080 VSS.n1871 VSS.n1846 3.59502
R9081 VSS.n1866 VSS.n1848 3.59502
R9082 VSS.n2139 VSS.n2138 3.57367
R9083 VSS.n3862 VSS.n3861 3.51386
R9084 VSS.n5190 VSS.n5189 3.50735
R9085 VSS.n5152 VSS.n5151 3.50735
R9086 VSS.n4983 VSS.n4982 3.50735
R9087 VSS.n938 VSS.n321 3.50735
R9088 VSS.n5431 VSS.n5389 3.50735
R9089 VSS.n3416 VSS.n3415 3.50735
R9090 VSS.n3318 VSS.n3317 3.50735
R9091 VSS.n1308 VSS.n1307 3.44377
R9092 VSS.n7 VSS.n0 3.43925
R9093 VSS.n5488 VSS.n5487 3.43925
R9094 VSS.n1936 VSS.n1930 3.43925
R9095 VSS.n2741 VSS.n2740 3.43925
R9096 VSS.n1238 VSS.n1237 3.43925
R9097 VSS.n1225 VSS.n1224 3.43925
R9098 VSS.n4644 VSS.n4643 3.43925
R9099 VSS.n4641 VSS.n4640 3.43925
R9100 VSS.n4825 VSS.n1770 3.43394
R9101 VSS.n4824 VSS.n4823 3.43394
R9102 VSS.n3860 VSS.n3859 3.43394
R9103 VSS.n3821 VSS.n1769 3.43394
R9104 VSS.n4287 VSS.n3903 3.42526
R9105 VSS.n5345 VSS.n5344 3.4105
R9106 VSS.n5344 VSS.n5343 3.4105
R9107 VSS.n5346 VSS.n5345 3.4105
R9108 VSS.n5343 VSS.n5342 3.4105
R9109 VSS.n5338 VSS.n107 3.4105
R9110 VSS.n105 VSS.n103 3.4105
R9111 VSS.n4 VSS.n2 3.4105
R9112 VSS.n5482 VSS.n5481 3.4105
R9113 VSS.n1933 VSS.n1931 3.4105
R9114 VSS.n2735 VSS.n2734 3.4105
R9115 VSS.n3541 VSS.n2745 3.4105
R9116 VSS.n3552 VSS.n3551 3.4105
R9117 VSS.n3537 VSS.n2743 3.4105
R9118 VSS.n3540 VSS.n3539 3.4105
R9119 VSS.n1193 VSS.n1192 3.4105
R9120 VSS.n1236 VSS.n1235 3.4105
R9121 VSS.n3557 VSS.n3555 3.4105
R9122 VSS.n4635 VSS.n1929 3.4105
R9123 VSS.n3553 VSS.n3552 3.4105
R9124 VSS.n3553 VSS.n2743 3.4105
R9125 VSS.n3263 VSS.n3262 3.4019
R9126 VSS.n1312 VSS.n1311 3.40077
R9127 VSS.n2440 VSS.n2439 3.38874
R9128 VSS.n2521 VSS.n1975 3.38874
R9129 VSS.n3512 VSS.n3511 3.38874
R9130 VSS.n3334 VSS.n3333 3.38874
R9131 VSS.n3159 VSS.n3157 3.38874
R9132 VSS.n1912 VSS.n1911 3.38874
R9133 VSS.n4075 VSS.n4074 3.38874
R9134 VSS.n1805 VSS.n1783 3.38874
R9135 VSS.n4548 VSS.n3591 3.38874
R9136 VSS.n4482 VSS.n4481 3.38874
R9137 VSS.n4415 VSS.n3655 3.38874
R9138 VSS.n4578 VSS.n3578 3.38874
R9139 VSS.n2883 VSS.n2879 3.31902
R9140 VSS.n3856 VSS.n3855 3.29357
R9141 VSS.n4805 VSS.n4804 3.29357
R9142 VSS.n1308 VSS.n1263 3.21921
R9143 VSS.n1305 VSS.n1265 3.21921
R9144 VSS.n5194 VSS.n168 3.2005
R9145 VSS.n5156 VSS.n183 3.2005
R9146 VSS.n4987 VSS.n268 3.2005
R9147 VSS.n935 VSS.n934 3.2005
R9148 VSS.n5430 VSS.n5390 3.2005
R9149 VSS.n3420 VSS.n2911 3.2005
R9150 VSS.n3322 VSS.n2960 3.2005
R9151 VSS.n1299 VSS.n1269 3.2005
R9152 VSS.n80 VSS.n79 3.13241
R9153 VSS.n15 VSS.n13 3.13241
R9154 VSS.n5455 VSS.n5454 3.13241
R9155 VSS.n2296 VSS.n2295 3.13241
R9156 VSS.n1229 VSS.n1228 3.13241
R9157 VSS.n1578 VSS.n1112 3.13241
R9158 VSS.n4510 VSS.n4509 3.13241
R9159 VSS.n3726 VSS.n1720 3.08333
R9160 VSS.n683 VSS.n682 3.04861
R9161 VSS.n1707 VSS.n986 3.04861
R9162 VSS.n5116 VSS.n5115 3.04861
R9163 VSS.n1706 VSS.n990 3.04861
R9164 VSS.n1313 VSS.n1261 3.04861
R9165 VSS.n1452 VSS.n1451 3.01226
R9166 VSS.n4292 VSS.n3890 3.01194
R9167 VSS.n4288 VSS.n4287 2.82936
R9168 VSS.n4829 VSS.n1766 2.8242
R9169 VSS.n4153 VSS.n3941 2.82286
R9170 VSS.n1301 VSS.n1300 2.76214
R9171 VSS.n3984 VSS.n3983 2.7505
R9172 VSS.n79 VSS.n78 2.7239
R9173 VSS.n393 VSS.n392 2.7239
R9174 VSS.n16 VSS.n15 2.7239
R9175 VSS.n5454 VSS.n5453 2.7239
R9176 VSS.n2295 VSS.n2294 2.7239
R9177 VSS.n1230 VSS.n1229 2.7239
R9178 VSS.n1114 VSS.n1112 2.7239
R9179 VSS.n4509 VSS.n3610 2.7239
R9180 VSS.t2925 VSS.t2923 2.72243
R9181 VSS.t3574 VSS.t3569 2.72243
R9182 VSS.n5042 VSS.n236 2.63579
R9183 VSS.n930 VSS.n929 2.63579
R9184 VSS.n904 VSS.n339 2.63579
R9185 VSS.n736 VSS.n735 2.63579
R9186 VSS.n709 VSS.n476 2.63579
R9187 VSS.n661 VSS.n660 2.63579
R9188 VSS.n573 VSS.n572 2.63579
R9189 VSS.n2123 VSS.n2122 2.63579
R9190 VSS.n2171 VSS.n2170 2.63579
R9191 VSS.n2695 VSS.n2694 2.63579
R9192 VSS.n2848 VSS.n2796 2.63579
R9193 VSS.n2855 VSS.n2853 2.63579
R9194 VSS.n3401 VSS.n3400 2.63579
R9195 VSS.n3365 VSS.n2935 2.63579
R9196 VSS.n3335 VSS.n2952 2.63579
R9197 VSS.n3121 VSS.n3005 2.63579
R9198 VSS.n3163 VSS.n3162 2.63579
R9199 VSS.n3269 VSS.n3232 2.63579
R9200 VSS.n1410 VSS.n1392 2.63579
R9201 VSS.n1059 VSS.n1058 2.63579
R9202 VSS.n1665 VSS.n1010 2.63579
R9203 VSS.n1703 VSS.n1700 2.63579
R9204 VSS.n4373 VSS.n3676 2.63579
R9205 VSS.n3988 VSS.n3972 2.63064
R9206 VSS.n3864 VSS.n3863 2.63064
R9207 VSS.n5193 VSS.n166 2.63064
R9208 VSS.n5155 VSS.n184 2.63064
R9209 VSS.n4986 VSS.n266 2.63064
R9210 VSS.n324 VSS.n322 2.63064
R9211 VSS.n5428 VSS.n5427 2.63064
R9212 VSS.n3419 VSS.n2909 2.63064
R9213 VSS.n3321 VSS.n2958 2.63064
R9214 VSS.n1297 VSS.n1296 2.63064
R9215 VSS.n1853 VSS.n1850 2.63064
R9216 VSS.n3246 VSS.n3245 2.5963
R9217 VSS.n5438 VSS.n5437 2.58773
R9218 VSS.n3409 VSS.n3408 2.58773
R9219 VSS.n4841 VSS.n4837 2.5605
R9220 VSS.n4142 VSS.n4141 2.5605
R9221 VSS.n4154 VSS.n4153 2.55728
R9222 VSS.n3103 VSS.n3009 2.53237
R9223 VSS.n2298 VSS.n2297 2.38348
R9224 VSS.n4293 VSS.n3889 2.341
R9225 VSS.n5457 VSS.n5456 2.31539
R9226 VSS.n989 VSS.n988 2.31539
R9227 VSS.n756 VSS.n755 2.2967
R9228 VSS.n5091 VSS.n5090 2.25932
R9229 VSS.n781 VSS.n780 2.25932
R9230 VSS.n2243 VSS.n2242 2.25932
R9231 VSS.n2359 VSS.n2006 2.25932
R9232 VSS.n2519 VSS.n2518 2.25932
R9233 VSS.n2569 VSS.n2567 2.25932
R9234 VSS.n2610 VSS.n2609 2.25932
R9235 VSS.n3899 VSS.n3898 2.1939
R9236 VSS.n4167 VSS.n4166 2.1851
R9237 VSS.n890 VSS.n349 2.13383
R9238 VSS.n813 VSS.n407 2.13383
R9239 VSS.n2421 VSS.n2420 2.13383
R9240 VSS.n2496 VSS.n1985 2.13383
R9241 VSS.n2880 VSS.n2860 2.13383
R9242 VSS.n3522 VSS.n2757 2.13383
R9243 VSS.n3082 VSS.n3081 2.13383
R9244 VSS.n3183 VSS.n3182 2.13383
R9245 VSS.n1346 VSS.n1162 2.13383
R9246 VSS.n3305 VSS.n2963 2.01789
R9247 VSS.n1871 VSS.n1870 2.01694
R9248 VSS.n1870 VSS.n1848 2.01694
R9249 VSS.n5464 VSS.n5463 1.97497
R9250 VSS.n1583 VSS.n1110 1.97497
R9251 VSS.n4899 VSS.n1720 1.91915
R9252 VSS.n3328 VSS.n3327 1.91116
R9253 VSS.n392 VSS.n391 1.90688
R9254 VSS.n2310 VSS.n2309 1.8968
R9255 VSS.n2457 VSS.n2456 1.8968
R9256 VSS.n2556 VSS.n2555 1.8968
R9257 VSS.n5049 VSS.n5048 1.88285
R9258 VSS.n920 VSS.n329 1.88285
R9259 VSS.n438 VSS.n435 1.88285
R9260 VSS.n700 VSS.n699 1.88285
R9261 VSS.n563 VSS.n562 1.88285
R9262 VSS.n2114 VSS.n2113 1.88285
R9263 VSS.n2177 VSS.n2150 1.88285
R9264 VSS.n2164 VSS.n2163 1.88285
R9265 VSS.n2694 VSS.n2693 1.88285
R9266 VSS.n2687 VSS.n2686 1.88285
R9267 VSS.n2672 VSS.n2671 1.88285
R9268 VSS.n2823 VSS.n2822 1.88285
R9269 VSS.n2840 VSS.n2839 1.88285
R9270 VSS.n2847 VSS.n2846 1.88285
R9271 VSS.n3372 VSS.n3371 1.88285
R9272 VSS.n3129 VSS.n3127 1.88285
R9273 VSS.n3172 VSS.n3171 1.88285
R9274 VSS.n1086 VSS.n1085 1.88285
R9275 VSS.n1067 VSS.n1066 1.88285
R9276 VSS.n4367 VSS.n4366 1.88285
R9277 VSS.n5363 VSS.n5362 1.8161
R9278 VSS.n5304 VSS.n122 1.8161
R9279 VSS.n5287 VSS.n128 1.8161
R9280 VSS.n5256 VSS.n143 1.8161
R9281 VSS.n925 VSS.n924 1.8161
R9282 VSS.n755 VSS.n450 1.8161
R9283 VSS.n704 VSS.n703 1.8161
R9284 VSS.n564 VSS.n560 1.8161
R9285 VSS.n2720 VSS.n2719 1.8161
R9286 VSS.n3475 VSS.n3471 1.8161
R9287 VSS.n1458 VSS.n1138 1.8161
R9288 VSS.n1601 VSS.n1103 1.8161
R9289 VSS.n1307 VSS.n1306 1.79699
R9290 VSS.n3251 VSS.n3250 1.79071
R9291 VSS.n4854 VSS.n4853 1.78349
R9292 VSS.n4133 VSS.n3942 1.78349
R9293 VSS.n3987 VSS.n3973 1.77828
R9294 VSS.n3866 VSS.n3865 1.77828
R9295 VSS.n5344 VSS.n106 1.69188
R9296 VSS.n4643 VSS.n4642 1.69188
R9297 VSS.n4642 VSS.n4641 1.69188
R9298 VSS.n3553 VSS.n2744 1.69188
R9299 VSS.n2742 VSS.n1930 1.69188
R9300 VSS.n2742 VSS.n2741 1.69188
R9301 VSS.n1237 VSS.n1 1.69188
R9302 VSS.n1224 VSS.n1 1.69188
R9303 VSS.n5489 VSS.n0 1.69188
R9304 VSS.n5489 VSS.n5488 1.69188
R9305 VSS.n2197 VSS.n2194 1.68471
R9306 VSS.n2811 VSS.n2810 1.6821
R9307 VSS.n293 VSS.n292 1.6819
R9308 VSS.n5407 VSS.n5406 1.6819
R9309 VSS.n2069 VSS.n2068 1.6819
R9310 VSS.n2662 VSS.n2661 1.6819
R9311 VSS.n3041 VSS.n3040 1.6819
R9312 VSS.n967 VSS.n966 1.6819
R9313 VSS.n1282 VSS.n1281 1.6819
R9314 VSS.n1350 VSS.n1349 1.6753
R9315 VSS.n3867 VSS.n3861 1.66667
R9316 VSS.n3186 VSS.n2983 1.65976
R9317 VSS.n1306 VSS.n1305 1.64728
R9318 VSS.n833 VSS.n832 1.63454
R9319 VSS.n4828 VSS.n1767 1.61027
R9320 VSS.n4121 VSS.n4120 1.54533
R9321 VSS.n898 VSS.n897 1.50638
R9322 VSS.n822 VSS.n821 1.50638
R9323 VSS.n821 VSS.n399 1.50638
R9324 VSS.n799 VSS.n798 1.50638
R9325 VSS.n742 VSS.n457 1.50638
R9326 VSS.n2078 VSS.n2077 1.50638
R9327 VSS.n2242 VSS.n2241 1.50638
R9328 VSS.n2481 VSS.n1987 1.50638
R9329 VSS.n2486 VSS.n2484 1.50638
R9330 VSS.n2524 VSS.n1975 1.50638
R9331 VSS.n2563 VSS.n1960 1.50638
R9332 VSS.n2588 VSS.n1950 1.50638
R9333 VSS.n2702 VSS.n2701 1.50638
R9334 VSS.n2830 VSS.n2801 1.50638
R9335 VSS.n3518 VSS.n3517 1.50638
R9336 VSS.n1218 VSS.n1199 1.50638
R9337 VSS.n1544 VSS.n1505 1.50638
R9338 VSS.n1649 VSS.n1017 1.50638
R9339 VSS.n1671 VSS.n1006 1.50638
R9340 VSS.n1228 VSS.n1196 1.49837
R9341 VSS.n940 VSS.n318 1.43682
R9342 VSS.n3889 VSS.n3886 1.43383
R9343 VSS.n2492 VSS.n2489 1.42272
R9344 VSS.n4204 VSS.n3903 1.41445
R9345 VSS.n4160 VSS.n4159 1.40119
R9346 VSS.n5469 VSS.n5468 1.3622
R9347 VSS.n3311 VSS.n3310 1.3622
R9348 VSS.n5452 VSS.n23 1.33898
R9349 VSS.n4289 VSS.n4288 1.32802
R9350 VSS.n4890 VSS.n1726 1.32464
R9351 VSS.n2812 VSS.n2811 1.30732
R9352 VSS.n296 VSS.n293 1.30718
R9353 VSS.n5410 VSS.n5407 1.30718
R9354 VSS.n2072 VSS.n2069 1.30718
R9355 VSS.n2663 VSS.n2662 1.30718
R9356 VSS.n3044 VSS.n3041 1.30718
R9357 VSS.n970 VSS.n967 1.30718
R9358 VSS.n1285 VSS.n1282 1.30718
R9359 VSS.n4828 VSS.n4827 1.28471
R9360 VSS.n4829 VSS.n4828 1.27382
R9361 VSS.n3327 VSS.n3325 1.24408
R9362 VSS.n4033 VSS.t3475 1.23959
R9363 VSS.n4961 VSS.n273 1.23559
R9364 VSS.n599 VSS.n598 1.23559
R9365 VSS.n2383 VSS.n2381 1.23559
R9366 VSS.n391 VSS.n388 1.22603
R9367 VSS.n2425 VSS.n2418 1.19136
R9368 VSS.n4814 VSS.n4811 1.18711
R9369 VSS.n4813 VSS.n4812 1.18711
R9370 VSS.n4806 VSS.n4803 1.18711
R9371 VSS.n4808 VSS.n4807 1.18711
R9372 VSS.n3848 VSS.n3842 1.18711
R9373 VSS.n3847 VSS.n3846 1.18711
R9374 VSS.n3854 VSS.n3826 1.18711
R9375 VSS.n3853 VSS.n3852 1.18711
R9376 VSS.n44 VSS.n43 1.18311
R9377 VSS.n5333 VSS.n5332 1.18311
R9378 VSS.n5246 VSS.n5245 1.18311
R9379 VSS.n5120 VSS.n196 1.18311
R9380 VSS.n5078 VSS.n5077 1.18311
R9381 VSS.n4924 VSS.n4923 1.18311
R9382 VSS.n633 VSS.n632 1.18311
R9383 VSS.n2323 VSS.n2322 1.18311
R9384 VSS.n3303 VSS.n3302 1.18311
R9385 VSS.n1837 VSS.n1836 1.18311
R9386 VSS.n3796 VSS.n3795 1.18311
R9387 VSS.n4688 VSS.n4687 1.18311
R9388 VSS.n5194 VSS.n5193 1.14023
R9389 VSS.n5156 VSS.n5155 1.14023
R9390 VSS.n4987 VSS.n4986 1.14023
R9391 VSS.n934 VSS.n322 1.14023
R9392 VSS.n5428 VSS.n5390 1.14023
R9393 VSS.n3420 VSS.n3419 1.14023
R9394 VSS.n3322 VSS.n3321 1.14023
R9395 VSS.n1297 VSS.n1269 1.14023
R9396 VSS.n1851 VSS.n1850 1.14023
R9397 VSS.n870 VSS.n869 1.12991
R9398 VSS.n2304 VSS.n2303 1.12991
R9399 VSS.n2449 VSS.n2448 1.12991
R9400 VSS.n1095 VSS.n1094 1.12991
R9401 VSS.n306 VSS.n305 1.11354
R9402 VSS.n3447 VSS.n3446 1.11354
R9403 VSS.n980 VSS.n979 1.11354
R9404 VSS.n4160 VSS.n3939 1.10883
R9405 VSS.n3087 VSS.n3086 1.06491
R9406 VSS.n3897 VSS.n3896 1.04229
R9407 VSS.n3979 VSS.n3978 1.01637
R9408 VSS.n3869 VSS.n3819 1.01637
R9409 VSS.n1302 VSS.n1301 1.00931
R9410 VSS.n3985 VSS.n1771 0.987643
R9411 VSS.n3984 VSS.n3940 0.987643
R9412 VSS.n4154 VSS.n3940 0.984154
R9413 VSS.n3986 VSS.n3985 0.973714
R9414 VSS.n201 VSS.n200 0.952566
R9415 VSS.n491 VSS.n490 0.952566
R9416 VSS.n989 VSS.n987 0.952566
R9417 VSS.n407 VSS.n404 0.948648
R9418 VSS.n4812 VSS.n4811 0.944548
R9419 VSS.n4814 VSS.n4813 0.944548
R9420 VSS.n4807 VSS.n4806 0.944548
R9421 VSS.n4808 VSS.n4803 0.944548
R9422 VSS.n3846 VSS.n3842 0.944548
R9423 VSS.n3848 VSS.n3847 0.944548
R9424 VSS.n3852 VSS.n3826 0.944548
R9425 VSS.n3854 VSS.n3853 0.944548
R9426 VSS.n688 VSS.n486 0.931411
R9427 VSS.n4889 VSS.n1728 0.883259
R9428 VSS.n4125 VSS.n4124 0.883259
R9429 VSS.n4118 VSS.n4117 0.848387
R9430 VSS.n1765 VSS.n1761 0.848386
R9431 VSS.n5189 VSS.n168 0.833377
R9432 VSS.n5151 VSS.n183 0.833377
R9433 VSS.n4982 VSS.n268 0.833377
R9434 VSS.n935 VSS.n321 0.833377
R9435 VSS.n5431 VSS.n5430 0.833377
R9436 VSS.n3415 VSS.n2911 0.833377
R9437 VSS.n3317 VSS.n2960 0.833377
R9438 VSS.n1300 VSS.n1299 0.833377
R9439 VSS.n3554 VSS.n1879 0.775551
R9440 VSS.n838 VSS.n383 0.753441
R9441 VSS.n424 VSS.n420 0.753441
R9442 VSS.n2077 VSS.n2076 0.753441
R9443 VSS.n2237 VSS.n2236 0.753441
R9444 VSS.n2260 VSS.n2259 0.753441
R9445 VSS.n2369 VSS.n2004 0.753441
R9446 VSS.n2475 VSS.n1991 0.753441
R9447 VSS.n2577 VSS.n2576 0.753441
R9448 VSS.n2578 VSS.n2577 0.753441
R9449 VSS.n2624 VSS.n2595 0.753441
R9450 VSS.n2673 VSS.n2672 0.753441
R9451 VSS.n3049 VSS.n3048 0.753441
R9452 VSS.n2824 VSS.n2823 0.753441
R9453 VSS.n3513 VSS.n3512 0.753441
R9454 VSS.n3500 VSS.n3499 0.753441
R9455 VSS.n3505 VSS.n3504 0.753441
R9456 VSS.n3491 VSS.n2774 0.753441
R9457 VSS.n3463 VSS.n3462 0.753441
R9458 VSS.n3464 VSS.n3463 0.753441
R9459 VSS.n3393 VSS.n3392 0.753441
R9460 VSS.n3387 VSS.n3386 0.753441
R9461 VSS.n3118 VSS.n3117 0.753441
R9462 VSS.n3123 VSS.n3002 0.753441
R9463 VSS.n3144 VSS.n2994 0.753441
R9464 VSS.n3195 VSS.n3194 0.753441
R9465 VSS.n1154 VSS.n1150 0.753441
R9466 VSS.n1435 VSS.n1434 0.753441
R9467 VSS.n1402 VSS.n1398 0.753441
R9468 VSS.n1566 VSS.n1565 0.753441
R9469 VSS.n1545 VSS.n1544 0.753441
R9470 VSS.n1534 VSS.n1512 0.753441
R9471 VSS.n1589 VSS.n1588 0.753441
R9472 VSS.n1657 VSS.n1656 0.753441
R9473 VSS.n4156 VSS.n1768 0.752461
R9474 VSS.n4836 VSS.n4834 0.750074
R9475 VSS.n4140 VSS.n4139 0.736693
R9476 VSS.n1824 VSS.n1822 0.732469
R9477 VSS.n1898 VSS.n1894 0.732469
R9478 VSS.n4061 VSS.n4059 0.732469
R9479 VSS.n1794 VSS.n1793 0.732469
R9480 VSS.n4855 VSS.n4854 0.728182
R9481 VSS.n4013 VSS.n3942 0.728182
R9482 VSS.n346 VSS.n344 0.711611
R9483 VSS.n816 VSS.n401 0.711611
R9484 VSS.n2425 VSS.n2424 0.711611
R9485 VSS.n2493 VSS.n2492 0.711611
R9486 VSS.n2884 VSS.n2883 0.711611
R9487 VSS.n3526 VSS.n3525 0.711611
R9488 VSS.n3086 VSS.n3085 0.711611
R9489 VSS.n3187 VSS.n3186 0.711611
R9490 VSS.n1349 VSS.n1158 0.711611
R9491 VSS.n4851 VSS.n4833 0.6935
R9492 VSS.n4135 VSS.n4132 0.6935
R9493 VSS.n4261 VSS.t3392 0.677631
R9494 VSS.n4854 VSS.n4830 0.661267
R9495 VSS.n4152 VSS.n3942 0.661267
R9496 VSS.n4852 VSS.n4832 0.627947
R9497 VSS.n4134 VSS.n3944 0.627947
R9498 VSS.n4845 VSS.n4832 0.598603
R9499 VSS.n4151 VSS.n3944 0.598603
R9500 VSS.n4847 VSS.n4833 0.596535
R9501 VSS.n4132 VSS.n3945 0.596535
R9502 VSS.n3444 VSS.n3443 0.578357
R9503 VSS.n3884 VSS.n3883 0.563
R9504 VSS.n3885 VSS.n3884 0.563
R9505 VSS.n4850 VSS.n4849 0.561264
R9506 VSS.n4136 VSS.n4131 0.561264
R9507 VSS.n1858 VSS.n1857 0.548538
R9508 VSS.n4743 VSS.n4739 0.548535
R9509 VSS.n4781 VSS.n4780 0.548535
R9510 VSS.n4094 VSS.n4091 0.548489
R9511 VSS.n4846 VSS.n1740 0.547559
R9512 VSS.n4150 VSS.n4149 0.547559
R9513 VSS.n3902 VSS.n3901 0.543
R9514 VSS.n3267 VSS.n3234 0.537563
R9515 VSS.n4155 VSS.n3554 0.533812
R9516 VSS.n5190 VSS.n5188 0.526527
R9517 VSS.n5152 VSS.n5150 0.526527
R9518 VSS.n4983 VSS.n4981 0.526527
R9519 VSS.n5389 VSS.n5387 0.526527
R9520 VSS.n3416 VSS.n3414 0.526527
R9521 VSS.n3318 VSS.n3316 0.526527
R9522 VSS.n4130 VSS.n3945 0.52524
R9523 VSS.n4848 VSS.n4847 0.523938
R9524 VSS.n4845 VSS.n4830 0.510917
R9525 VSS.n4152 VSS.n4151 0.510917
R9526 VSS.n4849 VSS.n4848 0.496683
R9527 VSS.n4131 VSS.n4130 0.496683
R9528 VSS.n939 VSS.n938 0.482692
R9529 VSS.n3900 VSS.n3899 0.4805
R9530 VSS.n2314 VSS.n2313 0.474574
R9531 VSS.n2461 VSS.n2460 0.474574
R9532 VSS.n2552 VSS.n2551 0.474574
R9533 VSS.n3898 VSS.n3897 0.472292
R9534 VSS.n4157 VSS.n4156 0.452653
R9535 VSS.n4291 VSS.n4290 0.449932
R9536 VSS.n4970 VSS.n4969 0.449623
R9537 VSS.n606 VSS.n605 0.449623
R9538 VSS.n2376 VSS.n2375 0.449623
R9539 VSS.n3100 VSS.n3098 0.449623
R9540 VSS.n3242 VSS.n3241 0.448052
R9541 VSS.n4885 VSS.n4884 0.441879
R9542 VSS.n4128 VSS.n4127 0.441879
R9543 VSS.n1874 VSS.n1846 0.438856
R9544 VSS.n1866 VSS.n1865 0.438856
R9545 VSS.n4186 VSS.n4185 0.438107
R9546 VSS.n47 VSS.n46 0.417891
R9547 VSS.n5330 VSS.n5329 0.417891
R9548 VSS.n5334 VSS.n5333 0.417891
R9549 VSS.n5243 VSS.n5242 0.417891
R9550 VSS.n5247 VSS.n5246 0.417891
R9551 VSS.n5119 VSS.n5118 0.417891
R9552 VSS.n5124 VSS.n196 0.417891
R9553 VSS.n5076 VSS.n5075 0.417891
R9554 VSS.n5077 VSS.n218 0.417891
R9555 VSS.n4928 VSS.n4922 0.417891
R9556 VSS.n302 VSS.n301 0.417891
R9557 VSS.n304 VSS.n284 0.417891
R9558 VSS.n632 VSS.n631 0.417891
R9559 VSS.n2268 VSS.n2266 0.417891
R9560 VSS.n2322 VSS.n2321 0.417891
R9561 VSS.n3445 VSS.n3444 0.417891
R9562 VSS.n3446 VSS.n2897 0.417891
R9563 VSS.n3300 VSS.n3299 0.417891
R9564 VSS.n976 VSS.n975 0.417891
R9565 VSS.n978 VSS.n959 0.417891
R9566 VSS.n1832 VSS.n1818 0.417891
R9567 VSS.n1838 VSS.n1837 0.417891
R9568 VSS.n3799 VSS.n3798 0.417891
R9569 VSS.n4692 VSS.n4686 0.417891
R9570 VSS.n29 VSS.n27 0.409011
R9571 VSS.n78 VSS.n77 0.409011
R9572 VSS.n5182 VSS.n5181 0.409011
R9573 VSS.n5144 VSS.n5143 0.409011
R9574 VSS.n5111 VSS.n5110 0.409011
R9575 VSS.n4975 VSS.n4974 0.409011
R9576 VSS.n316 VSS.n313 0.409011
R9577 VSS.n834 VSS.n833 0.409011
R9578 VSS.n827 VSS.n393 0.409011
R9579 VSS.n688 VSS.n687 0.409011
R9580 VSS.n5471 VSS.n5470 0.409011
R9581 VSS.n5460 VSS.n20 0.409011
R9582 VSS.n5453 VSS.n5452 0.409011
R9583 VSS.n5385 VSS.n5383 0.409011
R9584 VSS.n2301 VSS.n2276 0.409011
R9585 VSS.n2294 VSS.n2293 0.409011
R9586 VSS.n3407 VSS.n3406 0.409011
R9587 VSS.n3309 VSS.n3308 0.409011
R9588 VSS.n1220 VSS.n1219 0.409011
R9589 VSS.n1231 VSS.n1230 0.409011
R9590 VSS.n1575 VSS.n1114 0.409011
R9591 VSS.n1840 VSS.n1839 0.409011
R9592 VSS.n4507 VSS.n4506 0.409011
R9593 VSS.n4513 VSS.n3610 0.409011
R9594 VSS.n4156 VSS.n4155 0.406443
R9595 VSS.n4290 VSS.n1768 0.393625
R9596 VSS.n3979 VSS.n3974 0.388
R9597 VSS.n3983 VSS.n3972 0.388
R9598 VSS.n3863 VSS.n3862 0.388
R9599 VSS.n3869 VSS.n3868 0.388
R9600 VSS.n613 VSS.n612 0.376971
R9601 VSS.n2247 VSS.n2021 0.376971
R9602 VSS.n2502 VSS.n1983 0.376971
R9603 VSS.n2527 VSS.n2526 0.376971
R9604 VSS.n3332 VSS.n2956 0.376971
R9605 VSS.n3286 VSS.n3285 0.376971
R9606 VSS.n1320 VSS.n1319 0.376971
R9607 VSS.n1827 VSS.n1821 0.376971
R9608 VSS.n1901 VSS.n1893 0.376971
R9609 VSS.n1914 VSS.n1885 0.376971
R9610 VSS.n4064 VSS.n4058 0.376971
R9611 VSS.n4079 VSS.n4078 0.376971
R9612 VSS.n1810 VSS.n1809 0.376971
R9613 VSS.n1797 VSS.n1796 0.376971
R9614 VSS.n4547 VSS.n4546 0.376971
R9615 VSS.n4479 VSS.n4478 0.376971
R9616 VSS.n4417 VSS.n4416 0.376971
R9617 VSS.n4585 VSS.n4583 0.376971
R9618 VSS.n4223 VSS.n3880 0.376971
R9619 VSS.n4853 VSS.n4831 0.371802
R9620 VSS.n4133 VSS.n3943 0.371802
R9621 VSS.n1707 VSS.n1706 0.35916
R9622 VSS.n4852 VSS.n4851 0.343032
R9623 VSS.n4135 VSS.n4134 0.343032
R9624 VSS.n17 VSS.n16 0.340926
R9625 VSS.n1582 VSS.n1580 0.340926
R9626 VSS.n4293 VSS.n4292 0.338974
R9627 VSS.n4846 VSS.n4845 0.337621
R9628 VSS.n4151 VSS.n4150 0.337621
R9629 VSS.n4831 VSS.n4830 0.333523
R9630 VSS.n4152 VSS.n3943 0.333523
R9631 VSS.n3902 VSS.n3900 0.333
R9632 VSS.n4288 VSS.n3902 0.330857
R9633 VSS.n4847 VSS.n4846 0.328202
R9634 VSS.n4150 VSS.n3945 0.328202
R9635 VSS.n4136 VSS.n4135 0.32761
R9636 VSS.n4851 VSS.n4850 0.326799
R9637 VSS.n4871 VSS.n1740 0.3205
R9638 VSS.n4149 VSS.n3946 0.3205
R9639 VSS.n4853 VSS.n4852 0.318682
R9640 VSS.n4134 VSS.n4133 0.318682
R9641 VSS.n4006 VSS.n4003 0.311532
R9642 VSS.n3861 VSS.n3860 0.307193
R9643 VSS.n4766 VSS.n1879 0.301853
R9644 VSS.n4766 VSS.n4765 0.301853
R9645 VSS.n4158 VSS.n3932 0.3005
R9646 VSS.n3894 VSS.n3893 0.297375
R9647 VSS.n4827 VSS.n4826 0.290794
R9648 VSS.n4827 VSS.n1768 0.288701
R9649 VSS.n4904 VSS.n4903 0.283731
R9650 VSS.n523 VSS.n521 0.278761
R9651 VSS.n4161 VSS.n4160 0.267759
R9652 VSS.n5197 VSS.n166 0.263514
R9653 VSS.n184 VSS.n181 0.263514
R9654 VSS.n4990 VSS.n266 0.263514
R9655 VSS.n931 VSS.n324 0.263514
R9656 VSS.n5427 VSS.n5426 0.263514
R9657 VSS.n3423 VSS.n2909 0.263514
R9658 VSS.n3325 VSS.n2958 0.263514
R9659 VSS.n1296 VSS.n1295 0.263514
R9660 VSS.n1861 VSS.n1853 0.263514
R9661 VSS.n4815 VSS.n4810 0.248897
R9662 VSS.n3849 VSS.n3841 0.248897
R9663 VSS.n4848 VSS.n1729 0.242688
R9664 VSS.n4130 VSS.n4129 0.241385
R9665 VSS.n683 VSS.n489 0.239726
R9666 VSS.n5115 VSS.n5114 0.239726
R9667 VSS.n1315 VSS.n1261 0.239726
R9668 VSS.n5115 VSS.n198 0.239381
R9669 VSS.n684 VSS.n683 0.239381
R9670 VSS.n1708 VSS.n1707 0.239381
R9671 VSS.n1706 VSS.n1705 0.239381
R9672 VSS.n1310 VSS.n1261 0.239381
R9673 VSS.n3526 VSS.n3521 0.237537
R9674 VSS.n1311 VSS.n1263 0.225061
R9675 VSS.n1302 VSS.n1265 0.225061
R9676 VSS.n4287 VSS.n4286 0.216779
R9677 VSS.n3304 VSS.n3303 0.209196
R9678 VSS.n3305 VSS.n3304 0.209196
R9679 VSS.n4292 VSS.n4291 0.190841
R9680 VSS.n4809 VSS.n4802 0.179898
R9681 VSS.n3851 VSS.n3825 0.179898
R9682 VSS.n4642 VSS.n3554 0.171912
R9683 VSS.n3714 VSS.n3712 0.171884
R9684 VSS.n4289 VSS.n3895 0.164562
R9685 VSS.n4155 VSS.n4154 0.162788
R9686 VSS.n4823 VSS.n1770 0.15675
R9687 VSS.n3859 VSS.n3821 0.15675
R9688 VSS.n4824 VSS.n1771 0.153427
R9689 VSS.n5489 VSS.n1 0.1509
R9690 VSS.n2742 VSS.n1 0.1509
R9691 VSS.n3553 VSS.n2742 0.1509
R9692 VSS.n4642 VSS.n3553 0.1509
R9693 VSS.n2321 VSS.n2320 0.149858
R9694 VSS.n4162 VSS.n4161 0.145413
R9695 VSS.n4850 VSS.n4844 0.141388
R9696 VSS.n4138 VSS.n4136 0.140576
R9697 VSS.n301 VSS.n300 0.13963
R9698 VSS.n637 VSS.n521 0.13963
R9699 VSS.n975 VSS.n974 0.13963
R9700 VSS.n945 VSS.n944 0.13667
R9701 VSS.n685 VSS.n488 0.13667
R9702 VSS.n4290 VSS.n4289 0.122091
R9703 VSS.n4888 VSS.n1727 0.120292
R9704 VSS.n4888 VSS.n4887 0.120292
R9705 VSS.n4887 VSS.n1729 0.120292
R9706 VSS.n4927 VSS.n4926 0.120292
R9707 VSS.n4927 VSS.n4921 0.120292
R9708 VSS.n4921 VSS.n4919 0.120292
R9709 VSS.n4932 VSS.n4919 0.120292
R9710 VSS.n4933 VSS.n4932 0.120292
R9711 VSS.n4934 VSS.n4933 0.120292
R9712 VSS.n4934 VSS.n4916 0.120292
R9713 VSS.n4938 VSS.n4916 0.120292
R9714 VSS.n4939 VSS.n4938 0.120292
R9715 VSS.n4940 VSS.n4939 0.120292
R9716 VSS.n4940 VSS.n282 0.120292
R9717 VSS.n4944 VSS.n282 0.120292
R9718 VSS.n4945 VSS.n4944 0.120292
R9719 VSS.n4946 VSS.n4945 0.120292
R9720 VSS.n4946 VSS.n280 0.120292
R9721 VSS.n4950 VSS.n280 0.120292
R9722 VSS.n4951 VSS.n4950 0.120292
R9723 VSS.n4952 VSS.n4951 0.120292
R9724 VSS.n4952 VSS.n277 0.120292
R9725 VSS.n4956 VSS.n277 0.120292
R9726 VSS.n4957 VSS.n4956 0.120292
R9727 VSS.n4957 VSS.n274 0.120292
R9728 VSS.n4963 VSS.n274 0.120292
R9729 VSS.n4964 VSS.n4963 0.120292
R9730 VSS.n4965 VSS.n4964 0.120292
R9731 VSS.n4965 VSS.n272 0.120292
R9732 VSS.n4971 VSS.n272 0.120292
R9733 VSS.n4972 VSS.n4971 0.120292
R9734 VSS.n4973 VSS.n4972 0.120292
R9735 VSS.n4973 VSS.n270 0.120292
R9736 VSS.n4978 VSS.n270 0.120292
R9737 VSS.n4979 VSS.n4978 0.120292
R9738 VSS.n4980 VSS.n4979 0.120292
R9739 VSS.n4980 VSS.n267 0.120292
R9740 VSS.n4988 VSS.n267 0.120292
R9741 VSS.n4989 VSS.n4988 0.120292
R9742 VSS.n4989 VSS.n264 0.120292
R9743 VSS.n264 VSS.n262 0.120292
R9744 VSS.n4994 VSS.n262 0.120292
R9745 VSS.n4995 VSS.n4994 0.120292
R9746 VSS.n4996 VSS.n4995 0.120292
R9747 VSS.n4996 VSS.n259 0.120292
R9748 VSS.n259 VSS.n258 0.120292
R9749 VSS.n5001 VSS.n258 0.120292
R9750 VSS.n5002 VSS.n5001 0.120292
R9751 VSS.n5003 VSS.n5002 0.120292
R9752 VSS.n5003 VSS.n256 0.120292
R9753 VSS.n5007 VSS.n256 0.120292
R9754 VSS.n5008 VSS.n5007 0.120292
R9755 VSS.n5009 VSS.n5008 0.120292
R9756 VSS.n5009 VSS.n253 0.120292
R9757 VSS.n253 VSS.n252 0.120292
R9758 VSS.n5014 VSS.n252 0.120292
R9759 VSS.n5015 VSS.n5014 0.120292
R9760 VSS.n5016 VSS.n5015 0.120292
R9761 VSS.n5016 VSS.n248 0.120292
R9762 VSS.n5020 VSS.n248 0.120292
R9763 VSS.n5021 VSS.n5020 0.120292
R9764 VSS.n5022 VSS.n5021 0.120292
R9765 VSS.n5022 VSS.n245 0.120292
R9766 VSS.n5026 VSS.n245 0.120292
R9767 VSS.n5027 VSS.n5026 0.120292
R9768 VSS.n5028 VSS.n5027 0.120292
R9769 VSS.n5028 VSS.n242 0.120292
R9770 VSS.n242 VSS.n240 0.120292
R9771 VSS.n240 VSS.n239 0.120292
R9772 VSS.n5034 VSS.n239 0.120292
R9773 VSS.n5035 VSS.n5034 0.120292
R9774 VSS.n5036 VSS.n5035 0.120292
R9775 VSS.n5036 VSS.n237 0.120292
R9776 VSS.n5040 VSS.n237 0.120292
R9777 VSS.n5041 VSS.n5040 0.120292
R9778 VSS.n5041 VSS.n234 0.120292
R9779 VSS.n5045 VSS.n234 0.120292
R9780 VSS.n5046 VSS.n5045 0.120292
R9781 VSS.n5047 VSS.n5046 0.120292
R9782 VSS.n5047 VSS.n231 0.120292
R9783 VSS.n5052 VSS.n231 0.120292
R9784 VSS.n5053 VSS.n5052 0.120292
R9785 VSS.n5054 VSS.n5053 0.120292
R9786 VSS.n5054 VSS.n229 0.120292
R9787 VSS.n5058 VSS.n229 0.120292
R9788 VSS.n5059 VSS.n5058 0.120292
R9789 VSS.n5060 VSS.n5059 0.120292
R9790 VSS.n5060 VSS.n226 0.120292
R9791 VSS.n5064 VSS.n226 0.120292
R9792 VSS.n5065 VSS.n5064 0.120292
R9793 VSS.n5066 VSS.n5065 0.120292
R9794 VSS.n5066 VSS.n224 0.120292
R9795 VSS.n5070 VSS.n224 0.120292
R9796 VSS.n5071 VSS.n5070 0.120292
R9797 VSS.n5072 VSS.n5071 0.120292
R9798 VSS.n5072 VSS.n220 0.120292
R9799 VSS.n220 VSS.n219 0.120292
R9800 VSS.n5080 VSS.n219 0.120292
R9801 VSS.n5081 VSS.n5080 0.120292
R9802 VSS.n5082 VSS.n5081 0.120292
R9803 VSS.n5082 VSS.n216 0.120292
R9804 VSS.n216 VSS.n215 0.120292
R9805 VSS.n5087 VSS.n215 0.120292
R9806 VSS.n5088 VSS.n5087 0.120292
R9807 VSS.n5088 VSS.n212 0.120292
R9808 VSS.n5093 VSS.n212 0.120292
R9809 VSS.n5094 VSS.n5093 0.120292
R9810 VSS.n5095 VSS.n5094 0.120292
R9811 VSS.n5095 VSS.n208 0.120292
R9812 VSS.n5099 VSS.n208 0.120292
R9813 VSS.n5100 VSS.n5099 0.120292
R9814 VSS.n5101 VSS.n5100 0.120292
R9815 VSS.n5101 VSS.n206 0.120292
R9816 VSS.n206 VSS.n205 0.120292
R9817 VSS.n205 VSS.n204 0.120292
R9818 VSS.n5107 VSS.n204 0.120292
R9819 VSS.n5108 VSS.n5107 0.120292
R9820 VSS.n5109 VSS.n5108 0.120292
R9821 VSS.n5109 VSS.n202 0.120292
R9822 VSS.n5114 VSS.n202 0.120292
R9823 VSS.n198 VSS.n197 0.120292
R9824 VSS.n5122 VSS.n197 0.120292
R9825 VSS.n5123 VSS.n5122 0.120292
R9826 VSS.n5123 VSS.n195 0.120292
R9827 VSS.n5127 VSS.n195 0.120292
R9828 VSS.n5128 VSS.n5127 0.120292
R9829 VSS.n5129 VSS.n5128 0.120292
R9830 VSS.n5129 VSS.n191 0.120292
R9831 VSS.n5133 VSS.n191 0.120292
R9832 VSS.n5134 VSS.n5133 0.120292
R9833 VSS.n5135 VSS.n5134 0.120292
R9834 VSS.n5135 VSS.n188 0.120292
R9835 VSS.n5140 VSS.n188 0.120292
R9836 VSS.n5141 VSS.n5140 0.120292
R9837 VSS.n5142 VSS.n5141 0.120292
R9838 VSS.n5142 VSS.n186 0.120292
R9839 VSS.n5147 VSS.n186 0.120292
R9840 VSS.n5148 VSS.n5147 0.120292
R9841 VSS.n5149 VSS.n5148 0.120292
R9842 VSS.n5149 VSS.n182 0.120292
R9843 VSS.n5157 VSS.n182 0.120292
R9844 VSS.n5158 VSS.n5157 0.120292
R9845 VSS.n5159 VSS.n5158 0.120292
R9846 VSS.n5159 VSS.n180 0.120292
R9847 VSS.n5165 VSS.n180 0.120292
R9848 VSS.n5166 VSS.n5165 0.120292
R9849 VSS.n5167 VSS.n5166 0.120292
R9850 VSS.n5167 VSS.n177 0.120292
R9851 VSS.n5171 VSS.n177 0.120292
R9852 VSS.n5172 VSS.n5171 0.120292
R9853 VSS.n5173 VSS.n5172 0.120292
R9854 VSS.n5173 VSS.n174 0.120292
R9855 VSS.n174 VSS.n172 0.120292
R9856 VSS.n5178 VSS.n172 0.120292
R9857 VSS.n5179 VSS.n5178 0.120292
R9858 VSS.n5180 VSS.n5179 0.120292
R9859 VSS.n5180 VSS.n170 0.120292
R9860 VSS.n5185 VSS.n170 0.120292
R9861 VSS.n5186 VSS.n5185 0.120292
R9862 VSS.n5187 VSS.n5186 0.120292
R9863 VSS.n5187 VSS.n167 0.120292
R9864 VSS.n5195 VSS.n167 0.120292
R9865 VSS.n5196 VSS.n5195 0.120292
R9866 VSS.n5196 VSS.n165 0.120292
R9867 VSS.n5202 VSS.n165 0.120292
R9868 VSS.n5203 VSS.n5202 0.120292
R9869 VSS.n5204 VSS.n5203 0.120292
R9870 VSS.n5204 VSS.n163 0.120292
R9871 VSS.n5208 VSS.n163 0.120292
R9872 VSS.n5209 VSS.n5208 0.120292
R9873 VSS.n5210 VSS.n5209 0.120292
R9874 VSS.n5210 VSS.n160 0.120292
R9875 VSS.n5214 VSS.n160 0.120292
R9876 VSS.n5215 VSS.n5214 0.120292
R9877 VSS.n5216 VSS.n5215 0.120292
R9878 VSS.n5216 VSS.n156 0.120292
R9879 VSS.n5220 VSS.n156 0.120292
R9880 VSS.n5221 VSS.n5220 0.120292
R9881 VSS.n5222 VSS.n5221 0.120292
R9882 VSS.n5222 VSS.n154 0.120292
R9883 VSS.n154 VSS.n153 0.120292
R9884 VSS.n5227 VSS.n153 0.120292
R9885 VSS.n5228 VSS.n5227 0.120292
R9886 VSS.n5229 VSS.n5228 0.120292
R9887 VSS.n5229 VSS.n151 0.120292
R9888 VSS.n5233 VSS.n151 0.120292
R9889 VSS.n5234 VSS.n5233 0.120292
R9890 VSS.n5235 VSS.n5234 0.120292
R9891 VSS.n5235 VSS.n147 0.120292
R9892 VSS.n5239 VSS.n147 0.120292
R9893 VSS.n5240 VSS.n5239 0.120292
R9894 VSS.n5241 VSS.n5240 0.120292
R9895 VSS.n5241 VSS.n145 0.120292
R9896 VSS.n5248 VSS.n145 0.120292
R9897 VSS.n5249 VSS.n5248 0.120292
R9898 VSS.n5251 VSS.n5249 0.120292
R9899 VSS.n5251 VSS.n5250 0.120292
R9900 VSS.n5250 VSS.n142 0.120292
R9901 VSS.n5259 VSS.n142 0.120292
R9902 VSS.n5260 VSS.n5259 0.120292
R9903 VSS.n5261 VSS.n5260 0.120292
R9904 VSS.n5261 VSS.n139 0.120292
R9905 VSS.n139 VSS.n137 0.120292
R9906 VSS.n5266 VSS.n137 0.120292
R9907 VSS.n5267 VSS.n5266 0.120292
R9908 VSS.n5268 VSS.n5267 0.120292
R9909 VSS.n5268 VSS.n134 0.120292
R9910 VSS.n5272 VSS.n134 0.120292
R9911 VSS.n5273 VSS.n5272 0.120292
R9912 VSS.n5274 VSS.n5273 0.120292
R9913 VSS.n5274 VSS.n131 0.120292
R9914 VSS.n131 VSS.n130 0.120292
R9915 VSS.n5279 VSS.n130 0.120292
R9916 VSS.n5280 VSS.n5279 0.120292
R9917 VSS.n5282 VSS.n5280 0.120292
R9918 VSS.n5282 VSS.n5281 0.120292
R9919 VSS.n5281 VSS.n127 0.120292
R9920 VSS.n5290 VSS.n127 0.120292
R9921 VSS.n5291 VSS.n5290 0.120292
R9922 VSS.n5292 VSS.n5291 0.120292
R9923 VSS.n5292 VSS.n124 0.120292
R9924 VSS.n5296 VSS.n124 0.120292
R9925 VSS.n5297 VSS.n5296 0.120292
R9926 VSS.n5299 VSS.n5297 0.120292
R9927 VSS.n5299 VSS.n5298 0.120292
R9928 VSS.n5298 VSS.n121 0.120292
R9929 VSS.n5307 VSS.n121 0.120292
R9930 VSS.n5308 VSS.n5307 0.120292
R9931 VSS.n5309 VSS.n5308 0.120292
R9932 VSS.n5309 VSS.n118 0.120292
R9933 VSS.n118 VSS.n116 0.120292
R9934 VSS.n5314 VSS.n116 0.120292
R9935 VSS.n5315 VSS.n5314 0.120292
R9936 VSS.n5316 VSS.n5315 0.120292
R9937 VSS.n5316 VSS.n113 0.120292
R9938 VSS.n5320 VSS.n113 0.120292
R9939 VSS.n5321 VSS.n5320 0.120292
R9940 VSS.n5322 VSS.n5321 0.120292
R9941 VSS.n5322 VSS.n110 0.120292
R9942 VSS.n5326 VSS.n110 0.120292
R9943 VSS.n5327 VSS.n5326 0.120292
R9944 VSS.n5328 VSS.n5327 0.120292
R9945 VSS.n5328 VSS.n108 0.120292
R9946 VSS.n5335 VSS.n108 0.120292
R9947 VSS.n5354 VSS.n97 0.120292
R9948 VSS.n5355 VSS.n5354 0.120292
R9949 VSS.n5356 VSS.n5355 0.120292
R9950 VSS.n5356 VSS.n95 0.120292
R9951 VSS.n5364 VSS.n95 0.120292
R9952 VSS.n5365 VSS.n5364 0.120292
R9953 VSS.n5366 VSS.n5365 0.120292
R9954 VSS.n5366 VSS.n93 0.120292
R9955 VSS.n5370 VSS.n93 0.120292
R9956 VSS.n5371 VSS.n5370 0.120292
R9957 VSS.n5372 VSS.n5371 0.120292
R9958 VSS.n5372 VSS.n90 0.120292
R9959 VSS.n90 VSS.n89 0.120292
R9960 VSS.n89 VSS.n88 0.120292
R9961 VSS.n88 VSS.n26 0.120292
R9962 VSS.n84 VSS.n26 0.120292
R9963 VSS.n84 VSS.n83 0.120292
R9964 VSS.n83 VSS.n82 0.120292
R9965 VSS.n82 VSS.n28 0.120292
R9966 VSS.n76 VSS.n28 0.120292
R9967 VSS.n76 VSS.n75 0.120292
R9968 VSS.n75 VSS.n74 0.120292
R9969 VSS.n74 VSS.n31 0.120292
R9970 VSS.n69 VSS.n31 0.120292
R9971 VSS.n69 VSS.n68 0.120292
R9972 VSS.n68 VSS.n67 0.120292
R9973 VSS.n67 VSS.n34 0.120292
R9974 VSS.n63 VSS.n34 0.120292
R9975 VSS.n63 VSS.n62 0.120292
R9976 VSS.n62 VSS.n61 0.120292
R9977 VSS.n61 VSS.n37 0.120292
R9978 VSS.n57 VSS.n37 0.120292
R9979 VSS.n57 VSS.n56 0.120292
R9980 VSS.n56 VSS.n55 0.120292
R9981 VSS.n55 VSS.n40 0.120292
R9982 VSS.n50 VSS.n40 0.120292
R9983 VSS.n50 VSS.n49 0.120292
R9984 VSS.n49 VSS.n48 0.120292
R9985 VSS.n48 VSS.n42 0.120292
R9986 VSS.n297 VSS.n296 0.120292
R9987 VSS.n298 VSS.n297 0.120292
R9988 VSS.n298 VSS.n286 0.120292
R9989 VSS.n308 VSS.n286 0.120292
R9990 VSS.n309 VSS.n308 0.120292
R9991 VSS.n955 VSS.n309 0.120292
R9992 VSS.n955 VSS.n954 0.120292
R9993 VSS.n954 VSS.n953 0.120292
R9994 VSS.n953 VSS.n310 0.120292
R9995 VSS.n949 VSS.n310 0.120292
R9996 VSS.n949 VSS.n948 0.120292
R9997 VSS.n948 VSS.n947 0.120292
R9998 VSS.n947 VSS.n314 0.120292
R9999 VSS.n942 VSS.n314 0.120292
R10000 VSS.n942 VSS.n941 0.120292
R10001 VSS.n941 VSS.n319 0.120292
R10002 VSS.n933 VSS.n319 0.120292
R10003 VSS.n933 VSS.n932 0.120292
R10004 VSS.n932 VSS.n323 0.120292
R10005 VSS.n927 VSS.n323 0.120292
R10006 VSS.n927 VSS.n926 0.120292
R10007 VSS.n926 VSS.n327 0.120292
R10008 VSS.n919 VSS.n327 0.120292
R10009 VSS.n919 VSS.n918 0.120292
R10010 VSS.n918 VSS.n330 0.120292
R10011 VSS.n331 VSS.n330 0.120292
R10012 VSS.n913 VSS.n331 0.120292
R10013 VSS.n913 VSS.n912 0.120292
R10014 VSS.n912 VSS.n911 0.120292
R10015 VSS.n911 VSS.n334 0.120292
R10016 VSS.n907 VSS.n334 0.120292
R10017 VSS.n907 VSS.n906 0.120292
R10018 VSS.n906 VSS.n905 0.120292
R10019 VSS.n905 VSS.n337 0.120292
R10020 VSS.n901 VSS.n337 0.120292
R10021 VSS.n901 VSS.n900 0.120292
R10022 VSS.n900 VSS.n899 0.120292
R10023 VSS.n899 VSS.n342 0.120292
R10024 VSS.n893 VSS.n342 0.120292
R10025 VSS.n893 VSS.n892 0.120292
R10026 VSS.n892 VSS.n891 0.120292
R10027 VSS.n891 VSS.n345 0.120292
R10028 VSS.n887 VSS.n345 0.120292
R10029 VSS.n887 VSS.n886 0.120292
R10030 VSS.n886 VSS.n885 0.120292
R10031 VSS.n885 VSS.n351 0.120292
R10032 VSS.n881 VSS.n351 0.120292
R10033 VSS.n881 VSS.n880 0.120292
R10034 VSS.n880 VSS.n879 0.120292
R10035 VSS.n879 VSS.n355 0.120292
R10036 VSS.n875 VSS.n355 0.120292
R10037 VSS.n875 VSS.n874 0.120292
R10038 VSS.n874 VSS.n358 0.120292
R10039 VSS.n868 VSS.n358 0.120292
R10040 VSS.n868 VSS.n867 0.120292
R10041 VSS.n867 VSS.n866 0.120292
R10042 VSS.n866 VSS.n361 0.120292
R10043 VSS.n860 VSS.n361 0.120292
R10044 VSS.n860 VSS.n859 0.120292
R10045 VSS.n859 VSS.n858 0.120292
R10046 VSS.n858 VSS.n366 0.120292
R10047 VSS.n367 VSS.n366 0.120292
R10048 VSS.n369 VSS.n367 0.120292
R10049 VSS.n370 VSS.n369 0.120292
R10050 VSS.n371 VSS.n370 0.120292
R10051 VSS.n850 VSS.n371 0.120292
R10052 VSS.n850 VSS.n849 0.120292
R10053 VSS.n849 VSS.n848 0.120292
R10054 VSS.n848 VSS.n375 0.120292
R10055 VSS.n844 VSS.n375 0.120292
R10056 VSS.n844 VSS.n843 0.120292
R10057 VSS.n843 VSS.n842 0.120292
R10058 VSS.n842 VSS.n380 0.120292
R10059 VSS.n837 VSS.n380 0.120292
R10060 VSS.n837 VSS.n836 0.120292
R10061 VSS.n836 VSS.n384 0.120292
R10062 VSS.n830 VSS.n384 0.120292
R10063 VSS.n830 VSS.n829 0.120292
R10064 VSS.n829 VSS.n828 0.120292
R10065 VSS.n828 VSS.n389 0.120292
R10066 VSS.n396 VSS.n389 0.120292
R10067 VSS.n397 VSS.n396 0.120292
R10068 VSS.n398 VSS.n397 0.120292
R10069 VSS.n820 VSS.n398 0.120292
R10070 VSS.n820 VSS.n819 0.120292
R10071 VSS.n819 VSS.n400 0.120292
R10072 VSS.n815 VSS.n400 0.120292
R10073 VSS.n815 VSS.n814 0.120292
R10074 VSS.n814 VSS.n402 0.120292
R10075 VSS.n409 VSS.n402 0.120292
R10076 VSS.n809 VSS.n409 0.120292
R10077 VSS.n809 VSS.n808 0.120292
R10078 VSS.n808 VSS.n807 0.120292
R10079 VSS.n807 VSS.n411 0.120292
R10080 VSS.n803 VSS.n411 0.120292
R10081 VSS.n803 VSS.n802 0.120292
R10082 VSS.n802 VSS.n801 0.120292
R10083 VSS.n801 VSS.n417 0.120292
R10084 VSS.n419 VSS.n417 0.120292
R10085 VSS.n796 VSS.n419 0.120292
R10086 VSS.n796 VSS.n795 0.120292
R10087 VSS.n795 VSS.n794 0.120292
R10088 VSS.n794 VSS.n421 0.120292
R10089 VSS.n790 VSS.n421 0.120292
R10090 VSS.n790 VSS.n789 0.120292
R10091 VSS.n789 VSS.n788 0.120292
R10092 VSS.n788 VSS.n428 0.120292
R10093 VSS.n429 VSS.n428 0.120292
R10094 VSS.n783 VSS.n429 0.120292
R10095 VSS.n783 VSS.n782 0.120292
R10096 VSS.n782 VSS.n432 0.120292
R10097 VSS.n434 VSS.n432 0.120292
R10098 VSS.n776 VSS.n434 0.120292
R10099 VSS.n776 VSS.n775 0.120292
R10100 VSS.n775 VSS.n774 0.120292
R10101 VSS.n774 VSS.n436 0.120292
R10102 VSS.n770 VSS.n436 0.120292
R10103 VSS.n770 VSS.n769 0.120292
R10104 VSS.n769 VSS.n768 0.120292
R10105 VSS.n768 VSS.n440 0.120292
R10106 VSS.n441 VSS.n440 0.120292
R10107 VSS.n442 VSS.n441 0.120292
R10108 VSS.n444 VSS.n442 0.120292
R10109 VSS.n445 VSS.n444 0.120292
R10110 VSS.n760 VSS.n445 0.120292
R10111 VSS.n760 VSS.n759 0.120292
R10112 VSS.n759 VSS.n758 0.120292
R10113 VSS.n758 VSS.n449 0.120292
R10114 VSS.n452 VSS.n449 0.120292
R10115 VSS.n750 VSS.n452 0.120292
R10116 VSS.n750 VSS.n749 0.120292
R10117 VSS.n749 VSS.n748 0.120292
R10118 VSS.n748 VSS.n453 0.120292
R10119 VSS.n744 VSS.n453 0.120292
R10120 VSS.n744 VSS.n743 0.120292
R10121 VSS.n743 VSS.n456 0.120292
R10122 VSS.n739 VSS.n456 0.120292
R10123 VSS.n739 VSS.n738 0.120292
R10124 VSS.n738 VSS.n737 0.120292
R10125 VSS.n737 VSS.n460 0.120292
R10126 VSS.n462 VSS.n460 0.120292
R10127 VSS.n731 VSS.n462 0.120292
R10128 VSS.n731 VSS.n730 0.120292
R10129 VSS.n730 VSS.n729 0.120292
R10130 VSS.n729 VSS.n465 0.120292
R10131 VSS.n468 VSS.n465 0.120292
R10132 VSS.n724 VSS.n468 0.120292
R10133 VSS.n724 VSS.n723 0.120292
R10134 VSS.n723 VSS.n722 0.120292
R10135 VSS.n722 VSS.n471 0.120292
R10136 VSS.n472 VSS.n471 0.120292
R10137 VSS.n717 VSS.n472 0.120292
R10138 VSS.n717 VSS.n716 0.120292
R10139 VSS.n716 VSS.n715 0.120292
R10140 VSS.n715 VSS.n474 0.120292
R10141 VSS.n711 VSS.n474 0.120292
R10142 VSS.n711 VSS.n710 0.120292
R10143 VSS.n710 VSS.n477 0.120292
R10144 VSS.n706 VSS.n477 0.120292
R10145 VSS.n706 VSS.n705 0.120292
R10146 VSS.n705 VSS.n479 0.120292
R10147 VSS.n697 VSS.n479 0.120292
R10148 VSS.n697 VSS.n696 0.120292
R10149 VSS.n696 VSS.n695 0.120292
R10150 VSS.n695 VSS.n482 0.120292
R10151 VSS.n691 VSS.n482 0.120292
R10152 VSS.n691 VSS.n690 0.120292
R10153 VSS.n690 VSS.n689 0.120292
R10154 VSS.n689 VSS.n485 0.120292
R10155 VSS.n684 VSS.n485 0.120292
R10156 VSS.n678 VSS.n489 0.120292
R10157 VSS.n678 VSS.n677 0.120292
R10158 VSS.n677 VSS.n676 0.120292
R10159 VSS.n676 VSS.n495 0.120292
R10160 VSS.n672 VSS.n495 0.120292
R10161 VSS.n672 VSS.n671 0.120292
R10162 VSS.n671 VSS.n670 0.120292
R10163 VSS.n670 VSS.n499 0.120292
R10164 VSS.n500 VSS.n499 0.120292
R10165 VSS.n665 VSS.n500 0.120292
R10166 VSS.n665 VSS.n664 0.120292
R10167 VSS.n664 VSS.n663 0.120292
R10168 VSS.n663 VSS.n503 0.120292
R10169 VSS.n505 VSS.n503 0.120292
R10170 VSS.n657 VSS.n505 0.120292
R10171 VSS.n657 VSS.n656 0.120292
R10172 VSS.n656 VSS.n655 0.120292
R10173 VSS.n655 VSS.n507 0.120292
R10174 VSS.n650 VSS.n507 0.120292
R10175 VSS.n650 VSS.n649 0.120292
R10176 VSS.n649 VSS.n648 0.120292
R10177 VSS.n648 VSS.n512 0.120292
R10178 VSS.n644 VSS.n512 0.120292
R10179 VSS.n644 VSS.n643 0.120292
R10180 VSS.n643 VSS.n642 0.120292
R10181 VSS.n642 VSS.n515 0.120292
R10182 VSS.n518 VSS.n515 0.120292
R10183 VSS.n520 VSS.n518 0.120292
R10184 VSS.n636 VSS.n520 0.120292
R10185 VSS.n636 VSS.n635 0.120292
R10186 VSS.n635 VSS.n522 0.120292
R10187 VSS.n629 VSS.n522 0.120292
R10188 VSS.n629 VSS.n628 0.120292
R10189 VSS.n628 VSS.n627 0.120292
R10190 VSS.n627 VSS.n525 0.120292
R10191 VSS.n623 VSS.n525 0.120292
R10192 VSS.n623 VSS.n622 0.120292
R10193 VSS.n622 VSS.n528 0.120292
R10194 VSS.n618 VSS.n528 0.120292
R10195 VSS.n618 VSS.n617 0.120292
R10196 VSS.n617 VSS.n616 0.120292
R10197 VSS.n616 VSS.n533 0.120292
R10198 VSS.n610 VSS.n533 0.120292
R10199 VSS.n610 VSS.n609 0.120292
R10200 VSS.n609 VSS.n608 0.120292
R10201 VSS.n608 VSS.n537 0.120292
R10202 VSS.n602 VSS.n537 0.120292
R10203 VSS.n602 VSS.n601 0.120292
R10204 VSS.n601 VSS.n600 0.120292
R10205 VSS.n600 VSS.n539 0.120292
R10206 VSS.n594 VSS.n539 0.120292
R10207 VSS.n594 VSS.n593 0.120292
R10208 VSS.n593 VSS.n592 0.120292
R10209 VSS.n592 VSS.n542 0.120292
R10210 VSS.n546 VSS.n542 0.120292
R10211 VSS.n547 VSS.n546 0.120292
R10212 VSS.n586 VSS.n547 0.120292
R10213 VSS.n586 VSS.n585 0.120292
R10214 VSS.n585 VSS.n550 0.120292
R10215 VSS.n579 VSS.n550 0.120292
R10216 VSS.n579 VSS.n578 0.120292
R10217 VSS.n578 VSS.n577 0.120292
R10218 VSS.n577 VSS.n553 0.120292
R10219 VSS.n555 VSS.n553 0.120292
R10220 VSS.n571 VSS.n555 0.120292
R10221 VSS.n571 VSS.n570 0.120292
R10222 VSS.n570 VSS.n569 0.120292
R10223 VSS.n569 VSS.n559 0.120292
R10224 VSS.n5475 VSS.n5474 0.120292
R10225 VSS.n5474 VSS.n5473 0.120292
R10226 VSS.n5473 VSS.n12 0.120292
R10227 VSS.n5467 VSS.n12 0.120292
R10228 VSS.n5467 VSS.n5466 0.120292
R10229 VSS.n5466 VSS.n5465 0.120292
R10230 VSS.n5465 VSS.n14 0.120292
R10231 VSS.n5459 VSS.n14 0.120292
R10232 VSS.n5459 VSS.n5458 0.120292
R10233 VSS.n5458 VSS.n21 0.120292
R10234 VSS.n5451 VSS.n21 0.120292
R10235 VSS.n5451 VSS.n5450 0.120292
R10236 VSS.n5450 VSS.n24 0.120292
R10237 VSS.n5446 VSS.n24 0.120292
R10238 VSS.n5446 VSS.n5445 0.120292
R10239 VSS.n5445 VSS.n5380 0.120292
R10240 VSS.n5441 VSS.n5380 0.120292
R10241 VSS.n5441 VSS.n5440 0.120292
R10242 VSS.n5440 VSS.n5439 0.120292
R10243 VSS.n5439 VSS.n5384 0.120292
R10244 VSS.n5434 VSS.n5384 0.120292
R10245 VSS.n5434 VSS.n5433 0.120292
R10246 VSS.n5433 VSS.n5432 0.120292
R10247 VSS.n5432 VSS.n5388 0.120292
R10248 VSS.n5425 VSS.n5388 0.120292
R10249 VSS.n5425 VSS.n5424 0.120292
R10250 VSS.n5424 VSS.n5423 0.120292
R10251 VSS.n5423 VSS.n5393 0.120292
R10252 VSS.n5396 VSS.n5393 0.120292
R10253 VSS.n5418 VSS.n5396 0.120292
R10254 VSS.n5418 VSS.n5417 0.120292
R10255 VSS.n5417 VSS.n5416 0.120292
R10256 VSS.n5416 VSS.n5400 0.120292
R10257 VSS.n5412 VSS.n5400 0.120292
R10258 VSS.n5412 VSS.n5411 0.120292
R10259 VSS.n5411 VSS.n5410 0.120292
R10260 VSS.n2073 VSS.n2072 0.120292
R10261 VSS.n2074 VSS.n2073 0.120292
R10262 VSS.n2074 VSS.n2062 0.120292
R10263 VSS.n2080 VSS.n2062 0.120292
R10264 VSS.n2081 VSS.n2080 0.120292
R10265 VSS.n2082 VSS.n2081 0.120292
R10266 VSS.n2082 VSS.n2058 0.120292
R10267 VSS.n2087 VSS.n2058 0.120292
R10268 VSS.n2088 VSS.n2087 0.120292
R10269 VSS.n2089 VSS.n2088 0.120292
R10270 VSS.n2089 VSS.n2055 0.120292
R10271 VSS.n2093 VSS.n2055 0.120292
R10272 VSS.n2094 VSS.n2093 0.120292
R10273 VSS.n2095 VSS.n2094 0.120292
R10274 VSS.n2095 VSS.n2053 0.120292
R10275 VSS.n2100 VSS.n2053 0.120292
R10276 VSS.n2101 VSS.n2100 0.120292
R10277 VSS.n2102 VSS.n2101 0.120292
R10278 VSS.n2102 VSS.n2051 0.120292
R10279 VSS.n2107 VSS.n2051 0.120292
R10280 VSS.n2108 VSS.n2107 0.120292
R10281 VSS.n2109 VSS.n2108 0.120292
R10282 VSS.n2109 VSS.n2048 0.120292
R10283 VSS.n2115 VSS.n2048 0.120292
R10284 VSS.n2116 VSS.n2115 0.120292
R10285 VSS.n2117 VSS.n2116 0.120292
R10286 VSS.n2117 VSS.n2046 0.120292
R10287 VSS.n2124 VSS.n2046 0.120292
R10288 VSS.n2125 VSS.n2124 0.120292
R10289 VSS.n2126 VSS.n2125 0.120292
R10290 VSS.n2126 VSS.n2044 0.120292
R10291 VSS.n2131 VSS.n2044 0.120292
R10292 VSS.n2132 VSS.n2131 0.120292
R10293 VSS.n2133 VSS.n2132 0.120292
R10294 VSS.n2134 VSS.n2133 0.120292
R10295 VSS.n2201 VSS.n2134 0.120292
R10296 VSS.n2201 VSS.n2200 0.120292
R10297 VSS.n2200 VSS.n2199 0.120292
R10298 VSS.n2199 VSS.n2136 0.120292
R10299 VSS.n2192 VSS.n2136 0.120292
R10300 VSS.n2192 VSS.n2191 0.120292
R10301 VSS.n2191 VSS.n2190 0.120292
R10302 VSS.n2190 VSS.n2143 0.120292
R10303 VSS.n2186 VSS.n2143 0.120292
R10304 VSS.n2186 VSS.n2185 0.120292
R10305 VSS.n2185 VSS.n2184 0.120292
R10306 VSS.n2184 VSS.n2145 0.120292
R10307 VSS.n2180 VSS.n2145 0.120292
R10308 VSS.n2180 VSS.n2179 0.120292
R10309 VSS.n2179 VSS.n2178 0.120292
R10310 VSS.n2178 VSS.n2148 0.120292
R10311 VSS.n2174 VSS.n2148 0.120292
R10312 VSS.n2174 VSS.n2173 0.120292
R10313 VSS.n2173 VSS.n2172 0.120292
R10314 VSS.n2172 VSS.n2153 0.120292
R10315 VSS.n2167 VSS.n2153 0.120292
R10316 VSS.n2167 VSS.n2166 0.120292
R10317 VSS.n2166 VSS.n2165 0.120292
R10318 VSS.n2165 VSS.n2156 0.120292
R10319 VSS.n2160 VSS.n2156 0.120292
R10320 VSS.n2160 VSS.n2159 0.120292
R10321 VSS.n2159 VSS.n2042 0.120292
R10322 VSS.n2042 VSS.n2039 0.120292
R10323 VSS.n2210 VSS.n2039 0.120292
R10324 VSS.n2211 VSS.n2210 0.120292
R10325 VSS.n2212 VSS.n2211 0.120292
R10326 VSS.n2212 VSS.n2036 0.120292
R10327 VSS.n2217 VSS.n2036 0.120292
R10328 VSS.n2218 VSS.n2217 0.120292
R10329 VSS.n2219 VSS.n2218 0.120292
R10330 VSS.n2219 VSS.n2033 0.120292
R10331 VSS.n2224 VSS.n2033 0.120292
R10332 VSS.n2225 VSS.n2224 0.120292
R10333 VSS.n2225 VSS.n2030 0.120292
R10334 VSS.n2231 VSS.n2030 0.120292
R10335 VSS.n2232 VSS.n2231 0.120292
R10336 VSS.n2232 VSS.n2026 0.120292
R10337 VSS.n2238 VSS.n2026 0.120292
R10338 VSS.n2239 VSS.n2238 0.120292
R10339 VSS.n2239 VSS.n2022 0.120292
R10340 VSS.n2245 VSS.n2022 0.120292
R10341 VSS.n2246 VSS.n2245 0.120292
R10342 VSS.n2246 VSS.n2019 0.120292
R10343 VSS.n2252 VSS.n2019 0.120292
R10344 VSS.n2253 VSS.n2252 0.120292
R10345 VSS.n2254 VSS.n2253 0.120292
R10346 VSS.n2254 VSS.n2017 0.120292
R10347 VSS.n2261 VSS.n2017 0.120292
R10348 VSS.n2262 VSS.n2261 0.120292
R10349 VSS.n2263 VSS.n2262 0.120292
R10350 VSS.n2333 VSS.n2263 0.120292
R10351 VSS.n2333 VSS.n2332 0.120292
R10352 VSS.n2332 VSS.n2331 0.120292
R10353 VSS.n2331 VSS.n2265 0.120292
R10354 VSS.n2327 VSS.n2265 0.120292
R10355 VSS.n2327 VSS.n2326 0.120292
R10356 VSS.n2326 VSS.n2325 0.120292
R10357 VSS.n2325 VSS.n2267 0.120292
R10358 VSS.n2317 VSS.n2267 0.120292
R10359 VSS.n2317 VSS.n2316 0.120292
R10360 VSS.n2316 VSS.n2315 0.120292
R10361 VSS.n2315 VSS.n2271 0.120292
R10362 VSS.n2307 VSS.n2271 0.120292
R10363 VSS.n2307 VSS.n2306 0.120292
R10364 VSS.n2306 VSS.n2305 0.120292
R10365 VSS.n2305 VSS.n2273 0.120292
R10366 VSS.n2300 VSS.n2273 0.120292
R10367 VSS.n2300 VSS.n2299 0.120292
R10368 VSS.n2299 VSS.n2277 0.120292
R10369 VSS.n2292 VSS.n2277 0.120292
R10370 VSS.n2292 VSS.n2291 0.120292
R10371 VSS.n2291 VSS.n2290 0.120292
R10372 VSS.n2290 VSS.n2280 0.120292
R10373 VSS.n2282 VSS.n2280 0.120292
R10374 VSS.n2285 VSS.n2282 0.120292
R10375 VSS.n2285 VSS.n2284 0.120292
R10376 VSS.n2284 VSS.n2014 0.120292
R10377 VSS.n2339 VSS.n2014 0.120292
R10378 VSS.n2340 VSS.n2339 0.120292
R10379 VSS.n2341 VSS.n2340 0.120292
R10380 VSS.n2341 VSS.n2012 0.120292
R10381 VSS.n2346 VSS.n2012 0.120292
R10382 VSS.n2347 VSS.n2346 0.120292
R10383 VSS.n2348 VSS.n2347 0.120292
R10384 VSS.n2348 VSS.n2010 0.120292
R10385 VSS.n2353 VSS.n2010 0.120292
R10386 VSS.n2354 VSS.n2353 0.120292
R10387 VSS.n2355 VSS.n2354 0.120292
R10388 VSS.n2355 VSS.n2007 0.120292
R10389 VSS.n2361 VSS.n2007 0.120292
R10390 VSS.n2362 VSS.n2361 0.120292
R10391 VSS.n2363 VSS.n2362 0.120292
R10392 VSS.n2363 VSS.n2005 0.120292
R10393 VSS.n2367 VSS.n2005 0.120292
R10394 VSS.n2368 VSS.n2367 0.120292
R10395 VSS.n2368 VSS.n2002 0.120292
R10396 VSS.n2377 VSS.n2002 0.120292
R10397 VSS.n2378 VSS.n2377 0.120292
R10398 VSS.n2379 VSS.n2378 0.120292
R10399 VSS.n2379 VSS.n2000 0.120292
R10400 VSS.n2385 VSS.n2000 0.120292
R10401 VSS.n2386 VSS.n2385 0.120292
R10402 VSS.n2387 VSS.n2386 0.120292
R10403 VSS.n2387 VSS.n1998 0.120292
R10404 VSS.n2393 VSS.n1998 0.120292
R10405 VSS.n2470 VSS.n2393 0.120292
R10406 VSS.n2470 VSS.n2469 0.120292
R10407 VSS.n2469 VSS.n2468 0.120292
R10408 VSS.n2468 VSS.n2394 0.120292
R10409 VSS.n2464 VSS.n2394 0.120292
R10410 VSS.n2464 VSS.n2463 0.120292
R10411 VSS.n2463 VSS.n2462 0.120292
R10412 VSS.n2462 VSS.n2398 0.120292
R10413 VSS.n2400 VSS.n2398 0.120292
R10414 VSS.n2453 VSS.n2400 0.120292
R10415 VSS.n2453 VSS.n2452 0.120292
R10416 VSS.n2452 VSS.n2451 0.120292
R10417 VSS.n2451 VSS.n2403 0.120292
R10418 VSS.n2445 VSS.n2403 0.120292
R10419 VSS.n2445 VSS.n2444 0.120292
R10420 VSS.n2444 VSS.n2443 0.120292
R10421 VSS.n2443 VSS.n2407 0.120292
R10422 VSS.n2438 VSS.n2407 0.120292
R10423 VSS.n2438 VSS.n2437 0.120292
R10424 VSS.n2437 VSS.n2412 0.120292
R10425 VSS.n2433 VSS.n2412 0.120292
R10426 VSS.n2433 VSS.n2432 0.120292
R10427 VSS.n2432 VSS.n2431 0.120292
R10428 VSS.n2431 VSS.n2415 0.120292
R10429 VSS.n2427 VSS.n2415 0.120292
R10430 VSS.n2427 VSS.n2426 0.120292
R10431 VSS.n2426 VSS.n2419 0.120292
R10432 VSS.n2419 VSS.n1992 0.120292
R10433 VSS.n2476 VSS.n1992 0.120292
R10434 VSS.n2477 VSS.n2476 0.120292
R10435 VSS.n2477 VSS.n1988 0.120292
R10436 VSS.n2482 VSS.n1988 0.120292
R10437 VSS.n2483 VSS.n2482 0.120292
R10438 VSS.n2483 VSS.n1986 0.120292
R10439 VSS.n2494 VSS.n1986 0.120292
R10440 VSS.n2495 VSS.n2494 0.120292
R10441 VSS.n2495 VSS.n1984 0.120292
R10442 VSS.n2500 VSS.n1984 0.120292
R10443 VSS.n2501 VSS.n2500 0.120292
R10444 VSS.n2501 VSS.n1981 0.120292
R10445 VSS.n2506 VSS.n1981 0.120292
R10446 VSS.n2507 VSS.n2506 0.120292
R10447 VSS.n2508 VSS.n2507 0.120292
R10448 VSS.n2508 VSS.n1978 0.120292
R10449 VSS.n2513 VSS.n1978 0.120292
R10450 VSS.n2514 VSS.n2513 0.120292
R10451 VSS.n2515 VSS.n2514 0.120292
R10452 VSS.n2515 VSS.n1976 0.120292
R10453 VSS.n2522 VSS.n1976 0.120292
R10454 VSS.n2523 VSS.n2522 0.120292
R10455 VSS.n2523 VSS.n1974 0.120292
R10456 VSS.n2529 VSS.n1974 0.120292
R10457 VSS.n2530 VSS.n2529 0.120292
R10458 VSS.n2531 VSS.n2530 0.120292
R10459 VSS.n2531 VSS.n1971 0.120292
R10460 VSS.n2535 VSS.n1971 0.120292
R10461 VSS.n2536 VSS.n2535 0.120292
R10462 VSS.n2537 VSS.n2536 0.120292
R10463 VSS.n2537 VSS.n1969 0.120292
R10464 VSS.n2541 VSS.n1969 0.120292
R10465 VSS.n2542 VSS.n2541 0.120292
R10466 VSS.n2543 VSS.n2542 0.120292
R10467 VSS.n2543 VSS.n1967 0.120292
R10468 VSS.n2548 VSS.n1967 0.120292
R10469 VSS.n2549 VSS.n2548 0.120292
R10470 VSS.n2550 VSS.n2549 0.120292
R10471 VSS.n2550 VSS.n1965 0.120292
R10472 VSS.n2558 VSS.n1965 0.120292
R10473 VSS.n2559 VSS.n2558 0.120292
R10474 VSS.n2560 VSS.n2559 0.120292
R10475 VSS.n2560 VSS.n1962 0.120292
R10476 VSS.n2564 VSS.n1962 0.120292
R10477 VSS.n2565 VSS.n2564 0.120292
R10478 VSS.n2565 VSS.n1959 0.120292
R10479 VSS.n2572 VSS.n1959 0.120292
R10480 VSS.n2573 VSS.n2572 0.120292
R10481 VSS.n2574 VSS.n2573 0.120292
R10482 VSS.n2574 VSS.n1956 0.120292
R10483 VSS.n2580 VSS.n1956 0.120292
R10484 VSS.n2581 VSS.n2580 0.120292
R10485 VSS.n2582 VSS.n2581 0.120292
R10486 VSS.n2582 VSS.n1953 0.120292
R10487 VSS.n2590 VSS.n1953 0.120292
R10488 VSS.n2591 VSS.n2590 0.120292
R10489 VSS.n2632 VSS.n2591 0.120292
R10490 VSS.n2632 VSS.n2631 0.120292
R10491 VSS.n2631 VSS.n2592 0.120292
R10492 VSS.n2626 VSS.n2592 0.120292
R10493 VSS.n2626 VSS.n2625 0.120292
R10494 VSS.n2625 VSS.n2596 0.120292
R10495 VSS.n2599 VSS.n2596 0.120292
R10496 VSS.n2619 VSS.n2599 0.120292
R10497 VSS.n2619 VSS.n2618 0.120292
R10498 VSS.n2618 VSS.n2617 0.120292
R10499 VSS.n2617 VSS.n2602 0.120292
R10500 VSS.n2613 VSS.n2602 0.120292
R10501 VSS.n2613 VSS.n2612 0.120292
R10502 VSS.n2728 VSS.n2727 0.120292
R10503 VSS.n2727 VSS.n2726 0.120292
R10504 VSS.n2726 VSS.n1940 0.120292
R10505 VSS.n2722 VSS.n1940 0.120292
R10506 VSS.n2722 VSS.n2721 0.120292
R10507 VSS.n2721 VSS.n1944 0.120292
R10508 VSS.n2713 VSS.n1944 0.120292
R10509 VSS.n2713 VSS.n2712 0.120292
R10510 VSS.n2712 VSS.n2711 0.120292
R10511 VSS.n2711 VSS.n1946 0.120292
R10512 VSS.n2707 VSS.n1946 0.120292
R10513 VSS.n2707 VSS.n2706 0.120292
R10514 VSS.n2706 VSS.n2705 0.120292
R10515 VSS.n2705 VSS.n2637 0.120292
R10516 VSS.n2699 VSS.n2637 0.120292
R10517 VSS.n2699 VSS.n2698 0.120292
R10518 VSS.n2698 VSS.n2697 0.120292
R10519 VSS.n2697 VSS.n2640 0.120292
R10520 VSS.n2691 VSS.n2640 0.120292
R10521 VSS.n2691 VSS.n2690 0.120292
R10522 VSS.n2690 VSS.n2689 0.120292
R10523 VSS.n2689 VSS.n2644 0.120292
R10524 VSS.n2684 VSS.n2644 0.120292
R10525 VSS.n2684 VSS.n2683 0.120292
R10526 VSS.n2683 VSS.n2682 0.120292
R10527 VSS.n2682 VSS.n2647 0.120292
R10528 VSS.n2648 VSS.n2647 0.120292
R10529 VSS.n2677 VSS.n2648 0.120292
R10530 VSS.n2677 VSS.n2676 0.120292
R10531 VSS.n2676 VSS.n2675 0.120292
R10532 VSS.n2675 VSS.n2651 0.120292
R10533 VSS.n2669 VSS.n2651 0.120292
R10534 VSS.n2669 VSS.n2668 0.120292
R10535 VSS.n2668 VSS.n2667 0.120292
R10536 VSS.n2667 VSS.n2655 0.120292
R10537 VSS.n2663 VSS.n2655 0.120292
R10538 VSS.n3045 VSS.n3044 0.120292
R10539 VSS.n3046 VSS.n3045 0.120292
R10540 VSS.n3046 VSS.n3034 0.120292
R10541 VSS.n3051 VSS.n3034 0.120292
R10542 VSS.n3052 VSS.n3051 0.120292
R10543 VSS.n3053 VSS.n3052 0.120292
R10544 VSS.n3053 VSS.n3030 0.120292
R10545 VSS.n3057 VSS.n3030 0.120292
R10546 VSS.n3058 VSS.n3057 0.120292
R10547 VSS.n3059 VSS.n3058 0.120292
R10548 VSS.n3059 VSS.n3026 0.120292
R10549 VSS.n3063 VSS.n3026 0.120292
R10550 VSS.n3064 VSS.n3063 0.120292
R10551 VSS.n3065 VSS.n3064 0.120292
R10552 VSS.n3065 VSS.n3023 0.120292
R10553 VSS.n3070 VSS.n3023 0.120292
R10554 VSS.n3071 VSS.n3070 0.120292
R10555 VSS.n3072 VSS.n3071 0.120292
R10556 VSS.n3072 VSS.n3020 0.120292
R10557 VSS.n3078 VSS.n3020 0.120292
R10558 VSS.n3079 VSS.n3078 0.120292
R10559 VSS.n3080 VSS.n3079 0.120292
R10560 VSS.n3080 VSS.n3017 0.120292
R10561 VSS.n3089 VSS.n3017 0.120292
R10562 VSS.n3090 VSS.n3089 0.120292
R10563 VSS.n3091 VSS.n3090 0.120292
R10564 VSS.n3091 VSS.n3015 0.120292
R10565 VSS.n3095 VSS.n3015 0.120292
R10566 VSS.n3096 VSS.n3095 0.120292
R10567 VSS.n3097 VSS.n3096 0.120292
R10568 VSS.n3097 VSS.n3012 0.120292
R10569 VSS.n3105 VSS.n3012 0.120292
R10570 VSS.n3106 VSS.n3105 0.120292
R10571 VSS.n3107 VSS.n3106 0.120292
R10572 VSS.n3107 VSS.n3008 0.120292
R10573 VSS.n3112 VSS.n3008 0.120292
R10574 VSS.n3113 VSS.n3112 0.120292
R10575 VSS.n3114 VSS.n3113 0.120292
R10576 VSS.n3114 VSS.n3006 0.120292
R10577 VSS.n3119 VSS.n3006 0.120292
R10578 VSS.n3120 VSS.n3119 0.120292
R10579 VSS.n3120 VSS.n3003 0.120292
R10580 VSS.n3124 VSS.n3003 0.120292
R10581 VSS.n3125 VSS.n3124 0.120292
R10582 VSS.n3125 VSS.n3000 0.120292
R10583 VSS.n3132 VSS.n3000 0.120292
R10584 VSS.n3133 VSS.n3132 0.120292
R10585 VSS.n3134 VSS.n3133 0.120292
R10586 VSS.n3134 VSS.n2998 0.120292
R10587 VSS.n3138 VSS.n2998 0.120292
R10588 VSS.n3139 VSS.n3138 0.120292
R10589 VSS.n3140 VSS.n3139 0.120292
R10590 VSS.n3140 VSS.n2995 0.120292
R10591 VSS.n3145 VSS.n2995 0.120292
R10592 VSS.n3146 VSS.n3145 0.120292
R10593 VSS.n3146 VSS.n2991 0.120292
R10594 VSS.n3154 VSS.n2991 0.120292
R10595 VSS.n3155 VSS.n3154 0.120292
R10596 VSS.n3156 VSS.n3155 0.120292
R10597 VSS.n3156 VSS.n2989 0.120292
R10598 VSS.n3164 VSS.n2989 0.120292
R10599 VSS.n3165 VSS.n3164 0.120292
R10600 VSS.n3166 VSS.n3165 0.120292
R10601 VSS.n3166 VSS.n2987 0.120292
R10602 VSS.n3173 VSS.n2987 0.120292
R10603 VSS.n3174 VSS.n3173 0.120292
R10604 VSS.n3175 VSS.n3174 0.120292
R10605 VSS.n3175 VSS.n2985 0.120292
R10606 VSS.n3179 VSS.n2985 0.120292
R10607 VSS.n3180 VSS.n3179 0.120292
R10608 VSS.n3181 VSS.n3180 0.120292
R10609 VSS.n3181 VSS.n2982 0.120292
R10610 VSS.n3189 VSS.n2982 0.120292
R10611 VSS.n3190 VSS.n3189 0.120292
R10612 VSS.n3191 VSS.n3190 0.120292
R10613 VSS.n3191 VSS.n2978 0.120292
R10614 VSS.n3196 VSS.n2978 0.120292
R10615 VSS.n3197 VSS.n3196 0.120292
R10616 VSS.n3197 VSS.n2976 0.120292
R10617 VSS.n3202 VSS.n2976 0.120292
R10618 VSS.n3203 VSS.n3202 0.120292
R10619 VSS.n3204 VSS.n3203 0.120292
R10620 VSS.n3204 VSS.n2974 0.120292
R10621 VSS.n3209 VSS.n2974 0.120292
R10622 VSS.n3210 VSS.n3209 0.120292
R10623 VSS.n3211 VSS.n3210 0.120292
R10624 VSS.n3211 VSS.n2971 0.120292
R10625 VSS.n3215 VSS.n2971 0.120292
R10626 VSS.n3216 VSS.n3215 0.120292
R10627 VSS.n3217 VSS.n3216 0.120292
R10628 VSS.n3218 VSS.n3217 0.120292
R10629 VSS.n3289 VSS.n3218 0.120292
R10630 VSS.n3289 VSS.n3288 0.120292
R10631 VSS.n3288 VSS.n3221 0.120292
R10632 VSS.n3283 VSS.n3221 0.120292
R10633 VSS.n3283 VSS.n3282 0.120292
R10634 VSS.n3282 VSS.n3225 0.120292
R10635 VSS.n3228 VSS.n3225 0.120292
R10636 VSS.n3276 VSS.n3228 0.120292
R10637 VSS.n3276 VSS.n3275 0.120292
R10638 VSS.n3275 VSS.n3230 0.120292
R10639 VSS.n3271 VSS.n3230 0.120292
R10640 VSS.n3271 VSS.n3270 0.120292
R10641 VSS.n3270 VSS.n3233 0.120292
R10642 VSS.n3266 VSS.n3233 0.120292
R10643 VSS.n3266 VSS.n3265 0.120292
R10644 VSS.n3265 VSS.n3235 0.120292
R10645 VSS.n3260 VSS.n3235 0.120292
R10646 VSS.n3260 VSS.n3259 0.120292
R10647 VSS.n3259 VSS.n3258 0.120292
R10648 VSS.n3258 VSS.n3238 0.120292
R10649 VSS.n3254 VSS.n3238 0.120292
R10650 VSS.n3254 VSS.n3253 0.120292
R10651 VSS.n3253 VSS.n3240 0.120292
R10652 VSS.n3248 VSS.n3240 0.120292
R10653 VSS.n3248 VSS.n3247 0.120292
R10654 VSS.n3247 VSS.n2968 0.120292
R10655 VSS.n3296 VSS.n2968 0.120292
R10656 VSS.n3297 VSS.n3296 0.120292
R10657 VSS.n3298 VSS.n3297 0.120292
R10658 VSS.n3298 VSS.n2964 0.120292
R10659 VSS.n3306 VSS.n2964 0.120292
R10660 VSS.n3307 VSS.n3306 0.120292
R10661 VSS.n3307 VSS.n2962 0.120292
R10662 VSS.n3313 VSS.n2962 0.120292
R10663 VSS.n3314 VSS.n3313 0.120292
R10664 VSS.n3315 VSS.n3314 0.120292
R10665 VSS.n3315 VSS.n2959 0.120292
R10666 VSS.n3323 VSS.n2959 0.120292
R10667 VSS.n3324 VSS.n3323 0.120292
R10668 VSS.n3324 VSS.n2957 0.120292
R10669 VSS.n3330 VSS.n2957 0.120292
R10670 VSS.n3331 VSS.n3330 0.120292
R10671 VSS.n3331 VSS.n2953 0.120292
R10672 VSS.n3336 VSS.n2953 0.120292
R10673 VSS.n3337 VSS.n3336 0.120292
R10674 VSS.n3337 VSS.n2950 0.120292
R10675 VSS.n3341 VSS.n2950 0.120292
R10676 VSS.n3342 VSS.n3341 0.120292
R10677 VSS.n3342 VSS.n2948 0.120292
R10678 VSS.n2948 VSS.n2945 0.120292
R10679 VSS.n3349 VSS.n2945 0.120292
R10680 VSS.n3350 VSS.n3349 0.120292
R10681 VSS.n3351 VSS.n3350 0.120292
R10682 VSS.n3351 VSS.n2943 0.120292
R10683 VSS.n2943 VSS.n2939 0.120292
R10684 VSS.n3357 VSS.n2939 0.120292
R10685 VSS.n3358 VSS.n3357 0.120292
R10686 VSS.n3359 VSS.n3358 0.120292
R10687 VSS.n3359 VSS.n2936 0.120292
R10688 VSS.n3363 VSS.n2936 0.120292
R10689 VSS.n3364 VSS.n3363 0.120292
R10690 VSS.n3364 VSS.n2932 0.120292
R10691 VSS.n3368 VSS.n2932 0.120292
R10692 VSS.n3369 VSS.n3368 0.120292
R10693 VSS.n3370 VSS.n3369 0.120292
R10694 VSS.n3370 VSS.n2928 0.120292
R10695 VSS.n3375 VSS.n2928 0.120292
R10696 VSS.n3376 VSS.n3375 0.120292
R10697 VSS.n3377 VSS.n3376 0.120292
R10698 VSS.n3377 VSS.n2926 0.120292
R10699 VSS.n3381 VSS.n2926 0.120292
R10700 VSS.n3382 VSS.n3381 0.120292
R10701 VSS.n3383 VSS.n3382 0.120292
R10702 VSS.n3383 VSS.n2923 0.120292
R10703 VSS.n3389 VSS.n2923 0.120292
R10704 VSS.n3390 VSS.n3389 0.120292
R10705 VSS.n3390 VSS.n2919 0.120292
R10706 VSS.n3396 VSS.n2919 0.120292
R10707 VSS.n3397 VSS.n3396 0.120292
R10708 VSS.n3398 VSS.n3397 0.120292
R10709 VSS.n3398 VSS.n2916 0.120292
R10710 VSS.n3403 VSS.n2916 0.120292
R10711 VSS.n3404 VSS.n3403 0.120292
R10712 VSS.n3405 VSS.n3404 0.120292
R10713 VSS.n3405 VSS.n2913 0.120292
R10714 VSS.n3411 VSS.n2913 0.120292
R10715 VSS.n3412 VSS.n3411 0.120292
R10716 VSS.n3413 VSS.n3412 0.120292
R10717 VSS.n3413 VSS.n2910 0.120292
R10718 VSS.n3421 VSS.n2910 0.120292
R10719 VSS.n3422 VSS.n3421 0.120292
R10720 VSS.n3422 VSS.n2907 0.120292
R10721 VSS.n3426 VSS.n2907 0.120292
R10722 VSS.n3427 VSS.n3426 0.120292
R10723 VSS.n3428 VSS.n3427 0.120292
R10724 VSS.n3428 VSS.n2904 0.120292
R10725 VSS.n3432 VSS.n2904 0.120292
R10726 VSS.n3433 VSS.n3432 0.120292
R10727 VSS.n3434 VSS.n3433 0.120292
R10728 VSS.n3434 VSS.n2901 0.120292
R10729 VSS.n3438 VSS.n2901 0.120292
R10730 VSS.n3439 VSS.n3438 0.120292
R10731 VSS.n3440 VSS.n3439 0.120292
R10732 VSS.n3440 VSS.n2899 0.120292
R10733 VSS.n2899 VSS.n2898 0.120292
R10734 VSS.n3450 VSS.n2898 0.120292
R10735 VSS.n3451 VSS.n3450 0.120292
R10736 VSS.n3452 VSS.n3451 0.120292
R10737 VSS.n3452 VSS.n2896 0.120292
R10738 VSS.n2896 VSS.n2790 0.120292
R10739 VSS.n3458 VSS.n2790 0.120292
R10740 VSS.n3459 VSS.n3458 0.120292
R10741 VSS.n3460 VSS.n3459 0.120292
R10742 VSS.n3460 VSS.n2787 0.120292
R10743 VSS.n3466 VSS.n2787 0.120292
R10744 VSS.n3467 VSS.n3466 0.120292
R10745 VSS.n3468 VSS.n3467 0.120292
R10746 VSS.n3468 VSS.n2785 0.120292
R10747 VSS.n3476 VSS.n2785 0.120292
R10748 VSS.n3477 VSS.n3476 0.120292
R10749 VSS.n3478 VSS.n3477 0.120292
R10750 VSS.n3478 VSS.n2781 0.120292
R10751 VSS.n3482 VSS.n2781 0.120292
R10752 VSS.n3483 VSS.n3482 0.120292
R10753 VSS.n3484 VSS.n3483 0.120292
R10754 VSS.n3484 VSS.n2778 0.120292
R10755 VSS.n2778 VSS.n2775 0.120292
R10756 VSS.n3489 VSS.n2775 0.120292
R10757 VSS.n3490 VSS.n3489 0.120292
R10758 VSS.n3490 VSS.n2772 0.120292
R10759 VSS.n3494 VSS.n2772 0.120292
R10760 VSS.n3495 VSS.n3494 0.120292
R10761 VSS.n3496 VSS.n3495 0.120292
R10762 VSS.n3496 VSS.n2770 0.120292
R10763 VSS.n3501 VSS.n2770 0.120292
R10764 VSS.n3502 VSS.n3501 0.120292
R10765 VSS.n3502 VSS.n2766 0.120292
R10766 VSS.n3507 VSS.n2766 0.120292
R10767 VSS.n3508 VSS.n3507 0.120292
R10768 VSS.n3509 VSS.n3508 0.120292
R10769 VSS.n3509 VSS.n2761 0.120292
R10770 VSS.n3515 VSS.n2761 0.120292
R10771 VSS.n3516 VSS.n3515 0.120292
R10772 VSS.n3516 VSS.n2759 0.120292
R10773 VSS.n2759 VSS.n2758 0.120292
R10774 VSS.n3527 VSS.n2758 0.120292
R10775 VSS.n3528 VSS.n3527 0.120292
R10776 VSS.n3529 VSS.n3528 0.120292
R10777 VSS.n3529 VSS.n2755 0.120292
R10778 VSS.n2755 VSS.n2753 0.120292
R10779 VSS.n3534 VSS.n2753 0.120292
R10780 VSS.n3549 VSS.n2748 0.120292
R10781 VSS.n2867 VSS.n2748 0.120292
R10782 VSS.n2867 VSS.n2866 0.120292
R10783 VSS.n2866 VSS.n2863 0.120292
R10784 VSS.n2872 VSS.n2863 0.120292
R10785 VSS.n2873 VSS.n2872 0.120292
R10786 VSS.n2874 VSS.n2873 0.120292
R10787 VSS.n2874 VSS.n2861 0.120292
R10788 VSS.n2885 VSS.n2861 0.120292
R10789 VSS.n2886 VSS.n2885 0.120292
R10790 VSS.n2887 VSS.n2886 0.120292
R10791 VSS.n2887 VSS.n2859 0.120292
R10792 VSS.n2859 VSS.n2858 0.120292
R10793 VSS.n2858 VSS.n2857 0.120292
R10794 VSS.n2857 VSS.n2792 0.120292
R10795 VSS.n2851 VSS.n2792 0.120292
R10796 VSS.n2851 VSS.n2850 0.120292
R10797 VSS.n2850 VSS.n2849 0.120292
R10798 VSS.n2849 VSS.n2794 0.120292
R10799 VSS.n2843 VSS.n2794 0.120292
R10800 VSS.n2843 VSS.n2842 0.120292
R10801 VSS.n2842 VSS.n2841 0.120292
R10802 VSS.n2841 VSS.n2798 0.120292
R10803 VSS.n2835 VSS.n2798 0.120292
R10804 VSS.n2835 VSS.n2834 0.120292
R10805 VSS.n2834 VSS.n2833 0.120292
R10806 VSS.n2833 VSS.n2800 0.120292
R10807 VSS.n2828 VSS.n2800 0.120292
R10808 VSS.n2828 VSS.n2827 0.120292
R10809 VSS.n2827 VSS.n2826 0.120292
R10810 VSS.n2826 VSS.n2802 0.120292
R10811 VSS.n2820 VSS.n2802 0.120292
R10812 VSS.n2820 VSS.n2819 0.120292
R10813 VSS.n2819 VSS.n2818 0.120292
R10814 VSS.n2818 VSS.n2806 0.120292
R10815 VSS.n2812 VSS.n2806 0.120292
R10816 VSS.n971 VSS.n970 0.120292
R10817 VSS.n972 VSS.n971 0.120292
R10818 VSS.n972 VSS.n960 0.120292
R10819 VSS.n982 VSS.n960 0.120292
R10820 VSS.n983 VSS.n982 0.120292
R10821 VSS.n1716 VSS.n983 0.120292
R10822 VSS.n1716 VSS.n1715 0.120292
R10823 VSS.n1715 VSS.n1714 0.120292
R10824 VSS.n1714 VSS.n984 0.120292
R10825 VSS.n1708 VSS.n984 0.120292
R10826 VSS.n1705 VSS.n991 0.120292
R10827 VSS.n1699 VSS.n991 0.120292
R10828 VSS.n1699 VSS.n1698 0.120292
R10829 VSS.n1698 VSS.n1697 0.120292
R10830 VSS.n1697 VSS.n993 0.120292
R10831 VSS.n1692 VSS.n993 0.120292
R10832 VSS.n1692 VSS.n1691 0.120292
R10833 VSS.n1691 VSS.n997 0.120292
R10834 VSS.n1687 VSS.n997 0.120292
R10835 VSS.n1687 VSS.n1686 0.120292
R10836 VSS.n1686 VSS.n1685 0.120292
R10837 VSS.n1685 VSS.n1000 0.120292
R10838 VSS.n1681 VSS.n1000 0.120292
R10839 VSS.n1681 VSS.n1680 0.120292
R10840 VSS.n1680 VSS.n1679 0.120292
R10841 VSS.n1679 VSS.n1002 0.120292
R10842 VSS.n1674 VSS.n1002 0.120292
R10843 VSS.n1674 VSS.n1673 0.120292
R10844 VSS.n1673 VSS.n1672 0.120292
R10845 VSS.n1672 VSS.n1005 0.120292
R10846 VSS.n1668 VSS.n1005 0.120292
R10847 VSS.n1668 VSS.n1667 0.120292
R10848 VSS.n1667 VSS.n1666 0.120292
R10849 VSS.n1666 VSS.n1008 0.120292
R10850 VSS.n1662 VSS.n1008 0.120292
R10851 VSS.n1662 VSS.n1661 0.120292
R10852 VSS.n1661 VSS.n1660 0.120292
R10853 VSS.n1660 VSS.n1013 0.120292
R10854 VSS.n1654 VSS.n1013 0.120292
R10855 VSS.n1654 VSS.n1653 0.120292
R10856 VSS.n1653 VSS.n1652 0.120292
R10857 VSS.n1652 VSS.n1016 0.120292
R10858 VSS.n1647 VSS.n1016 0.120292
R10859 VSS.n1647 VSS.n1646 0.120292
R10860 VSS.n1646 VSS.n1645 0.120292
R10861 VSS.n1645 VSS.n1018 0.120292
R10862 VSS.n1639 VSS.n1018 0.120292
R10863 VSS.n1639 VSS.n1638 0.120292
R10864 VSS.n1638 VSS.n1637 0.120292
R10865 VSS.n1637 VSS.n1021 0.120292
R10866 VSS.n1632 VSS.n1021 0.120292
R10867 VSS.n1632 VSS.n1631 0.120292
R10868 VSS.n1631 VSS.n1630 0.120292
R10869 VSS.n1630 VSS.n1024 0.120292
R10870 VSS.n1026 VSS.n1024 0.120292
R10871 VSS.n1051 VSS.n1026 0.120292
R10872 VSS.n1053 VSS.n1051 0.120292
R10873 VSS.n1054 VSS.n1053 0.120292
R10874 VSS.n1055 VSS.n1054 0.120292
R10875 VSS.n1055 VSS.n1047 0.120292
R10876 VSS.n1060 VSS.n1047 0.120292
R10877 VSS.n1061 VSS.n1060 0.120292
R10878 VSS.n1062 VSS.n1061 0.120292
R10879 VSS.n1062 VSS.n1044 0.120292
R10880 VSS.n1068 VSS.n1044 0.120292
R10881 VSS.n1069 VSS.n1068 0.120292
R10882 VSS.n1070 VSS.n1069 0.120292
R10883 VSS.n1070 VSS.n1042 0.120292
R10884 VSS.n1074 VSS.n1042 0.120292
R10885 VSS.n1075 VSS.n1074 0.120292
R10886 VSS.n1076 VSS.n1075 0.120292
R10887 VSS.n1076 VSS.n1039 0.120292
R10888 VSS.n1039 VSS.n1036 0.120292
R10889 VSS.n1081 VSS.n1036 0.120292
R10890 VSS.n1082 VSS.n1081 0.120292
R10891 VSS.n1083 VSS.n1082 0.120292
R10892 VSS.n1083 VSS.n1033 0.120292
R10893 VSS.n1089 VSS.n1033 0.120292
R10894 VSS.n1090 VSS.n1089 0.120292
R10895 VSS.n1091 VSS.n1090 0.120292
R10896 VSS.n1091 VSS.n1030 0.120292
R10897 VSS.n1096 VSS.n1030 0.120292
R10898 VSS.n1623 VSS.n1096 0.120292
R10899 VSS.n1623 VSS.n1622 0.120292
R10900 VSS.n1622 VSS.n1621 0.120292
R10901 VSS.n1621 VSS.n1097 0.120292
R10902 VSS.n1616 VSS.n1097 0.120292
R10903 VSS.n1616 VSS.n1615 0.120292
R10904 VSS.n1615 VSS.n1614 0.120292
R10905 VSS.n1614 VSS.n1100 0.120292
R10906 VSS.n1609 VSS.n1100 0.120292
R10907 VSS.n1609 VSS.n1608 0.120292
R10908 VSS.n1608 VSS.n1607 0.120292
R10909 VSS.n1607 VSS.n1102 0.120292
R10910 VSS.n1599 VSS.n1102 0.120292
R10911 VSS.n1599 VSS.n1598 0.120292
R10912 VSS.n1598 VSS.n1597 0.120292
R10913 VSS.n1597 VSS.n1105 0.120292
R10914 VSS.n1592 VSS.n1105 0.120292
R10915 VSS.n1592 VSS.n1591 0.120292
R10916 VSS.n1591 VSS.n1590 0.120292
R10917 VSS.n1590 VSS.n1107 0.120292
R10918 VSS.n1585 VSS.n1107 0.120292
R10919 VSS.n1585 VSS.n1584 0.120292
R10920 VSS.n1584 VSS.n1111 0.120292
R10921 VSS.n1577 VSS.n1111 0.120292
R10922 VSS.n1577 VSS.n1576 0.120292
R10923 VSS.n1576 VSS.n1113 0.120292
R10924 VSS.n1572 VSS.n1113 0.120292
R10925 VSS.n1572 VSS.n1571 0.120292
R10926 VSS.n1571 VSS.n1570 0.120292
R10927 VSS.n1570 VSS.n1117 0.120292
R10928 VSS.n1520 VSS.n1117 0.120292
R10929 VSS.n1521 VSS.n1520 0.120292
R10930 VSS.n1521 VSS.n1517 0.120292
R10931 VSS.n1525 VSS.n1517 0.120292
R10932 VSS.n1526 VSS.n1525 0.120292
R10933 VSS.n1527 VSS.n1526 0.120292
R10934 VSS.n1527 VSS.n1515 0.120292
R10935 VSS.n1515 VSS.n1513 0.120292
R10936 VSS.n1532 VSS.n1513 0.120292
R10937 VSS.n1533 VSS.n1532 0.120292
R10938 VSS.n1533 VSS.n1510 0.120292
R10939 VSS.n1538 VSS.n1510 0.120292
R10940 VSS.n1539 VSS.n1538 0.120292
R10941 VSS.n1540 VSS.n1539 0.120292
R10942 VSS.n1540 VSS.n1507 0.120292
R10943 VSS.n1507 VSS.n1506 0.120292
R10944 VSS.n1546 VSS.n1506 0.120292
R10945 VSS.n1547 VSS.n1546 0.120292
R10946 VSS.n1547 VSS.n1503 0.120292
R10947 VSS.n1551 VSS.n1503 0.120292
R10948 VSS.n1552 VSS.n1551 0.120292
R10949 VSS.n1553 VSS.n1552 0.120292
R10950 VSS.n1553 VSS.n1498 0.120292
R10951 VSS.n1561 VSS.n1498 0.120292
R10952 VSS.n1562 VSS.n1561 0.120292
R10953 VSS.n1563 VSS.n1562 0.120292
R10954 VSS.n1563 VSS.n1495 0.120292
R10955 VSS.n1495 VSS.n1494 0.120292
R10956 VSS.n1494 VSS.n1493 0.120292
R10957 VSS.n1493 VSS.n1121 0.120292
R10958 VSS.n1488 VSS.n1121 0.120292
R10959 VSS.n1488 VSS.n1487 0.120292
R10960 VSS.n1487 VSS.n1124 0.120292
R10961 VSS.n1482 VSS.n1124 0.120292
R10962 VSS.n1482 VSS.n1481 0.120292
R10963 VSS.n1481 VSS.n1480 0.120292
R10964 VSS.n1480 VSS.n1127 0.120292
R10965 VSS.n1476 VSS.n1127 0.120292
R10966 VSS.n1476 VSS.n1475 0.120292
R10967 VSS.n1475 VSS.n1130 0.120292
R10968 VSS.n1471 VSS.n1130 0.120292
R10969 VSS.n1471 VSS.n1470 0.120292
R10970 VSS.n1470 VSS.n1469 0.120292
R10971 VSS.n1469 VSS.n1135 0.120292
R10972 VSS.n1465 VSS.n1135 0.120292
R10973 VSS.n1465 VSS.n1464 0.120292
R10974 VSS.n1464 VSS.n1463 0.120292
R10975 VSS.n1463 VSS.n1137 0.120292
R10976 VSS.n1456 VSS.n1137 0.120292
R10977 VSS.n1456 VSS.n1455 0.120292
R10978 VSS.n1455 VSS.n1454 0.120292
R10979 VSS.n1454 VSS.n1141 0.120292
R10980 VSS.n1449 VSS.n1141 0.120292
R10981 VSS.n1449 VSS.n1448 0.120292
R10982 VSS.n1448 VSS.n1447 0.120292
R10983 VSS.n1447 VSS.n1143 0.120292
R10984 VSS.n1400 VSS.n1143 0.120292
R10985 VSS.n1401 VSS.n1400 0.120292
R10986 VSS.n1401 VSS.n1396 0.120292
R10987 VSS.n1406 VSS.n1396 0.120292
R10988 VSS.n1407 VSS.n1406 0.120292
R10989 VSS.n1407 VSS.n1393 0.120292
R10990 VSS.n1411 VSS.n1393 0.120292
R10991 VSS.n1412 VSS.n1411 0.120292
R10992 VSS.n1412 VSS.n1390 0.120292
R10993 VSS.n1416 VSS.n1390 0.120292
R10994 VSS.n1417 VSS.n1416 0.120292
R10995 VSS.n1418 VSS.n1417 0.120292
R10996 VSS.n1418 VSS.n1388 0.120292
R10997 VSS.n1388 VSS.n1386 0.120292
R10998 VSS.n1386 VSS.n1385 0.120292
R10999 VSS.n1424 VSS.n1385 0.120292
R11000 VSS.n1425 VSS.n1424 0.120292
R11001 VSS.n1426 VSS.n1425 0.120292
R11002 VSS.n1426 VSS.n1381 0.120292
R11003 VSS.n1431 VSS.n1381 0.120292
R11004 VSS.n1432 VSS.n1431 0.120292
R11005 VSS.n1433 VSS.n1432 0.120292
R11006 VSS.n1433 VSS.n1377 0.120292
R11007 VSS.n1439 VSS.n1377 0.120292
R11008 VSS.n1440 VSS.n1439 0.120292
R11009 VSS.n1441 VSS.n1440 0.120292
R11010 VSS.n1441 VSS.n1374 0.120292
R11011 VSS.n1374 VSS.n1373 0.120292
R11012 VSS.n1373 VSS.n1372 0.120292
R11013 VSS.n1372 VSS.n1146 0.120292
R11014 VSS.n1368 VSS.n1146 0.120292
R11015 VSS.n1368 VSS.n1367 0.120292
R11016 VSS.n1367 VSS.n1366 0.120292
R11017 VSS.n1366 VSS.n1149 0.120292
R11018 VSS.n1362 VSS.n1149 0.120292
R11019 VSS.n1362 VSS.n1361 0.120292
R11020 VSS.n1361 VSS.n1360 0.120292
R11021 VSS.n1360 VSS.n1151 0.120292
R11022 VSS.n1355 VSS.n1151 0.120292
R11023 VSS.n1355 VSS.n1354 0.120292
R11024 VSS.n1354 VSS.n1353 0.120292
R11025 VSS.n1353 VSS.n1157 0.120292
R11026 VSS.n1348 VSS.n1157 0.120292
R11027 VSS.n1348 VSS.n1347 0.120292
R11028 VSS.n1347 VSS.n1159 0.120292
R11029 VSS.n1343 VSS.n1159 0.120292
R11030 VSS.n1343 VSS.n1342 0.120292
R11031 VSS.n1342 VSS.n1341 0.120292
R11032 VSS.n1341 VSS.n1165 0.120292
R11033 VSS.n1337 VSS.n1165 0.120292
R11034 VSS.n1337 VSS.n1336 0.120292
R11035 VSS.n1336 VSS.n1168 0.120292
R11036 VSS.n1332 VSS.n1168 0.120292
R11037 VSS.n1332 VSS.n1331 0.120292
R11038 VSS.n1331 VSS.n1330 0.120292
R11039 VSS.n1330 VSS.n1172 0.120292
R11040 VSS.n1204 VSS.n1172 0.120292
R11041 VSS.n1204 VSS.n1203 0.120292
R11042 VSS.n1209 VSS.n1203 0.120292
R11043 VSS.n1210 VSS.n1209 0.120292
R11044 VSS.n1211 VSS.n1210 0.120292
R11045 VSS.n1211 VSS.n1201 0.120292
R11046 VSS.n1201 VSS.n1200 0.120292
R11047 VSS.n1216 VSS.n1200 0.120292
R11048 VSS.n1217 VSS.n1216 0.120292
R11049 VSS.n1217 VSS.n1197 0.120292
R11050 VSS.n1222 VSS.n1197 0.120292
R11051 VSS.n1240 VSS.n1187 0.120292
R11052 VSS.n1244 VSS.n1187 0.120292
R11053 VSS.n1245 VSS.n1244 0.120292
R11054 VSS.n1246 VSS.n1245 0.120292
R11055 VSS.n1246 VSS.n1183 0.120292
R11056 VSS.n1183 VSS.n1181 0.120292
R11057 VSS.n1251 VSS.n1181 0.120292
R11058 VSS.n1252 VSS.n1251 0.120292
R11059 VSS.n1253 VSS.n1252 0.120292
R11060 VSS.n1253 VSS.n1178 0.120292
R11061 VSS.n1257 VSS.n1178 0.120292
R11062 VSS.n1325 VSS.n1257 0.120292
R11063 VSS.n1325 VSS.n1324 0.120292
R11064 VSS.n1324 VSS.n1323 0.120292
R11065 VSS.n1323 VSS.n1258 0.120292
R11066 VSS.n1317 VSS.n1258 0.120292
R11067 VSS.n1317 VSS.n1316 0.120292
R11068 VSS.n1316 VSS.n1315 0.120292
R11069 VSS.n1310 VSS.n1309 0.120292
R11070 VSS.n1309 VSS.n1264 0.120292
R11071 VSS.n1304 VSS.n1264 0.120292
R11072 VSS.n1304 VSS.n1303 0.120292
R11073 VSS.n1303 VSS.n1266 0.120292
R11074 VSS.n1271 VSS.n1266 0.120292
R11075 VSS.n1294 VSS.n1271 0.120292
R11076 VSS.n1294 VSS.n1293 0.120292
R11077 VSS.n1293 VSS.n1292 0.120292
R11078 VSS.n1292 VSS.n1272 0.120292
R11079 VSS.n1275 VSS.n1272 0.120292
R11080 VSS.n1287 VSS.n1275 0.120292
R11081 VSS.n1287 VSS.n1286 0.120292
R11082 VSS.n1286 VSS.n1285 0.120292
R11083 VSS.n4007 VSS.n4006 0.120292
R11084 VSS.n4008 VSS.n4007 0.120292
R11085 VSS.n1828 VSS.n1822 0.120292
R11086 VSS.n1829 VSS.n1828 0.120292
R11087 VSS.n1829 VSS.n1819 0.120292
R11088 VSS.n1833 VSS.n1819 0.120292
R11089 VSS.n1834 VSS.n1833 0.120292
R11090 VSS.n1834 VSS.n1817 0.120292
R11091 VSS.n1841 VSS.n1817 0.120292
R11092 VSS.n1842 VSS.n1841 0.120292
R11093 VSS.n1843 VSS.n1842 0.120292
R11094 VSS.n1843 VSS.n1814 0.120292
R11095 VSS.n1877 VSS.n1815 0.120292
R11096 VSS.n1873 VSS.n1815 0.120292
R11097 VSS.n1873 VSS.n1872 0.120292
R11098 VSS.n1872 VSS.n1847 0.120292
R11099 VSS.n1864 VSS.n1847 0.120292
R11100 VSS.n1864 VSS.n1863 0.120292
R11101 VSS.n1863 VSS.n1862 0.120292
R11102 VSS.n1862 VSS.n1852 0.120292
R11103 VSS.n1858 VSS.n1852 0.120292
R11104 VSS.n1902 VSS.n1894 0.120292
R11105 VSS.n1903 VSS.n1902 0.120292
R11106 VSS.n1903 VSS.n1890 0.120292
R11107 VSS.n1908 VSS.n1890 0.120292
R11108 VSS.n1909 VSS.n1908 0.120292
R11109 VSS.n1910 VSS.n1909 0.120292
R11110 VSS.n1910 VSS.n1886 0.120292
R11111 VSS.n1915 VSS.n1886 0.120292
R11112 VSS.n1916 VSS.n1915 0.120292
R11113 VSS.n1916 VSS.n1881 0.120292
R11114 VSS.n4763 VSS.n1882 0.120292
R11115 VSS.n4759 VSS.n1882 0.120292
R11116 VSS.n4759 VSS.n4758 0.120292
R11117 VSS.n4758 VSS.n4757 0.120292
R11118 VSS.n4757 VSS.n4737 0.120292
R11119 VSS.n4751 VSS.n4737 0.120292
R11120 VSS.n4751 VSS.n4750 0.120292
R11121 VSS.n4750 VSS.n4749 0.120292
R11122 VSS.n4749 VSS.n4739 0.120292
R11123 VSS.n4065 VSS.n4059 0.120292
R11124 VSS.n4066 VSS.n4065 0.120292
R11125 VSS.n4066 VSS.n4056 0.120292
R11126 VSS.n4071 VSS.n4056 0.120292
R11127 VSS.n4072 VSS.n4071 0.120292
R11128 VSS.n4073 VSS.n4072 0.120292
R11129 VSS.n4073 VSS.n4053 0.120292
R11130 VSS.n4080 VSS.n4053 0.120292
R11131 VSS.n4081 VSS.n4080 0.120292
R11132 VSS.n4082 VSS.n4081 0.120292
R11133 VSS.n4085 VSS.n4084 0.120292
R11134 VSS.n4106 VSS.n4085 0.120292
R11135 VSS.n4106 VSS.n4105 0.120292
R11136 VSS.n4105 VSS.n4104 0.120292
R11137 VSS.n4104 VSS.n4088 0.120292
R11138 VSS.n4100 VSS.n4088 0.120292
R11139 VSS.n4100 VSS.n4099 0.120292
R11140 VSS.n4099 VSS.n4098 0.120292
R11141 VSS.n4098 VSS.n4091 0.120292
R11142 VSS.n1794 VSS.n1786 0.120292
R11143 VSS.n1799 VSS.n1786 0.120292
R11144 VSS.n1800 VSS.n1799 0.120292
R11145 VSS.n1801 VSS.n1800 0.120292
R11146 VSS.n1801 VSS.n1784 0.120292
R11147 VSS.n1806 VSS.n1784 0.120292
R11148 VSS.n1807 VSS.n1806 0.120292
R11149 VSS.n1807 VSS.n1778 0.120292
R11150 VSS.n1812 VSS.n1778 0.120292
R11151 VSS.n1813 VSS.n1812 0.120292
R11152 VSS.n4796 VSS.n4795 0.120292
R11153 VSS.n4795 VSS.n4794 0.120292
R11154 VSS.n4794 VSS.n4768 0.120292
R11155 VSS.n4788 VSS.n4768 0.120292
R11156 VSS.n4788 VSS.n4787 0.120292
R11157 VSS.n4787 VSS.n4786 0.120292
R11158 VSS.n4786 VSS.n4772 0.120292
R11159 VSS.n4782 VSS.n4772 0.120292
R11160 VSS.n4782 VSS.n4781 0.120292
R11161 VSS.n4905 VSS.n4904 0.120292
R11162 VSS.n3800 VSS.n3794 0.120292
R11163 VSS.n3801 VSS.n3800 0.120292
R11164 VSS.n3802 VSS.n3801 0.120292
R11165 VSS.n3802 VSS.n3792 0.120292
R11166 VSS.n3792 VSS.n3789 0.120292
R11167 VSS.n3807 VSS.n3789 0.120292
R11168 VSS.n3808 VSS.n3807 0.120292
R11169 VSS.n3809 VSS.n3808 0.120292
R11170 VSS.n3809 VSS.n3787 0.120292
R11171 VSS.n3787 VSS.n3786 0.120292
R11172 VSS.n3786 VSS.n3785 0.120292
R11173 VSS.n3785 VSS.n3730 0.120292
R11174 VSS.n3781 VSS.n3730 0.120292
R11175 VSS.n3781 VSS.n3780 0.120292
R11176 VSS.n3780 VSS.n3779 0.120292
R11177 VSS.n3779 VSS.n3732 0.120292
R11178 VSS.n3775 VSS.n3732 0.120292
R11179 VSS.n3775 VSS.n3774 0.120292
R11180 VSS.n3774 VSS.n3773 0.120292
R11181 VSS.n3773 VSS.n3736 0.120292
R11182 VSS.n3767 VSS.n3736 0.120292
R11183 VSS.n3767 VSS.n3766 0.120292
R11184 VSS.n3766 VSS.n3765 0.120292
R11185 VSS.n3765 VSS.n3738 0.120292
R11186 VSS.n3761 VSS.n3738 0.120292
R11187 VSS.n3761 VSS.n3760 0.120292
R11188 VSS.n3760 VSS.n3759 0.120292
R11189 VSS.n3759 VSS.n3740 0.120292
R11190 VSS.n3754 VSS.n3740 0.120292
R11191 VSS.n3754 VSS.n3753 0.120292
R11192 VSS.n3753 VSS.n3752 0.120292
R11193 VSS.n3752 VSS.n3742 0.120292
R11194 VSS.n3748 VSS.n3742 0.120292
R11195 VSS.n3748 VSS.n3747 0.120292
R11196 VSS.n3747 VSS.n3746 0.120292
R11197 VSS.n3746 VSS.n3710 0.120292
R11198 VSS.n4304 VSS.n3710 0.120292
R11199 VSS.n4305 VSS.n4304 0.120292
R11200 VSS.n4306 VSS.n4305 0.120292
R11201 VSS.n4306 VSS.n3708 0.120292
R11202 VSS.n3708 VSS.n3706 0.120292
R11203 VSS.n4311 VSS.n3706 0.120292
R11204 VSS.n4312 VSS.n4311 0.120292
R11205 VSS.n4313 VSS.n4312 0.120292
R11206 VSS.n4313 VSS.n3703 0.120292
R11207 VSS.n3703 VSS.n3701 0.120292
R11208 VSS.n4318 VSS.n3701 0.120292
R11209 VSS.n4319 VSS.n4318 0.120292
R11210 VSS.n4320 VSS.n4319 0.120292
R11211 VSS.n4320 VSS.n3699 0.120292
R11212 VSS.n4324 VSS.n3699 0.120292
R11213 VSS.n4325 VSS.n4324 0.120292
R11214 VSS.n4326 VSS.n4325 0.120292
R11215 VSS.n4326 VSS.n3697 0.120292
R11216 VSS.n4330 VSS.n3697 0.120292
R11217 VSS.n4331 VSS.n4330 0.120292
R11218 VSS.n4332 VSS.n4331 0.120292
R11219 VSS.n4332 VSS.n3695 0.120292
R11220 VSS.n3695 VSS.n3693 0.120292
R11221 VSS.n4337 VSS.n3693 0.120292
R11222 VSS.n4338 VSS.n4337 0.120292
R11223 VSS.n4339 VSS.n4338 0.120292
R11224 VSS.n4339 VSS.n3690 0.120292
R11225 VSS.n4343 VSS.n3690 0.120292
R11226 VSS.n4344 VSS.n4343 0.120292
R11227 VSS.n4345 VSS.n4344 0.120292
R11228 VSS.n4345 VSS.n3687 0.120292
R11229 VSS.n4349 VSS.n3687 0.120292
R11230 VSS.n4350 VSS.n4349 0.120292
R11231 VSS.n4351 VSS.n4350 0.120292
R11232 VSS.n4351 VSS.n3684 0.120292
R11233 VSS.n4355 VSS.n3684 0.120292
R11234 VSS.n4356 VSS.n4355 0.120292
R11235 VSS.n4357 VSS.n4356 0.120292
R11236 VSS.n4357 VSS.n3682 0.120292
R11237 VSS.n4361 VSS.n3682 0.120292
R11238 VSS.n4362 VSS.n4361 0.120292
R11239 VSS.n4363 VSS.n4362 0.120292
R11240 VSS.n4363 VSS.n3679 0.120292
R11241 VSS.n4368 VSS.n3679 0.120292
R11242 VSS.n4369 VSS.n4368 0.120292
R11243 VSS.n4370 VSS.n4369 0.120292
R11244 VSS.n4370 VSS.n3677 0.120292
R11245 VSS.n4374 VSS.n3677 0.120292
R11246 VSS.n4375 VSS.n4374 0.120292
R11247 VSS.n4375 VSS.n3674 0.120292
R11248 VSS.n4380 VSS.n3674 0.120292
R11249 VSS.n4381 VSS.n4380 0.120292
R11250 VSS.n4382 VSS.n4381 0.120292
R11251 VSS.n4382 VSS.n3671 0.120292
R11252 VSS.n4387 VSS.n3671 0.120292
R11253 VSS.n4388 VSS.n4387 0.120292
R11254 VSS.n4388 VSS.n3669 0.120292
R11255 VSS.n3669 VSS.n3666 0.120292
R11256 VSS.n4393 VSS.n3666 0.120292
R11257 VSS.n4394 VSS.n4393 0.120292
R11258 VSS.n4395 VSS.n4394 0.120292
R11259 VSS.n4395 VSS.n3663 0.120292
R11260 VSS.n4399 VSS.n3663 0.120292
R11261 VSS.n4400 VSS.n4399 0.120292
R11262 VSS.n4401 VSS.n4400 0.120292
R11263 VSS.n4401 VSS.n3661 0.120292
R11264 VSS.n3661 VSS.n3659 0.120292
R11265 VSS.n4406 VSS.n3659 0.120292
R11266 VSS.n4407 VSS.n4406 0.120292
R11267 VSS.n4408 VSS.n4407 0.120292
R11268 VSS.n4408 VSS.n3657 0.120292
R11269 VSS.n3657 VSS.n3656 0.120292
R11270 VSS.n4413 VSS.n3656 0.120292
R11271 VSS.n4414 VSS.n4413 0.120292
R11272 VSS.n4414 VSS.n3652 0.120292
R11273 VSS.n4419 VSS.n3652 0.120292
R11274 VSS.n4420 VSS.n4419 0.120292
R11275 VSS.n4421 VSS.n4420 0.120292
R11276 VSS.n4421 VSS.n3650 0.120292
R11277 VSS.n4425 VSS.n3650 0.120292
R11278 VSS.n4426 VSS.n4425 0.120292
R11279 VSS.n4427 VSS.n4426 0.120292
R11280 VSS.n4427 VSS.n3647 0.120292
R11281 VSS.n4431 VSS.n3647 0.120292
R11282 VSS.n4432 VSS.n4431 0.120292
R11283 VSS.n4433 VSS.n4432 0.120292
R11284 VSS.n4433 VSS.n3644 0.120292
R11285 VSS.n4437 VSS.n3644 0.120292
R11286 VSS.n4438 VSS.n4437 0.120292
R11287 VSS.n4439 VSS.n4438 0.120292
R11288 VSS.n4439 VSS.n3642 0.120292
R11289 VSS.n4443 VSS.n3642 0.120292
R11290 VSS.n4444 VSS.n4443 0.120292
R11291 VSS.n4445 VSS.n4444 0.120292
R11292 VSS.n4445 VSS.n3639 0.120292
R11293 VSS.n4449 VSS.n3639 0.120292
R11294 VSS.n4450 VSS.n4449 0.120292
R11295 VSS.n4451 VSS.n4450 0.120292
R11296 VSS.n4451 VSS.n3637 0.120292
R11297 VSS.n4455 VSS.n3637 0.120292
R11298 VSS.n4456 VSS.n4455 0.120292
R11299 VSS.n4457 VSS.n4456 0.120292
R11300 VSS.n4457 VSS.n3634 0.120292
R11301 VSS.n4461 VSS.n3634 0.120292
R11302 VSS.n4462 VSS.n4461 0.120292
R11303 VSS.n4463 VSS.n4462 0.120292
R11304 VSS.n4463 VSS.n3632 0.120292
R11305 VSS.n3632 VSS.n3630 0.120292
R11306 VSS.n4468 VSS.n3630 0.120292
R11307 VSS.n4469 VSS.n4468 0.120292
R11308 VSS.n4470 VSS.n4469 0.120292
R11309 VSS.n4470 VSS.n3627 0.120292
R11310 VSS.n4474 VSS.n3627 0.120292
R11311 VSS.n4475 VSS.n4474 0.120292
R11312 VSS.n4476 VSS.n4475 0.120292
R11313 VSS.n4476 VSS.n3624 0.120292
R11314 VSS.n4483 VSS.n3624 0.120292
R11315 VSS.n4484 VSS.n4483 0.120292
R11316 VSS.n4485 VSS.n4484 0.120292
R11317 VSS.n4485 VSS.n3622 0.120292
R11318 VSS.n3622 VSS.n3620 0.120292
R11319 VSS.n4490 VSS.n3620 0.120292
R11320 VSS.n4491 VSS.n4490 0.120292
R11321 VSS.n4492 VSS.n4491 0.120292
R11322 VSS.n4492 VSS.n3617 0.120292
R11323 VSS.n4496 VSS.n3617 0.120292
R11324 VSS.n4497 VSS.n4496 0.120292
R11325 VSS.n4498 VSS.n4497 0.120292
R11326 VSS.n4498 VSS.n3615 0.120292
R11327 VSS.n3615 VSS.n3613 0.120292
R11328 VSS.n4503 VSS.n3613 0.120292
R11329 VSS.n4504 VSS.n4503 0.120292
R11330 VSS.n4505 VSS.n4504 0.120292
R11331 VSS.n4505 VSS.n3611 0.120292
R11332 VSS.n4511 VSS.n3611 0.120292
R11333 VSS.n4512 VSS.n4511 0.120292
R11334 VSS.n4512 VSS.n3609 0.120292
R11335 VSS.n4516 VSS.n3609 0.120292
R11336 VSS.n4517 VSS.n4516 0.120292
R11337 VSS.n4518 VSS.n4517 0.120292
R11338 VSS.n4518 VSS.n3606 0.120292
R11339 VSS.n3606 VSS.n3604 0.120292
R11340 VSS.n4523 VSS.n3604 0.120292
R11341 VSS.n4524 VSS.n4523 0.120292
R11342 VSS.n4525 VSS.n4524 0.120292
R11343 VSS.n4525 VSS.n3602 0.120292
R11344 VSS.n3602 VSS.n3601 0.120292
R11345 VSS.n4530 VSS.n3601 0.120292
R11346 VSS.n4531 VSS.n4530 0.120292
R11347 VSS.n4532 VSS.n4531 0.120292
R11348 VSS.n4532 VSS.n3598 0.120292
R11349 VSS.n4536 VSS.n3598 0.120292
R11350 VSS.n4537 VSS.n4536 0.120292
R11351 VSS.n4538 VSS.n4537 0.120292
R11352 VSS.n4538 VSS.n3595 0.120292
R11353 VSS.n4542 VSS.n3595 0.120292
R11354 VSS.n4543 VSS.n4542 0.120292
R11355 VSS.n4544 VSS.n4543 0.120292
R11356 VSS.n4544 VSS.n3592 0.120292
R11357 VSS.n4549 VSS.n3592 0.120292
R11358 VSS.n4550 VSS.n4549 0.120292
R11359 VSS.n4550 VSS.n3589 0.120292
R11360 VSS.n4554 VSS.n3589 0.120292
R11361 VSS.n4555 VSS.n4554 0.120292
R11362 VSS.n4556 VSS.n4555 0.120292
R11363 VSS.n4556 VSS.n3587 0.120292
R11364 VSS.n4560 VSS.n3587 0.120292
R11365 VSS.n4561 VSS.n4560 0.120292
R11366 VSS.n4562 VSS.n4561 0.120292
R11367 VSS.n4562 VSS.n3584 0.120292
R11368 VSS.n4566 VSS.n3584 0.120292
R11369 VSS.n4567 VSS.n4566 0.120292
R11370 VSS.n4568 VSS.n4567 0.120292
R11371 VSS.n4568 VSS.n3581 0.120292
R11372 VSS.n4572 VSS.n3581 0.120292
R11373 VSS.n4573 VSS.n4572 0.120292
R11374 VSS.n4574 VSS.n4573 0.120292
R11375 VSS.n4574 VSS.n3579 0.120292
R11376 VSS.n4580 VSS.n3579 0.120292
R11377 VSS.n4581 VSS.n4580 0.120292
R11378 VSS.n4582 VSS.n4581 0.120292
R11379 VSS.n4582 VSS.n3577 0.120292
R11380 VSS.n4588 VSS.n3577 0.120292
R11381 VSS.n4589 VSS.n4588 0.120292
R11382 VSS.n4590 VSS.n4589 0.120292
R11383 VSS.n4590 VSS.n3575 0.120292
R11384 VSS.n4595 VSS.n3575 0.120292
R11385 VSS.n4596 VSS.n4595 0.120292
R11386 VSS.n4597 VSS.n4596 0.120292
R11387 VSS.n4597 VSS.n3573 0.120292
R11388 VSS.n4601 VSS.n3573 0.120292
R11389 VSS.n4602 VSS.n4601 0.120292
R11390 VSS.n4603 VSS.n4602 0.120292
R11391 VSS.n4603 VSS.n3570 0.120292
R11392 VSS.n4608 VSS.n3570 0.120292
R11393 VSS.n4609 VSS.n4608 0.120292
R11394 VSS.n4610 VSS.n4609 0.120292
R11395 VSS.n4610 VSS.n3567 0.120292
R11396 VSS.n4614 VSS.n3567 0.120292
R11397 VSS.n4615 VSS.n4614 0.120292
R11398 VSS.n4616 VSS.n4615 0.120292
R11399 VSS.n4616 VSS.n3564 0.120292
R11400 VSS.n4620 VSS.n3564 0.120292
R11401 VSS.n4621 VSS.n4620 0.120292
R11402 VSS.n4622 VSS.n4621 0.120292
R11403 VSS.n4622 VSS.n3561 0.120292
R11404 VSS.n4627 VSS.n3561 0.120292
R11405 VSS.n4628 VSS.n4627 0.120292
R11406 VSS.n4629 VSS.n4628 0.120292
R11407 VSS.n4646 VSS.n1925 0.120292
R11408 VSS.n4651 VSS.n1925 0.120292
R11409 VSS.n4652 VSS.n4651 0.120292
R11410 VSS.n4653 VSS.n4652 0.120292
R11411 VSS.n4653 VSS.n1923 0.120292
R11412 VSS.n4657 VSS.n1923 0.120292
R11413 VSS.n4658 VSS.n4657 0.120292
R11414 VSS.n4659 VSS.n4658 0.120292
R11415 VSS.n4659 VSS.n1921 0.120292
R11416 VSS.n4664 VSS.n1921 0.120292
R11417 VSS.n4665 VSS.n4664 0.120292
R11418 VSS.n4666 VSS.n4665 0.120292
R11419 VSS.n4667 VSS.n4666 0.120292
R11420 VSS.n4727 VSS.n4667 0.120292
R11421 VSS.n4727 VSS.n4726 0.120292
R11422 VSS.n4726 VSS.n4725 0.120292
R11423 VSS.n4725 VSS.n4670 0.120292
R11424 VSS.n4721 VSS.n4670 0.120292
R11425 VSS.n4721 VSS.n4720 0.120292
R11426 VSS.n4720 VSS.n4719 0.120292
R11427 VSS.n4719 VSS.n4673 0.120292
R11428 VSS.n4715 VSS.n4673 0.120292
R11429 VSS.n4715 VSS.n4714 0.120292
R11430 VSS.n4714 VSS.n4713 0.120292
R11431 VSS.n4713 VSS.n4676 0.120292
R11432 VSS.n4709 VSS.n4676 0.120292
R11433 VSS.n4709 VSS.n4708 0.120292
R11434 VSS.n4708 VSS.n4707 0.120292
R11435 VSS.n4707 VSS.n4679 0.120292
R11436 VSS.n4703 VSS.n4679 0.120292
R11437 VSS.n4703 VSS.n4702 0.120292
R11438 VSS.n4702 VSS.n4701 0.120292
R11439 VSS.n4701 VSS.n4682 0.120292
R11440 VSS.n4697 VSS.n4682 0.120292
R11441 VSS.n4697 VSS.n4696 0.120292
R11442 VSS.n4696 VSS.n4695 0.120292
R11443 VSS.n4695 VSS.n4685 0.120292
R11444 VSS.n4691 VSS.n4685 0.120292
R11445 VSS.n4691 VSS.n4690 0.120292
R11446 VSS.n4129 VSS.n4114 0.120292
R11447 VSS.n4123 VSS.n4114 0.120292
R11448 VSS.n4123 VSS.n4122 0.120292
R11449 VSS.n4166 VSS.n3935 0.120292
R11450 VSS.n4162 VSS.n3935 0.120292
R11451 VSS.n4830 VSS.n4829 0.119329
R11452 VSS.n4153 VSS.n4152 0.119329
R11453 VSS.n2198 VSS.n2139 0.112781
R11454 VSS.n4008 VSS.n3998 0.108833
R11455 VSS.n4820 VSS.n1772 0.104667
R11456 VSS.n4822 VSS.n1772 0.104667
R11457 VSS.n3858 VSS.n3857 0.104667
R11458 VSS.n3857 VSS.n3823 0.104667
R11459 VSS VSS.n5489 0.101274
R11460 VSS.n3940 VSS.n1771 0.101002
R11461 VSS.n3998 VSS.n3939 0.0963333
R11462 VSS.n5342 VSS.n5341 0.0950946
R11463 VSS.n5347 VSS.n5346 0.0950946
R11464 VSS.n5487 VSS.n5486 0.0950946
R11465 VSS.n5480 VSS.n7 0.0950946
R11466 VSS.n2740 VSS.n2739 0.0950946
R11467 VSS.n2733 VSS.n1936 0.0950946
R11468 VSS.n3538 VSS.n3537 0.0950946
R11469 VSS.n3551 VSS.n2746 0.0950946
R11470 VSS.n1225 VSS.n1223 0.0950946
R11471 VSS.n1238 VSS.n1191 0.0950946
R11472 VSS.n4640 VSS.n4639 0.0950946
R11473 VSS.n4644 VSS.n1928 0.0950946
R11474 VSS.n1878 VSS.n1877 0.09425
R11475 VSS.n4764 VSS.n4763 0.09425
R11476 VSS.n4084 VSS.n1880 0.09425
R11477 VSS.n4796 VSS.n4767 0.09425
R11478 VSS.n104 VSS.n97 0.0916458
R11479 VSS.n5475 VSS.n8 0.0916458
R11480 VSS.n2728 VSS.n1937 0.0916458
R11481 VSS.n3550 VSS.n3549 0.0916458
R11482 VSS.n1240 VSS.n1239 0.0916458
R11483 VSS.n4646 VSS.n4645 0.0916458
R11484 VSS.n3246 VSS.n3242 0.0900105
R11485 VSS.n3982 VSS.n3981 0.0882358
R11486 VSS.n3987 VSS.n3986 0.0882358
R11487 VSS.n3820 VSS.n3818 0.0882358
R11488 VSS.n3867 VSS.n3866 0.0882358
R11489 VSS.n4805 VSS.n4802 0.0840129
R11490 VSS.n3855 VSS.n3825 0.0840129
R11491 VSS.n5340 VSS.n102 0.0838333
R11492 VSS.n5485 VSS.n5484 0.0838333
R11493 VSS.n2738 VSS.n2737 0.0838333
R11494 VSS.n3543 VSS.n2752 0.0838333
R11495 VSS.n1233 VSS.n1194 0.0838333
R11496 VSS.n4638 VSS.n4637 0.0838333
R11497 VSS.n1766 VSS.n1765 0.0812292
R11498 VSS.n4118 VSS.n3941 0.0812292
R11499 VSS.n4810 VSS.n1775 0.0744504
R11500 VSS.n3845 VSS.n3841 0.0744504
R11501 VSS.n305 VSS.n304 0.0700652
R11502 VSS.n3448 VSS.n3447 0.0700652
R11503 VSS.n979 VSS.n978 0.0700652
R11504 VSS.n317 VSS.n316 0.0685851
R11505 VSS.n5464 VSS.n17 0.0685851
R11506 VSS.n1583 VSS.n1582 0.0685851
R11507 VSS.n5338 VSS.n5337 0.0680676
R11508 VSS.n5337 VSS.n103 0.0680676
R11509 VSS.n5483 VSS.n4 0.0680676
R11510 VSS.n5483 VSS.n5482 0.0680676
R11511 VSS.n2736 VSS.n1933 0.0680676
R11512 VSS.n2736 VSS.n2735 0.0680676
R11513 VSS.n3542 VSS.n3540 0.0680676
R11514 VSS.n3542 VSS.n3541 0.0680676
R11515 VSS.n1234 VSS.n1193 0.0680676
R11516 VSS.n1235 VSS.n1234 0.0680676
R11517 VSS.n4636 VSS.n3557 0.0680676
R11518 VSS.n4636 VSS.n4635 0.0680676
R11519 VSS.n3726 VSS.n3725 0.0677515
R11520 VSS.n3725 VSS.n3724 0.0677515
R11521 VSS.n3724 VSS.n3720 0.0677515
R11522 VSS.n5339 VSS.n5336 0.0656042
R11523 VSS.n5349 VSS.n5348 0.0656042
R11524 VSS.n5 VSS.n3 0.0656042
R11525 VSS.n5479 VSS.n6 0.0656042
R11526 VSS.n1934 VSS.n1932 0.0656042
R11527 VSS.n2732 VSS.n1935 0.0656042
R11528 VSS.n3536 VSS.n3535 0.0656042
R11529 VSS.n3545 VSS.n3544 0.0656042
R11530 VSS.n1227 VSS.n1226 0.0656042
R11531 VSS.n1232 VSS.n1195 0.0656042
R11532 VSS.n3558 VSS.n3556 0.0656042
R11533 VSS.n4634 VSS.n3559 0.0656042
R11534 VSS.n4294 VSS.n4293 0.0620894
R11535 VSS.n5343 VSS.n107 0.0574697
R11536 VSS.n5345 VSS.n105 0.0574697
R11537 VSS.n5481 VSS.n2 0.0574697
R11538 VSS.n2734 VSS.n1931 0.0574697
R11539 VSS.n3539 VSS.n2743 0.0574697
R11540 VSS.n3552 VSS.n2745 0.0574697
R11541 VSS.n1236 VSS.n1192 0.0574697
R11542 VSS.n3555 VSS.n1929 0.0574697
R11543 VSS.n5336 VSS.n5335 0.0551875
R11544 VSS.n5348 VSS.n99 0.0551875
R11545 VSS.n559 VSS.n3 0.0551875
R11546 VSS.n5479 VSS.n5478 0.0551875
R11547 VSS.n2612 VSS.n1932 0.0551875
R11548 VSS.n2732 VSS.n2731 0.0551875
R11549 VSS.n3536 VSS.n3534 0.0551875
R11550 VSS.n3544 VSS.n2747 0.0551875
R11551 VSS.n1226 VSS.n1222 0.0551875
R11552 VSS.n1195 VSS.n1190 0.0551875
R11553 VSS.n4629 VSS.n3556 0.0551875
R11554 VSS.n3559 VSS.n1927 0.0551875
R11555 VSS.n4844 VSS.n4834 0.0550024
R11556 VSS.n4139 VSS.n4138 0.0550024
R11557 VSS.n4804 VSS.n1773 0.052157
R11558 VSS.n3856 VSS.n3824 0.052157
R11559 VSS.n4826 VSS.n4825 0.046482
R11560 VSS.n940 VSS.n939 0.0443356
R11561 VSS.n4826 VSS.n1769 0.0437119
R11562 VSS.n5341 VSS.n5338 0.0410405
R11563 VSS.n5347 VSS.n103 0.0410405
R11564 VSS.n5486 VSS.n4 0.0410405
R11565 VSS.n5482 VSS.n5480 0.0410405
R11566 VSS.n2739 VSS.n1933 0.0410405
R11567 VSS.n2735 VSS.n2733 0.0410405
R11568 VSS.n3540 VSS.n3538 0.0410405
R11569 VSS.n3541 VSS.n2746 0.0410405
R11570 VSS.n1223 VSS.n1193 0.0410405
R11571 VSS.n1235 VSS.n1191 0.0410405
R11572 VSS.n4639 VSS.n3557 0.0410405
R11573 VSS.n4635 VSS.n1928 0.0410405
R11574 VSS.n1766 VSS.n1727 0.0395625
R11575 VSS.n4122 VSS.n3941 0.0395625
R11576 VSS.n106 VSS.n105 0.0292489
R11577 VSS.n107 VSS.n106 0.0292489
R11578 VSS.n2745 VSS.n2744 0.0292489
R11579 VSS.n4641 VSS.n3555 0.0292489
R11580 VSS.n4643 VSS.n1929 0.0292489
R11581 VSS.n3539 VSS.n2744 0.0292489
R11582 VSS.n2741 VSS.n1931 0.0292489
R11583 VSS.n2734 VSS.n1930 0.0292489
R11584 VSS.n1224 VSS.n1192 0.0292489
R11585 VSS.n1237 VSS.n1236 0.0292489
R11586 VSS.n5488 VSS.n2 0.0292489
R11587 VSS.n5481 VSS.n0 0.0292489
R11588 VSS.n104 VSS.n99 0.0291458
R11589 VSS.n5478 VSS.n8 0.0291458
R11590 VSS.n2731 VSS.n1937 0.0291458
R11591 VSS.n3550 VSS.n2747 0.0291458
R11592 VSS.n1239 VSS.n1190 0.0291458
R11593 VSS.n4645 VSS.n1927 0.0291458
R11594 VSS.n1878 VSS.n1814 0.0265417
R11595 VSS.n4764 VSS.n1881 0.0265417
R11596 VSS.n4082 VSS.n1880 0.0265417
R11597 VSS.n4767 VSS.n1813 0.0265417
R11598 VSS.n5490 VSS 0.025175
R11599 VSS VSS.n5490 0.0237235
R11600 VSS.n4158 VSS.n4157 0.0200312
R11601 VSS.n3720 VSS.n1767 0.0187749
R11602 VSS.n5340 VSS.n5339 0.0187292
R11603 VSS.n5349 VSS.n102 0.0187292
R11604 VSS.n5485 VSS.n5 0.0187292
R11605 VSS.n5484 VSS.n6 0.0187292
R11606 VSS.n2738 VSS.n1934 0.0187292
R11607 VSS.n2737 VSS.n1935 0.0187292
R11608 VSS.n3535 VSS.n2752 0.0187292
R11609 VSS.n3545 VSS.n3543 0.0187292
R11610 VSS.n1227 VSS.n1194 0.0187292
R11611 VSS.n1233 VSS.n1232 0.0187292
R11612 VSS.n4638 VSS.n3558 0.0187292
R11613 VSS.n4637 VSS.n4634 0.0187292
R11614 VSS.n5490 VSS 0.0146
R11615 VSS.n5344 VSS 0.0144531
R11616 VSS.n5490 VSS 0.0137706
R11617 VSS.n4159 VSS.n4158 0.0122188
R11618 VSS.n4905 VSS.n4900 0.00701042
R11619 VSS.n3886 VSS.n3881 0.00675
R11620 VSS.n4825 VSS.n4824 0.00609092
R11621 VSS.n3860 VSS.n1769 0.00605668
R11622 VDAC_P.n3 VDAC_P.t19 946.489
R11623 VDAC_P.n0 VDAC_P.t16 946.489
R11624 VDAC_P.n7 VDAC_P.t13 946.345
R11625 VDAC_P.n13 VDAC_P.t10 945.764
R11626 VDAC_P.n12 VDAC_P.t8 945.755
R11627 VDAC_P.n11 VDAC_P.t20 945.755
R11628 VDAC_P.n10 VDAC_P.t9 945.755
R11629 VDAC_P.n9 VDAC_P.t18 945.755
R11630 VDAC_P.n8 VDAC_P.t23 945.755
R11631 VDAC_P.n7 VDAC_P.t12 945.755
R11632 VDAC_P.n5 VDAC_P.t14 945.755
R11633 VDAC_P.n4 VDAC_P.t17 945.755
R11634 VDAC_P.n3 VDAC_P.t21 945.755
R11635 VDAC_P.n2 VDAC_P.t15 945.755
R11636 VDAC_P.n1 VDAC_P.t11 945.755
R11637 VDAC_P.n0 VDAC_P.t22 945.755
R11638 VDAC_P.n20 VDAC_P.n18 14.894
R11639 VDAC_P.n17 VDAC_P.n15 14.894
R11640 VDAC_P.n20 VDAC_P.n19 14.394
R11641 VDAC_P.n17 VDAC_P.n16 14.394
R11642 VDAC_P.n22 VDAC_P.n14 13.3642
R11643 VDAC_P.n22 VDAC_P.n21 13.0284
R11644 VDAC_P.n10 VDAC_P.n9 6.67373
R11645 VDAC_P.n6 VDAC_P.n2 6.20847
R11646 VDAC_P.n14 VDAC_P.n6 5.45883
R11647 VDAC_P.n14 VDAC_P.n13 4.5005
R11648 VDAC_P.n19 VDAC_P.t5 2.4755
R11649 VDAC_P.n19 VDAC_P.t2 2.4755
R11650 VDAC_P.n18 VDAC_P.t1 2.4755
R11651 VDAC_P.n18 VDAC_P.t3 2.4755
R11652 VDAC_P.n15 VDAC_P.t7 2.4755
R11653 VDAC_P.n15 VDAC_P.t4 2.4755
R11654 VDAC_P.n16 VDAC_P.t6 2.4755
R11655 VDAC_P.n16 VDAC_P.t0 2.4755
R11656 VDAC_P VDAC_P.n22 1.91687
R11657 VDAC_P.n11 VDAC_P.n10 0.733109
R11658 VDAC_P.n12 VDAC_P.n11 0.733109
R11659 VDAC_P.n4 VDAC_P.n3 0.733109
R11660 VDAC_P.n5 VDAC_P.n4 0.733109
R11661 VDAC_P.n1 VDAC_P.n0 0.733109
R11662 VDAC_P.n2 VDAC_P.n1 0.733109
R11663 VDAC_P.n13 VDAC_P.n12 0.675138
R11664 VDAC_P.n8 VDAC_P.n7 0.589359
R11665 VDAC_P.n9 VDAC_P.n8 0.589359
R11666 VDAC_P.n6 VDAC_P.n5 0.491804
R11667 VDAC_P.n21 VDAC_P.n20 0.21925
R11668 VDAC_P.n21 VDAC_P.n17 0.188
R11669 a_5088_37509.n8 a_5088_37509.t19 120.862
R11670 a_5088_37509.n9 a_5088_37509.t17 120.564
R11671 a_5088_37509.n8 a_5088_37509.n7 104.312
R11672 a_5088_37509.n2 a_5088_37509.n0 40.84
R11673 a_5088_37509.n6 a_5088_37509.n5 40.5431
R11674 a_5088_37509.n4 a_5088_37509.n3 40.5431
R11675 a_5088_37509.n2 a_5088_37509.n1 40.5431
R11676 a_5088_37509.n17 a_5088_37509.n16 40.4813
R11677 a_5088_37509.n12 a_5088_37509.n11 40.1844
R11678 a_5088_37509.n14 a_5088_37509.n13 40.1844
R11679 a_5088_37509.n16 a_5088_37509.n15 40.1844
R11680 a_5088_37509.n10 a_5088_37509.n9 24.9745
R11681 a_5088_37509.n7 a_5088_37509.t18 16.253
R11682 a_5088_37509.n7 a_5088_37509.t16 16.253
R11683 a_5088_37509.n12 a_5088_37509.n10 13.188
R11684 a_5088_37509.n11 a_5088_37509.t7 4.76133
R11685 a_5088_37509.n11 a_5088_37509.t15 4.76133
R11686 a_5088_37509.n13 a_5088_37509.t12 4.76133
R11687 a_5088_37509.n13 a_5088_37509.t3 4.76133
R11688 a_5088_37509.n15 a_5088_37509.t10 4.76133
R11689 a_5088_37509.n15 a_5088_37509.t5 4.76133
R11690 a_5088_37509.n5 a_5088_37509.t6 4.76133
R11691 a_5088_37509.n5 a_5088_37509.t9 4.76133
R11692 a_5088_37509.n3 a_5088_37509.t11 4.76133
R11693 a_5088_37509.n3 a_5088_37509.t13 4.76133
R11694 a_5088_37509.n1 a_5088_37509.t2 4.76133
R11695 a_5088_37509.n1 a_5088_37509.t14 4.76133
R11696 a_5088_37509.n0 a_5088_37509.t4 4.76133
R11697 a_5088_37509.n0 a_5088_37509.t1 4.76133
R11698 a_5088_37509.t0 a_5088_37509.n17 4.76133
R11699 a_5088_37509.n17 a_5088_37509.t8 4.76133
R11700 a_5088_37509.n4 a_5088_37509.n2 0.313
R11701 a_5088_37509.n6 a_5088_37509.n4 0.313
R11702 a_5088_37509.n16 a_5088_37509.n14 0.313
R11703 a_5088_37509.n14 a_5088_37509.n12 0.313
R11704 a_5088_37509.n9 a_5088_37509.n8 0.297375
R11705 a_5088_37509.n10 a_5088_37509.n6 0.297375
R11706 a_8912_37509.n14 a_8912_37509.t14 45.8845
R11707 a_8912_37509.n33 a_8912_37509.t31 45.6616
R11708 a_8912_37509.n19 a_8912_37509.t9 45.6572
R11709 a_8912_37509.n20 a_8912_37509.t27 45.6572
R11710 a_8912_37509.n27 a_8912_37509.t16 45.6572
R11711 a_8912_37509.n38 a_8912_37509.t23 45.4344
R11712 a_8912_37509.n39 a_8912_37509.t4 45.4344
R11713 a_8912_37509.n31 a_8912_37509.t5 45.4344
R11714 a_8912_37509.n14 a_8912_37509.n13 40.8964
R11715 a_8912_37509.n16 a_8912_37509.n15 40.8964
R11716 a_8912_37509.n18 a_8912_37509.n17 40.8964
R11717 a_8912_37509.n22 a_8912_37509.n21 40.8964
R11718 a_8912_37509.n24 a_8912_37509.n23 40.8964
R11719 a_8912_37509.n26 a_8912_37509.n25 40.8964
R11720 a_8912_37509.n33 a_8912_37509.n32 40.6735
R11721 a_8912_37509.n35 a_8912_37509.n34 40.6735
R11722 a_8912_37509.n37 a_8912_37509.n36 40.6735
R11723 a_8912_37509.n41 a_8912_37509.n40 40.6735
R11724 a_8912_37509.n43 a_8912_37509.n42 40.6735
R11725 a_8912_37509.n45 a_8912_37509.n44 40.6735
R11726 a_8912_37509.n2 a_8912_37509.t33 30.0869
R11727 a_8912_37509.n29 a_8912_37509.t32 30.0869
R11728 a_8912_37509.n11 a_8912_37509.t36 30.0869
R11729 a_8912_37509.n9 a_8912_37509.t34 30.0869
R11730 a_8912_37509.n6 a_8912_37509.t35 30.0869
R11731 a_8912_37509.n4 a_8912_37509.t37 30.0869
R11732 a_8912_37509.n3 a_8912_37509.n2 5.95542
R11733 a_8912_37509.n29 a_8912_37509.n28 5.6486
R11734 a_8912_37509.n12 a_8912_37509.n11 5.6486
R11735 a_8912_37509.n10 a_8912_37509.n9 5.6486
R11736 a_8912_37509.n6 a_8912_37509.n1 5.6486
R11737 a_8912_37509.n4 a_8912_37509.n3 5.6486
R11738 a_8912_37509.n5 a_8912_37509.n2 4.80732
R11739 a_8912_37509.n32 a_8912_37509.t29 4.76133
R11740 a_8912_37509.n32 a_8912_37509.t28 4.76133
R11741 a_8912_37509.n34 a_8912_37509.t25 4.76133
R11742 a_8912_37509.n34 a_8912_37509.t24 4.76133
R11743 a_8912_37509.n36 a_8912_37509.t30 4.76133
R11744 a_8912_37509.n36 a_8912_37509.t20 4.76133
R11745 a_8912_37509.n40 a_8912_37509.t8 4.76133
R11746 a_8912_37509.n40 a_8912_37509.t12 4.76133
R11747 a_8912_37509.n42 a_8912_37509.t10 4.76133
R11748 a_8912_37509.n42 a_8912_37509.t1 4.76133
R11749 a_8912_37509.n13 a_8912_37509.t2 4.76133
R11750 a_8912_37509.n13 a_8912_37509.t11 4.76133
R11751 a_8912_37509.n15 a_8912_37509.t3 4.76133
R11752 a_8912_37509.n15 a_8912_37509.t0 4.76133
R11753 a_8912_37509.n17 a_8912_37509.t6 4.76133
R11754 a_8912_37509.n17 a_8912_37509.t7 4.76133
R11755 a_8912_37509.n21 a_8912_37509.t21 4.76133
R11756 a_8912_37509.n21 a_8912_37509.t17 4.76133
R11757 a_8912_37509.n23 a_8912_37509.t19 4.76133
R11758 a_8912_37509.n23 a_8912_37509.t22 4.76133
R11759 a_8912_37509.n25 a_8912_37509.t18 4.76133
R11760 a_8912_37509.n25 a_8912_37509.t26 4.76133
R11761 a_8912_37509.n45 a_8912_37509.t13 4.76133
R11762 a_8912_37509.t15 a_8912_37509.n45 4.76133
R11763 a_8912_37509.n5 a_8912_37509.n4 4.5005
R11764 a_8912_37509.n7 a_8912_37509.n6 4.5005
R11765 a_8912_37509.n9 a_8912_37509.n8 4.5005
R11766 a_8912_37509.n11 a_8912_37509.n0 4.5005
R11767 a_8912_37509.n30 a_8912_37509.n29 4.5005
R11768 a_8912_37509.n28 a_8912_37509.n27 1.19141
R11769 a_8912_37509.n31 a_8912_37509.n30 1.18686
R11770 a_8912_37509.n10 a_8912_37509.n1 0.614136
R11771 a_8912_37509.n8 a_8912_37509.n7 0.614136
R11772 a_8912_37509.n12 a_8912_37509.n10 0.318682
R11773 a_8912_37509.n8 a_8912_37509.n0 0.318682
R11774 a_8912_37509.n3 a_8912_37509.n1 0.307318
R11775 a_8912_37509.n28 a_8912_37509.n12 0.307318
R11776 a_8912_37509.n7 a_8912_37509.n5 0.307318
R11777 a_8912_37509.n30 a_8912_37509.n0 0.307318
R11778 a_8912_37509.n20 a_8912_37509.n19 0.261864
R11779 a_8912_37509.n39 a_8912_37509.n38 0.261864
R11780 a_8912_37509.n27 a_8912_37509.n26 0.227773
R11781 a_8912_37509.n24 a_8912_37509.n22 0.227773
R11782 a_8912_37509.n19 a_8912_37509.n18 0.227773
R11783 a_8912_37509.n18 a_8912_37509.n16 0.227773
R11784 a_8912_37509.n44 a_8912_37509.n43 0.227773
R11785 a_8912_37509.n43 a_8912_37509.n41 0.227773
R11786 a_8912_37509.n38 a_8912_37509.n37 0.227773
R11787 a_8912_37509.n37 a_8912_37509.n35 0.227773
R11788 a_8912_37509.n26 a_8912_37509.n24 0.216409
R11789 a_8912_37509.n22 a_8912_37509.n20 0.216409
R11790 a_8912_37509.n16 a_8912_37509.n14 0.216409
R11791 a_8912_37509.n44 a_8912_37509.n31 0.216409
R11792 a_8912_37509.n41 a_8912_37509.n39 0.216409
R11793 a_8912_37509.n35 a_8912_37509.n33 0.216409
R11794 VDD.n193 VDD.t1766 187509
R11795 VDD.n295 VDD.n193 135375
R11796 VDD.t69 VDD.n295 115781
R11797 VDD.n176 VDD.n99 15352.9
R11798 VDD.n176 VDD.n96 15352.9
R11799 VDD.n97 VDD.n95 15352.9
R11800 VDD.n167 VDD.n95 15352.9
R11801 VDD.n58 VDD.n50 13260
R11802 VDD.n55 VDD.n51 13260
R11803 VDD.n21 VDD.n14 13260
R11804 VDD.n18 VDD.n15 13260
R11805 VDD.n55 VDD.n50 13154.1
R11806 VDD.n58 VDD.n51 13154.1
R11807 VDD.n18 VDD.n14 13154.1
R11808 VDD.n21 VDD.n15 13154.1
R11809 VDD.n177 VDD.n93 11297.6
R11810 VDD.n177 VDD.n94 11297.6
R11811 VDD.n294 VDD.n293 9790.59
R11812 VDD.n171 VDD.n170 8029.09
R11813 VDD.n293 VDD.n195 8022.35
R11814 VDD.n325 VDD.n298 6963.53
R11815 VDD.n310 VDD.n298 6963.53
R11816 VDD.n294 VDD.n191 6374.12
R11817 VDD.n200 VDD.n192 5516.47
R11818 VDD.n107 VDD.n92 5440
R11819 VDD.n308 VDD.n192 5379.02
R11820 VDD.n326 VDD.n297 5177.65
R11821 VDD.n309 VDD.n297 5177.65
R11822 VDD.n106 VDD.n103 4253.52
R11823 VDD.n99 VDD.n94 4055.29
R11824 VDD.n96 VDD.n93 4055.29
R11825 VDD.n97 VDD.n94 4055.29
R11826 VDD.n330 VDD.n191 3220
R11827 VDD.n330 VDD.n192 3220
R11828 VDD.n233 VDD.n230 2311.76
R11829 VDD.n235 VDD.n230 2311.76
R11830 VDD.n241 VDD.n227 2311.76
R11831 VDD.n239 VDD.n227 2311.76
R11832 VDD.n173 VDD.n100 2291.2
R11833 VDD.n203 VDD.n202 2068.24
R11834 VDD.n202 VDD.n201 2068.24
R11835 VDD.n370 VDD.n364 1937.65
R11836 VDD.n371 VDD.n370 1937.65
R11837 VDD.n327 VDD.n326 1785.88
R11838 VDD.n326 VDD.n325 1785.88
R11839 VDD.n309 VDD.n308 1785.88
R11840 VDD.n310 VDD.n309 1785.88
R11841 VDD.n195 VDD.n194 1768.24
R11842 VDD.n376 VDD.n369 1757.65
R11843 VDD.n415 VDD.n360 1757.65
R11844 VDD.n376 VDD.n367 1757.65
R11845 VDD.n116 VDD.n110 1754.12
R11846 VDD.n121 VDD.n118 1754.12
R11847 VDD.n415 VDD.n361 1750.59
R11848 VDD.n327 VDD.n191 1718.82
R11849 VDD.n420 VDD.n355 1436.47
R11850 VDD.n388 VDD.n354 1436.47
R11851 VDD.n385 VDD.n374 1436.47
R11852 VDD.n384 VDD.n379 1436.47
R11853 VDD.n321 VDD.n302 1312.94
R11854 VDD.n317 VDD.n302 1312.94
R11855 VDD.n321 VDD.n303 1312.94
R11856 VDD.n231 VDD.n226 1231.76
R11857 VDD.n231 VDD.n228 1231.76
R11858 VDD.n178 VDD.n92 1195.67
R11859 VDD.n179 VDD.n178 1187.39
R11860 VDD.n233 VDD.n226 1080
R11861 VDD.n241 VDD.n226 1080
R11862 VDD.n235 VDD.n228 1080
R11863 VDD.n239 VDD.n228 1080
R11864 VDD.n111 VDD.n109 1080
R11865 VDD.n110 VDD.n108 1020
R11866 VDD.n121 VDD.n120 1020
R11867 VDD.n119 VDD.n109 1020
R11868 VDD.n120 VDD.n119 924.444
R11869 VDD.n119 VDD.n108 924.444
R11870 VDD.n434 VDD.t358 879.831
R11871 VDD.n356 VDD.n354 878.823
R11872 VDD.n379 VDD.n378 878.823
R11873 VDD.n378 VDD.n374 878.823
R11874 VDD.n67 VDD.t1659 877.016
R11875 VDD.n29 VDD.t2408 877.016
R11876 VDD.n2699 VDD.t56 873.438
R11877 VDD.n353 VDD.t1206 871.962
R11878 VDD.n72 VDD.t3071 871.962
R11879 VDD.n32 VDD.t3060 871.962
R11880 VDD.n420 VDD.n356 871.765
R11881 VDD.n4589 VDD.t943 871.529
R11882 VDD.n4245 VDD.t2377 871.529
R11883 VDD.n2384 VDD.t2260 870.221
R11884 VDD.n4237 VDD.t1546 869.669
R11885 VDD.n3229 VDD.t2365 867.614
R11886 VDD.n1915 VDD.t2750 866.47
R11887 VDD.n54 VDD.n52 861.352
R11888 VDD.n17 VDD.n12 861.268
R11889 VDD.n200 VDD.n194 857.648
R11890 VDD.n54 VDD.n53 857.359
R11891 VDD.n17 VDD.n16 857.183
R11892 VDD.n1043 VDD.t833 842.073
R11893 VDD.n4263 VDD.t2252 840.826
R11894 VDD.n106 VDD.n105 839.439
R11895 VDD.n2936 VDD.t1114 838.817
R11896 VDD.n2049 VDD.t3525 838.817
R11897 VDD.n2115 VDD.t3536 838.817
R11898 VDD.n2127 VDD.t3542 838.817
R11899 VDD.n4301 VDD.t1188 836.124
R11900 VDD.n3603 VDD.t955 836.124
R11901 VDD.n3552 VDD.t839 836.124
R11902 VDD.n2389 VDD.t1315 836.124
R11903 VDD.n1410 VDD.t2499 836.124
R11904 VDD.n3524 VDD.t2486 832.876
R11905 VDD.n3414 VDD.t2186 832.876
R11906 VDD.n3006 VDD.t679 832.876
R11907 VDD.n4629 VDD.t2256 807.261
R11908 VDD.n4566 VDD.t2784 806.511
R11909 VDD.n4322 VDD.t1723 806.511
R11910 VDD.n4203 VDD.t2856 806.511
R11911 VDD.n3685 VDD.t472 806.511
R11912 VDD.n3448 VDD.t3323 806.511
R11913 VDD.n3367 VDD.t2478 806.511
R11914 VDD.n2482 VDD.t2788 806.511
R11915 VDD.n1556 VDD.t1605 806.511
R11916 VDD.n1808 VDD.t992 806.511
R11917 VDD.n2182 VDD.t2422 806.511
R11918 VDD.n802 VDD.t1524 806.511
R11919 VDD.n1015 VDD.t2813 806.511
R11920 VDD.n3116 VDD.t3348 806.367
R11921 VDD.n4628 VDD.t100 804.731
R11922 VDD.n4008 VDD.t115 804.731
R11923 VDD.n4020 VDD.t103 804.731
R11924 VDD.n4444 VDD.t117 804.731
R11925 VDD.n4414 VDD.t152 804.731
R11926 VDD.n4066 VDD.t217 804.731
R11927 VDD.n4090 VDD.t84 804.731
R11928 VDD.n4164 VDD.t106 804.731
R11929 VDD.n4167 VDD.t195 804.731
R11930 VDD.n3970 VDD.t204 804.731
R11931 VDD.n3975 VDD.t193 804.731
R11932 VDD.t192 VDD.n3913 804.731
R11933 VDD.n3933 VDD.t139 804.731
R11934 VDD.n3936 VDD.t184 804.731
R11935 VDD.n3309 VDD.t226 804.731
R11936 VDD.n3312 VDD.t75 804.731
R11937 VDD.n3322 VDD.t220 804.731
R11938 VDD.n3330 VDD.t109 804.731
R11939 VDD.n3333 VDD.t207 804.731
R11940 VDD.n3114 VDD.t162 804.731
R11941 VDD.n3136 VDD.t156 804.731
R11942 VDD.n3139 VDD.t229 804.731
R11943 VDD.n2571 VDD.t142 804.731
R11944 VDD.n2580 VDD.t190 804.731
R11945 VDD.n2583 VDD.t211 804.731
R11946 VDD.t145 VDD.n2295 804.731
R11947 VDD.n2315 VDD.t78 804.731
R11948 VDD.n2318 VDD.t187 804.731
R11949 VDD.n1537 VDD.t159 804.731
R11950 VDD.n1696 VDD.t123 804.731
R11951 VDD.n1699 VDD.t93 804.731
R11952 VDD.n1899 VDD.t168 804.731
R11953 VDD.n1885 VDD.t167 804.731
R11954 VDD.n1870 VDD.t112 804.731
R11955 VDD.n1585 VDD.t90 804.731
R11956 VDD.n1910 VDD.t81 804.731
R11957 VDD.n2199 VDD.t232 804.731
R11958 VDD.n2202 VDD.t179 804.731
R11959 VDD.n859 VDD.t173 804.731
R11960 VDD.n862 VDD.t149 804.731
R11961 VDD.n1435 VDD.t202 804.731
R11962 VDD.n1438 VDD.t209 804.731
R11963 VDD.n611 VDD.t132 804.731
R11964 VDD.n2347 VDD.t330 804.216
R11965 VDD.n4022 VDD.t1190 804.135
R11966 VDD.n4446 VDD.t412 803.572
R11967 VDD.n4050 VDD.t570 803.572
R11968 VDD.n4072 VDD.t1428 803.572
R11969 VDD.n3525 VDD.t996 803.572
R11970 VDD.n3278 VDD.t540 803.572
R11971 VDD.n3461 VDD.t2121 803.572
R11972 VDD.n2511 VDD.t1182 803.572
R11973 VDD.n2180 VDD.t446 803.572
R11974 VDD.n968 VDD.t2544 803.572
R11975 VDD.n777 VDD.t2247 803.572
R11976 VDD.n1178 VDD.t2883 803.572
R11977 VDD.n1468 VDD.t1264 803.572
R11978 VDD.n2398 VDD.t1096 789.686
R11979 VDD.n2720 VDD.t3670 789.686
R11980 VDD.n1853 VDD.t3678 789.686
R11981 VDD.n1778 VDD.t3120 789.686
R11982 VDD.n1879 VDD.t1363 789.686
R11983 VDD.n1562 VDD.t1110 789.686
R11984 VDD.n1070 VDD.t2996 789.686
R11985 VDD.n731 VDD.t444 789.686
R11986 VDD.n744 VDD.t1106 789.686
R11987 VDD.n1281 VDD.t1804 789.686
R11988 VDD.n763 VDD.t526 789.686
R11989 VDD.n1191 VDD.t3635 789.686
R11990 VDD.n1373 VDD.t3442 789.686
R11991 VDD.n100 VDD.n92 787.201
R11992 VDD.n1486 VDD.t1920 786.62
R11993 VDD.n1101 VDD.t241 786.62
R11994 VDD.n1153 VDD.t3264 786.62
R11995 VDD.n3471 VDD.t1060 783.403
R11996 VDD.n2860 VDD.t1025 783.403
R11997 VDD.n2829 VDD.t492 783.403
R11998 VDD.n1807 VDD.t622 783.403
R11999 VDD.n3041 VDD.t20 779.372
R12000 VDD.n203 VDD.n200 755.294
R12001 VDD.n201 VDD.n195 755.294
R12002 VDD.t117 VDD.n4443 751.692
R12003 VDD.t152 VDD.n4048 751.692
R12004 VDD.t204 VDD.n3969 751.692
R12005 VDD.t193 VDD.n3974 751.692
R12006 VDD.n3972 VDD.t192 751.692
R12007 VDD.t226 VDD.n3308 751.692
R12008 VDD.n2297 VDD.t145 751.692
R12009 VDD.t90 VDD.n1584 751.692
R12010 VDD.n312 VDD.n311 742.777
R12011 VDD.t1205 VDD.n353 731.598
R12012 VDD.n104 VDD.n91 728.284
R12013 VDD.t100 VDD.n4627 725.173
R12014 VDD.t115 VDD.n4007 725.173
R12015 VDD.t103 VDD.n4019 725.173
R12016 VDD.t217 VDD.n4065 725.173
R12017 VDD.t84 VDD.n4089 725.173
R12018 VDD.t106 VDD.n4163 725.173
R12019 VDD.t195 VDD.n4166 725.173
R12020 VDD.t139 VDD.n3932 725.173
R12021 VDD.t184 VDD.n3935 725.173
R12022 VDD.t75 VDD.n3311 725.173
R12023 VDD.t220 VDD.n3321 725.173
R12024 VDD.t109 VDD.n3329 725.173
R12025 VDD.t207 VDD.n3332 725.173
R12026 VDD.t162 VDD.n3113 725.173
R12027 VDD.t156 VDD.n3135 725.173
R12028 VDD.t229 VDD.n3138 725.173
R12029 VDD.t142 VDD.n2570 725.173
R12030 VDD.t190 VDD.n2579 725.173
R12031 VDD.t211 VDD.n2582 725.173
R12032 VDD.t78 VDD.n2314 725.173
R12033 VDD.t187 VDD.n2317 725.173
R12034 VDD.t159 VDD.n1536 725.173
R12035 VDD.t123 VDD.n1695 725.173
R12036 VDD.t93 VDD.n1698 725.173
R12037 VDD.t112 VDD.n1869 725.173
R12038 VDD.t81 VDD.n1909 725.173
R12039 VDD.t232 VDD.n2198 725.173
R12040 VDD.t179 VDD.n2201 725.173
R12041 VDD.t173 VDD.n858 725.173
R12042 VDD.t149 VDD.n861 725.173
R12043 VDD.t202 VDD.n1434 725.173
R12044 VDD.t209 VDD.n1437 725.173
R12045 VDD.t132 VDD.n610 725.173
R12046 VDD.t2049 VDD.t1207 725.078
R12047 VDD.n1834 VDD.n1613 721.278
R12048 VDD.n2015 VDD.n2014 716.76
R12049 VDD.n3519 VDD.t246 700.506
R12050 VDD.n2871 VDD.t1879 700.506
R12051 VDD.n3073 VDD.t3445 700.506
R12052 VDD.n2485 VDD.t3123 700.506
R12053 VDD.n1384 VDD.t2991 700.506
R12054 VDD.n1379 VDD.t3715 700.506
R12055 VDD.n2720 VDD.t1521 699.386
R12056 VDD.n3195 VDD.t1916 696.322
R12057 VDD.n2650 VDD.t1961 685.97
R12058 VDD.n3976 VDD.t1887 677.846
R12059 VDD.n4470 VDD.t3240 675.293
R12060 VDD.n4051 VDD.t3752 675.293
R12061 VDD.n4365 VDD.t2842 675.293
R12062 VDD.n3721 VDD.t1499 675.293
R12063 VDD.n883 VDD.t1530 675.293
R12064 VDD.n118 VDD.n111 674.119
R12065 VDD.n116 VDD.n111 674.119
R12066 VDD.n152 VDD.t2540 672.854
R12067 VDD.n152 VDD.t2392 672.77
R12068 VDD.n154 VDD.t1244 671.888
R12069 VDD.n151 VDD.t1243 671.888
R12070 VDD.n4424 VDD.t1874 671.408
R12071 VDD.n3768 VDD.t320 671.408
R12072 VDD.n2915 VDD.t3570 671.408
R12073 VDD.n2289 VDD.t1250 671.408
R12074 VDD.n2597 VDD.t3201 671.408
R12075 VDD.n2139 VDD.t691 671.408
R12076 VDD.n923 VDD.t3423 671.408
R12077 VDD.n4614 VDD.t763 667.778
R12078 VDD.n3991 VDD.t749 667.778
R12079 VDD.n4014 VDD.t1673 667.778
R12080 VDD.n4452 VDD.t2633 667.778
R12081 VDD.n4406 VDD.t1583 667.778
R12082 VDD.n2620 VDD.t294 667.778
R12083 VDD.n1550 VDD.t1491 667.778
R12084 VDD.n2226 VDD.t2578 667.778
R12085 VDD.n2220 VDD.t583 667.778
R12086 VDD.n1122 VDD.t2322 667.778
R12087 VDD.n986 VDD.t2862 667.778
R12088 VDD.n1133 VDD.t2584 667.778
R12089 VDD.n4635 VDD.t1468 667.751
R12090 VDD.n4557 VDD.t1687 667.751
R12091 VDD.n4270 VDD.t887 667.751
R12092 VDD.n4139 VDD.t1353 667.751
R12093 VDD.n3733 VDD.t2586 667.751
R12094 VDD.n3262 VDD.t798 667.751
R12095 VDD.n3459 VDD.t2617 667.751
R12096 VDD.n3384 VDD.t2304 667.751
R12097 VDD.n2522 VDD.t2703 667.751
R12098 VDD.n2354 VDD.t2720 667.751
R12099 VDD.n2643 VDD.t2200 667.751
R12100 VDD.n2241 VDD.t2330 667.751
R12101 VDD.n1037 VDD.t2482 667.751
R12102 VDD.n960 VDD.t2133 667.751
R12103 VDD.n1210 VDD.t1156 667.751
R12104 VDD.n3270 VDD.t3506 667.611
R12105 VDD.n3448 VDD.t1414 666.366
R12106 VDD.n4308 VDD.t1180 665.736
R12107 VDD.n1846 VDD.t3177 665.307
R12108 VDD.n4030 VDD.t1222 664.455
R12109 VDD.n4440 VDD.t2158 664.455
R12110 VDD.n4043 VDD.t2654 664.455
R12111 VDD.n4373 VDD.t3485 664.455
R12112 VDD.n3477 VDD.t2819 664.455
R12113 VDD.n3355 VDD.t1736 664.455
R12114 VDD.n3178 VDD.t1456 664.455
R12115 VDD.n1981 VDD.t1184 664.455
R12116 VDD.n1800 VDD.t2647 664.455
R12117 VDD.n2248 VDD.t544 664.455
R12118 VDD.n1100 VDD.t1671 664.455
R12119 VDD.n1145 VDD.t3327 664.455
R12120 VDD.n1478 VDD.t1327 664.455
R12121 VDD.n4394 VDD.t1202 664.326
R12122 VDD.n4372 VDD.t2954 663.636
R12123 VDD.n4216 VDD.t2289 663.426
R12124 VDD.n3678 VDD.t2574 663.426
R12125 VDD.n3539 VDD.t292 663.426
R12126 VDD.n3435 VDD.t2786 663.426
R12127 VDD.n3294 VDD.t873 663.426
R12128 VDD.n3121 VDD.t2353 663.426
R12129 VDD.n2504 VDD.t2782 663.426
R12130 VDD.n2303 VDD.t646 663.426
R12131 VDD.n1619 VDD.t2324 663.426
R12132 VDD.n1010 VDD.t903 663.426
R12133 VDD.n771 VDD.t1519 663.426
R12134 VDD.n1421 VDD.t587 663.426
R12135 VDD.n1596 VDD.t2772 662.841
R12136 VDD.n1588 VDD.t3108 662.841
R12137 VDD.n1998 VDD.t514 659.593
R12138 VDD.n60 VDD.n48 657.715
R12139 VDD.n24 VDD.n23 657.715
R12140 VDD.n59 VDD.n49 647.111
R12141 VDD.n22 VDD.n13 647.111
R12142 VDD.n4092 VDD.n4091 630.699
R12143 VDD.n3900 VDD.n3899 629.801
R12144 VDD.n4582 VDD.n3990 629.801
R12145 VDD.n4565 VDD.n3997 629.801
R12146 VDD.n4535 VDD.n4016 629.801
R12147 VDD.n4505 VDD.n4037 629.801
R12148 VDD.n4328 VDD.n4273 629.801
R12149 VDD.n3695 VDD.n3694 629.801
R12150 VDD.n3691 VDD.n3690 629.801
R12151 VDD.n3656 VDD.n3212 629.801
R12152 VDD.n3226 VDD.n3225 629.801
R12153 VDD.n3614 VDD.n3577 629.801
R12154 VDD.n3365 VDD.n3302 629.801
R12155 VDD.n3182 VDD.n3181 629.801
R12156 VDD.n3844 VDD.n3821 629.801
R12157 VDD.n3097 VDD.n3096 629.801
R12158 VDD.n2838 VDD.n2837 629.801
R12159 VDD.n2281 VDD.n2280 629.801
R12160 VDD.n2460 VDD.n2459 629.801
R12161 VDD.n2669 VDD.n2668 629.801
R12162 VDD.n1318 VDD.n1317 629.801
R12163 VDD.t1643 VDD.t88 621.025
R12164 VDD.n1839 VDD.n1609 613.89
R12165 VDD.n2012 VDD.n2011 611.178
R12166 VDD.n3483 VDD.n3281 611.122
R12167 VDD.n2827 VDD.n2826 611.122
R12168 VDD.n2418 VDD.n2417 611.122
R12169 VDD.n1817 VDD.n1622 611.122
R12170 VDD.n2853 VDD.n2842 610.861
R12171 VDD.n2844 VDD.n2843 610.861
R12172 VDD.n2413 VDD.n2412 610.861
R12173 VDD.n3051 VDD.n3011 610.861
R12174 VDD.n3049 VDD.n3014 610.307
R12175 VDD.n2880 VDD.n2879 610.098
R12176 VDD.n1809 VDD.n1627 610.098
R12177 VDD.n2855 VDD.n2840 609.847
R12178 VDD.n3016 VDD.n3015 609.847
R12179 VDD.n3498 VDD.n3272 609.615
R12180 VDD.n3274 VDD.n3273 609.615
R12181 VDD.n3490 VDD.n3277 609.615
R12182 VDD.n2815 VDD.n2814 609.615
R12183 VDD.n1833 VDD.n1614 609.615
R12184 VDD.n1824 VDD.n1618 609.615
R12185 VDD.n2907 VDD.n2407 609.37
R12186 VDD.n2999 VDD.n2998 609.37
R12187 VDD.n2821 VDD.n2420 608.178
R12188 VDD.n622 VDD.n618 607.212
R12189 VDD.n622 VDD.n619 607.212
R12190 VDD.n634 VDD.n608 607.212
R12191 VDD.n539 VDD.n535 607.212
R12192 VDD.n539 VDD.n536 607.212
R12193 VDD.n551 VDD.n527 607.212
R12194 VDD.n551 VDD.n528 607.212
R12195 VDD.n459 VDD.n455 607.212
R12196 VDD.n459 VDD.n456 607.212
R12197 VDD.n471 VDD.n447 607.212
R12198 VDD.n471 VDD.n448 607.212
R12199 VDD.n1866 VDD.n1593 607.155
R12200 VDD.n823 VDD.n822 607.155
R12201 VDD.n1326 VDD.n1325 607.155
R12202 VDD.n1289 VDD.n746 607.155
R12203 VDD.n422 VDD.t2049 606.698
R12204 VDD.n4252 VDD.n4106 606.505
R12205 VDD.n4250 VDD.n4109 606.505
R12206 VDD.n3479 VDD.n3286 606.42
R12207 VDD.n3485 VDD.n3280 606.42
R12208 VDD.n2886 VDD.n2825 606.42
R12209 VDD.n3053 VDD.n3008 606.42
R12210 VDD.n1625 VDD.n1624 606.42
R12211 VDD.n1819 VDD.n1621 606.42
R12212 VDD.n4257 VDD.n4102 605.971
R12213 VDD.n3476 VDD.n3287 605.581
R12214 VDD.n2409 VDD.n2408 605.186
R12215 VDD.n2898 VDD.n2411 605.186
R12216 VDD.n2362 VDD.n2361 605.186
R12217 VDD.n3058 VDD.n3005 605.186
R12218 VDD.n2416 VDD.n2415 605.186
R12219 VDD.n1616 VDD.n1615 605.186
R12220 VDD.n4604 VDD.n4603 604.457
R12221 VDD.n4559 VDD.n4000 604.457
R12222 VDD.n4526 VDD.n4028 604.457
R12223 VDD.n4375 VDD.n4076 604.457
R12224 VDD.n4197 VDD.n4138 604.457
R12225 VDD.n3688 VDD.n3687 604.457
R12226 VDD.n3517 VDD.n3260 604.457
R12227 VDD.n3455 VDD.n3454 604.457
R12228 VDD.n2525 VDD.n2524 604.457
R12229 VDD.n2658 VDD.n2657 604.457
R12230 VDD.n1979 VDD.n1978 604.457
R12231 VDD.n1802 VDD.n1633 604.457
R12232 VDD.n2174 VDD.n2173 604.457
R12233 VDD.n805 VDD.n804 604.457
R12234 VDD.n1020 VDD.n1019 604.457
R12235 VDD.n782 VDD.n781 604.457
R12236 VDD.n1170 VDD.n1143 604.457
R12237 VDD.n1475 VDD.n1406 604.457
R12238 VDD.n4671 VDD.n4670 604.394
R12239 VDD.n4584 VDD.n3989 604.394
R12240 VDD.n4543 VDD.n4013 604.394
R12241 VDD.n4463 VDD.n4462 604.394
R12242 VDD.n4396 VDD.n4062 604.394
R12243 VDD.n4286 VDD.n4285 604.394
R12244 VDD.n3249 VDD.n3248 604.394
R12245 VDD.n3505 VDD.n3267 604.394
R12246 VDD.n3408 VDD.n3407 604.394
R12247 VDD.n2611 VDD.n2610 604.394
R12248 VDD.n2048 VDD.n1547 604.394
R12249 VDD.n2221 VDD.n2188 604.394
R12250 VDD.n1125 VDD.n793 604.394
R12251 VDD.n1066 VDD.n1065 604.394
R12252 VDD.n1237 VDD.n768 604.394
R12253 VDD.n1192 VDD.n1130 604.394
R12254 VDD.n1454 VDD.n1423 604.394
R12255 VDD.n4527 VDD.n4025 604.076
R12256 VDD.n4397 VDD.n4059 604.076
R12257 VDD.n4104 VDD.n4103 604.076
R12258 VDD.n1930 VDD.n1569 603.859
R12259 VDD.n1114 VDD.n801 603.859
R12260 VDD.n1208 VDD.n784 603.859
R12261 VDD.n840 VDD.n838 603.402
R12262 VDD.n3652 VDD.n3217 603.231
R12263 VDD.n3429 VDD.n3428 603.231
R12264 VDD.n3854 VDD.n3814 603.231
R12265 VDD.n3838 VDD.n3824 603.231
R12266 VDD.n2735 VDD.n2466 603.231
R12267 VDD.n1950 VDD.n1949 603.231
R12268 VDD.n1302 VDD.n739 603.231
R12269 VDD.n4463 VDD.n4455 603.106
R12270 VDD.n3783 VDD.n3781 603.106
R12271 VDD.n2795 VDD.n2433 602.456
R12272 VDD.n2777 VDD.n2443 602.456
R12273 VDD.n1739 VDD.n1667 602.456
R12274 VDD.n4022 VDD.n4021 602.326
R12275 VDD.n1766 VDD.n1650 601.943
R12276 VDD.n4569 VDD.n4568 601.679
R12277 VDD.n4477 VDD.n4476 601.679
R12278 VDD.n3748 VDD.n3747 601.679
R12279 VDD.n3492 VDD.n3276 601.679
R12280 VDD.n3396 VDD.n3395 601.679
R12281 VDD.n3372 VDD.n3299 601.679
R12282 VDD.n2629 VDD.n2628 601.679
R12283 VDD.n2234 VDD.n2181 601.679
R12284 VDD.n2227 VDD.n2184 601.679
R12285 VDD.n1052 VDD.n1051 601.679
R12286 VDD.n1138 VDD.n1137 601.679
R12287 VDD.n1414 VDD.n1413 601.679
R12288 VDD.n3359 VDD.n3358 601.317
R12289 VDD.n4400 VDD.n4057 601.097
R12290 VDD.n4223 VDD.n4125 601.097
R12291 VDD.n3670 VDD.n3669 601.097
R12292 VDD.n3442 VDD.n3403 601.097
R12293 VDD.n3389 VDD.n3386 601.097
R12294 VDD.n3123 VDD.n3122 601.097
R12295 VDD.n2502 VDD.n2501 601.097
R12296 VDD.n2306 VDD.n2305 601.097
R12297 VDD.n1827 VDD.n1826 601.097
R12298 VDD.n2214 VDD.n2191 601.097
R12299 VDD.n990 VDD.n989 601.097
R12300 VDD.n3566 VDD.n3231 600.904
R12301 VDD.n3553 VDD.n3241 600.904
R12302 VDD.n4440 VDD.n4439 600.105
R12303 VDD.n4421 VDD.n4045 600.105
R12304 VDD.n4329 VDD.n4272 600.105
R12305 VDD.n3284 VDD.n3283 600.105
R12306 VDD.n3388 VDD.n3387 600.105
R12307 VDD.n3110 VDD.n3109 600.105
R12308 VDD.n2349 VDD.n2294 600.105
R12309 VDD.n2480 VDD.n2479 600.105
R12310 VDD.n2704 VDD.n2661 600.105
R12311 VDD.n1759 VDD.n1656 600.105
R12312 VDD.n2179 VDD.n2178 600.105
R12313 VDD.n1783 VDD.n1641 599.966
R12314 VDD.n1752 VDD.n1660 599.966
R12315 VDD.n3253 VDD.n3252 599.933
R12316 VDD.n2982 VDD.n2373 599.933
R12317 VDD.n2706 VDD.n2660 599.933
R12318 VDD.n4620 VDD.n4610 599.808
R12319 VDD.n4643 VDD.n4598 599.808
R12320 VDD.n4005 VDD.n4004 599.808
R12321 VDD.n4437 VDD.n4436 599.808
R12322 VDD.n4264 VDD.n4098 599.808
R12323 VDD.n3927 VDD.n3926 599.808
R12324 VDD.n2983 VDD.n2372 599.808
R12325 VDD.n853 VDD.n852 599.808
R12326 VDD.n3584 VDD.n3583 599.74
R12327 VDD.n3571 VDD.n3570 599.74
R12328 VDD.n3558 VDD.n3237 599.74
R12329 VDD.n3546 VDD.n3247 599.74
R12330 VDD.n1965 VDD.n1964 599.74
R12331 VDD.n1854 VDD.n1600 599.74
R12332 VDD.n1524 VDD.n1523 599.74
R12333 VDD.n1878 VDD.n1877 599.74
R12334 VDD.n987 VDD.n829 599.74
R12335 VDD.n3116 VDD.n3115 599.212
R12336 VDD.n2687 VDD.n2671 599.159
R12337 VDD.n980 VDD.n833 599.159
R12338 VDD.n2544 VDD.n2506 598.986
R12339 VDD.n1635 VDD.n1634 598.986
R12340 VDD.n1776 VDD.n1644 598.986
R12341 VDD.n1745 VDD.n1663 598.986
R12342 VDD.n3662 VDD.n3209 598.965
R12343 VDD.n3579 VDD.n3578 598.965
R12344 VDD.n2832 VDD.n2831 598.965
R12345 VDD.n3034 VDD.n3025 598.965
R12346 VDD.n2754 VDD.n2454 598.965
R12347 VDD.n2742 VDD.n2462 598.965
R12348 VDD.n2019 VDD.n1958 598.965
R12349 VDD.n4609 VDD.n4608 598.383
R12350 VDD.n4050 VDD.n4049 598.383
R12351 VDD.n4387 VDD.n4071 598.383
R12352 VDD.n4281 VDD.n4278 598.383
R12353 VDD.n4208 VDD.n4130 598.383
R12354 VDD.n3528 VDD.n3527 598.383
R12355 VDD.n3401 VDD.n3400 598.383
R12356 VDD.n2537 VDD.n2509 598.383
R12357 VDD.n2343 VDD.n2299 598.383
R12358 VDD.n2036 VDD.n1555 598.383
R12359 VDD.n1811 VDD.n1810 598.383
R12360 VDD.n1115 VDD.n800 598.383
R12361 VDD.n978 VDD.n834 598.383
R12362 VDD.n1224 VDD.n776 598.383
R12363 VDD.n3796 VDD.n3185 596.97
R12364 VDD.n2821 VDD.n2421 596.97
R12365 VDD.n2536 VDD.n2510 596.619
R12366 VDD.n1787 VDD.n1785 596.619
R12367 VDD.n2084 VDD.n2083 596.442
R12368 VDD.n3709 VDD.n3703 595.668
R12369 VDD.n2997 VDD.n2364 595.668
R12370 VDD.n2085 VDD.n2082 595.668
R12371 VDD.n4132 VDD.n4131 594.144
R12372 VDD.n2813 VDD.n2424 594.144
R12373 VDD.n205 VDD.n190 588.424
R12374 VDD.n4135 VDD.n4134 585
R12375 VDD.n4196 VDD.n4195 585
R12376 VDD.n3791 VDD.n3790 585
R12377 VDD.n3803 VDD.n3802 585
R12378 VDD.n2805 VDD.n2804 585
R12379 VDD.n2613 VDD.n2612 585
R12380 VDD.n2615 VDD.n2614 585
R12381 VDD.n970 VDD.n969 585
R12382 VDD.n972 VDD.n971 585
R12383 VDD.n307 VDD.n190 573.763
R12384 VDD.n646 VDD.t3822 571.745
R12385 VDD.n385 VDD.n369 557.648
R12386 VDD.n394 VDD.n369 557.648
R12387 VDD.n394 VDD.n371 557.648
R12388 VDD.n371 VDD.n363 557.648
R12389 VDD.n363 VDD.n360 557.648
R12390 VDD.n388 VDD.n360 557.648
R12391 VDD.n384 VDD.n367 557.648
R12392 VDD.n395 VDD.n367 557.648
R12393 VDD.n395 VDD.n364 557.648
R12394 VDD.n413 VDD.n364 557.648
R12395 VDD.n413 VDD.n361 557.648
R12396 VDD.n361 VDD.n355 557.648
R12397 VDD.n175 VDD.n90 557.184
R12398 VDD.n305 VDD.n304 552.283
R12399 VDD.n306 VDD.n305 552.283
R12400 VDD.n313 VDD.n312 552.283
R12401 VDD.n201 VDD.t1757 545.926
R12402 VDD.n203 VDD.t3431 545.926
R12403 VDD.n2895 VDD.t315 543.817
R12404 VDD.n1200 VDD.t2959 543.817
R12405 VDD.n167 VDD.n108 542.485
R12406 VDD.n120 VDD.n93 531.895
R12407 VDD.n169 VDD.n100 514.134
R12408 VDD.n173 VDD.n172 477.44
R12409 VDD.t1411 VDD.t3103 473.322
R12410 VDD.t3462 VDD.t1967 471.644
R12411 VDD.t841 VDD.t3130 469.966
R12412 VDD.t2749 VDD.t169 464.93
R12413 VDD.t191 VDD.t203 463.252
R12414 VDD.t582 VDD.t3051 441.432
R12415 VDD.t2946 VDD.n422 440.348
R12416 VDD.n174 VDD.n173 435.346
R12417 VDD.t343 VDD.t2624 433.039
R12418 VDD.n341 VDD.t2050 431.428
R12419 VDD.t3339 VDD.n1658 421.291
R12420 VDD.t3261 VDD.t79 416.255
R12421 VDD.t1753 VDD.t1755 409.875
R12422 VDD.t1753 VDD.t1758 409.875
R12423 VDD.n648 VDD.t176 402.748
R12424 VDD.t215 VDD.t639 396.113
R12425 VDD.t361 VDD.t2015 396.113
R12426 VDD.n2081 VDD.t3039 395.495
R12427 VDD.n2097 VDD.t3037 395.495
R12428 VDD.n644 VDD.t175 394.139
R12429 VDD.t3237 VDD.n4502 392.757
R12430 VDD.t1703 VDD.t876 392.757
R12431 VDD.t3510 VDD.t349 392.757
R12432 VDD.t946 VDD.t104 391.079
R12433 VDD.t2517 VDD.t2545 391.079
R12434 VDD.t1133 VDD.t137 391.079
R12435 VDD.t473 VDD.t107 391.079
R12436 VDD.t1405 VDD.t154 391.079
R12437 VDD.t393 VDD.t188 391.079
R12438 VDD.t259 VDD.t76 391.079
R12439 VDD.t1167 VDD.t91 391.079
R12440 VDD.t287 VDD.t177 391.079
R12441 VDD.t3334 VDD.t147 391.079
R12442 VDD.t925 VDD.t200 391.079
R12443 VDD.t2086 VDD.t73 389.399
R12444 VDD.t3314 VDD.n3634 389.399
R12445 VDD.t865 VDD.n1199 389.399
R12446 VDD.n4448 VDD.t118 388.656
R12447 VDD.n4422 VDD.t153 388.656
R12448 VDD.n4381 VDD.t86 388.656
R12449 VDD.n4388 VDD.t87 388.656
R12450 VDD.n4128 VDD.t135 388.656
R12451 VDD.n4224 VDD.t136 388.656
R12452 VDD.n3671 VDD.t198 388.656
R12453 VDD.n3679 VDD.t199 388.656
R12454 VDD.n3357 VDD.t227 388.656
R12455 VDD.n3831 VDD.t125 388.656
R12456 VDD.n3886 VDD.t126 388.656
R12457 VDD.n2500 VDD.t128 388.656
R12458 VDD.n2550 VDD.t129 388.656
R12459 VDD.n3043 VDD.t234 388.656
R12460 VDD.n3023 VDD.t235 388.656
R12461 VDD.n2761 VDD.t164 388.656
R12462 VDD.n2764 VDD.t165 388.656
R12463 VDD.n2300 VDD.t146 388.656
R12464 VDD.n1272 VDD.t214 388.656
R12465 VDD.n1257 VDD.t213 388.656
R12466 VDD.n4659 VDD.t95 388.656
R12467 VDD.n3907 VDD.t96 388.656
R12468 VDD.n4315 VDD.t181 388.656
R12469 VDD.n4284 VDD.t182 388.656
R12470 VDD.n3962 VDD.t205 388.656
R12471 VDD.n3164 VDD.t120 388.656
R12472 VDD.n3125 VDD.t121 388.656
R12473 VDD.n1574 VDD.t170 388.656
R12474 VDD.n1923 VDD.t171 388.656
R12475 VDD.n1238 VDD.t222 388.656
R12476 VDD.n1245 VDD.t223 388.656
R12477 VDD.n1583 VDD.t89 387.682
R12478 VDD.t73 VDD.t225 386.043
R12479 VDD.t1245 VDD.t3481 384.365
R12480 VDD.t936 VDD.t1937 384.365
R12481 VDD.n4626 VDD.t99 380.193
R12482 VDD.n4006 VDD.t114 380.193
R12483 VDD.n4018 VDD.t102 380.193
R12484 VDD.n4064 VDD.t216 380.193
R12485 VDD.n4088 VDD.t83 380.193
R12486 VDD.n4162 VDD.t105 380.193
R12487 VDD.n4165 VDD.t194 380.193
R12488 VDD.n3931 VDD.t138 380.193
R12489 VDD.n3934 VDD.t183 380.193
R12490 VDD.n3310 VDD.t74 380.193
R12491 VDD.n3320 VDD.t219 380.193
R12492 VDD.n3328 VDD.t108 380.193
R12493 VDD.n3331 VDD.t206 380.193
R12494 VDD.n3112 VDD.t161 380.193
R12495 VDD.n3134 VDD.t155 380.193
R12496 VDD.n3137 VDD.t228 380.193
R12497 VDD.n2569 VDD.t141 380.193
R12498 VDD.n2578 VDD.t189 380.193
R12499 VDD.n2581 VDD.t210 380.193
R12500 VDD.n2313 VDD.t77 380.193
R12501 VDD.n2316 VDD.t186 380.193
R12502 VDD.n1535 VDD.t158 380.193
R12503 VDD.n1694 VDD.t122 380.193
R12504 VDD.n1697 VDD.t92 380.193
R12505 VDD.n1868 VDD.t111 380.193
R12506 VDD.n1908 VDD.t80 380.193
R12507 VDD.n2197 VDD.t231 380.193
R12508 VDD.n2200 VDD.t178 380.193
R12509 VDD.n857 VDD.t172 380.193
R12510 VDD.n860 VDD.t148 380.193
R12511 VDD.n1433 VDD.t201 380.193
R12512 VDD.n1436 VDD.t208 380.193
R12513 VDD.n609 VDD.t131 380.193
R12514 VDD.t1886 VDD.t191 372.615
R12515 VDD.t723 VDD.t1876 367.579
R12516 VDD.t882 VDD.t2877 367.579
R12517 VDD.t281 VDD.t1761 367.579
R12518 VDD.t1509 VDD.t1352 360.866
R12519 VDD.t886 VDD.t888 360.866
R12520 VDD.t2157 VDD.t908 360.866
R12521 VDD.t1739 VDD.t1735 360.866
R12522 VDD.t931 VDD.t2585 360.866
R12523 VDD.n165 VDD.t936 360.866
R12524 VDD.t3641 VDD.t764 359.188
R12525 VDD.t3345 VDD.t1647 359.188
R12526 VDD.t648 VDD.t3110 359.188
R12527 VDD.t238 VDD.t3758 359.188
R12528 VDD.n3641 VDD.t877 353.774
R12529 VDD.t1610 VDD.n164 352.082
R12530 VDD.n165 VDD.t660 350.796
R12531 VDD.n4597 VDD.t1474 350.582
R12532 VDD.n1968 VDD.t856 350.582
R12533 VDD.n1786 VDD.t298 350.582
R12534 VDD.n1028 VDD.t1633 350.582
R12535 VDD.n3101 VDD.t2452 350.582
R12536 VDD.n1510 VDD.t550 350.582
R12537 VDD.n811 VDD.t2599 350.582
R12538 VDD.n1154 VDD.t919 350.582
R12539 VDD.n1155 VDD.t1460 350.582
R12540 VDD.n706 VDD.t819 350.582
R12541 VDD.n2888 VDD.t3046 349.507
R12542 VDD.n2437 VDD.t3705 349.507
R12543 VDD.n4637 VDD.t1472 347.572
R12544 VDD.n1973 VDD.t860 347.572
R12545 VDD.n1795 VDD.t304 347.572
R12546 VDD.n1035 VDD.t1637 347.572
R12547 VDD.n620 VDD.t1047 347.572
R12548 VDD.n612 VDD.t724 347.572
R12549 VDD.n537 VDD.t2649 347.572
R12550 VDD.n529 VDD.t883 347.572
R12551 VDD.n457 VDD.t1151 347.572
R12552 VDD.n449 VDD.t282 347.572
R12553 VDD.n3868 VDD.t2456 347.57
R12554 VDD.n2250 VDD.t546 347.57
R12555 VDD.n1098 VDD.t2601 347.57
R12556 VDD.n1165 VDD.t915 347.57
R12557 VDD.n1207 VDD.t1466 347.57
R12558 VDD.n710 VDD.t813 347.57
R12559 VDD.n620 VDD.t1375 347.57
R12560 VDD.n537 VDD.t404 347.57
R12561 VDD.n529 VDD.t2160 347.57
R12562 VDD.n457 VDD.t705 347.57
R12563 VDD.n449 VDD.t1616 347.57
R12564 VDD.n1901 VDD.t1041 346.693
R12565 VDD.n1738 VDD.t634 345.885
R12566 VDD.t1024 VDD.t3101 345.76
R12567 VDD.n4085 VDD.t790 344.887
R12568 VDD.n4625 VDD.t2314 344.06
R12569 VDD.n4529 VDD.t1345 344.06
R12570 VDD.n4465 VDD.t733 344.06
R12571 VDD.n4497 VDD.t1214 344.06
R12572 VDD.n4395 VDD.t462 344.06
R12573 VDD.n4257 VDD.t2174 344.06
R12574 VDD.n3187 VDD.t2226 344.06
R12575 VDD.n4520 VDD.t1497 343.579
R12576 VDD.n4488 VDD.t909 343.579
R12577 VDD.n4077 VDD.t2805 343.579
R12578 VDD.n4190 VDD.t1510 343.579
R12579 VDD.n3731 VDD.t932 343.579
R12580 VDD.n3288 VDD.t2347 343.579
R12581 VDD.n2517 VDD.t2672 343.579
R12582 VDD.n2476 VDD.t986 343.579
R12583 VDD.n2243 VDD.t2738 343.579
R12584 VDD.n4335 VDD.t889 343.577
R12585 VDD.n331 VDD.n190 343.467
R12586 VDD.n958 VDD.t2135 343.308
R12587 VDD.n3411 VDD.t1825 342.841
R12588 VDD.n2152 VDD.t2998 342.841
R12589 VDD.n1341 VDD.t3532 342.839
R12590 VDD.n4096 VDD.t2127 342.772
R12591 VDD.t3543 VDD.t3428 342.404
R12592 VDD.n2398 VDD.t1506 341.553
R12593 VDD.n1664 VDD.t2940 341.154
R12594 VDD.n2985 VDD.t667 340.243
R12595 VDD.n866 VDD.t1239 340.243
R12596 VDD.n4596 VDD.t2113 340.241
R12597 VDD.n4005 VDD.t2396 340.241
R12598 VDD.n3940 VDD.t420 340.241
R12599 VDD.n2920 VDD.t3205 340.212
R12600 VDD.n2990 VDD.t3225 340.212
R12601 VDD.n3265 VDD.t3171 340.211
R12602 VDD.n2803 VDD.t3695 340.211
R12603 VDD.n4550 VDD.t1058 340.012
R12604 VDD.n4430 VDD.t2512 340.012
R12605 VDD.n3394 VDD.t2387 340.012
R12606 VDD.n3306 VDD.t1740 340.012
R12607 VDD.n2291 VDD.t1176 340.012
R12608 VDD.n3510 VDD.t802 340.01
R12609 VDD.n3379 VDD.t770 340.01
R12610 VDD.t872 VDD.t2303 339.046
R12611 VDD.t212 VDD.t3716 339.046
R12612 VDD.n1521 VDD.t3254 338.555
R12613 VDD.n2964 VDD.t434 338.11
R12614 VDD.n2756 VDD.t237 338.082
R12615 VDD.n2746 VDD.t1301 338.082
R12616 VDD.n2091 VDD.t2372 338.08
R12617 VDD.n2015 VDD.t3491 338.08
R12618 VDD.n2938 VDD.t1112 337.952
R12619 VDD.n1397 VDD.t697 337.95
R12620 VDD.n332 VDD.n331 337.423
R12621 VDD.n1771 VDD.t1692 337.096
R12622 VDD.n4237 VDD.t1412 336.567
R12623 VDD.n3788 VDD.t3487 336.567
R12624 VDD.n2158 VDD.t6 336.567
R12625 VDD.n2042 VDD.t52 336.567
R12626 VDD.n1975 VDD.t743 336.567
R12627 VDD.n918 VDD.t2558 336.567
R12628 VDD.n1606 VDD.t3223 336.522
R12629 VDD.n1526 VDD.t3003 335.257
R12630 VDD.n660 VDD.t1890 334.784
R12631 VDD.n671 VDD.t2919 334.784
R12632 VDD.n564 VDD.t3615 334.784
R12633 VDD.n567 VDD.t2876 334.784
R12634 VDD.n484 VDD.t2894 334.784
R12635 VDD.n487 VDD.t3706 334.784
R12636 VDD.n3560 VDD.t3504 334.784
R12637 VDD.n660 VDD.t2106 334.784
R12638 VDD.n564 VDD.t2890 334.784
R12639 VDD.n567 VDD.t1984 334.784
R12640 VDD.n484 VDD.t2026 334.784
R12641 VDD.n487 VDD.t2044 334.784
R12642 VDD.n4096 VDD.t2254 334.108
R12643 VDD.t2918 VDD.t333 334.012
R12644 VDD.t2889 VDD.t779 334.012
R12645 VDD.t2025 VDD.t1711 334.012
R12646 VDD.n654 VDD.t334 334.009
R12647 VDD.n593 VDD.t2521 334.009
R12648 VDD.n580 VDD.t1554 334.009
R12649 VDD.n513 VDD.t2547 334.009
R12650 VDD.n500 VDD.t1712 334.009
R12651 VDD.n654 VDD.t2320 334.007
R12652 VDD.n593 VDD.t368 334.007
R12653 VDD.n580 VDD.t780 334.007
R12654 VDD.n513 VDD.t1382 334.007
R12655 VDD.n500 VDD.t2362 334.007
R12656 VDD.n4292 VDD.t2576 333.368
R12657 VDD.n1515 VDD.t2643 333.368
R12658 VDD.n1059 VDD.t1446 333.366
R12659 VDD.n639 VDD.t1576 333.212
R12660 VDD.t2451 VDD.t3252 332.332
R12661 VDD.t1841 VDD.t569 330.654
R12662 VDD.t2980 VDD.t411 330.654
R12663 VDD.t2477 VDD.t3408 330.654
R12664 VDD.t3410 VDD.t3322 330.654
R12665 VDD.t1604 VDD.t3377 330.654
R12666 VDD.t2882 VDD.t1845 330.654
R12667 VDD.t3347 VDD.t160 328.976
R12668 VDD.n76 VDD.n71 326.158
R12669 VDD.n37 VDD.n36 326.158
R12670 VDD.n2909 VDD.n2908 325.82
R12671 VDD.n4450 VDD.n4449 325.627
R12672 VDD.n4407 VDD.n4053 325.627
R12673 VDD.n3698 VDD.n3697 325.627
R12674 VDD.n3193 VDD.n3192 325.627
R12675 VDD.n2145 VDD.n2137 325.627
R12676 VDD.n939 VDD.n938 325.627
R12677 VDD.n1018 VDD.n1017 324.74
R12678 VDD.n4642 VDD.n4599 323.988
R12679 VDD.n1988 VDD.n1970 323.988
R12680 VDD.n1793 VDD.n1637 323.988
R12681 VDD.n1027 VDD.n1026 323.988
R12682 VDD.n3873 VDD.n3102 323.986
R12683 VDD.n2255 VDD.n1514 323.986
R12684 VDD.n1093 VDD.n810 323.986
R12685 VDD.n1162 VDD.n1150 323.986
R12686 VDD.n789 VDD.n788 323.986
R12687 VDD.n1484 VDD.n707 323.986
R12688 VDD.n3911 VDD.n3910 322.329
R12689 VDD.n4431 VDD.n4042 322.329
R12690 VDD.n4359 VDD.n4358 322.329
R12691 VDD.n3067 VDD.n2288 322.329
R12692 VDD.n2604 VDD.n2491 322.329
R12693 VDD.n888 VDD.n887 322.329
R12694 VDD.t457 VDD.t2948 322.262
R12695 VDD.t2189 VDD.t345 322.262
R12696 VDD.t1409 VDD.t966 322.262
R12697 VDD.t3004 VDD.t2916 322.262
R12698 VDD.t1902 VDD.t1123 322.262
R12699 VDD.n2970 VDD.n2967 320.976
R12700 VDD.n352 VDD.n351 320.976
R12701 VDD.n717 VDD.n716 320.976
R12702 VDD.n1353 VDD.n715 320.976
R12703 VDD.n1346 VDD.n720 320.976
R12704 VDD.n432 VDD.n346 320.976
R12705 VDD.n69 VDD.n65 320.976
R12706 VDD.n40 VDD.n39 320.976
R12707 VDD.t2763 VDD.t1187 320.584
R12708 VDD.t429 VDD.t1872 320.584
R12709 VDD.t3643 VDD.t750 320.584
R12710 VDD.t3253 VDD.t2801 320.584
R12711 VDD.n616 VDD.n615 320.224
R12712 VDD.n688 VDD.n635 320.224
R12713 VDD.n533 VDD.n532 320.224
R12714 VDD.n600 VDD.n553 320.224
R12715 VDD.n453 VDD.n452 320.224
R12716 VDD.n520 VDD.n473 320.224
R12717 VDD.n616 VDD.n614 320.223
R12718 VDD.n533 VDD.n531 320.223
R12719 VDD.n600 VDD.n552 320.223
R12720 VDD.n453 VDD.n451 320.223
R12721 VDD.n520 VDD.n472 320.223
R12722 VDD.t134 VDD.t1196 318.906
R12723 VDD.t954 VDD.t3276 318.906
R12724 VDD.t119 VDD.t1586 318.906
R12725 VDD.t3136 VDD.t347 318.906
R12726 VDD.t1484 VDD.t3142 318.906
R12727 VDD.t163 VDD.t1749 318.906
R12728 VDD.t1826 VDD.t317 318.906
R12729 VDD.t1502 VDD.t2307 318.906
R12730 VDD.t1445 VDD.t1690 318.906
R12731 VDD.n1740 VDD.n1666 318.305
R12732 VDD.n136 VDD.n134 318.303
R12733 VDD.n4355 VDD.n4082 318.293
R12734 VDD.n3985 VDD.n3984 317.943
R12735 VDD.n4243 VDD.n4114 317.943
R12736 VDD.n4118 VDD.n4117 317.942
R12737 VDD.n2944 VDD.n2386 317.942
R12738 VDD.n898 VDD.n897 317.755
R12739 VDD.n2622 VDD.n2621 317.478
R12740 VDD.t2286 VDD.t3099 317.226
R12741 VDD.t1732 VDD.t2761 317.226
R12742 VDD.t595 VDD.t1891 317.226
R12743 VDD.t1157 VDD.t1163 317.226
R12744 VDD.t2532 VDD.t1165 317.226
R12745 VDD.t2029 VDD.t2141 317.226
R12746 VDD.t2213 VDD.t1762 317.226
R12747 VDD.t2968 VDD.t2791 317.226
R12748 VDD.t1423 VDD.t1441 317.226
R12749 VDD.t2449 VDD.t1981 317.226
R12750 VDD.n3776 VDD.n3775 317.104
R12751 VDD.n2835 VDD.n2834 317.104
R12752 VDD.n2123 VDD.n2122 317.104
R12753 VDD.n2635 VDD.n2483 317.103
R12754 VDD.n2713 VDD.n2655 317.103
R12755 VDD.t3572 VDD.t1977 315.548
R12756 VDD.t2847 VDD.t1496 315.548
R12757 VDD.t1933 VDD.t2109 315.548
R12758 VDD.t3166 VDD.t801 315.548
R12759 VDD.t3728 VDD.t1915 315.548
R12760 VDD.t1817 VDD.t3486 315.548
R12761 VDD.t373 VDD.t1385 315.548
R12762 VDD.t3743 VDD.t2021 315.548
R12763 VDD.t2425 VDD.t267 315.548
R12764 VDD.t2634 VDD.t3488 315.548
R12765 VDD.t2031 VDD.t2419 315.548
R12766 VDD.t1691 VDD.t2433 315.548
R12767 VDD.t3176 VDD.t822 315.548
R12768 VDD.t2755 VDD.t1813 315.548
R12769 VDD.t2965 VDD.t2766 315.548
R12770 VDD.t2969 VDD.t1415 315.548
R12771 VDD.t1717 VDD.t1559 315.548
R12772 VDD.t2306 VDD.t2967 315.548
R12773 VDD.t1354 VDD.t2966 315.548
R12774 VDD.t3747 VDD.t1985 315.548
R12775 VDD.n2878 VDD.n2877 315.406
R12776 VDD.n3029 VDD.n3027 315.406
R12777 VDD.n1366 VDD.n1365 315.406
R12778 VDD.n2367 VDD.n2366 315.334
R12779 VDD.n3504 VDD.n3268 315.334
R12780 VDD.n3270 VDD.n3269 315.334
R12781 VDD.n2427 VDD.n2426 315.334
R12782 VDD.n1611 VDD.n1610 315.334
R12783 VDD.n2104 VDD.n2103 315.301
R12784 VDD.n2152 VDD.n2132 315.301
R12785 VDD.n1943 VDD.n1942 315.221
R12786 VDD.n1310 VDD.n734 315.221
R12787 VDD.n1193 VDD.n1129 315.221
R12788 VDD.n1163 VDD.n1149 315.221
R12789 VDD.n1483 VDD.n709 315.221
R12790 VDD.n2928 VDD.n2396 315.221
R12791 VDD.n1876 VDD.n1591 315.221
R12792 VDD.n1288 VDD.n747 315.221
R12793 VDD.n1497 VDD.n702 315.221
R12794 VDD.n2405 VDD.n2404 315.089
R12795 VDD.n1911 VDD.n1907 314.49
R12796 VDD.n4357 VDD.n4081 313.94
R12797 VDD.t3630 VDD.t110 313.87
R12798 VDD.t3040 VDD.t1145 313.87
R12799 VDD.n3171 VDD.n3170 313.337
R12800 VDD.n1991 VDD.n1990 313.336
R12801 VDD.n1565 VDD.n1564 312.978
R12802 VDD.n4306 VDD.n4305 312.829
R12803 VDD.n2943 VDD.n2388 312.829
R12804 VDD.n3601 VDD.n3585 312.827
R12805 VDD.n3420 VDD.n3419 312.827
R12806 VDD.n433 VDD.n345 312.699
R12807 VDD.t3119 VDD.t2678 312.192
R12808 VDD.t1897 VDD.t3634 312.192
R12809 VDD.t3128 VDD.t221 312.192
R12810 VDD.n4145 VDD.n4144 312.053
R12811 VDD.n4181 VDD.n4149 312.053
R12812 VDD.n4178 VDD.n4155 312.053
R12813 VDD.n4161 VDD.n4160 312.053
R12814 VDD.n3919 VDD.n3918 312.053
R12815 VDD.n3923 VDD.n3922 312.053
R12816 VDD.n3348 VDD.n3316 312.053
R12817 VDD.n3763 VDD.n3762 312.053
R12818 VDD.n3327 VDD.n3326 312.053
R12819 VDD.n3150 VDD.n3128 312.053
R12820 VDD.n3144 VDD.n3132 312.053
R12821 VDD.n2565 VDD.n2564 312.053
R12822 VDD.n2577 VDD.n2576 312.053
R12823 VDD.n2312 VDD.n2311 312.053
R12824 VDD.n2069 VDD.n1534 312.053
R12825 VDD.n1731 VDD.n1676 312.053
R12826 VDD.n1685 VDD.n1684 312.053
R12827 VDD.n1688 VDD.n1687 312.053
R12828 VDD.n1693 VDD.n1692 312.053
R12829 VDD.n1955 VDD.n1954 312.053
R12830 VDD.n2196 VDD.n2195 312.053
R12831 VDD.n1123 VDD.n795 312.053
R12832 VDD.n1001 VDD.n821 312.053
R12833 VDD.n840 VDD.n839 312.053
R12834 VDD.n958 VDD.n843 312.053
R12835 VDD.n901 VDD.n900 312.053
R12836 VDD.n1354 VDD.n714 312.053
R12837 VDD.n724 VDD.n723 312.053
R12838 VDD.n1283 VDD.n750 312.053
R12839 VDD.n1251 VDD.n762 312.053
R12840 VDD.n1236 VDD.n770 312.053
R12841 VDD.n1184 VDD.n1136 312.053
R12842 VDD.n1172 VDD.n1142 312.053
R12843 VDD.n1398 VDD.n1360 312.053
R12844 VDD.n1369 VDD.n1368 312.053
R12845 VDD.n1372 VDD.n1371 312.053
R12846 VDD.n1474 VDD.n1409 312.053
R12847 VDD.n1461 VDD.n1417 312.053
R12848 VDD.n1455 VDD.n1422 312.053
R12849 VDD.n1428 VDD.n1427 312.053
R12850 VDD.n1432 VDD.n1431 312.053
R12851 VDD.n4348 VDD.n4087 312.051
R12852 VDD.n4244 VDD.n4112 312.051
R12853 VDD.n4230 VDD.n4121 312.051
R12854 VDD.n4189 VDD.n4141 312.051
R12855 VDD.n4182 VDD.n4147 312.051
R12856 VDD.n4177 VDD.n4156 312.051
R12857 VDD.n4161 VDD.n4159 312.051
R12858 VDD.n3953 VDD.n3921 312.051
R12859 VDD.n3348 VDD.n3315 312.051
R12860 VDD.n3327 VDD.n3325 312.051
R12861 VDD.n3150 VDD.n3126 312.051
R12862 VDD.n3144 VDD.n3131 312.051
R12863 VDD.n2393 VDD.n2392 312.051
R12864 VDD.n2529 VDD.n2515 312.051
R12865 VDD.n2563 VDD.n2562 312.051
R12866 VDD.n2577 VDD.n2575 312.051
R12867 VDD.n2312 VDD.n2310 312.051
R12868 VDD.n2047 VDD.n1548 312.051
R12869 VDD.n1685 VDD.n1683 312.051
R12870 VDD.n1693 VDD.n1691 312.051
R12871 VDD.n2118 VDD.n2117 312.051
R12872 VDD.n2157 VDD.n2129 312.051
R12873 VDD.n2196 VDD.n2194 312.051
R12874 VDD.n932 VDD.n931 312.051
R12875 VDD.n944 VDD.n881 312.051
R12876 VDD.n1428 VDD.n1426 312.051
R12877 VDD.n1432 VDD.n1430 312.051
R12878 VDD.n1541 VDD.n1540 312.005
R12879 VDD.n2375 VDD.n2374 311.659
R12880 VDD.n4618 VDD.n4612 311.659
R12881 VDD.n4458 VDD.n4457 311.659
R12882 VDD.n4490 VDD.n4489 311.659
R12883 VDD.n4100 VDD.n4099 311.659
R12884 VDD.n4251 VDD.n4107 311.659
R12885 VDD.n3947 VDD.n3925 311.659
R12886 VDD.n3190 VDD.n3189 311.659
R12887 VDD.n3512 VDD.n3264 311.521
R12888 VDD.n1391 VDD.n1364 311.521
R12889 VDD.n2641 VDD.n2478 311.519
R12890 VDD.n2006 VDD.n1962 311.519
R12891 VDD.n1334 VDD.n726 311.519
R12892 VDD.n2402 VDD.n2401 311.151
R12893 VDD.n1841 VDD.n1608 311.149
R12894 VDD.n3239 VDD.n3238 310.974
R12895 VDD.n2996 VDD.n2365 310.904
R12896 VDD.n2811 VDD.n2425 310.902
R12897 VDD.n2473 VDD.n2472 310.87
R12898 VDD.n808 VDD.n807 310.87
R12899 VDD.n1848 VDD.n1605 310.868
R12900 VDD.n1646 VDD.n1645 310.868
R12901 VDD.n1006 VDD.n1005 310.868
R12902 VDD.n1275 VDD.n1274 310.868
R12903 VDD.n1243 VDD.n765 310.868
R12904 VDD.t1496 VDD.t2976 310.512
R12905 VDD.n3594 VDD.n3593 310.502
R12906 VDD.n3621 VDD.n3620 310.502
R12907 VDD.n2930 VDD.n2395 310.502
R12908 VDD.n2136 VDD.n2135 310.502
R12909 VDD.n3565 VDD.n3232 310.5
R12910 VDD.n4299 VDD.n4298 309.726
R12911 VDD.n4232 VDD.n4120 309.726
R12912 VDD.n3783 VDD.n3782 309.726
R12913 VDD.n2163 VDD.n2126 309.726
R12914 VDD.n1013 VDD.n1012 309.724
R12915 VDD.n3960 VDD.n3959 309.647
R12916 VDD.n3529 VDD.n3257 309.531
R12917 VDD.n1467 VDD.n1412 309.531
R12918 VDD.n3548 VDD.n3245 309.531
R12919 VDD.n3059 VDD.n3004 309.531
R12920 VDD.n3852 VDD.n3815 309.519
R12921 VDD.n2969 VDD.n2968 309.517
R12922 VDD.n2680 VDD.n2674 309.517
R12923 VDD.n1579 VDD.n1578 309.517
R12924 VDD.n1872 VDD.n1871 309.476
R12925 VDD.n1886 VDD.t3774 309.034
R12926 VDD.n4342 VDD.t82 308.834
R12927 VDD.t985 VDD.t1960 308.834
R12928 VDD.t1175 VDD.t2961 308.834
R12929 VDD.t88 VDD.t166 308.834
R12930 VDD.n3942 VDD.n3929 308.755
R12931 VDD.n3324 VDD.n3323 308.755
R12932 VDD.n2574 VDD.n2573 308.755
R12933 VDD.n1654 VDD.n1653 308.755
R12934 VDD.n1734 VDD.n1673 308.755
R12935 VDD.n1724 VDD.n1681 308.755
R12936 VDD.n2140 VDD.n2138 308.755
R12937 VDD.n1348 VDD.n719 308.755
R12938 VDD.n753 VDD.n752 308.755
R12939 VDD.n1225 VDD.n775 308.755
R12940 VDD.n1086 VDD.n813 308.755
R12941 VDD.n1072 VDD.n1007 308.755
R12942 VDD.n912 VDD.n896 308.755
R12943 VDD.n1218 VDD.n779 308.755
R12944 VDD.n3967 VDD.n3915 308.755
R12945 VDD.n4293 VDD.n4290 308.755
R12946 VDD.n3708 VDD.n3704 308.755
R12947 VDD.n2336 VDD.n2302 308.755
R12948 VDD.n2309 VDD.n2308 308.755
R12949 VDD.n2213 VDD.n2192 308.755
R12950 VDD.n1085 VDD.n814 308.755
R12951 VDD.n1034 VDD.n1022 308.755
R12952 VDD.n925 VDD.n889 308.755
R12953 VDD.n868 VDD.n855 308.755
R12954 VDD.n873 VDD.n851 308.151
R12955 VDD.n4601 VDD.n4600 308.149
R12956 VDD.n4551 VDD.n4549 308.149
R12957 VDD.n4525 VDD.n4029 308.149
R12958 VDD.n4399 VDD.n4058 308.149
R12959 VDD.n3415 VDD.n3413 307.204
R12960 VDD.n2005 VDD.n1963 307.204
R12961 VDD.n1603 VDD.n1602 307.204
R12962 VDD.n826 VDD.n825 307.204
R12963 VDD.n431 VDD.n347 307.204
R12964 VDD.t2616 VDD.t2120 307.156
R12965 VDD.n847 VDD.n846 306.896
R12966 VDD.n2257 VDD.n1513 306.428
R12967 VDD.n664 VDD.n656 306.428
R12968 VDD.n659 VDD.n658 306.428
R12969 VDD.n651 VDD.n650 306.428
R12970 VDD.n677 VDD.n641 306.428
R12971 VDD.n561 VDD.n560 306.428
R12972 VDD.n587 VDD.n563 306.428
R12973 VDD.n571 VDD.n570 306.428
R12974 VDD.n574 VDD.n573 306.428
R12975 VDD.n481 VDD.n480 306.428
R12976 VDD.n507 VDD.n483 306.428
R12977 VDD.n491 VDD.n490 306.428
R12978 VDD.n494 VDD.n493 306.428
R12979 VDD.n1553 VDD.n1552 306.428
R12980 VDD.n1982 VDD.n1974 306.428
R12981 VDD.n895 VDD.n894 306.428
R12982 VDD.n664 VDD.n655 306.428
R12983 VDD.n659 VDD.n657 306.428
R12984 VDD.n561 VDD.n559 306.428
R12985 VDD.n587 VDD.n562 306.428
R12986 VDD.n571 VDD.n569 306.428
R12987 VDD.n574 VDD.n572 306.428
R12988 VDD.n481 VDD.n479 306.428
R12989 VDD.n507 VDD.n482 306.428
R12990 VDD.n491 VDD.n489 306.428
R12991 VDD.n494 VDD.n492 306.428
R12992 VDD.t3147 VDD.t2995 305.478
R12993 VDD.t732 VDD.t2632 302.12
R12994 VDD.t746 VDD.t3244 302.12
R12995 VDD.t3524 VDD.t1815 302.12
R12996 VDD.t914 VDD.t519 302.12
R12997 VDD.t3124 VDD.t2163 298.764
R12998 VDD.t2445 VDD.t1095 298.764
R12999 VDD.n133 VDD.t2282 293.685
R13000 VDD.t2700 VDD.t694 292.05
R13001 VDD.t1490 VDD.t2822 292.05
R13002 VDD.t3272 VDD.t3316 290.372
R13003 VDD.t1995 VDD.t1179 288.693
R13004 VDD.t3520 VDD.t2785 288.693
R13005 VDD.t1181 VDD.t1255 287.014
R13006 VDD.t1518 VDD.t1259 287.014
R13007 VDD.t586 VDD.t3053 287.014
R13008 VDD.t1824 VDD.t3764 285.337
R13009 VDD.t197 VDD.t2573 283.658
R13010 VDD.t1888 VDD.t2602 281.979
R13011 VDD.n423 VDD.t2682 281.979
R13012 VDD.t2565 VDD.t3280 278.623
R13013 VDD.t1535 VDD.t2747 275.265
R13014 VDD.t2313 VDD.t2255 270.231
R13015 VDD.t328 VDD.t561 268.551
R13016 VDD.t1757 VDD.n193 265.26
R13017 VDD.t3431 VDD.n193 265.26
R13018 VDD.n322 VDD.t1770 264.262
R13019 VDD.t1300 VDD.t1640 263.517
R13020 VDD.t1310 VDD.t251 263.517
R13021 VDD.t3739 VDD.t1871 261.837
R13022 VDD.t3242 VDD.t3737 261.837
R13023 VDD.t3625 VDD.t1632 261.837
R13024 VDD.n3234 VDD.n3233 260.031
R13025 VDD.n3243 VDD.n3242 260.031
R13026 VDD.n2431 VDD.n2430 259.697
R13027 VDD.n2780 VDD.n2441 259.697
R13028 VDD.n2693 VDD.n2667 259.697
R13029 VDD.n1671 VDD.n1670 259.697
R13030 VDD.n350 VDD.t2947 259.577
R13031 VDD.t1038 VDD.t2630 258.481
R13032 VDD.n844 VDD.t408 257.913
R13033 VDD.n3426 VDD.t1347 257.474
R13034 VDD.n2922 VDD.t2446 257.474
R13035 VDD.n2130 VDD.t2631 257.474
R13036 VDD.n3792 VDD.t3685 255.905
R13037 VDD.n2380 VDD.t322 255.905
R13038 VDD.n2796 VDD.t510 255.905
R13039 VDD.n2064 VDD.t1503 255.905
R13040 VDD.n135 VDD.t1609 255.905
R13041 VDD.n143 VDD.t661 255.905
R13042 VDD.n125 VDD.t937 255.905
R13043 VDD.n4630 VDD.t2357 255.904
R13044 VDD.n4560 VDD.t1620 255.904
R13045 VDD.n4032 VDD.t2442 255.904
R13046 VDD.n4035 VDD.t2237 255.904
R13047 VDD.n4074 VDD.t3757 255.904
R13048 VDD.n3581 VDD.t3277 255.904
R13049 VDD.n3009 VDD.t384 255.904
R13050 VDD.n2772 VDD.t3637 255.904
R13051 VDD.n2070 VDD.t3010 255.904
R13052 VDD.n1730 VDD.t3083 255.904
R13053 VDD.n2075 VDD.t2917 255.904
R13054 VDD.n141 VDD.t3482 255.904
R13055 VDD.n125 VDD.t2390 255.904
R13056 VDD.n76 VDD.t1655 255.904
R13057 VDD.n37 VDD.t2194 255.904
R13058 VDD.n638 VDD.t3093 255.125
R13059 VDD.n556 VDD.t1962 255.125
R13060 VDD.n476 VDD.t1772 255.125
R13061 VDD.n3727 VDD.t2016 255.075
R13062 VDD.n1396 VDD.t3708 254.907
R13063 VDD.n4497 VDD.t3238 254.541
R13064 VDD.n4340 VDD.t3181 254.475
R13065 VDD.n4336 VDD.t3203 252.95
R13066 VDD.n2958 VDD.t318 252.95
R13067 VDD.n2794 VDD.t512 252.95
R13068 VDD.n2698 VDD.t2839 252.95
R13069 VDD.n3982 VDD.t3496 252.948
R13070 VDD.n4634 VDD.t2355 252.948
R13071 VDD.n4558 VDD.t1618 252.948
R13072 VDD.n4512 VDD.t2444 252.948
R13073 VDD.n4511 VDD.t2239 252.948
R13074 VDD.n4374 VDD.t3755 252.948
R13075 VDD.n3608 VDD.t3273 252.948
R13076 VDD.n3440 VDD.t1394 252.948
R13077 VDD.n3012 VDD.t380 252.948
R13078 VDD.n2770 VDD.t3628 252.948
R13079 VDD.n2489 VDD.t1485 252.948
R13080 VDD.n1732 VDD.t3085 252.948
R13081 VDD.n2074 VDD.t3005 252.948
R13082 VDD.n1530 VDD.t2910 252.948
R13083 VDD.n3731 VDD.t2014 251.786
R13084 VDD.t1427 VDD.t85 251.768
R13085 VDD.t3444 VDD.t1883 251.768
R13086 VDD.t329 VDD.t144 251.768
R13087 VDD.n556 VDD.t367 251.768
R13088 VDD.n476 VDD.t1381 251.768
R13089 VDD.n1688 VDD.t632 251.516
R13090 VDD.n3796 VDD.t3692 251.044
R13091 VDD.n2499 VDD.t3137 250.724
R13092 VDD.n2665 VDD.t2846 250.724
R13093 VDD.n208 VDD.t1767 250.724
R13094 VDD.n3912 VDD.t3498 250.722
R13095 VDD.n3406 VDD.t1400 250.722
R13096 VDD.n2603 VDD.t1488 250.722
R13097 VDD.n1710 VDD.t630 250.722
R13098 VDD.n4491 VDD.t907 250.464
R13099 VDD.n4040 VDD.t2516 250.464
R13100 VDD.n3727 VDD.t934 250.464
R13101 VDD.n4095 VDD.t891 250.463
R13102 VDD.n4341 VDD.t2126 250.089
R13103 VDD.n4010 VDD.t2395 250.089
R13104 VDD.t2112 VDD.n4650 250.089
R13105 VDD.t834 VDD.t1855 250.089
R13106 VDD.n3045 VDD.t701 249.972
R13107 VDD.n712 VDD.t3453 249.901
R13108 VDD.n133 VDD.t2283 249.387
R13109 VDD.n4188 VDD.t1268 249.363
R13110 VDD.n4176 VDD.t1681 249.363
R13111 VDD.n4170 VDD.t947 249.363
R13112 VDD.n3317 VDD.t1434 249.363
R13113 VDD.n3197 VDD.t2693 249.363
R13114 VDD.n3859 VDD.t374 249.363
R13115 VDD.n3336 VDD.t474 249.363
R13116 VDD.n3129 VDD.t2525 249.363
R13117 VDD.n3133 VDD.t2567 249.363
R13118 VDD.n2975 VDD.t3463 249.363
R13119 VDD.n2771 VDD.t1282 249.363
R13120 VDD.n2468 VDD.t3759 249.363
R13121 VDD.n2714 VDD.t2844 249.363
R13122 VDD.n2586 VDD.t394 249.363
R13123 VDD.n2321 VDD.t2167 249.363
R13124 VDD.n2055 VDD.t1501 249.363
R13125 VDD.n2054 VDD.t1108 249.363
R13126 VDD.n1764 VDD.t747 249.363
R13127 VDD.n1729 VDD.t951 249.363
R13128 VDD.n1722 VDD.t2142 249.363
R13129 VDD.n1716 VDD.t1562 249.363
R13130 VDD.n1702 VDD.t2432 249.363
R13131 VDD.n2080 VDD.t1426 249.363
R13132 VDD.n2111 VDD.t3247 249.363
R13133 VDD.n2020 VDD.t897 249.363
R13134 VDD.n2268 VDD.t1124 249.363
R13135 VDD.n2205 VDD.t288 249.363
R13136 VDD.n1121 VDD.t452 249.363
R13137 VDD.n1088 VDD.t2769 249.363
R13138 VDD.n966 VDD.t2180 249.363
R13139 VDD.n905 VDD.t2218 249.363
R13140 VDD.n910 VDD.t1729 249.363
R13141 VDD.n1216 VDD.t1404 249.363
R13142 VDD.n1396 VDD.t274 249.363
R13143 VDD.n1378 VDD.t982 249.363
R13144 VDD.n701 VDD.t772 249.363
R13145 VDD.n1453 VDD.t312 249.363
R13146 VDD.n1447 VDD.t2450 249.363
R13147 VDD.n1441 VDD.t926 249.363
R13148 VDD.n161 VDD.t2638 249.363
R13149 VDD.n4288 VDD.t809 249.362
R13150 VDD.n4110 VDD.t458 249.362
R13151 VDD.n4180 VDD.t2268 249.362
R13152 VDD.n4170 VDD.t2561 249.362
R13153 VDD.n3199 VDD.t1337 249.362
R13154 VDD.n3653 VDD.t961 249.362
R13155 VDD.n3629 VDD.t3315 249.362
R13156 VDD.n3317 VDD.t1333 249.362
R13157 VDD.n3761 VDD.t1894 249.362
R13158 VDD.n3336 VDD.t2212 249.362
R13159 VDD.n3129 VDD.t1733 249.362
R13160 VDD.n3133 VDD.t1406 249.362
R13161 VDD.n2861 VDD.t3102 249.362
R13162 VDD.n2495 VDD.t1227 249.362
R13163 VDD.n3033 VDD.t2104 249.362
R13164 VDD.n2757 VDD.t2190 249.362
R13165 VDD.n2586 VDD.t578 249.362
R13166 VDD.n2327 VDD.t1158 249.362
R13167 VDD.n2321 VDD.t260 249.362
R13168 VDD.n1867 VDD.t1483 249.362
R13169 VDD.n1861 VDD.t1390 249.362
R13170 VDD.n1716 VDD.t1275 249.362
R13171 VDD.n1702 VDD.t1168 249.362
R13172 VDD.n2211 VDD.t2214 249.362
R13173 VDD.n2205 VDD.t459 249.362
R13174 VDD.n936 VDD.t2807 249.362
R13175 VDD.n727 VDD.t2048 249.362
R13176 VDD.n1447 VDD.t2825 249.362
R13177 VDD.n1441 VDD.t1357 249.362
R13178 VDD.n161 VDD.t1938 249.362
R13179 VDD.n2445 VDD.t3648 248.929
R13180 VDD.n844 VDD.t262 248.865
R13181 VDD.n70 VDD.t3062 248.843
R13182 VDD.n41 VDD.t3058 248.843
R13183 VDD.n77 VDD.t1661 248.843
R13184 VDD.n38 VDD.t2410 248.843
R13185 VDD.n3947 VDD.t574 248.688
R13186 VDD.t1207 VDD.t1209 248.599
R13187 VDD.t1209 VDD.t1203 248.599
R13188 VDD.t1203 VDD.t1205 248.599
R13189 VDD.n3953 VDD.t3331 248.475
R13190 VDD.n3919 VDD.t1174 248.475
R13191 VDD.n3923 VDD.t844 248.475
R13192 VDD.n4502 VDD.t2515 248.411
R13193 VDD.n1070 VDD.t560 248.243
R13194 VDD.n1281 VDD.t2860 248.243
R13195 VDD.n763 VDD.t913 248.243
R13196 VDD.n4495 VDD.t3236 248.219
R13197 VDD.n2556 VDD.t3150 248.219
R13198 VDD.n2062 VDD.t1508 248.219
R13199 VDD.n1362 VDD.t3723 248.219
R13200 VDD.n73 VDD.t1657 248.219
R13201 VDD.n33 VDD.t2196 248.219
R13202 VDD.n3812 VDD.t3260 247.394
R13203 VDD.n2802 VDD.t310 247.394
R13204 VDD.n2778 VDD.t3608 247.394
R13205 VDD.n2734 VDD.t1449 247.394
R13206 VDD.n2712 VDD.t806 247.394
R13207 VDD.n1545 VDD.t1816 247.394
R13208 VDD.n2076 VDD.t2713 247.394
R13209 VDD.n123 VDD.t1611 247.394
R13210 VDD.n3651 VDD.t3564 247.394
R13211 VDD.n3642 VDD.t2623 247.394
R13212 VDD.n3627 VDD.t1870 247.394
R13213 VDD.n3757 VDD.t2389 247.394
R13214 VDD.n2865 VDD.t2831 247.394
R13215 VDD.n2957 VDD.t563 247.394
R13216 VDD.n3013 VDD.t3440 247.394
R13217 VDD.n3035 VDD.t2531 247.394
R13218 VDD.n2793 VDD.t1410 247.394
R13219 VDD.n2755 VDD.t2232 247.394
R13220 VDD.n1594 VDD.t1002 247.394
R13221 VDD.n1324 VDD.t2732 247.394
R13222 VDD.n123 VDD.t1612 247.394
R13223 VDD.n238 VDD.n225 247.387
R13224 VDD.n236 VDD.n229 247.316
R13225 VDD.n1572 VDD.t3041 247.292
R13226 VDD.n1859 VDD.t2864 247.261
R13227 VDD.n2777 VDD.t2351 246.805
R13228 VDD.t3451 VDD.t2502 246.732
R13229 VDD.n2115 VDD.t829 246.573
R13230 VDD.n169 VDD.n168 245.761
R13231 VDD.n4627 VDD.t3770 245.667
R13232 VDD.n4007 VDD.t3773 245.667
R13233 VDD.n4019 VDD.t3815 245.667
R13234 VDD.n4065 VDD.t3800 245.667
R13235 VDD.n4089 VDD.t3780 245.667
R13236 VDD.n4163 VDD.t3794 245.667
R13237 VDD.n4166 VDD.t3792 245.667
R13238 VDD.n3932 VDD.t3767 245.667
R13239 VDD.n3935 VDD.t3806 245.667
R13240 VDD.n3311 VDD.t3789 245.667
R13241 VDD.n3321 VDD.t3802 245.667
R13242 VDD.n3329 VDD.t3797 245.667
R13243 VDD.n3332 VDD.t3816 245.667
R13244 VDD.n3113 VDD.t3769 245.667
R13245 VDD.n3135 VDD.t3813 245.667
R13246 VDD.n3138 VDD.t3777 245.667
R13247 VDD.n2570 VDD.t3810 245.667
R13248 VDD.n2579 VDD.t3827 245.667
R13249 VDD.n2582 VDD.t3807 245.667
R13250 VDD.n2314 VDD.t3795 245.667
R13251 VDD.n2317 VDD.t3801 245.667
R13252 VDD.n1536 VDD.t3781 245.667
R13253 VDD.n1695 VDD.t3791 245.667
R13254 VDD.n1698 VDD.t3782 245.667
R13255 VDD.n1869 VDD.t3778 245.667
R13256 VDD.n1909 VDD.t3826 245.667
R13257 VDD.n2198 VDD.t3821 245.667
R13258 VDD.n2201 VDD.t3803 245.667
R13259 VDD.n858 VDD.t3818 245.667
R13260 VDD.n861 VDD.t3796 245.667
R13261 VDD.n1434 VDD.t3808 245.667
R13262 VDD.n1437 VDD.t3814 245.667
R13263 VDD.n610 VDD.t3819 245.667
R13264 VDD.n3930 VDD.t1134 245.178
R13265 VDD.n3324 VDD.t2287 245.178
R13266 VDD.n2797 VDD.t1866 245.178
R13267 VDD.n2781 VDD.t3043 245.178
R13268 VDD.n2765 VDD.t1976 245.178
R13269 VDD.n2574 VDD.t596 245.178
R13270 VDD.n1708 VDD.t2533 245.178
R13271 VDD.n1332 VDD.t46 245.178
R13272 VDD.n1177 VDD.t2412 245.178
R13273 VDD.n1477 VDD.t2554 245.178
R13274 VDD.n1420 VDD.t899 245.178
R13275 VDD.n3645 VDD.t3243 245.178
R13276 VDD.n2513 VDD.t2152 245.178
R13277 VDD.n2899 VDD.t3561 245.178
R13278 VDD.n2951 VDD.t316 245.178
R13279 VDD.n2788 VDD.t2835 245.178
R13280 VDD.n890 VDD.t2792 245.178
R13281 VDD.n848 VDD.t1438 245.178
R13282 VDD.n856 VDD.t3335 245.178
R13283 VDD.t2543 VDD.t1999 245.054
R13284 VDD.n341 VDD.t1208 244.737
R13285 VDD.n348 VDD.t354 244.737
R13286 VDD.n3714 VDD.t342 244.498
R13287 VDD.n3657 VDD.t973 244.498
R13288 VDD.n3616 VDD.t1581 244.498
R13289 VDD.n2873 VDD.t530 244.496
R13290 VDD.n2991 VDD.t687 244.496
R13291 VDD.n2881 VDD.t3568 244.192
R13292 VDD.n2439 VDD.t3113 244.192
R13293 VDD.n1906 VDD.t3262 243.512
R13294 VDD.n917 VDD.t1398 243.512
R13295 VDD.n1301 VDD.t2012 243.512
R13296 VDD.n2494 VDD.t3734 243.512
R13297 VDD.n2609 VDD.t1544 243.512
R13298 VDD.n817 VDD.t3626 243.512
R13299 VDD.n2448 VDD.t1750 243.508
R13300 VDD.n2450 VDD.t346 243.508
R13301 VDD.n2057 VDD.t1557 243.508
R13302 VDD.n2905 VDD.t3342 243.508
R13303 VDD.t2855 VDD.t2659 243.375
R13304 VDD.n1929 VDD.t1043 242.76
R13305 VDD.n1928 VDD.t1868 242.268
R13306 VDD.n170 VDD.n169 242.036
R13307 VDD.n169 VDD.n103 242.036
R13308 VDD.n3755 VDD.t2388 241.696
R13309 VDD.t1895 VDD.t918 241.696
R13310 VDD.t818 VDD.t1905 241.696
R13311 VDD.n3022 VDD.t975 241.201
R13312 VDD.n1538 VDD.t3544 241.113
R13313 VDD.n3644 VDD.t344 240.792
R13314 VDD.n2952 VDD.t2897 240.215
R13315 VDD.n946 VDD.t256 240.215
R13316 VDD.n721 VDD.t3438 240.215
R13317 VDD.n755 VDD.t3717 240.215
R13318 VDD.n1266 VDD.t2904 240.215
R13319 VDD.n1231 VDD.t1806 240.215
R13320 VDD.n1147 VDD.t520 240.215
R13321 VDD.n426 VDD.t2683 240.215
R13322 VDD.n2292 VDD.t2993 240.214
R13323 VDD.n2492 VDD.t868 240.214
R13324 VDD.n1679 VDD.t3191 240.214
R13325 VDD.n2096 VDD.t3540 240.214
R13326 VDD.n875 VDD.t1992 240.214
R13327 VDD.t1867 VDD.t527 240.018
R13328 VDD.n3827 VDD.n3825 239.6
R13329 VDD.n1310 VDD.n733 239.6
R13330 VDD.n4543 VDD.n4012 238.544
R13331 VDD.n3714 VDD.n3701 238.544
R13332 VDD.n4651 VDD.t3495 238.339
R13333 VDD.t3636 VDD.n2726 238.339
R13334 VDD.n317 VDD.n316 237.584
R13335 VDD.n4503 VDD.t2240 236.661
R13336 VDD.n3319 VDD.t1332 236.661
R13337 VDD.n3755 VDD.t1336 236.661
R13338 VDD.n1689 VDD.t1274 236.661
R13339 VDD.t1437 VDD.n951 236.661
R13340 VDD.t2768 VDD.t2598 236.661
R13341 VDD.t2579 VDD.t3391 236.661
R13342 VDD.n3905 VDD.n3904 235.248
R13343 VDD.n4591 VDD.n4590 235.248
R13344 VDD.n4576 VDD.n3993 235.248
R13345 VDD.n4514 VDD.n4513 235.248
R13346 VDD.n4354 VDD.n4084 235.248
R13347 VDD.n4280 VDD.n4279 235.248
R13348 VDD.n3745 VDD.n3684 235.248
R13349 VDD.n3206 VDD.n3205 235.248
R13350 VDD.n3596 VDD.n3587 235.248
R13351 VDD.n3574 VDD.n3573 235.248
R13352 VDD.n3297 VDD.n3296 235.248
R13353 VDD.n3810 VDD.n3809 235.248
R13354 VDD.n3104 VDD.n3103 235.248
R13355 VDD.n2847 VDD.n2846 235.248
R13356 VDD.n2286 VDD.n2285 235.248
R13357 VDD.n2753 VDD.n2455 235.248
R13358 VDD.n2678 VDD.n2675 235.248
R13359 VDD.n4152 VDD.t2869 234.982
R13360 VDD.t2563 VDD.t1198 234.982
R13361 VDD.t3151 VDD.n4151 234.982
R13362 VDD.n4151 VDD.t2873 234.982
R13363 VDD.t1720 VDD.t2275 234.982
R13364 VDD.n4342 VDD.t2972 234.982
R13365 VDD.t1429 VDD.t642 234.982
R13366 VDD.t710 VDD.t275 234.982
R13367 VDD.t1592 VDD.n4010 234.982
R13368 VDD.n4651 VDD.t1547 234.982
R13369 VDD.n3469 VDD.t2346 234.982
R13370 VDD.t2155 VDD.t1626 234.982
R13371 VDD.n3634 VDD.t40 234.982
R13372 VDD.t2733 VDD.t2753 234.982
R13373 VDD.t2710 VDD.t1588 234.982
R13374 VDD.t2242 VDD.n2594 234.982
R13375 VDD.n2595 VDD.t2671 234.982
R13376 VDD.t331 VDD.t1317 234.982
R13377 VDD.n1658 VDD.t714 234.982
R13378 VDD.t649 VDD.n1598 234.982
R13379 VDD.t1453 VDD.t2691 234.982
R13380 VDD.n951 VDD.t835 234.982
R13381 VDD.t1147 VDD.t1435 234.982
R13382 VDD.t2290 VDD.t2559 234.982
R13383 VDD.n1078 VDD.t2924 234.982
R13384 VDD.t555 VDD.n1078 234.982
R13385 VDD.t1525 VDD.t1667 234.982
R13386 VDD.n1199 VDD.t3138 234.982
R13387 VDD.t1877 VDD.n1200 234.982
R13388 VDD.n1404 VDD.t2851 234.982
R13389 VDD.t2500 VDD.n1404 234.982
R13390 VDD.n406 VDD.t2055 234.042
R13391 VDD.n399 VDD.t2057 234.042
R13392 VDD.n5 VDD.t3645 233.44
R13393 VDD.n82 VDD.t3133 233.44
R13394 VDD.t1672 VDD.t3753 233.304
R13395 VDD.n406 VDD.t2058 232.798
R13396 VDD.n399 VDD.t2059 232.798
R13397 VDD.n638 VDD.t174 231.625
R13398 VDD.n336 VDD.t1771 230.201
R13399 VDD.n166 VDD.t1755 227.642
R13400 VDD.n98 VDD.t1758 227.642
R13401 VDD.t1688 VDD.t752 224.912
R13402 VDD.t1324 VDD.t43 224.912
R13403 VDD.n3820 VDD.n3819 224.139
R13404 VDD.n3654 VDD.n3214 223.869
R13405 VDD.n3541 VDD.n3251 223.869
R13406 VDD.n3827 VDD.n3826 223.869
R13407 VDD.n2663 VDD.n2662 223.869
R13408 VDD.n3433 VDD.n3409 223.868
R13409 VDD.n2464 VDD.n2463 223.868
R13410 VDD.t2429 VDD.t1646 223.233
R13411 VDD.n292 VDD.n188 222.655
R13412 VDD.n204 VDD.n199 220.613
R13413 VDD.n199 VDD.n198 220.613
R13414 VDD.n3111 VDD.n3108 219.787
R13415 VDD.n2965 VDD.n2379 219.787
R13416 VDD.n2471 VDD.n2470 219.787
R13417 VDD.n1996 VDD.n1967 219.787
R13418 VDD.n1893 VDD.n1581 219.787
R13419 VDD.n3851 VDD.n3816 219.516
R13420 VDD.n2370 VDD.n2369 219.516
R13421 VDD.n1560 VDD.n1559 219.516
R13422 VDD.n1304 VDD.n738 219.516
R13423 VDD.t1040 VDD.t2960 218.198
R13424 VDD.t2721 VDD.t1549 218.198
R13425 VDD.t543 VDD.t2642 216.519
R13426 VDD.n168 VDD.n107 215.041
R13427 VDD.t1621 VDD.t1686 214.841
R13428 VDD.t1467 VDD.t2358 214.841
R13429 VDD.t385 VDD.t375 214.841
R13430 VDD.t2953 VDD.t3484 213.163
R13431 VDD.t1309 VDD.t2702 213.163
R13432 VDD.t3558 VDD.t2132 213.163
R13433 VDD.t2884 VDD.t2481 213.163
R13434 VDD.n1584 VDD.t3799 213.148
R13435 VDD.n4341 VDD.n4340 213.119
R13436 VDD.n4393 VDD.n4069 213.119
R13437 VDD.n4504 VDD.n4503 213.119
R13438 VDD.n4650 VDD.n4649 213.119
R13439 VDD.n4179 VDD.n4152 213.119
R13440 VDD.n3470 VDD.n3469 213.119
R13441 VDD.n3634 VDD.n3633 213.119
R13442 VDD.n3754 VDD.n3753 213.119
R13443 VDD.n3865 VDD.n3864 213.119
R13444 VDD.n3343 VDD.n3319 213.119
R13445 VDD.n2726 VDD.n2445 213.119
R13446 VDD.n2594 VDD.n2593 213.119
R13447 VDD.n1715 VDD.n1689 213.119
R13448 VDD.n1806 VDD.n1631 213.119
R13449 VDD.n1597 VDD.n1576 213.119
R13450 VDD.n2030 VDD.n2029 213.119
R13451 VDD.n2171 VDD.n2170 213.119
R13452 VDD.n3756 VDD.n3755 213.119
R13453 VDD.n3636 VDD.n3635 213.119
R13454 VDD.n3468 VDD.n3258 213.119
R13455 VDD.n3467 VDD.n3466 213.119
R13456 VDD.n2895 VDD.n2384 213.119
R13457 VDD.n2596 VDD.n2595 213.119
R13458 VDD.n2028 VDD.n1532 213.119
R13459 VDD.n1859 VDD.n1598 213.119
R13460 VDD.n1757 VDD.n1658 213.119
R13461 VDD.n1080 VDD.n1079 213.119
R13462 VDD.n953 VDD.n952 213.119
R13463 VDD.n4658 VDD.t3784 210.964
R13464 VDD.n4314 VDD.t3787 210.964
R13465 VDD.n3830 VDD.t3768 210.964
R13466 VDD.n3042 VDD.t3793 210.964
R13467 VDD.n2762 VDD.t3772 210.964
R13468 VDD.n766 VDD.t3776 210.964
R13469 VDD.n246 VDD.n245 209.963
R13470 VDD.t748 VDD.t1917 209.806
R13471 VDD.t1921 VDD.t762 209.806
R13472 VDD.n3867 VDD.n3866 209.368
R13473 VDD.n3066 VDD.n3065 209.368
R13474 VDD.n2894 VDD.n2893 209.368
R13475 VDD.n2728 VDD.n2727 209.368
R13476 VDD.n2725 VDD.n2724 209.368
R13477 VDD.n2897 VDD.n2896 209.368
R13478 VDD.n3064 VDD.n3063 209.368
R13479 VDD.n2247 VDD.n2172 209.368
R13480 VDD.n2027 VDD.n2026 209.368
R13481 VDD.n1479 VDD.n1405 209.368
R13482 VDD.n1305 VDD.n737 209.368
R13483 VDD.n1202 VDD.n1201 209.368
R13484 VDD.n683 VDD.n638 209.368
R13485 VDD.n424 VDD.n423 209.368
R13486 VDD.n3973 VDD.t3811 208.409
R13487 VDD.t321 VDD.t1911 208.127
R13488 VDD.t185 VDD.n230 206.778
R13489 VDD.t133 VDD.n227 206.778
R13490 VDD.n410 VDD.n365 206.683
R13491 VDD.n392 VDD.n365 206.683
R13492 VDD.n171 VDD.n100 205.227
R13493 VDD.n81 VDD.t3785 204.754
R13494 VDD.n9 VDD.t3783 204.751
R13495 VDD.t1644 VDD.t2951 203.093
R13496 VDD.n1260 VDD.n1258 202.66
R13497 VDD.n6 VDD.t3824 202.582
R13498 VDD.n83 VDD.t3786 202.581
R13499 VDD.n84 VDD.t3825 202.576
R13500 VDD.n7 VDD.t3805 202.573
R13501 VDD.t3029 VDD.t531 201.413
R13502 VDD.t166 VDD.t3182 201.413
R13503 VDD.t2982 VDD.t3015 201.413
R13504 VDD.n67 VDD.n66 201.373
R13505 VDD.n29 VDD.n28 201.373
R13506 VDD.t1539 VDD.t2187 199.736
R13507 VDD.t2380 VDD.t2273 199.736
R13508 VDD.t716 VDD.t1397 198.058
R13509 VDD.t752 VDD.t297 196.379
R13510 VDD.n3866 VDD.t2455 194.701
R13511 VDD.n1405 VDD.t812 194.701
R13512 VDD.t3002 VDD.t3539 193.022
R13513 VDD.n307 VDD.n306 190.494
R13514 VDD.n311 VDD.n306 190.494
R13515 VDD.n1259 VDD.n757 190.165
R13516 VDD.t233 VDD.t19 187.987
R13517 VDD.n372 VDD.n366 187.482
R13518 VDD.n387 VDD.n372 187.482
R13519 VDD.n390 VDD.n359 187.482
R13520 VDD.n112 VDD.n101 187.107
R13521 VDD.n115 VDD.n114 187.107
R13522 VDD.n411 VDD.n359 186.73
R13523 VDD.n378 VDD.n377 185.882
R13524 VDD.n377 VDD.n376 185.882
R13525 VDD.n207 VDD.n206 184.056
R13526 VDD.t196 VDD.n232 183.653
R13527 VDD.n232 VDD.t224 183.653
R13528 VDD.t2063 VDD.t2489 182.952
R13529 VDD.t1141 VDD.t841 182.952
R13530 VDD.t2007 VDD.t2382 182.952
R13531 VDD.t588 VDD.t359 182.952
R13532 VDD.t1385 VDD.t377 182.952
R13533 VDD.t1230 VDD.t3652 182.952
R13534 VDD.t407 VDD.t261 182.952
R13535 VDD.n416 VDD.n415 182.309
R13536 VDD.n416 VDD.n356 182.309
R13537 VDD.t2513 VDD.t1827 181.273
R13538 VDD.t904 VDD.t2970 181.273
R13539 VDD.t3361 VDD.t1737 181.273
R13540 VDD.t1839 VDD.t799 181.273
R13541 VDD.t3316 VDD.t3296 181.273
R13542 VDD.t755 VDD.t1348 181.273
R13543 VDD.t1135 VDD.t1787 181.273
R13544 VDD.t3476 VDD.t3258 181.273
R13545 VDD.t3426 VDD.t2673 181.273
R13546 VDD.t3047 VDD.t3704 181.273
R13547 VDD.t3286 VDD.t3565 181.273
R13548 VDD.t3464 VDD.t1251 181.273
R13549 VDD.t3393 VDD.t1177 181.273
R13550 VDD.t3404 VDD.t299 181.273
R13551 VDD.t2935 VDD.t1040 181.273
R13552 VDD.t1146 VDD.t1823 181.273
R13553 VDD.t863 VDD.t3397 181.273
R13554 VDD.t1253 VDD.t3518 181.273
R13555 VDD.t3516 VDD.t1147 181.273
R13556 VDD.t1831 VDD.t1628 181.273
R13557 VDD.t1853 VDD.t920 181.273
R13558 VDD.t1479 VDD.t3385 179.595
R13559 VDD.t1641 VDD.t2231 179.595
R13560 VDD.t3320 VDD.t2935 179.595
R13561 VDD.n419 VDD.n357 178.008
R13562 VDD.n383 VDD.n382 178.008
R13563 VDD.t2111 VDD.t788 177.916
R13564 VDD.t956 VDD.t1878 176.238
R13565 VDD.t1189 VDD.t101 174.559
R13566 VDD.t1279 VDD.t1225 174.559
R13567 VDD.t1764 VDD.t1302 174.559
R13568 VDD.t656 VDD.t3642 172.881
R13569 VDD.t1881 VDD.t2620 172.881
R13570 VDD.t2840 VDD.t1931 172.881
R13571 VDD.t3753 VDD.t2019 172.881
R13572 VDD.t1884 VDD.t2608 172.881
R13573 VDD.t1871 VDD.t1923 172.881
R13574 VDD.t1909 VDD.t3242 172.881
R13575 VDD.t359 VDD.t1880 172.881
R13576 VDD.t3652 VDD.t2264 172.881
R13577 VDD.t2439 VDD.t756 172.881
R13578 VDD.t1783 VDD.t413 171.202
R13579 VDD.t2343 VDD.t3153 171.202
R13580 VDD.t2655 VDD.t3122 171.202
R13581 VDD.t1820 VDD.t389 171.202
R13582 VDD.t2217 VDD.t1308 171.202
R13583 VDD.t2988 VDD.t1118 171.202
R13584 VDD.t3687 VDD.t1677 171.202
R13585 VDD.t3537 VDD.t2587 171.202
R13586 VDD.t1745 VDD.t1997 169.524
R13587 VDD.t1161 VDD.t3690 169.524
R13588 VDD.t2922 VDD.t1048 169.524
R13589 VDD.t2891 VDD.t719 169.524
R13590 VDD.t1571 VDD.t3611 169.524
R13591 VDD.t337 VDD.t2078 169.524
R13592 VDD.t2036 VDD.t399 169.524
R13593 VDD.t2023 VDD.t884 169.524
R13594 VDD.t369 VDD.t3228 169.524
R13595 VDD.t777 VDD.t1970 169.524
R13596 VDD.t2027 VDD.t708 169.524
R13597 VDD.t2887 VDD.t285 169.524
R13598 VDD.t1379 VDD.t2956 169.524
R13599 VDD.t1707 VDD.t3094 169.524
R13600 VDD.t788 VDD.t2804 167.845
R13601 VDD.t3288 VDD.t1099 167.845
R13602 VDD.t3107 VDD.t1450 167.845
R13603 VDD.t513 VDD.t3448 167.845
R13604 VDD.t3000 VDD.t653 167.845
R13605 VDD.t2493 VDD.t2165 167.845
R13606 VDD.t684 VDD.t3458 167.845
R13607 VDD.t449 VDD.t1668 167.845
R13608 VDD.t3545 VDD.t590 167.845
R13609 VDD.n242 VDD.n225 166.901
R13610 VDD.n229 VDD.n223 166.611
R13611 VDD.t1198 VDD.t1350 166.167
R13612 VDD.t2795 VDD.t2066 166.167
R13613 VDD.t1722 VDD.t1719 166.167
R13614 VDD.t641 VDD.t1427 166.167
R13615 VDD.t411 VDD.t1093 166.167
R13616 VDD.t2469 VDD.t1189 166.167
R13617 VDD.t2475 VDD.t2611 166.167
R13618 VDD.t3290 VDD.t2299 166.167
R13619 VDD.t3298 VDD.t2590 166.167
R13620 VDD.t3508 VDD.t727 166.167
R13621 VDD.t1588 VDD.t1590 166.167
R13622 VDD.t1646 VDD.t2415 166.167
R13623 VDD.t3730 VDD.t2849 166.167
R13624 VDD.t3468 VDD.t565 166.167
R13625 VDD.t1316 VDD.t329 166.167
R13626 VDD.t1317 VDD.t2491 166.167
R13627 VDD.t2435 VDD.t2332 166.167
R13628 VDD.t2630 VDD.t2494 166.167
R13629 VDD.t445 VDD.t2739 166.167
R13630 VDD.t1603 VDD.t542 166.167
R13631 VDD.t1666 VDD.t1523 166.167
R13632 VDD.t1667 VDD.t1285 166.167
R13633 VDD.t2696 VDD.t3324 166.167
R13634 VDD.t3707 VDD.t273 166.167
R13635 VDD.t580 VDD.t1358 164.488
R13636 VDD.t2751 VDD.t197 164.488
R13637 VDD.t431 VDD.t760 164.488
R13638 VDD.t2838 VDD.t55 164.488
R13639 VDD.t3310 VDD.t2612 164.488
R13640 VDD.t565 VDD.t3224 164.488
R13641 VDD.t381 VDD.t2700 164.488
R13642 VDD.t1103 VDD.t2277 164.488
R13643 VDD.t1223 VDD.t3009 164.488
R13644 VDD.t2165 VDD.t3550 164.488
R13645 VDD.t688 VDD.t786 164.488
R13646 VDD.t692 VDD.t591 164.488
R13647 VDD.n117 VDD.t2391 164.072
R13648 VDD.t1267 VDD.t2871 162.81
R13649 VDD.t1835 VDD.t1429 162.81
R13650 VDD.t275 VDD.t1841 162.81
R13651 VDD.t3367 VDD.t1191 162.81
R13652 VDD.t3385 VDD.t2325 162.81
R13653 VDD.t2978 VDD.t2733 162.81
R13654 VDD.t3712 VDD.t371 162.81
R13655 VDD.t3446 VDD.t682 162.81
R13656 VDD.t3371 VDD.t2710 162.81
R13657 VDD.t3349 VDD.t2604 162.81
R13658 VDD.t2201 VDD.t3406 162.81
R13659 VDD.t3204 VDD.t3606 162.81
R13660 VDD.t2017 VDD.t2905 162.81
R13661 VDD.t3365 VDD.t331 162.81
R13662 VDD.t2950 VDD.t950 162.81
R13663 VDD.t3182 VDD.t3278 162.81
R13664 VDD.t3308 VDD.t523 162.81
R13665 VDD.t1859 VDD.t295 162.81
R13666 VDD.t1101 VDD.t1809 162.81
R13667 VDD.t1149 VDD.t3682 162.81
R13668 VDD.t1425 VDD.t3528 162.81
R13669 VDD.t3021 VDD.t1728 162.81
R13670 VDD.t251 VDD.t3659 162.81
R13671 VDD.t1855 VDD.t2814 162.81
R13672 VDD.t1845 VDD.t2337 162.81
R13673 VDD.t1811 VDD.t968 162.81
R13674 VDD.t3711 VDD.t981 162.81
R13675 VDD.t3363 VDD.t1324 162.81
R13676 VDD.t1283 VDD.t1989 161.131
R13677 VDD.t2618 VDD.t775 161.131
R13678 VDD.t2240 VDD.t738 161.131
R13679 VDD.t1907 VDD.t567 161.131
R13680 VDD.t1917 VDD.t1513 161.131
R13681 VDD.t2536 VDD.t1921 161.131
R13682 VDD.t2640 VDD.t421 161.131
R13683 VDD.t1693 VDD.t1193 161.131
R13684 VDD.t3157 VDD.t3196 161.131
R13685 VDD.t876 VDD.t2622 161.131
R13686 VDD.t2624 VDD.t958 161.131
R13687 VDD.t1139 VDD.t1143 161.131
R13688 VDD.t2729 VDD.t361 161.131
R13689 VDD.t3282 VDD.t2227 161.131
R13690 VDD.t375 VDD.t1127 161.131
R13691 VDD.t824 VDD.t1797 161.131
R13692 VDD.t1421 VDD.t1417 161.131
R13693 VDD.t2090 VDD.t3762 161.131
R13694 VDD.t127 VDD.t3149 161.131
R13695 VDD.t1960 VDD.t1638 161.131
R13696 VDD.t1000 VDD.t1520 161.131
R13697 VDD.t1364 VDD.t242 161.131
R13698 VDD.t2614 VDD.t3112 161.131
R13699 VDD.t3704 VDD.t2834 161.131
R13700 VDD.t2004 VDD.t964 161.131
R13701 VDD.t1823 VDD.t1807 161.131
R13702 VDD.t308 VDD.t962 161.131
R13703 VDD.t3492 VDD.t1500 161.131
R13704 VDD.t3535 VDD.t3248 161.131
R13705 VDD.t3550 VDD.t978 161.131
R13706 VDD.t3006 VDD.t3541 161.131
R13707 VDD.t2569 VDD.t1240 161.131
R13708 VDD.t425 VDD.t2907 161.131
R13709 VDD.t676 VDD.t3537 161.131
R13710 VDD.n971 VDD.n970 159.476
R13711 VDD.t1977 VDD.t944 159.452
R13712 VDD.t1989 VDD.t1265 159.452
R13713 VDD.t1185 VDD.t1995 159.452
R13714 VDD.t2109 VDD.t1171 159.452
R13715 VDD.t1987 VDD.t3328 159.452
R13716 VDD.t3650 VDD.t845 159.452
R13717 VDD.t2878 VDD.t575 159.452
R13718 VDD.t3099 VDD.t475 159.452
R13719 VDD.t2045 VDD.t2284 159.452
R13720 VDD.t1330 VDD.t2086 159.452
R13721 VDD.t2341 VDD.t3520 159.452
R13722 VDD.n3469 VDD.t1955 159.452
R13723 VDD.t1358 VDD.t3629 159.452
R13724 VDD.t247 VDD.t643 159.452
R13725 VDD.t1334 VDD.t1857 159.452
R13726 VDD.t2694 VDD.t3728 159.452
R13727 VDD.t3443 VDD.t431 159.452
R13728 VDD.t3337 VDD.t2828 159.452
R13729 VDD.t2826 VDD.t385 159.452
R13730 VDD.t2021 VDD.t1730 159.452
R13731 VDD.t2761 VDD.t1407 159.452
R13732 VDD.t1891 VDD.t395 159.452
R13733 VDD.t1965 VDD.t593 159.452
R13734 VDD.t2854 VDD.t3522 159.452
R13735 VDD.t1957 VDD.t2853 159.452
R13736 VDD.t1387 VDD.t42 159.452
R13737 VDD.t970 VDD.t2913 159.452
R13738 VDD.t1312 VDD.t2743 159.452
R13739 VDD.t974 VDD.t233 159.452
R13740 VDD.t1163 VDD.t257 159.452
R13741 VDD.t1165 VDD.t1169 159.452
R13742 VDD.t1276 VDD.t2029 159.452
R13743 VDD.t2143 VDD.t2041 159.452
R13744 VDD.t3518 VDD.t684 159.452
R13745 VDD.t1762 VDD.t289 159.452
R13746 VDD.t2559 VDD.t2808 159.452
R13747 VDD.t453 VDD.t449 159.452
R13748 VDD.t3336 VDD.t1461 159.452
R13749 VDD.t2765 VDD.t688 159.452
R13750 VDD.t773 VDD.t2203 159.452
R13751 VDD.t2496 VDD.t1935 159.452
R13752 VDD.t3053 VDD.t313 159.452
R13753 VDD.t1985 VDD.t2447 159.452
R13754 VDD.t1981 VDD.t927 159.452
R13755 VDD.t3622 VDD.t3290 157.774
R13756 VDD.t3140 VDD.t127 157.774
R13757 VDD.t3669 VDD.t3292 157.774
R13758 VDD.t242 VDD.t3730 157.774
R13759 VDD.t1801 VDD.t631 157.774
R13760 VDD.t3460 VDD.t1109 157.774
R13761 VDD.t3048 VDD.t3255 157.774
R13762 VDD.t3017 VDD.t240 157.774
R13763 VDD.t2092 VDD.t525 157.774
R13764 VDD.t2094 VDD.t1803 157.774
R13765 VDD.t2011 VDD.t425 157.774
R13766 VDD.t2907 VDD.t3472 157.774
R13767 VDD.n2430 VDD.t3266 157.014
R13768 VDD.n2441 VDD.t3619 157.014
R13769 VDD.n2667 VDD.t3125 156.998
R13770 VDD.n1670 VDD.t2929 156.998
R13771 VDD.t2401 VDD.t1511 156.095
R13772 VDD.t2575 VDD.t810 156.095
R13773 VDD.t101 VDD.t3367 156.095
R13774 VDD.t55 VDD.t1387 156.095
R13775 VDD.t2147 VDD.t2901 156.095
R13776 VDD.t2758 VDD.t3109 156.095
R13777 VDD.t1297 VDD.t1859 156.095
R13778 VDD.t2911 VDD.t2986 156.095
R13779 VDD.t2822 VDD.t2436 156.095
R13780 VDD.t3248 VDD.t1161 156.095
R13781 VDD.t2096 VDD.t771 156.095
R13782 VDD.t2836 VDD.t674 154.417
R13783 VDD.t1527 VDD.t1283 154.417
R13784 VDD.t1350 VDD.t2288 154.417
R13785 VDD.t3103 VDD.t1395 154.417
R13786 VDD.t1179 VDD.t2244 154.417
R13787 VDD.t1444 VDD.t1201 154.417
R13788 VDD.t2632 VDD.t1715 154.417
R13789 VDD.t1684 VDD.t748 154.417
R13790 VDD.t1713 VDD.t940 154.417
R13791 VDD.t762 VDD.t2727 154.417
R13792 VDD.t1863 VDD.t39 154.417
R13793 VDD.t2573 VDD.t469 154.417
R13794 VDD.t1590 VDD.t2352 154.417
R13795 VDD.t347 VDD.t3574 154.417
R13796 VDD.t1296 VDD.t3689 154.417
R13797 VDD.t3042 VDD.t2614 154.417
R13798 VDD.n3065 VDD.t2262 154.417
R13799 VDD.t822 VDD.t3300 154.417
R13800 VDD.t1549 VDD.t3460 154.417
R13801 VDD.t3528 VDD.t3038 154.417
R13802 VDD.t1435 VDD.t2962 154.417
R13803 VDD.t2098 VDD.t555 154.417
R13804 VDD.t2479 VDD.t902 154.417
R13805 VDD.t3011 VDD.t865 154.417
R13806 VDD.t1516 VDD.t2092 154.417
R13807 VDD.t1441 VDD.t3478 154.417
R13808 VDD.t584 VDD.t2096 154.417
R13809 VDD.n386 VDD.n373 153.225
R13810 VDD.n389 VDD.n358 153.225
R13811 VDD.t2541 VDD.t2980 152.739
R13812 VDD.t2828 VDD.t3684 152.739
R13813 VDD.t3109 VDD.t1691 152.739
R13814 VDD.t2494 VDD.t5 152.739
R13815 VDD.t525 VDD.t912 152.739
R13816 VDD.t1803 VDD.t2859 152.739
R13817 VDD.n1261 VDD.n1260 152
R13818 VDD.n647 VDD.n646 152
R13819 VDD.n643 VDD.n642 152
R13820 VDD.t1547 VDD.t94 151.06
R13821 VDD.n3635 VDD.t1703 151.06
R13822 VDD.t1520 VDD.t3669 151.06
R13823 VDD.t3265 VDD.t1865 151.06
R13824 VDD.t1137 VDD.t2928 151.06
R13825 VDD.t3541 VDD.t3507 151.06
R13826 VDD.t2691 VDD.t1600 151.06
R13827 VDD.t997 VDD.t3021 151.06
R13828 VDD.t1545 VDD.t1411 149.382
R13829 VDD.t2271 VDD.t1824 149.382
R13830 VDD.t2183 VDD.t1522 149.382
R13831 VDD.t838 VDD.t247 149.382
R13832 VDD.t2747 VDD.t293 149.382
R13833 VDD.t2502 VDD.t45 149.382
R13834 VDD.t1320 VDD.t900 149.382
R13835 VDD.n179 VDD.n91 149.249
R13836 VDD.t2871 VDD.t1052 147.703
R13837 VDD.t2873 VDD.t2795 147.703
R13838 VDD.t409 VDD.t1768 147.703
R13839 VDD.t2804 VDD.t2953 147.703
R13840 VDD.t1191 VDD.t2009 147.703
R13841 VDD.t2465 VDD.t1933 147.703
R13842 VDD.t1393 VDD.t2343 147.703
R13843 VDD.t2612 VDD.t3618 147.703
R13844 VDD.t2423 VDD.t3265 147.703
R13845 VDD.t2901 VDD.t1262 147.703
R13846 VDD.t2419 VDD.t1137 147.703
R13847 VDD.t2928 VDD.t2417 147.703
R13848 VDD.t3428 VDD.t1223 147.703
R13849 VDD.t828 VDD.t3535 147.703
R13850 VDD.t405 VDD.t3724 147.703
R13851 VDD.t2134 VDD.t3558 147.703
R13852 VDD.t2766 VDD.t2571 147.703
R13853 VDD.t1837 VDD.t3274 147.703
R13854 VDD.t2538 VDD.t2107 147.703
R13855 VDD.t1259 VDD.t3233 147.703
R13856 VDD.t1415 VDD.t2296 147.703
R13857 VDD.t3714 VDD.t3545 147.703
R13858 VDD.n180 VDD.n90 147.328
R13859 VDD.t1057 VDD.t1621 146.025
R13860 VDD.t3490 VDD.t2439 146.025
R13861 VDD.t1118 VDD.t571 146.025
R13862 VDD.t2066 VDD.t2663 144.346
R13863 VDD.t2171 VDD.t2169 144.346
R13864 VDD.t2169 VDD.t2173 144.346
R13865 VDD.t2130 VDD.t2124 144.346
R13866 VDD.t1719 VDD.t2245 144.346
R13867 VDD.t2669 VDD.t2763 144.346
R13868 VDD.t1443 VDD.t641 144.346
R13869 VDD.t467 VDD.t463 144.346
R13870 VDD.t463 VDD.t465 144.346
R13871 VDD.t713 VDD.t2295 144.346
R13872 VDD.t1217 VDD.t1215 144.346
R13873 VDD.t1211 VDD.t1217 144.346
R13874 VDD.t1093 VDD.t1716 144.346
R13875 VDD.t734 VDD.t732 144.346
R13876 VDD.t738 VDD.t736 144.346
R13877 VDD.t2399 VDD.t2393 144.346
R13878 VDD.t2393 VDD.t2397 144.346
R13879 VDD.t1685 VDD.t2800 144.346
R13880 VDD.t2207 VDD.t2728 144.346
R13881 VDD.t2309 VDD.t2311 144.346
R13882 VDD.t421 VDD.t415 144.346
R13883 VDD.t1059 VDD.t1081 144.346
R13884 VDD.t1081 VDD.t1063 144.346
R13885 VDD.t1079 VDD.t1069 144.346
R13886 VDD.t1071 VDD.t1073 144.346
R13887 VDD.t1087 VDD.t3168 144.346
R13888 VDD.t3168 VDD.t3212 144.346
R13889 VDD.t3212 VDD.t3216 144.346
R13890 VDD.t993 VDD.t1627 144.346
R13891 VDD.t1366 VDD.t1368 144.346
R13892 VDD.t2366 VDD.t2364 144.346
R13893 VDD.t470 VDD.t2754 144.346
R13894 VDD.t2227 VDD.t2223 144.346
R13895 VDD.t1591 VDD.t1589 144.346
R13896 VDD.t725 VDD.t3347 144.346
R13897 VDD.t3186 VDD.t2655 144.346
R13898 VDD.t3114 VDD.t1292 144.346
R13899 VDD.t3689 VDD.t3116 144.346
R13900 VDD.t3679 VDD.t249 144.346
R13901 VDD.t3694 VDD.t3700 144.346
R13902 VDD.t3698 VDD.t3696 144.346
R13903 VDD.t483 VDD.t507 144.346
R13904 VDD.t503 VDD.t489 144.346
R13905 VDD.t505 VDD.t493 144.346
R13906 VDD.t497 VDD.t485 144.346
R13907 VDD.t499 VDD.t481 144.346
R13908 VDD.t495 VDD.t487 144.346
R13909 VDD.t501 VDD.t495 144.346
R13910 VDD.t1028 VDD.t1022 144.346
R13911 VDD.t1006 VDD.t1030 144.346
R13912 VDD.t1020 VDD.t1034 144.346
R13913 VDD.t1014 VDD.t1012 144.346
R13914 VDD.t1012 VDD.t1018 144.346
R13915 VDD.t3208 VDD.t3218 144.346
R13916 VDD.t3218 VDD.t3204 144.346
R13917 VDD.t1911 VDD.t433 144.346
R13918 VDD.t672 VDD.t666 144.346
R13919 VDD.t3224 VDD.t3226 144.346
R13920 VDD.t3172 VDD.t3214 144.346
R13921 VDD.t11 VDD.t37 144.346
R13922 VDD.t21 VDD.t33 144.346
R13923 VDD.t17 VDD.t29 144.346
R13924 VDD.t25 VDD.t17 144.346
R13925 VDD.t19 VDD.t7 144.346
R13926 VDD.t2492 VDD.t1316 144.346
R13927 VDD.t635 VDD.t2926 144.346
R13928 VDD.t2926 VDD.t2939 144.346
R13929 VDD.t2065 VDD.t2062 144.346
R13930 VDD.t2062 VDD.t3121 144.346
R13931 VDD.t619 VDD.t599 144.346
R13932 VDD.t627 VDD.t605 144.346
R13933 VDD.t601 VDD.t603 144.346
R13934 VDD.t603 VDD.t615 144.346
R13935 VDD.t597 VDD.t623 144.346
R13936 VDD.t3174 VDD.t3210 144.346
R13937 VDD.t3210 VDD.t3222 144.346
R13938 VDD.t1362 VDD.t3107 144.346
R13939 VDD.t3267 VDD.t3686 144.346
R13940 VDD.t756 VDD.t3267 144.346
R13941 VDD.t3448 VDD.t1261 144.346
R13942 VDD.t740 VDD.t2145 144.346
R13943 VDD.t2438 VDD.t2331 144.346
R13944 VDD.t3038 VDD.t2914 144.346
R13945 VDD.t2914 VDD.t324 144.346
R13946 VDD.t652 VDD.t3002 144.346
R13947 VDD.t3036 VDD.t3048 144.346
R13948 VDD.t541 VDD.t1602 144.346
R13949 VDD.t1240 VDD.t1234 144.346
R13950 VDD.t1121 VDD.t1117 144.346
R13951 VDD.t2861 VDD.t2982 144.346
R13952 VDD.t1899 VDD.t2984 144.346
R13953 VDD.t1286 VDD.t1666 144.346
R13954 VDD.t1677 VDD.t2963 144.346
R13955 VDD.t2774 VDD.t1321 144.346
R13956 VDD.t1575 VDD.t1573 144.346
R13957 VDD.t1573 VDD.t1577 144.346
R13958 VDD.t1577 VDD.t1571 144.346
R13959 VDD.t3611 VDD.t2918 144.346
R13960 VDD.t333 VDD.t335 144.346
R13961 VDD.t335 VDD.t339 144.346
R13962 VDD.t339 VDD.t337 144.346
R13963 VDD.t2078 VDD.t1889 144.346
R13964 VDD.t367 VDD.t365 144.346
R13965 VDD.t365 VDD.t363 144.346
R13966 VDD.t363 VDD.t369 144.346
R13967 VDD.t3228 VDD.t2889 144.346
R13968 VDD.t779 VDD.t781 144.346
R13969 VDD.t781 VDD.t783 144.346
R13970 VDD.t783 VDD.t777 144.346
R13971 VDD.t1970 VDD.t1983 144.346
R13972 VDD.t1381 VDD.t1383 144.346
R13973 VDD.t1383 VDD.t1377 144.346
R13974 VDD.t1377 VDD.t1379 144.346
R13975 VDD.t2956 VDD.t2025 144.346
R13976 VDD.t1711 VDD.t1705 144.346
R13977 VDD.t1705 VDD.t1709 144.346
R13978 VDD.t1709 VDD.t1707 144.346
R13979 VDD.t3094 VDD.t2043 144.346
R13980 VDD.n1650 VDD.t1821 143.06
R13981 VDD.t892 VDD.t658 142.668
R13982 VDD.t1822 VDD.t2669 142.668
R13983 VDD.t2039 VDD.t417 142.668
R13984 VDD.t1368 VDD.t3194 142.668
R13985 VDD.t1199 VDD.t1279 142.668
R13986 VDD.t1419 VDD.t2723 142.668
R13987 VDD.t2745 VDD.t2197 142.668
R13988 VDD.t2229 VDD.t1641 142.668
R13989 VDD.t507 VDD.t1650 142.668
R13990 VDD.t485 VDD.t477 142.668
R13991 VDD.t15 VDD.t9 142.668
R13992 VDD.t1700 VDD.t621 142.668
R13993 VDD.t3566 VDD.t1515 142.668
R13994 VDD.t3507 VDD.t3250 142.668
R13995 VDD.t2034 VDD.t1236 142.668
R13996 VDD.t3027 VDD.t716 142.668
R13997 VDD.t3514 VDD.t2088 142.668
R13998 VDD.t1308 VDD.t997 142.668
R13999 VDD.t944 VDD.t946 140.989
R14000 VDD.t1682 VDD.t1680 140.989
R14001 VDD.t2267 VDD.t2269 140.989
R14002 VDD.t1265 VDD.t1267 140.989
R14003 VDD.t1511 VDD.t1351 140.989
R14004 VDD.t1196 VDD.t3151 140.989
R14005 VDD.t1594 VDD.t1545 140.989
R14006 VDD.t3667 VDD.t2376 140.989
R14007 VDD.t455 VDD.t457 140.989
R14008 VDD.t2948 VDD.t2937 140.989
R14009 VDD.t3178 VDD.t3188 140.989
R14010 VDD.t3188 VDD.t2934 140.989
R14011 VDD.t3202 VDD.t3180 140.989
R14012 VDD.t888 VDD.t890 140.989
R14013 VDD.t3414 VDD.t886 140.989
R14014 VDD.t180 VDD.t1720 140.989
R14015 VDD.t1187 VDD.t1185 140.989
R14016 VDD.t810 VDD.t808 140.989
R14017 VDD.t789 VDD.t791 140.989
R14018 VDD.t791 VDD.t793 140.989
R14019 VDD.t793 VDD.t795 140.989
R14020 VDD.t2802 VDD.t1443 140.989
R14021 VDD.t3162 VDD.t711 140.989
R14022 VDD.t2295 VDD.t2513 140.989
R14023 VDD.t1827 VDD.t2653 140.989
R14024 VDD.t1873 VDD.t1799 140.989
R14025 VDD.t2970 VDD.t2157 140.989
R14026 VDD.t3126 VDD.t1091 140.989
R14027 VDD.t2236 VDD.t2238 140.989
R14028 VDD.t2443 VDD.t2441 140.989
R14029 VDD.t2467 VDD.t1592 140.989
R14030 VDD.t1055 VDD.t1685 140.989
R14031 VDD.t942 VDD.t3033 140.989
R14032 VDD.t2728 VDD.t1475 140.989
R14033 VDD.t1785 VDD.t1886 140.989
R14034 VDD.t1171 VDD.t1173 140.989
R14035 VDD.t3328 VDD.t3330 140.989
R14036 VDD.t845 VDD.t843 140.989
R14037 VDD.t575 VDD.t573 140.989
R14038 VDD.t475 VDD.t473 140.989
R14039 VDD.t1332 VDD.t1330 140.989
R14040 VDD.t1735 VDD.t3361 140.989
R14041 VDD.t1737 VDD.t2610 140.989
R14042 VDD.t767 VDD.t2301 140.989
R14043 VDD.t2485 VDD.t2487 140.989
R14044 VDD.t1624 VDD.t3157 140.989
R14045 VDD.t3196 VDD.t1745 140.989
R14046 VDD.t3276 VDD.t3272 140.989
R14047 VDD.t960 VDD.t3298 140.989
R14048 VDD.t3130 VDD.t2751 140.989
R14049 VDD.t929 VDD.t470 140.989
R14050 VDD.t1787 VDD.t1498 140.989
R14051 VDD.t2388 VDD.t1893 140.989
R14052 VDD.t2692 VDD.t2694 140.989
R14053 VDD.t319 VDD.t1781 140.989
R14054 VDD.t3684 VDD.t3691 140.989
R14055 VDD.t1455 VDD.t3395 140.989
R14056 VDD.t1586 VDD.t3743 140.989
R14057 VDD.t1730 VDD.t1732 140.989
R14058 VDD.t1407 VDD.t1405 140.989
R14059 VDD.t395 VDD.t393 140.989
R14060 VDD.t1228 VDD.t1226 140.989
R14061 VDD.t3149 VDD.t3136 140.989
R14062 VDD.t1647 VDD.t3140 140.989
R14063 VDD.t2702 VDD.t3426 140.989
R14064 VDD.t3200 VDD.t2930 140.989
R14065 VDD.t2198 VDD.t987 140.989
R14066 VDD.t3111 VDD.t1000 140.989
R14067 VDD.t805 VDD.t2843 140.989
R14068 VDD.t2845 VDD.t2838 140.989
R14069 VDD.t345 VDD.t1975 140.989
R14070 VDD.t1749 VDD.t1281 140.989
R14071 VDD.t3627 VDD.t3636 140.989
R14072 VDD.t3647 VDD.t2350 140.989
R14073 VDD.t3607 VDD.t3042 140.989
R14074 VDD.t2834 VDD.t1409 140.989
R14075 VDD.t511 VDD.t509 140.989
R14076 VDD.t1865 VDD.t309 140.989
R14077 VDD.t3606 VDD.t3044 140.989
R14078 VDD.t1505 VDD.t1480 140.989
R14079 VDD.t2898 VDD.t1111 140.989
R14080 VDD.t852 VDD.t2261 140.989
R14081 VDD.t2261 VDD.t1819 140.989
R14082 VDD.t1314 VDD.t1312 140.989
R14083 VDD.t2905 VDD.t2259 140.989
R14084 VDD.t317 VDD.t321 140.989
R14085 VDD.t2103 VDD.t2530 140.989
R14086 VDD.t1795 VDD.t1249 140.989
R14087 VDD.t1177 VDD.t2492 140.989
R14088 VDD.t1318 VDD.t3749 140.989
R14089 VDD.t1159 VDD.t1157 140.989
R14090 VDD.t257 VDD.t259 140.989
R14091 VDD.t1169 VDD.t1167 140.989
R14092 VDD.t1274 VDD.t1276 140.989
R14093 VDD.t2141 VDD.t2143 140.989
R14094 VDD.t950 VDD.t948 140.989
R14095 VDD.t3082 VDD.t3084 140.989
R14096 VDD.t3118 VDD.t3339 140.989
R14097 VDD.t714 VDD.t869 140.989
R14098 VDD.t305 VDD.t301 140.989
R14099 VDD.t301 VDD.t303 140.989
R14100 VDD.t2646 VDD.t3404 140.989
R14101 VDD.t299 VDD.t989 140.989
R14102 VDD.t807 VDD.t649 140.989
R14103 VDD.t2863 VDD.t1389 140.989
R14104 VDD.t803 VDD.t731 140.989
R14105 VDD.t1450 VDD.t1643 140.989
R14106 VDD.t3278 VDD.t3320 140.989
R14107 VDD.t523 VDD.t2749 140.989
R14108 VDD.t1145 VDD.t1257 140.989
R14109 VDD.t1257 VDD.t1867 140.989
R14110 VDD.t1258 VDD.t307 140.989
R14111 VDD.t1807 VDD.t2721 140.989
R14112 VDD.t758 VDD.t3284 140.989
R14113 VDD.t896 VDD.t894 140.989
R14114 VDD.t1813 VDD.t2911 140.989
R14115 VDD.t521 VDD.t1101 140.989
R14116 VDD.t857 VDD.t855 140.989
R14117 VDD.t859 VDD.t861 140.989
R14118 VDD.t2436 VDD.t3097 140.989
R14119 VDD.t2794 VDD.t3492 140.989
R14120 VDD.t1500 VDD.t1556 140.989
R14121 VDD.t2916 VDD.t2909 140.989
R14122 VDD.t2712 VDD.t1425 140.989
R14123 VDD.t2801 VDD.t2250 140.989
R14124 VDD.t2250 VDD.t2138 140.989
R14125 VDD.t3246 VDD.t828 140.989
R14126 VDD.t654 VDD.t2493 140.989
R14127 VDD.t1123 VDD.t1125 140.989
R14128 VDD.t545 VDD.t553 140.989
R14129 VDD.t547 VDD.t541 140.989
R14130 VDD.t2329 VDD.t3381 140.989
R14131 VDD.t2739 VDD.t2328 140.989
R14132 VDD.t2688 VDD.t3741 140.989
R14133 VDD.t2215 VDD.t2213 140.989
R14134 VDD.t289 VDD.t287 140.989
R14135 VDD.t1529 VDD.t3516 140.989
R14136 VDD.t2808 VDD.t2806 140.989
R14137 VDD.t1728 VDD.t1726 140.989
R14138 VDD.t261 VDD.t263 140.989
R14139 VDD.t3659 VDD.t999 140.989
R14140 VDD.t559 VDD.t557 140.989
R14141 VDD.t1634 VDD.t1630 140.989
R14142 VDD.t1632 VDD.t1634 140.989
R14143 VDD.t2770 VDD.t2768 140.989
R14144 VDD.t2598 VDD.t2594 140.989
R14145 VDD.t2594 VDD.t2592 140.989
R14146 VDD.t1670 VDD.t1847 140.989
R14147 VDD.t1271 VDD.t2339 140.989
R14148 VDD.t2339 VDD.t3302 140.989
R14149 VDD.t1668 VDD.t3138 140.989
R14150 VDD.t2697 VDD.t3011 140.989
R14151 VDD.t515 VDD.t1895 140.989
R14152 VDD.t1463 VDD.t1459 140.989
R14153 VDD.t1457 VDD.t1465 140.989
R14154 VDD.t1461 VDD.t1678 140.989
R14155 VDD.t1675 VDD.t3128 140.989
R14156 VDD.t912 VDD.t910 140.989
R14157 VDD.t1898 VDD.t1877 140.989
R14158 VDD.t2859 VDD.t2857 140.989
R14159 VDD.t1901 VDD.t1717 140.989
R14160 VDD.t2298 VDD.t2793 140.989
R14161 VDD.t1558 VDD.t2306 140.989
R14162 VDD.t2587 VDD.t924 140.989
R14163 VDD.t3529 VDD.t3552 140.989
R14164 VDD.t3466 VDD.t3470 140.989
R14165 VDD.t3454 VDD.t2851 140.989
R14166 VDD.t976 VDD.t2500 140.989
R14167 VDD.t273 VDD.t271 140.989
R14168 VDD.t3722 VDD.t3707 140.989
R14169 VDD.t981 VDD.t983 140.989
R14170 VDD.t1904 VDD.t3711 140.989
R14171 VDD.t1905 VDD.t3450 140.989
R14172 VDD.t2447 VDD.t2449 140.989
R14173 VDD.t927 VDD.t925 140.989
R14174 VDD.t1044 VDD.t1046 140.989
R14175 VDD.t1050 VDD.t1044 140.989
R14176 VDD.t1048 VDD.t1050 140.989
R14177 VDD.t717 VDD.t721 140.989
R14178 VDD.t719 VDD.t717 140.989
R14179 VDD.t401 VDD.t403 140.989
R14180 VDD.t397 VDD.t401 140.989
R14181 VDD.t399 VDD.t397 140.989
R14182 VDD.t878 VDD.t882 140.989
R14183 VDD.t880 VDD.t878 140.989
R14184 VDD.t884 VDD.t880 140.989
R14185 VDD.t702 VDD.t704 140.989
R14186 VDD.t706 VDD.t702 140.989
R14187 VDD.t708 VDD.t706 140.989
R14188 VDD.t283 VDD.t281 140.989
R14189 VDD.t279 VDD.t283 140.989
R14190 VDD.t285 VDD.t279 140.989
R14191 VDD.t2282 VDD.t662 140.989
R14192 VDD.t1937 VDD.t1610 140.989
R14193 VDD.t1664 VDD.t1662 140.989
R14194 VDD.t1662 VDD.t1660 140.989
R14195 VDD.t3061 VDD.t3068 140.989
R14196 VDD.t3068 VDD.t3064 140.989
R14197 VDD.t3055 VDD.t3066 140.989
R14198 VDD.t3057 VDD.t3055 140.989
R14199 VDD.t2405 VDD.t2409 140.989
R14200 VDD.t2403 VDD.t2405 140.989
R14201 VDD.n319 VDD.n318 140.702
R14202 VDD.n320 VDD.n319 140.048
R14203 VDD.t536 VDD.t3170 139.311
R14204 VDD.t1645 VDD.t1724 139.311
R14205 VDD.t1869 VDD.t1579 139.311
R14206 VDD.t952 VDD.t1278 139.311
R14207 VDD.t2231 VDD.t236 139.311
R14208 VDD.t2 VDD.t956 139.311
R14209 VDD.t2335 VDD.t1026 139.311
R14210 VDD.t2534 VDD.t629 139.311
R14211 VDD.t3441 VDD.t773 139.311
R14212 VDD.t1322 VDD.t311 139.311
R14213 VDD.n1766 VDD.n1651 138.415
R14214 VDD.t1537 VDD.t871 137.633
R14215 VDD.t2799 VDD.t664 137.633
R14216 VDD.t3666 VDD.t1247 137.633
R14217 VDD.t1069 VDD.t3412 137.633
R14218 VDD.t3501 VDD.t3632 137.633
R14219 VDD.t1569 VDD.t2221 137.633
R14220 VDD.t2292 VDD.t2225 137.633
R14221 VDD.t1797 VDD.t3259 137.633
R14222 VDD.t2717 VDD.t648 137.633
R14223 VDD.t1448 VDD.t1364 137.633
R14224 VDD.t861 VDD.t2820 137.633
R14225 VDD.t653 VDD.t2371 137.633
R14226 VDD.n2667 VDD.t2164 137.095
R14227 VDD.n1670 VDD.t2420 137.095
R14228 VDD.n2430 VDD.t2426 137.079
R14229 VDD.n2441 VDD.t2615 137.079
R14230 VDD.t3499 VDD.t2210 135.954
R14231 VDD.t2384 VDD.t2122 135.954
R14232 VDD.t2714 VDD.t2628 135.954
R14233 VDD.t0 VDD.t2830 135.954
R14234 VDD.t854 VDD.t1115 135.954
R14235 VDD.t1861 VDD.t1849 134.276
R14236 VDD.t2255 VDD.t98 134.276
R14237 VDD.t1413 VDD.t2340 134.276
R14238 VDD.t3155 VDD.t2378 134.276
R14239 VDD.t1075 VDD.t3505 134.276
R14240 VDD.n3468 VDD.t995 134.276
R14241 VDD.t836 VDD.t3318 134.276
R14242 VDD.t3726 VDD.t3548 134.276
R14243 VDD.t7 VDD.t700 134.276
R14244 VDD.t3294 VDD.t253 134.276
R14245 VDD.n2029 VDD.t1604 134.276
R14246 VDD.t2506 VDD.t1906 134.276
R14247 VDD.t1285 VDD.t451 134.276
R14248 VDD.t3470 VDD.t3616 134.276
R14249 VDD.n3233 VDD.t2952 133.571
R14250 VDD.n3233 VDD.t3313 133.571
R14251 VDD.n3242 VDD.t2942 133.571
R14252 VDD.n3242 VDD.t3319 133.571
R14253 VDD.t461 VDD.t3159 132.597
R14254 VDD.t2191 VDD.t906 132.597
R14255 VDD.t2611 VDD.t769 132.597
R14256 VDD.t2816 VDD.t1089 132.597
R14257 VDD.n3866 VDD.t1455 132.597
R14258 VDD.n2727 VDD.t1370 132.597
R14259 VDD.t670 VDD.t1929 132.597
R14260 VDD.n3064 VDD.t37 132.597
R14261 VDD.t2491 VDD.t3091 132.597
R14262 VDD.t613 VDD.t2932 132.597
R14263 VDD.t3324 VDD.t3269 132.597
R14264 VDD.t2990 VDD.t692 132.597
R14265 VDD.n1405 VDD.t1326 132.597
R14266 VDD.n243 VDD.n224 131.388
R14267 VDD.n237 VDD.n224 131.388
R14268 VDD.t1596 VDD.t3192 130.919
R14269 VDD.t2606 VDD.t2783 130.919
R14270 VDD.t1346 VDD.t1693 130.919
R14271 VDD.t933 VDD.t2013 130.919
R14272 VDD.t3640 VDD.t2090 130.919
R14273 VDD.t265 VDD.t3698 130.919
R14274 VDD.t1973 VDD.t505 130.919
R14275 VDD.t3045 VDD.t497 130.919
R14276 VDD.t23 VDD.t3439 130.919
R14277 VDD.t3458 VDD.t1037 130.919
R14278 VDD.t3134 VDD.t1310 130.919
R14279 VDD.n165 VDD.t1242 130.65
R14280 VDD.n353 VDD.n352 129.506
R14281 VDD.n4382 VDD.t3804 129.344
R14282 VDD.n3203 VDD.t3788 129.344
R14283 VDD.n2557 VDD.t3771 129.344
R14284 VDD.t2288 VDD.t134 129.24
R14285 VDD.t1582 VDD.t1789 129.24
R14286 VDD.t3235 VDD.t1213 129.24
R14287 VDD.t2951 VDD.t3503 129.24
R14288 VDD.t3435 VDD.t53 129.24
R14289 VDD.t2352 VDD.t119 129.24
R14290 VDD.t3206 VDD.t49 129.24
R14291 VDD.t3533 VDD.t443 129.24
R14292 VDD.t1131 VDD.t419 127.562
R14293 VDD.n3865 VDD.t1872 127.562
R14294 VDD.t1417 VDD.t3712 127.562
R14295 VDD.t2453 VDD.t1927 127.562
R14296 VDD.t3675 VDD.t2658 127.562
R14297 VDD.t1113 VDD.t2898 127.562
R14298 VDD.t2280 VDD.t1107 127.562
R14299 VDD.t3332 VDD.t1238 127.562
R14300 VDD.t2508 VDD.t572 127.562
R14301 VDD.n1201 VDD.t1457 127.562
R14302 VDD.t696 VDD.t269 127.562
R14303 VDD.t1654 VDD.t3070 127.562
R14304 VDD.t2193 VDD.t3059 127.562
R14305 VDD.t3595 VDD.t3582 127.291
R14306 VDD.t3582 VDD.t3584 127.291
R14307 VDD.t3584 VDD.t3580 127.291
R14308 VDD.t3580 VDD.t3602 127.291
R14309 VDD.t3602 VDD.t3590 127.291
R14310 VDD.t3576 VDD.t3590 127.291
R14311 VDD.t3586 VDD.t3576 127.291
R14312 VDD.t3600 VDD.t3586 127.291
R14313 VDD.t3578 VDD.t3600 127.291
R14314 VDD.t3598 VDD.t3588 127.291
R14315 VDD.t3588 VDD.t3592 127.291
R14316 VDD.t3257 VDD.t1672 125.883
R14317 VDD.t3503 VDD.t3312 125.883
R14318 VDD.t477 VDD.n2894 125.883
R14319 VDD.n2896 VDD.t1016 125.883
R14320 VDD.t645 VDD.t2634 125.883
R14321 VDD.t2145 VDD.t859 125.883
R14322 VDD.t2327 VDD.t3745 125.883
R14323 VDD.t698 VDD.t47 125.883
R14324 VDD.t2302 VDD.t2344 124.206
R14325 VDD.t1067 VDD.t2483 124.206
R14326 VDD.t2706 VDD.t3023 124.206
R14327 VDD.t3563 VDD.t516 124.206
R14328 VDD.t1336 VDD.t423 124.206
R14329 VDD.t383 VDD.t15 124.206
R14330 VDD.t3300 VDD.t2867 124.206
R14331 VDD.t2625 VDD.t3270 124.206
R14332 VDD.t447 VDD.t2421 124.206
R14333 VDD.t1122 VDD.t1307 124.206
R14334 VDD.t2773 VDD.t898 124.206
R14335 VDD.t2682 VDD.t353 124.206
R14336 VDD.t2684 VDD.t355 124.206
R14337 VDD.t2680 VDD.t351 124.206
R14338 VDD.t2686 VDD.t357 124.206
R14339 VDD.n4513 VDD.t1932 123.507
R14340 VDD.n4084 VDD.t2621 123.507
R14341 VDD.n4279 VDD.t657 123.507
R14342 VDD.n3809 VDD.t378 123.507
R14343 VDD.n3103 VDD.t3513 123.507
R14344 VDD.n2285 VDD.t3653 123.507
R14345 VDD.n2675 VDD.t1293 123.507
R14346 VDD.n3904 VDD.t1910 123.507
R14347 VDD.n4590 VDD.t1924 123.507
R14348 VDD.n3993 VDD.t2609 123.507
R14349 VDD.n4012 VDD.t2020 123.507
R14350 VDD.n3701 VDD.t360 123.507
R14351 VDD.n3684 VDD.t2008 123.507
R14352 VDD.n3205 VDD.t1142 123.507
R14353 VDD.n3587 VDD.t1702 123.507
R14354 VDD.n3573 VDD.t2707 123.507
R14355 VDD.n3296 VDD.t2064 123.507
R14356 VDD.n3825 VDD.t1420 123.507
R14357 VDD.n2846 VDD.t2336 123.507
R14358 VDD.n2455 VDD.t1299 123.507
R14359 VDD.n733 VDD.t3534 123.507
R14360 VDD.t2463 VDD.n3467 122.526
R14361 VDD.t1399 VDD.t2345 122.526
R14362 VDD.t849 VDD.t2854 122.526
R14363 VDD.t441 VDD.t435 122.526
R14364 VDD.t2899 VDD.t3456 122.526
R14365 VDD.t633 VDD.t1598 122.526
R14366 VDD.t744 VDD.t2757 122.526
R14367 VDD.t754 VDD.t1688 122.526
R14368 VDD.n1631 VDD.t1700 122.526
R14369 VDD.t2332 VDD.t51 122.526
R14370 VDD.t3523 VDD.t826 122.526
R14371 VDD.t902 VDD.t1445 122.526
R14372 VDD.t1847 VDD.t1896 122.526
R14373 VDD.t2056 VDD.n375 121.245
R14374 VDD.t2056 VDD.n368 121.245
R14375 VDD.t2051 VDD.n368 121.245
R14376 VDD.t2051 VDD.n362 121.245
R14377 VDD.t2944 VDD.n362 121.245
R14378 VDD.n414 VDD.t2944 121.245
R14379 VDD.n414 VDD.t2054 121.245
R14380 VDD.n421 VDD.t2054 121.245
R14381 VDD.t1486 VDD.t2265 120.849
R14382 VDD.t775 VDD.t2529 120.849
R14383 VDD.t567 VDD.t323 120.849
R14384 VDD.t2509 VDD.t1479 120.849
R14385 VDD.t1751 VDD.t1054 120.849
R14386 VDD.t2941 VDD.t836 120.849
R14387 VDD.t1747 VDD.t3641 120.849
R14388 VDD.t3562 VDD.t343 120.849
R14389 VDD.t1565 VDD.t1504 120.849
R14390 VDD.t3483 VDD.t2729 120.849
R14391 VDD.t3258 VDD.t341 120.849
R14392 VDD.t1127 VDD.t3241 120.849
R14393 VDD.t3008 VDD.t1421 120.849
R14394 VDD.t3252 VDD.t2880 120.849
R14395 VDD.t3733 VDD.t1309 120.849
R14396 VDD.t3090 VDD.t867 120.849
R14397 VDD.t2368 VDD.t244 120.849
R14398 VDD.t244 VDD.t2787 120.849
R14399 VDD.t2853 VDD.t2504 120.849
R14400 VDD.t2715 VDD.t647 120.849
R14401 VDD.t3112 VDD.t3047 120.849
R14402 VDD.t487 VDD.t2279 120.849
R14403 VDD.t1959 VDD.t2004 120.849
R14404 VDD.t3565 VDD.t529 120.849
R14405 VDD.t2913 VDD.t2 120.849
R14406 VDD.t686 VDD.t326 120.849
R14407 VDD.t2775 VDD.t35 120.849
R14408 VDD.t379 VDD.t27 120.849
R14409 VDD.t1251 VDD.t974 120.849
R14410 VDD.t3190 VDD.t2950 120.849
R14411 VDD.t991 VDD.t619 120.849
R14412 VDD.t3539 VDD.t1306 120.849
R14413 VDD.t3389 VDD.t2690 120.849
R14414 VDD.t835 VDD.t1991 120.849
R14415 VDD.t2219 VDD.t3732 120.849
R14416 VDD.t3420 VDD.t2181 120.849
R14417 VDD.t2600 VDD.t3017 120.849
R14418 VDD.t2321 VDD.t453 120.849
R14419 VDD.t2959 VDD.t2903 120.849
R14420 VDD.t3716 VDD.t2969 120.849
R14421 VDD.t977 VDD.t2501 120.849
R14422 VDD.t785 VDD.t2765 120.849
R14423 VDD.t590 VDD.t2994 120.849
R14424 VDD.t1876 VDD.t2922 120.849
R14425 VDD.t3093 VDD.t2891 120.849
R14426 VDD.t2877 VDD.t2036 120.849
R14427 VDD.t1962 VDD.t2023 120.849
R14428 VDD.t1761 VDD.t2027 120.849
R14429 VDD.t1772 VDD.t2887 120.849
R14430 VDD.n4603 VDD.t1476 119.608
R14431 VDD.n4000 VDD.t1056 119.608
R14432 VDD.n4028 VDD.t1495 119.608
R14433 VDD.n4439 VDD.t905 119.608
R14434 VDD.n4045 VDD.t2514 119.608
R14435 VDD.n4076 VDD.t2803 119.608
R14436 VDD.n4272 VDD.t893 119.608
R14437 VDD.n4138 VDD.t1512 119.608
R14438 VDD.n3687 VDD.t930 119.608
R14439 VDD.n3260 VDD.t800 119.608
R14440 VDD.n3283 VDD.t2349 119.608
R14441 VDD.n3454 VDD.t2385 119.608
R14442 VDD.n3387 VDD.t768 119.608
R14443 VDD.n3358 VDD.t1738 119.608
R14444 VDD.n3109 VDD.t2454 119.608
R14445 VDD.n2524 VDD.t2674 119.608
R14446 VDD.n2294 VDD.t1178 119.608
R14447 VDD.n2479 VDD.t988 119.608
R14448 VDD.n1978 VDD.t864 119.608
R14449 VDD.n1633 VDD.t300 119.608
R14450 VDD.n2173 VDD.t548 119.608
R14451 VDD.n2178 VDD.t2740 119.608
R14452 VDD.n804 VDD.t2597 119.608
R14453 VDD.n1019 VDD.t1629 119.608
R14454 VDD.n838 VDD.t2137 119.608
R14455 VDD.n781 VDD.t1462 119.608
R14456 VDD.n1143 VDD.t921 119.608
R14457 VDD.n1406 VDD.t821 119.608
R14458 VDD.t2124 VDD.t2251 119.171
R14459 VDD.t2653 VDD.t1873 119.171
R14460 VDD.t2060 VDD.t2476 119.171
R14461 VDD.t1328 VDD.t305 119.171
R14462 VDD.n2172 VDD.t3399 119.171
R14463 VDD.t2583 VDD.t1897 119.171
R14464 VDD.t968 VDD.t1155 119.171
R14465 VDD.t2235 VDD.t3375 119.171
R14466 VDD.n4443 VDD.t3798 118.853
R14467 VDD.n4048 VDD.t3823 118.853
R14468 VDD.n3969 VDD.t3790 118.853
R14469 VDD.n3308 VDD.t3820 118.853
R14470 VDD.n2297 VDD.t3779 118.853
R14471 VDD.n645 VDD.n644 118.316
R14472 VDD.t2001 VDD.t2102 118.267
R14473 VDD.t3604 VDD.t2921 118.267
R14474 VDD.t3416 VDD.t3418 117.492
R14475 VDD.t1701 VDD.t2665 117.492
R14476 VDD.t3763 VDD.t373 117.492
R14477 VDD.t1543 VDD.t2656 117.492
R14478 VDD.t1003 VDD.t3643 117.492
R14479 VDD.t3664 VDD.t3025 117.492
R14480 VDD.t3105 VDD.t847 117.492
R14481 VDD.t3758 VDD.t804 117.492
R14482 VDD.t1289 VDD.t1298 117.492
R14483 VDD.t830 VDD.t3013 117.492
R14484 VDD.t611 VDD.t3718 117.492
R14485 VDD.t1556 VDD.t1149 117.492
R14486 VDD.t1304 VDD.t2140 117.492
R14487 VDD.t1397 VDD.t2557 117.492
R14488 VDD.t2967 VDD.t1555 117.492
R14489 VDD.n1963 VDD.t1926 117.451
R14490 VDD.n1602 VDD.t2868 117.451
R14491 VDD.n1871 VDD.t3281 117.451
R14492 VDD.n4214 VDD.t3775 117.294
R14493 VDD.n3162 VDD.t3809 117.294
R14494 VDD.n1916 VDD.t3812 117.294
R14495 VDD.t2102 VDD.t2893 116.82
R14496 VDD.t2893 VDD.t2033 116.82
R14497 VDD.t2033 VDD.t3702 116.82
R14498 VDD.t3702 VDD.t3663 116.82
R14499 VDD.t3663 VDD.t3547 116.82
R14500 VDD.t3761 VDD.t2955 116.82
R14501 VDD.t3766 VDD.t3761 116.82
R14502 VDD.t3096 VDD.t3766 116.82
R14503 VDD.t3231 VDD.t3096 116.82
R14504 VDD.t2921 VDD.t3231 116.82
R14505 VDD.n3910 VDD.t1786 116.341
R14506 VDD.n4449 VDD.t1784 116.341
R14507 VDD.n4042 VDD.t1800 116.341
R14508 VDD.n4053 VDD.t1790 116.341
R14509 VDD.n4358 VDD.t3089 116.341
R14510 VDD.n3697 VDD.t1788 116.341
R14511 VDD.n3192 VDD.t1782 116.341
R14512 VDD.n2908 VDD.t1792 116.341
R14513 VDD.n2288 VDD.t1796 116.341
R14514 VDD.n2491 VDD.t2931 116.341
R14515 VDD.n2137 VDD.t1254 116.341
R14516 VDD.n887 VDD.t1534 116.341
R14517 VDD.n938 VDD.t3517 116.341
R14518 VDD.t2128 VDD.t2253 115.814
R14519 VDD.t2294 VDD.t3751 115.814
R14520 VDD.t2002 VDD.t2974 115.814
R14521 VDD.t1967 VDD.t564 115.814
R14522 VDD.t668 VDD.t439 115.814
R14523 VDD.t3399 VDD.t2737 115.814
R14524 VDD.t1439 VDD.t255 115.814
R14525 VDD.t2481 VDD.t2652 115.814
R14526 VDD.n237 VDD.n236 115.201
R14527 VDD.n238 VDD.n237 115.201
R14528 VDD.n113 VDD.n102 115.201
R14529 VDD.t3383 VDD.t1340 114.135
R14530 VDD.t1781 VDD.t759 114.135
R14531 VDD.t2459 VDD.t3638 114.135
R14532 VDD.t2896 VDD.t562 114.135
R14533 VDD.t1699 VDD.t609 114.135
R14534 VDD.t277 VDD.t3620 114.135
R14535 VDD.t1109 VDD.t308 114.135
R14536 VDD.t1636 VDD.t2884 114.135
R14537 VDD.n323 VDD.n322 113.448
R14538 VDD.t2358 VDD.t1471 112.457
R14539 VDD.t2386 VDD.t2463 112.457
R14540 VDD.t1272 VDD.t1008 112.457
R14541 VDD.t3724 VDD.t1531 112.457
R14542 VDD.t1117 VDD.t1743 112.457
R14543 VDD.t1321 VDD.t2498 112.457
R14544 VDD.t2175 VDD.t3184 110.778
R14545 VDD.t3359 VDD.t656 110.778
R14546 VDD.t3198 VDD.t3088 110.778
R14547 VDD.t2886 VDD.t2841 110.778
R14548 VDD.t2238 VDD.t2840 110.778
R14549 VDD.t1221 VDD.t1338 110.778
R14550 VDD.t3497 VDD.t1785 110.778
R14551 VDD.t2427 VDD.t2781 110.778
R14552 VDD.t2930 VDD.t1487 110.778
R14553 VDD.t491 VDD.t874 110.778
R14554 VDD.t1882 VDD.t1028 110.778
R14555 VDD.t3677 VDD.t1764 110.778
R14556 VDD.t3306 VDD.t518 110.778
R14557 VDD.t2642 VDD.t545 110.778
R14558 VDD.t2421 VDD.t1603 110.778
R14559 VDD.t1851 VDD.t2943 109.1
R14560 VDD.t151 VDD.t713 109.1
R14561 VDD.t2303 VDD.t2473 109.1
R14562 VDD.t3424 VDD.t3164 109.1
R14563 VDD.t291 VDD.t3622 109.1
R14564 VDD.t1016 VDD.t3493 109.1
R14565 VDD.t2480 VDD.t3657 109.1
R14566 VDD.t1628 VDD.t832 109.1
R14567 VDD.t230 VDD.t185 108.832
R14568 VDD.t150 VDD.t196 108.832
R14569 VDD.t224 VDD.t143 108.832
R14570 VDD.t97 VDD.t133 108.832
R14571 VDD.n170 VDD.n101 108.8
R14572 VDD.n169 VDD.n102 108.8
R14573 VDD.n114 VDD.n103 108.8
R14574 VDD.t3822 VDD.n645 107.793
R14575 VDD.t1768 VDD.t1881 107.421
R14576 VDD.t795 VDD.t2527 107.421
R14577 VDD.t323 VDD.t2236 107.421
R14578 VDD.t1626 VDD.t1447 107.421
R14579 VDD.t1489 VDD.t471 107.421
R14580 VDD.t2588 VDD.t824 107.421
R14581 VDD.t2416 VDD.t2149 107.421
R14582 VDD.t2369 VDD.t2198 107.421
R14583 VDD.t2264 VDD.t3444 107.421
R14584 VDD.t1925 VDD.t1103 107.421
R14585 VDD.t1630 VDD.t729 107.421
R14586 VDD.t2592 VDD.t1652 107.421
R14587 VDD.t3325 VDD.t2413 107.421
R14588 VDD.t3437 VDD.t3529 107.421
R14589 VDD.n1404 VDD.n1403 106.561
R14590 VDD.n4652 VDD.n4651 106.559
R14591 VDD.n4547 VDD.n4010 106.559
R14592 VDD.n4502 VDD.n4501 106.559
R14593 VDD.n4343 VDD.n4342 106.559
R14594 VDD.n4151 VDD.n4123 106.559
R14595 VDD.n1200 VDD.n760 106.559
R14596 VDD.n1199 VDD.n1198 106.559
R14597 VDD.n1078 VDD.n1077 106.559
R14598 VDD.n951 VDD.n950 106.559
R14599 VDD.t3484 VDD.t3754 105.743
R14600 VDD.t1829 VDD.t3756 105.743
R14601 VDD.t1686 VDD.t1617 105.743
R14602 VDD.t3379 VDD.t1619 105.743
R14603 VDD.t2354 VDD.t1467 105.743
R14604 VDD.t2356 VDD.t3387 105.743
R14605 VDD.t3353 VDD.t1083 105.743
R14606 VDD.t1348 VDD.t1885 105.743
R14607 VDD.t3680 VDD.t2997 105.743
R14608 VDD.t2505 VDD.t3671 105.743
R14609 VDD.n595 VDD.n556 104.684
R14610 VDD.n515 VDD.n476 104.684
R14611 VDD.t2529 VDD.t409 104.064
R14612 VDD.t371 VDD.t2471 104.064
R14613 VDD.t1649 VDD.t2151 104.064
R14614 VDD.t850 VDD.t3351 104.064
R14615 VDD.t2205 VDD.t479 104.064
R14616 VDD.t1022 VDD.t2679 104.064
R14617 VDD.t2699 VDD.t2411 104.064
R14618 VDD.t1678 VDD.t1403 104.064
R14619 VDD.t1326 VDD.t2553 104.064
R14620 VDD.t3373 VDD.t2555 104.064
R14621 VDD.n4069 VDD.t1444 102.385
R14622 VDD.t2818 VDD.t1085 102.385
R14623 VDD.t1089 VDD.t535 102.385
R14624 VDD.t994 VDD.t3304 102.385
R14625 VDD.t2704 VDD.t1875 102.385
R14626 VDD.n3754 VDD.t469 102.385
R14627 VDD.t1370 VDD.t533 102.385
R14628 VDD.t650 VDD.t2715 102.385
R14629 VDD.t623 VDD.t3 102.385
R14630 VDD.t2132 VDD.t2177 102.385
R14631 VDD.t3015 VDD.t1119 102.385
R14632 VDD.t1799 VDD.t2511 100.707
R14633 VDD.t995 VDD.t2485 100.707
R14634 VDD.t2810 VDD.t2457 100.707
R14635 VDD.t979 VDD.t1431 100.707
R14636 VDD.t3369 VDD.t2577 100.707
R14637 VDD.t1533 VDD.t2865 100.707
R14638 VDD.t1741 VDD.t2626 100.707
R14639 VDD.t916 VDD.t2581 100.707
R14640 VDD.t1674 VDD.t1401 100.707
R14641 VDD.t2793 VDD.t1558 100.707
R14642 VDD.t3526 VDD.t1979 100.707
R14643 VDD.t1451 VDD.t814 100.707
R14644 VDD.t2464 VDD.t2384 99.0288
R14645 VDD.t391 VDD.t1820 99.0288
R14646 VDD.t1269 VDD.t3253 99.0288
R14647 VDD.t1679 VDD.t1805 99.0288
R14648 VDD.t721 VDD.t130 99.0288
R14649 VDD.n3775 VDD.t432 98.5005
R14650 VDD.n2834 VDD.t971 98.5005
R14651 VDD.n2621 VDD.t3187 98.5005
R14652 VDD.n2483 VDD.t3676 98.5005
R14653 VDD.n2655 VDD.t1958 98.5005
R14654 VDD.n2122 VDD.t3551 98.5005
R14655 VDD.n293 VDD.t3595 97.4361
R14656 VDD.t2999 VDD.t3739 97.3503
R14657 VDD.t3737 VDD.t1252 97.3503
R14658 VDD.t1492 VDD.t1141 97.3503
R14659 VDD.t1010 VDD.t2333 97.3503
R14660 VDD.t3710 VDD.t3654 97.3503
R14661 VDD.t2391 VDD.t935 97.2286
R14662 VDD.t1242 VDD.t3480 97.2286
R14663 VDD.n3984 VDD.t941 96.1553
R14664 VDD.n4114 VDD.t3104 96.1553
R14665 VDD.n4117 VDD.t1538 96.1553
R14666 VDD.n3264 VDD.t1359 96.1553
R14667 VDD.n2386 VDD.t2018 96.1553
R14668 VDD.n2877 VDD.t965 96.1553
R14669 VDD.n3027 VDD.t382 96.1553
R14670 VDD.n2433 VDD.t2424 96.1553
R14671 VDD.n2443 VDD.t2613 96.1553
R14672 VDD.n2478 VDD.t3674 96.1553
R14673 VDD.n2671 VDD.t1432 96.1553
R14674 VDD.n1540 VDD.t3683 96.1553
R14675 VDD.n1962 VDD.t1104 96.1553
R14676 VDD.n1593 VDD.t3631 96.1553
R14677 VDD.n1667 VDD.t2418 96.1553
R14678 VDD.n2103 VDD.t1305 96.1553
R14679 VDD.n1907 VDD.t3309 96.1553
R14680 VDD.n1569 VDD.t528 96.1553
R14681 VDD.n2132 VDD.t3681 96.1553
R14682 VDD.n801 VDD.t3275 96.1553
R14683 VDD.n822 VDD.t252 96.1553
R14684 VDD.n833 VDD.t1742 96.1553
R14685 VDD.n726 VDD.t699 96.1553
R14686 VDD.n1325 VDD.t3452 96.1553
R14687 VDD.n746 VDD.t2006 96.1553
R14688 VDD.n784 VDD.t1812 96.1553
R14689 VDD.n1364 VDD.t689 96.1553
R14690 VDD.n1365 VDD.t693 96.1553
R14691 VDD.t3547 VDD.n55 95.7389
R14692 VDD.t2955 VDD.n18 95.7389
R14693 VDD.t765 VDD.t3029 95.6719
R14694 VDD.t1129 VDD.t1701 95.6719
R14695 VDD.t647 VDD.t1300 95.6719
R14696 VDD.t680 VDD.t13 95.6719
R14697 VDD.t2519 VDD.t754 95.6719
R14698 VDD.t2273 VDD.t2646 95.6719
R14699 VDD.t3326 VDD.t2964 95.6719
R14700 VDD.n3108 VDD.t3447 95.3969
R14701 VDD.n3819 VDD.t3713 95.3969
R14702 VDD.n2379 VDD.t1912 95.3969
R14703 VDD.n2470 VDD.t239 95.3969
R14704 VDD.n1967 VDD.t1810 95.3969
R14705 VDD.n1581 VDD.t3183 95.3969
R14706 VDD.n318 VDD.n315 95.0755
R14707 VDD.t1195 VDD.t1391 93.9934
R14708 VDD.t1065 VDD.t539 93.9934
R14709 VDD.t867 VDD.t3200 93.9934
R14710 VDD.t1389 VDD.t803 93.9934
R14711 VDD.n2027 VDD.t3284 93.9934
R14712 VDD.t655 VDD.t2139 93.9934
R14713 VDD.t2246 VDD.t2579 93.9934
R14714 VDD.t3472 VDD.n737 93.9934
R14715 VDD.t3552 VDD.t1695 93.9934
R14716 VDD.n4608 VDD.t2258 93.81
R14717 VDD.n4568 VDD.t2326 93.81
R14718 VDD.n4021 VDD.t1192 93.81
R14719 VDD.n4476 VDD.t414 93.81
R14720 VDD.n4049 VDD.t276 93.81
R14721 VDD.n4071 VDD.t1430 93.81
R14722 VDD.n4278 VDD.t2276 93.81
R14723 VDD.n4130 VDD.t2564 93.81
R14724 VDD.n3747 VDD.t2734 93.81
R14725 VDD.n3527 VDD.t2156 93.81
R14726 VDD.n3276 VDD.t2817 93.81
R14727 VDD.n3400 VDD.t1564 93.81
R14728 VDD.n3395 VDD.t2123 93.81
R14729 VDD.n3299 VDD.t1248 93.81
R14730 VDD.n3115 VDD.t2711 93.81
R14731 VDD.n2509 VDD.t2605 93.81
R14732 VDD.n2628 VDD.t2202 93.81
R14733 VDD.n2299 VDD.t332 93.81
R14734 VDD.n1555 VDD.t1607 93.81
R14735 VDD.n1613 VDD.t3719 93.81
R14736 VDD.n1810 VDD.t2645 93.81
R14737 VDD.n2014 VDD.t2987 93.81
R14738 VDD.n2181 VDD.t448 93.81
R14739 VDD.n2184 VDD.t1454 93.81
R14740 VDD.n800 VDD.t1526 93.81
R14741 VDD.n1051 VDD.t2815 93.81
R14742 VDD.n834 VDD.t2627 93.81
R14743 VDD.n776 VDD.t2249 93.81
R14744 VDD.n1137 VDD.t2338 93.81
R14745 VDD.n1413 VDD.t1325 93.81
R14746 VDD.n381 VDD.n373 93.7417
R14747 VDD.n418 VDD.n358 93.7417
R14748 VDD.n382 VDD.n381 93.7417
R14749 VDD.n58 VDD.t1941 93.3253
R14750 VDD.n21 VDD.t2068 93.3253
R14751 VDD.n419 VDD.n418 92.9887
R14752 VDD.n417 VDD.n416 92.5005
R14753 VDD.n416 VDD.t2054 92.5005
R14754 VDD.n389 VDD.n388 92.5005
R14755 VDD.n388 VDD.t2054 92.5005
R14756 VDD.n391 VDD.n363 92.5005
R14757 VDD.t2944 VDD.n363 92.5005
R14758 VDD.n394 VDD.n393 92.5005
R14759 VDD.t2051 VDD.n394 92.5005
R14760 VDD.n386 VDD.n385 92.5005
R14761 VDD.n385 VDD.t2056 92.5005
R14762 VDD.n380 VDD.n377 92.5005
R14763 VDD.t2056 VDD.n377 92.5005
R14764 VDD.n384 VDD.n383 92.5005
R14765 VDD.t2056 VDD.n384 92.5005
R14766 VDD.n396 VDD.n395 92.5005
R14767 VDD.n395 VDD.t2051 92.5005
R14768 VDD.n413 VDD.n412 92.5005
R14769 VDD.t2944 VDD.n413 92.5005
R14770 VDD.n357 VDD.n355 92.5005
R14771 VDD.n355 VDD.t2054 92.5005
R14772 VDD.n319 VDD.n303 92.5005
R14773 VDD.n315 VDD.n302 92.5005
R14774 VDD.n302 VDD.t1770 92.5005
R14775 VDD.t2153 VDD.t1220 92.315
R14776 VDD.t2114 VDD.t1477 92.315
R14777 VDD.t2185 VDD.t1793 92.315
R14778 VDD.t3086 VDD.t2155 92.315
R14779 VDD.t678 VDD.t31 92.315
R14780 VDD.t990 VDD.t617 92.315
R14781 VDD.t662 VDD.t1608 92.315
R14782 VDD.n206 VDD.n205 91.4829
R14783 VDD.n295 VDD.t3578 91.2567
R14784 VDD.t2661 VDD.t2563 90.6365
R14785 VDD.t2275 VDD.t1584 90.6365
R14786 VDD.t1099 VDD.t2147 90.6365
R14787 VDD.t3720 VDD.t2895 90.6365
R14788 VDD.t561 VDD.t2305 90.6365
R14789 VDD.n329 VDD.t3592 90.3207
R14790 VDD.n291 VDD.n196 90.2911
R14791 VDD.t1715 VDD.t3239 88.9581
R14792 VDD.t2118 VDD.t1469 88.9581
R14793 VDD.t797 VDD.t579 88.9581
R14794 VDD.t2487 VDD.t1843 88.9581
R14795 VDD.t2781 VDD.t3345 88.9581
R14796 VDD.t2673 VDD.t1541 88.9581
R14797 VDD.t3406 VDD.t2368 88.9581
R14798 VDD.t1294 VDD.t483 88.9581
R14799 VDD.t920 VDD.t2777 88.9581
R14800 VDD.t2659 VDD.t1833 87.2797
R14801 VDD.t2009 VDD.t2470 87.2797
R14802 VDD.t2880 VDD.t124 87.2797
R14803 VDD.t1287 VDD.t3124 87.2797
R14804 VDD.n1598 VDD.t2863 87.2797
R14805 VDD.t731 VDD.t1001 87.2797
R14806 VDD.t1360 VDD.t1482 87.2797
R14807 VDD.t690 VDD.t2741 87.2797
R14808 VDD.n952 VDD.t405 87.2797
R14809 VDD.t2281 VDD.t2924 87.2797
R14810 VDD.t922 VDD.t3019 87.2797
R14811 VDD.t3474 VDD.t1097 87.2797
R14812 VDD.t924 VDD.t2731 87.2797
R14813 VDD.t427 VDD.t2047 87.2797
R14814 VDD.t2966 VDD.t3531 87.2797
R14815 VDD.t2100 VDD.t816 87.2797
R14816 VDD.t1263 VDD.t2496 87.2797
R14817 VDD.n3899 VDD.t2537 86.7743
R14818 VDD.n3990 VDD.t1514 86.7743
R14819 VDD.n3997 VDD.t2510 86.7743
R14820 VDD.n4016 VDD.t2154 86.7743
R14821 VDD.n4037 VDD.t568 86.7743
R14822 VDD.n4091 VDD.t776 86.7743
R14823 VDD.n4273 VDD.t2266 86.7743
R14824 VDD.n3694 VDD.t2730 86.7743
R14825 VDD.n3690 VDD.t1566 86.7743
R14826 VDD.n3212 VDD.t1144 86.7743
R14827 VDD.n3225 VDD.t1748 86.7743
R14828 VDD.n3577 VDD.t2709 86.7743
R14829 VDD.n3302 VDD.t1752 86.7743
R14830 VDD.n3181 VDD.t1128 86.7743
R14831 VDD.n3821 VDD.t1422 86.7743
R14832 VDD.n3096 VDD.t2881 86.7743
R14833 VDD.n2837 VDD.t2833 86.7743
R14834 VDD.n2280 VDD.t2736 86.7743
R14835 VDD.n2459 VDD.t2716 86.7743
R14836 VDD.n2668 VDD.t980 86.7743
R14837 VDD.n1964 VDD.t3721 86.7743
R14838 VDD.n1964 VDD.t3449 86.7743
R14839 VDD.n1600 VDD.t1765 86.7743
R14840 VDD.n1600 VDD.t1303 86.7743
R14841 VDD.n1877 VDD.t3621 86.7743
R14842 VDD.n1877 VDD.t254 86.7743
R14843 VDD.n970 VDD.t2000 86.7743
R14844 VDD.n1317 VDD.t677 86.7743
R14845 VDD.t116 VDD.t904 85.6012
R14846 VDD.t113 VDD.t2399 85.6012
R14847 VDD.t2116 VDD.t1473 85.6012
R14848 VDD.t2461 VDD.t3410 85.6012
R14849 VDD.t2590 VDD.t1139 85.6012
R14850 VDD.t3116 VDD.t1290 85.6012
R14851 VDD.t527 VDD.t1042 85.6012
R14852 VDD.t1818 VDD.t1183 85.6012
R14853 VDD.t1999 VDD.t3355 85.6012
R14854 VDD.n333 VDD.n188 85.5545
R14855 VDD.n383 VDD.n366 84.2672
R14856 VDD.n396 VDD.n366 84.2672
R14857 VDD.n410 VDD.n396 84.2672
R14858 VDD.n412 VDD.n410 84.2672
R14859 VDD.n412 VDD.n411 84.2672
R14860 VDD.n411 VDD.n357 84.2672
R14861 VDD.t3180 VDD.n4341 83.9228
R14862 VDD.t2315 VDD.t3401 83.9228
R14863 VDD.t1567 VDD.t3462 83.9228
R14864 VDD.t387 VDD.t11 83.9228
R14865 VDD.t607 VDD.t2644 83.9228
R14866 VDD.t3377 VDD.t3343 83.9228
R14867 VDD.t2233 VDD.t2248 83.9228
R14868 VDD.t1935 VDD.t3363 83.9228
R14869 VDD.t799 VDD.t245 82.2443
R14870 VDD.t2382 VDD.t2978 82.2443
R14871 VDD.t2457 VDD.t3512 82.2443
R14872 VDD.t3013 VDD.t938 82.2443
R14873 VDD.t3422 VDD.t2789 82.2443
R14874 VDD.t3735 VDD.t3134 82.2443
R14875 VDD.t2596 VDD.t3624 82.2443
R14876 VDD.t820 VDD.t2551 82.2443
R14877 VDD.n4152 VDD.t2836 80.5659
R14878 VDD.t2511 VDD.t1232 80.5659
R14879 VDD.t1219 VDD.t1344 80.5659
R14880 VDD.n4650 VDD.t940 80.5659
R14881 VDD.n3319 VDD.t2045 80.5659
R14882 VDD.n2594 VDD.t1965 80.5659
R14883 VDD.n2595 VDD.t3090 80.5659
R14884 VDD.t3673 VDD.t2199 80.5659
R14885 VDD.t3292 VDD.n2725 80.5659
R14886 VDD.n2726 VDD.t3647 80.5659
R14887 VDD.t1004 VDD.t2832 80.5659
R14888 VDD.t437 VDD.t21 80.5659
R14889 VDD.t2262 VDD.t1230 80.5659
R14890 VDD.n1689 VDD.t1801 80.5659
R14891 VDD.t2323 VDD.t601 80.5659
R14892 VDD.t110 VDD.t2565 80.5659
R14893 VDD.t79 VDD.t3308 80.5659
R14894 VDD.t2865 VDD.t2290 80.5659
R14895 VDD.t2136 VDD.t2179 80.5659
R14896 VDD.t999 VDD.t2373 80.5659
R14897 VDD.t2812 VDD.t834 80.5659
R14898 VDD.t1459 VDD.t515 80.5659
R14899 VDD.n320 VDD.n314 80.5652
R14900 VDD.n205 VDD.n204 80.5652
R14901 VDD.t1351 VDD.t1993 78.8874
R14902 VDD.t85 VDD.t1835 78.8874
R14903 VDD.t2257 VDD.t2315 78.8874
R14904 VDD.t3296 VDD.t2704 78.8874
R14905 VDD.t3569 VDD.t3208 78.8874
R14906 VDD.t2259 VDD.n2895 78.8874
R14907 VDD.t144 VDD.t3365 78.8874
R14908 VDD.t3357 VDD.t607 78.8874
R14909 VDD.t615 VDD.t1697 78.8874
R14910 VDD.t742 VDD.t863 78.8874
R14911 VDD.t3343 VDD.t1606 78.8874
R14912 VDD.t3391 VDD.t2233 78.8874
R14913 VDD.t1559 VDD.t2005 78.8874
R14914 VDD.n66 VDD.t1664 78.8874
R14915 VDD.n28 VDD.t2403 78.8874
R14916 VDD.n4195 VDD.t1862 77.3934
R14917 VDD.n4134 VDD.t1994 77.3934
R14918 VDD.n4131 VDD.t2660 77.3934
R14919 VDD.n3231 VDD.t3633 77.3934
R14920 VDD.n3241 VDD.t248 77.3934
R14921 VDD.n3802 VDD.t430 77.3934
R14922 VDD.n3790 VDD.t2829 77.3934
R14923 VDD.n3185 VDD.t386 77.3934
R14924 VDD.n2804 VDD.t266 77.3934
R14925 VDD.n2421 VDD.t1974 77.3934
R14926 VDD.n2424 VDD.t1295 77.3934
R14927 VDD.t3239 VDD.t1094 77.209
R14928 VDD.t1494 VDD.t1342 77.209
R14929 VDD.t1513 VDD.t2797 77.209
R14930 VDD.t2208 VDD.t2536 77.209
R14931 VDD.t1563 VDD.t2461 77.209
R14932 VDD.t2602 VDD.t2714 77.209
R14933 VDD.t764 VDD.t1129 77.209
R14934 VDD.t987 VDD.t850 77.209
R14935 VDD.t2187 VDD.t2065 77.209
R14936 VDD.t2667 VDD.t3118 77.209
R14937 VDD.t1042 VDD.t3306 77.209
R14938 VDD.t2639 VDD.t551 77.209
R14939 VDD.t2555 VDD.t820 77.209
R14940 VDD.t72 VDD.n323 76.2813
R14941 VDD.t3756 VDD.t2802 75.5305
R14942 VDD.t1619 VDD.t1055 75.5305
R14943 VDD.t1475 VDD.t2356 75.5305
R14944 VDD.t1955 VDD.t2185 75.5305
R14945 VDD.t1083 VDD.t2348 75.5305
R14946 VDD.t1885 VDD.t1492 75.5305
R14947 VDD.t3341 VDD.t1014 75.5305
R14948 VDD.t1791 VDD.t3220 75.5305
R14949 VDD.t938 VDD.t3119 75.5305
R14950 VDD.t625 VDD.t3145 75.5305
R14951 VDD.t1482 VDD.t3630 75.5305
R14952 VDD.t1507 VDD.t853 75.5305
R14953 VDD.t1913 VDD.t549 75.5305
R14954 VDD.t2814 VDD.t1899 75.5305
R14955 VDD.t2005 VDD.t3474 75.5305
R14956 VDD.t2047 VDD.t3451 75.5305
R14957 VDD.n329 VDD.t69 75.3453
R14958 VDD.n2510 VDD.t2430 75.0481
R14959 VDD.n1785 VDD.t1329 75.0481
R14960 VDD.n1641 VDD.t2520 75.0481
R14961 VDD.n1660 VDD.t2668 75.0481
R14962 VDD.t2470 VDD.t2153 73.8521
R14963 VDD.t124 VDD.t3510 73.8521
R14964 VDD.n2725 VDD.t1638 73.8521
R14965 VDD.t2960 VDD.n1597 73.8521
R14966 VDD.t2307 VDD.t157 73.8521
R14967 VDD.t3255 VDD.t655 73.8521
R14968 VDD.n1079 VDD.t2965 73.8521
R14969 VDD.t1391 VDD.t2855 72.1736
R14970 VDD.t1833 VDD.t2661 72.1736
R14971 VDD.t1584 VDD.t3359 72.1736
R14972 VDD.t218 VDD.t2286 72.1736
R14973 VDD.t3164 VDD.t767 72.1736
R14974 VDD.t1061 VDD.t2484 72.1736
R14975 VDD.t2484 VDD.t1077 72.1736
R14976 VDD.t1077 VDD.t538 72.1736
R14977 VDD.t538 VDD.t1065 72.1736
R14978 VDD.t1143 VDD.t972 72.1736
R14979 VDD.t840 VDD.t755 72.1736
R14980 VDD.t140 VDD.t595 72.1736
R14981 VDD.t2199 VDD.t849 72.1736
R14982 VDD.t1034 VDD.t3560 72.1736
R14983 VDD.t3560 VDD.t1032 72.1736
R14984 VDD.t2992 VDD.t3393 72.1736
R14985 VDD.t295 VDD.n2027 72.1736
R14986 VDD.t1125 VDD.t690 72.1736
R14987 VDD.n737 VDD.t1423 72.1736
R14988 VDD.n113 VDD.n112 71.9064
R14989 VDD.n115 VDD.n113 71.9064
R14990 VDD.n316 VDD.n303 70.7763
R14991 VDD.t2527 VDD.t3198 70.4952
R14992 VDD.t3495 VDD.t637 70.4952
R14993 VDD.t637 VDD.t3497 70.4952
R14994 VDD.t1843 VDD.t3086 70.4952
R14995 VDD.t1487 VDD.t2675 70.4952
R14996 VDD.t2675 VDD.t1484 70.4952
R14997 VDD.t3009 VDD.n2028 70.4952
R14998 VDD.n2028 VDD.t3004 70.4952
R14999 VDD.n2171 VDD.t3690 70.4952
R15000 VDD.t2337 VDD.t2538 70.4952
R15001 VDD.t3263 VDD.t922 70.4952
R15002 VDD.t918 VDD.t3263 70.4952
R15003 VDD.t1097 VDD.t1105 70.4952
R15004 VDD.t1105 VDD.t2298 70.4952
R15005 VDD.t327 VDD.t676 70.4952
R15006 VDD.t1919 VDD.t818 70.4952
R15007 VDD.t816 VDD.t1919 70.4952
R15008 VDD.n846 VDD.t1532 69.9355
R15009 VDD.n352 VDD.n342 69.2711
R15010 VDD.t2284 VDD.t218 68.8168
R15011 VDD.t2348 VDD.t1061 68.8168
R15012 VDD.t593 VDD.t140 68.8168
R15013 VDD.t1032 VDD.t3341 68.8168
R15014 VDD.t1008 VDD.t1791 68.8168
R15015 VDD.t2719 VDD.t2992 68.8168
R15016 VDD.t3145 VDD.t597 68.8168
R15017 VDD.t549 VDD.t1902 68.8168
R15018 VDD.t2806 VDD.t1529 68.8168
R15019 VDD.t1608 VDD.t1245 68.8168
R15020 VDD.n3899 VDD.t1922 68.0124
R15021 VDD.n3990 VDD.t1918 68.0124
R15022 VDD.n3997 VDD.t2607 68.0124
R15023 VDD.n4016 VDD.t2010 68.0124
R15024 VDD.n4037 VDD.t1908 68.0124
R15025 VDD.n4091 VDD.t2619 68.0124
R15026 VDD.n4273 VDD.t659 68.0124
R15027 VDD.n3694 VDD.t362 68.0124
R15028 VDD.n3690 VDD.t2003 68.0124
R15029 VDD.n3212 VDD.t1140 68.0124
R15030 VDD.n3225 VDD.t1704 68.0124
R15031 VDD.n3577 VDD.t2705 68.0124
R15032 VDD.n3302 VDD.t2061 68.0124
R15033 VDD.n3181 VDD.t376 68.0124
R15034 VDD.n3821 VDD.t1418 68.0124
R15035 VDD.n3096 VDD.t3511 68.0124
R15036 VDD.n2837 VDD.t2334 68.0124
R15037 VDD.n2280 VDD.t3655 68.0124
R15038 VDD.n2459 VDD.t1291 68.0124
R15039 VDD.n2668 VDD.t1288 68.0124
R15040 VDD.n1317 VDD.t3538 68.0124
R15041 VDD.t1340 VDD.t1494 67.1383
R15042 VDD.t759 VDD.t2725 67.1383
R15043 VDD.t3762 VDD.t3008 67.1383
R15044 VDD.t1249 VDD.t1175 67.1383
R15045 VDD.t3121 VDD.t2667 67.1383
R15046 VDD.t1037 VDD.t1036 67.1383
R15047 VDD.n2614 VDD.n2613 66.9805
R15048 VDD.n971 VDD.t1744 66.8398
R15049 VDD.t1993 VDD.t1195 65.4599
R15050 VDD.t2311 VDD.t2257 65.4599
R15051 VDD.t2665 VDD.t765 65.4599
R15052 VDD.t471 VDD.t2007 65.4599
R15053 VDD.t3220 VDD.t3569 65.4599
R15054 VDD.t599 VDD.t3357 65.4599
R15055 VDD.t1697 VDD.t625 65.4599
R15056 VDD.t1606 VDD.t3566 65.4599
R15057 VDD.t853 VDD.t1502 65.4599
R15058 VDD.t551 VDD.t1913 65.4599
R15059 VDD.t2737 VDD.t547 65.4599
R15060 VDD.t1401 VDD.t2246 65.4599
R15061 VDD.n342 VDD.n341 64.0005
R15062 VDD.n404 VDD.t2945 63.8266
R15063 VDD.t642 VDD.n4069 63.7814
R15064 VDD.t1094 VDD.t1783 63.7814
R15065 VDD.t1342 VDD.t1219 63.7814
R15066 VDD.t1344 VDD.t2469 63.7814
R15067 VDD.t3153 VDD.t1563 63.7814
R15068 VDD.t2753 VDD.n3754 63.7814
R15069 VDD.t3122 VDD.t2201 63.7814
R15070 VDD.t3661 VDD.t979 63.7814
R15071 VDD.t2832 VDD.t1010 63.7814
R15072 VDD.t13 VDD.t437 63.7814
R15073 VDD.t2735 VDD.t3710 63.7814
R15074 VDD.t1883 VDD.t2779 63.7814
R15075 VDD.t553 VDD.t2639 63.7814
R15076 VDD.t2626 VDD.t2988 63.7814
R15077 VDD.t2248 VDD.t3687 63.7814
R15078 VDD.n398 VDD.t2052 63.7312
R15079 VDD.n4608 VDD.t3402 63.3219
R15080 VDD.n4603 VDD.t3388 63.3219
R15081 VDD.n4568 VDD.t3386 63.3219
R15082 VDD.n4000 VDD.t3380 63.3219
R15083 VDD.n4021 VDD.t3368 63.3219
R15084 VDD.n4028 VDD.t3384 63.3219
R15085 VDD.n4476 VDD.t2981 63.3219
R15086 VDD.n4439 VDD.t2971 63.3219
R15087 VDD.n4045 VDD.t1828 63.3219
R15088 VDD.n4049 VDD.t1842 63.3219
R15089 VDD.n4071 VDD.t1836 63.3219
R15090 VDD.n4076 VDD.t1830 63.3219
R15091 VDD.n4278 VDD.t3360 63.3219
R15092 VDD.n4272 VDD.t3415 63.3219
R15093 VDD.n4130 VDD.t1834 63.3219
R15094 VDD.n4138 VDD.t1850 63.3219
R15095 VDD.n3687 VDD.t2975 63.3219
R15096 VDD.n3747 VDD.t2979 63.3219
R15097 VDD.n3237 VDD.t3195 63.3219
R15098 VDD.n3237 VDD.t1725 63.3219
R15099 VDD.n3247 VDD.t3197 63.3219
R15100 VDD.n3247 VDD.t1746 63.3219
R15101 VDD.n3527 VDD.t1844 63.3219
R15102 VDD.n3260 VDD.t1840 63.3219
R15103 VDD.n3276 VDD.t3413 63.3219
R15104 VDD.n3283 VDD.t3354 63.3219
R15105 VDD.n3400 VDD.t3411 63.3219
R15106 VDD.n3454 VDD.t3417 63.3219
R15107 VDD.n3395 VDD.t3419 63.3219
R15108 VDD.n3387 VDD.t3425 63.3219
R15109 VDD.n3299 VDD.t3409 63.3219
R15110 VDD.n3358 VDD.t3362 63.3219
R15111 VDD.n3109 VDD.t3396 63.3219
R15112 VDD.n3115 VDD.t3372 63.3219
R15113 VDD.n2524 VDD.t3427 63.3219
R15114 VDD.n2509 VDD.t3350 63.3219
R15115 VDD.n2506 VDD.t3346 63.3219
R15116 VDD.n2506 VDD.t2428 63.3219
R15117 VDD.n2294 VDD.t3394 63.3219
R15118 VDD.n2433 VDD.t967 63.3219
R15119 VDD.n2443 VDD.t3311 63.3219
R15120 VDD.n2628 VDD.t3407 63.3219
R15121 VDD.n2479 VDD.t3352 63.3219
R15122 VDD.n2671 VDD.t3662 63.3219
R15123 VDD.n2299 VDD.t3366 63.3219
R15124 VDD.n1555 VDD.t3378 63.3219
R15125 VDD.n1978 VDD.t3398 63.3219
R15126 VDD.n2011 VDD.t2912 63.3219
R15127 VDD.n2011 VDD.t1814 63.3219
R15128 VDD.n1609 VDD.t2933 63.3219
R15129 VDD.n1609 VDD.t50 63.3219
R15130 VDD.n1810 VDD.t3358 63.3219
R15131 VDD.n1633 VDD.t3405 63.3219
R15132 VDD.n1634 VDD.t2381 63.3219
R15133 VDD.n1634 VDD.t2274 63.3219
R15134 VDD.n1644 VDD.t831 63.3219
R15135 VDD.n1644 VDD.t939 63.3219
R15136 VDD.n1656 VDD.t715 63.3219
R15137 VDD.n1656 VDD.t870 63.3219
R15138 VDD.n1663 VDD.t1540 63.3219
R15139 VDD.n1663 VDD.t2188 63.3219
R15140 VDD.n1667 VDD.t1599 63.3219
R15141 VDD.n2173 VDD.t3400 63.3219
R15142 VDD.n2178 VDD.t3382 63.3219
R15143 VDD.n2181 VDD.t3390 63.3219
R15144 VDD.n2184 VDD.t3370 63.3219
R15145 VDD.n800 VDD.t1838 63.3219
R15146 VDD.n804 VDD.t1848 63.3219
R15147 VDD.n1019 VDD.t1832 63.3219
R15148 VDD.n1051 VDD.t1856 63.3219
R15149 VDD.n834 VDD.t3356 63.3219
R15150 VDD.n833 VDD.t2989 63.3219
R15151 VDD.n838 VDD.t3421 63.3219
R15152 VDD.n776 VDD.t3392 63.3219
R15153 VDD.n781 VDD.t3376 63.3219
R15154 VDD.n1137 VDD.t1846 63.3219
R15155 VDD.n1143 VDD.t1854 63.3219
R15156 VDD.n1406 VDD.t3374 63.3219
R15157 VDD.n1413 VDD.t3364 63.3219
R15158 VDD.n646 VDD.n643 62.9556
R15159 VDD.t2708 VDD.t1580 62.103
R15160 VDD.t2151 VDD.t1181 62.103
R15161 VDD.t1115 VDD.t3288 62.103
R15162 VDD.t3654 VDD.t381 62.103
R15163 VDD.t617 VDD.t2323 62.103
R15164 VDD.t2331 VDD.t742 62.103
R15165 VDD.t2577 VDD.t1453 62.103
R15166 VDD.t3355 VDD.t1741 62.103
R15167 VDD.t2411 VDD.t2882 62.103
R15168 VDD.n66 VDD.t1658 62.103
R15169 VDD.n28 VDD.t2407 62.103
R15170 VDD.t1941 VDD.t1940 61.7891
R15171 VDD.t1940 VDD.t1953 61.7891
R15172 VDD.t1953 VDD.t1948 61.7891
R15173 VDD.t1948 VDD.t1944 61.7891
R15174 VDD.t1944 VDD.t1947 61.7891
R15175 VDD.t1947 VDD.t1954 61.7891
R15176 VDD.t1954 VDD.t1950 61.7891
R15177 VDD.t1950 VDD.t1942 61.7891
R15178 VDD.t1942 VDD.t1952 61.7891
R15179 VDD.t1952 VDD.t1946 61.7891
R15180 VDD.t1946 VDD.t1939 61.7891
R15181 VDD.t1939 VDD.t1949 61.7891
R15182 VDD.t1949 VDD.t1951 61.7891
R15183 VDD.t1951 VDD.t1943 61.7891
R15184 VDD.t1943 VDD.t1945 61.7891
R15185 VDD.t1945 VDD.t1775 61.7891
R15186 VDD.t1775 VDD.t1774 61.7891
R15187 VDD.t1774 VDD.t1779 61.7891
R15188 VDD.t1779 VDD.t1778 61.7891
R15189 VDD.t1778 VDD.t1776 61.7891
R15190 VDD.t1780 VDD.t1773 61.7891
R15191 VDD.t1773 VDD.t1777 61.7891
R15192 VDD.t1777 VDD.t3557 61.7891
R15193 VDD.t3557 VDD.t3556 61.7891
R15194 VDD.t3556 VDD.t3554 61.7891
R15195 VDD.t3554 VDD.t3555 61.7891
R15196 VDD.t3555 VDD.t1964 61.7891
R15197 VDD.t1964 VDD.t1963 61.7891
R15198 VDD.t1963 VDD.t2001 61.7891
R15199 VDD.t1972 VDD.t3604 61.7891
R15200 VDD.t1969 VDD.t1972 61.7891
R15201 VDD.t3609 VDD.t1969 61.7891
R15202 VDD.t3613 VDD.t3609 61.7891
R15203 VDD.t3610 VDD.t3613 61.7891
R15204 VDD.t3614 VDD.t3610 61.7891
R15205 VDD.t3072 VDD.t3614 61.7891
R15206 VDD.t3079 VDD.t3072 61.7891
R15207 VDD.t3073 VDD.t3079 61.7891
R15208 VDD.t3075 VDD.t3080 61.7891
R15209 VDD.t3076 VDD.t3075 61.7891
R15210 VDD.t3078 VDD.t3076 61.7891
R15211 VDD.t3074 VDD.t3078 61.7891
R15212 VDD.t2072 VDD.t3074 61.7891
R15213 VDD.t2073 VDD.t2072 61.7891
R15214 VDD.t2074 VDD.t2073 61.7891
R15215 VDD.t2069 VDD.t2074 61.7891
R15216 VDD.t2084 VDD.t2069 61.7891
R15217 VDD.t2071 VDD.t2084 61.7891
R15218 VDD.t2085 VDD.t2071 61.7891
R15219 VDD.t2081 VDD.t2085 61.7891
R15220 VDD.t2075 VDD.t2081 61.7891
R15221 VDD.t2083 VDD.t2075 61.7891
R15222 VDD.t2077 VDD.t2083 61.7891
R15223 VDD.t2070 VDD.t2077 61.7891
R15224 VDD.t2076 VDD.t2070 61.7891
R15225 VDD.t2082 VDD.t2076 61.7891
R15226 VDD.t2080 VDD.t2082 61.7891
R15227 VDD.t2068 VDD.t2080 61.7891
R15228 VDD.n1651 VDD.t392 60.9739
R15229 VDD.t1232 VDD.t2515 60.4245
R15230 VDD.t3401 VDD.t2313 60.4245
R15231 VDD.t1915 VDD.t319 60.4245
R15232 VDD.t3351 VDD.t3673 60.4245
R15233 VDD.t1431 VDD.t1287 60.4245
R15234 VDD.t35 VDD.t387 60.4245
R15235 VDD.t2644 VDD.t627 60.4245
R15236 VDD.t2181 VDD.t2136 60.4245
R15237 VDD.t2179 VDD.t1121 60.4245
R15238 VDD.t2373 VDD.t2281 60.4245
R15239 VDD.t3671 VDD.t2812 60.4245
R15240 VDD.n1651 VDD.t390 59.9892
R15241 VDD.n387 VDD.n386 59.4829
R15242 VDD.n393 VDD.n387 59.4829
R15243 VDD.n393 VDD.n392 59.4829
R15244 VDD.n392 VDD.n391 59.4829
R15245 VDD.n391 VDD.n390 59.4829
R15246 VDD.n390 VDD.n389 59.4829
R15247 VDD.t2395 VDD.t113 58.7461
R15248 VDD.t1473 VDD.t2112 58.7461
R15249 VDD.t245 VDD.t993 58.7461
R15250 VDD.t1447 VDD.t994 58.7461
R15251 VDD.t3023 VDD.t1199 58.7461
R15252 VDD.t1580 VDD.t1888 58.7461
R15253 VDD.t1875 VDD.t2708 58.7461
R15254 VDD.t2754 VDD.t1489 58.7461
R15255 VDD.t3512 VDD.t2459 58.7461
R15256 VDD.t1290 VDD.t650 58.7461
R15257 VDD.t2789 VDD.t1533 58.7461
R15258 VDD.t2791 VDD.t3422 58.7461
R15259 VDD.t1119 VDD.t3735 58.7461
R15260 VDD.t1896 VDD.t2596 58.7461
R15261 VDD.t3624 VDD.t1286 58.7461
R15262 VDD.t2551 VDD.t2774 58.7461
R15263 VDD.t569 VDD.t151 57.0676
R15264 VDD.t3110 VDD.t3661 57.0676
R15265 VDD.t3456 VDD.t1567 57.0676
R15266 VDD.t2779 VDD.t2735 57.0676
R15267 VDD.t1183 VDD.t740 57.0676
R15268 VDD.t2997 VDD.t1038 57.0676
R15269 VDD.n4290 VDD.t2973 55.4067
R15270 VDD.n4112 VDD.t1396 55.4067
R15271 VDD.n4144 VDD.t1990 55.4067
R15272 VDD.n4147 VDD.t1284 55.4067
R15273 VDD.n4155 VDD.t2837 55.4067
R15274 VDD.n4159 VDD.t3703 55.4067
R15275 VDD.n4160 VDD.t1978 55.4067
R15276 VDD.n3959 VDD.t2110 55.4067
R15277 VDD.n3918 VDD.t1988 55.4067
R15278 VDD.n3921 VDD.t3651 55.4067
R15279 VDD.n3922 VDD.t2879 55.4067
R15280 VDD.n3929 VDD.t2040 55.4067
R15281 VDD.n3704 VDD.t1858 55.4067
R15282 VDD.n3315 VDD.t2087 55.4067
R15283 VDD.n3316 VDD.t3245 55.4067
R15284 VDD.n3762 VDD.t3729 55.4067
R15285 VDD.n3323 VDD.t2046 55.4067
R15286 VDD.n3325 VDD.t3646 55.4067
R15287 VDD.n3326 VDD.t3100 55.4067
R15288 VDD.n3126 VDD.t2875 55.4067
R15289 VDD.n3128 VDD.t2022 55.4067
R15290 VDD.n3131 VDD.t2762 55.4067
R15291 VDD.n3132 VDD.t3693 55.4067
R15292 VDD.n2515 VDD.t1542 55.4067
R15293 VDD.n2562 VDD.t348 55.4067
R15294 VDD.n2573 VDD.t1966 55.4067
R15295 VDD.n2575 VDD.t1892 55.4067
R15296 VDD.n2576 VDD.t2105 55.4067
R15297 VDD.n2308 VDD.t3489 55.4067
R15298 VDD.n2310 VDD.t1164 55.4067
R15299 VDD.n2311 VDD.t3709 55.4067
R15300 VDD.n1653 VDD.t2677 55.4067
R15301 VDD.n1676 VDD.t2032 55.4067
R15302 VDD.n1681 VDD.t2042 55.4067
R15303 VDD.n1683 VDD.t3656 55.4067
R15304 VDD.n1684 VDD.t2030 55.4067
R15305 VDD.n1687 VDD.t1802 55.4067
R15306 VDD.n1691 VDD.t1166 55.4067
R15307 VDD.n1692 VDD.t2958 55.4067
R15308 VDD.n1954 VDD.t1860 55.4067
R15309 VDD.n2138 VDD.t2742 55.4067
R15310 VDD.n2192 VDD.t3052 55.4067
R15311 VDD.n2194 VDD.t1763 55.4067
R15312 VDD.n2195 VDD.t3035 55.4067
R15313 VDD.n795 VDD.t450 55.4067
R15314 VDD.n813 VDD.t2767 55.4067
R15315 VDD.n1007 VDD.t556 55.4067
R15316 VDD.n839 VDD.t2178 55.4067
R15317 VDD.n843 VDD.t3559 55.4067
R15318 VDD.n900 VDD.t3725 55.4067
R15319 VDD.n896 VDD.t2089 55.4067
R15320 VDD.n889 VDD.t2866 55.4067
R15321 VDD.n931 VDD.t2560 55.4067
R15322 VDD.n881 VDD.t1436 55.4067
R15323 VDD.n855 VDD.t2035 55.4067
R15324 VDD.n723 VDD.t1355 55.4067
R15325 VDD.n750 VDD.t1718 55.4067
R15326 VDD.n762 VDD.t2760 55.4067
R15327 VDD.n779 VDD.t2580 55.4067
R15328 VDD.n1142 VDD.t2778 55.4067
R15329 VDD.n1360 VDD.t270 55.4067
R15330 VDD.n1368 VDD.t3546 55.4067
R15331 VDD.n1371 VDD.t2204 55.4067
R15332 VDD.n1409 VDD.t2552 55.4067
R15333 VDD.n1417 VDD.t44 55.4067
R15334 VDD.n1422 VDD.t3054 55.4067
R15335 VDD.n1426 VDD.t1986 55.4067
R15336 VDD.n1427 VDD.t2780 55.4067
R15337 VDD.n1430 VDD.t1982 55.4067
R15338 VDD.n1431 VDD.t3649 55.4067
R15339 VDD.t1716 VDD.t116 55.3892
R15340 VDD.t1469 VDD.t2116 55.3892
R15341 VDD.t1640 VDD.t1289 55.3892
R15342 VDD.t479 VDD.t1294 55.3892
R15343 VDD.t3397 VDD.t1818 55.3892
R15344 VDD.t1805 VDD.t1518 55.3892
R15345 VDD.n234 VDD.t230 54.4158
R15346 VDD.n234 VDD.t150 54.4158
R15347 VDD.n240 VDD.t143 54.4158
R15348 VDD.n240 VDD.t97 54.4158
R15349 VDD.t2120 VDD.t2386 53.7107
R15350 VDD.t2725 VDD.t3443 53.7107
R15351 VDD.t964 VDD.t491 53.7107
R15352 VDD.t1001 VDD.t1360 53.7107
R15353 VDD.t2895 VDD.t1925 53.7107
R15354 VDD.t1036 VDD.t3680 53.7107
R15355 VDD.t2741 VDD.t1253 53.7107
R15356 VDD.t542 VDD.t3369 53.7107
R15357 VDD.n952 VDD.t407 53.7107
R15358 VDD.t1743 VDD.t2543 53.7107
R15359 VDD.t3019 VDD.t916 53.7107
R15360 VDD.t2731 VDD.t427 53.7107
R15361 VDD.t814 VDD.t2100 53.7107
R15362 VDD.t2498 VDD.t1263 53.7107
R15363 VDD.n846 VDD.t406 53.1905
R15364 VDD.t2943 VDD.t2130 52.0323
R15365 VDD.t1201 VDD.t215 52.0323
R15366 VDD.t2545 VDD.t1582 52.0323
R15367 VDD.t1477 VDD.t2118 52.0323
R15368 VDD.t579 VDD.t1839 52.0323
R15369 VDD.t3304 VDD.t291 52.0323
R15370 VDD.t1541 VDD.t2416 52.0323
R15371 VDD.t9 VDD.t678 52.0323
R15372 VDD.t2961 VDD.t2719 52.0323
R15373 VDD.t609 VDD.t990 52.0323
R15374 VDD.t2777 VDD.t3325 52.0323
R15375 VDD.n3593 VDD.t2666 51.2205
R15376 VDD.n3620 VDD.t2629 51.2205
R15377 VDD.n825 VDD.t3736 51.2205
R15378 VDD.n1259 VDD.t3817 50.5057
R15379 VDD.t67 VDD.n300 50.3751
R15380 VDD.n300 VDD.t71 50.3751
R15381 VDD.t3751 VDD.t710 50.3539
R15382 VDD.t2976 VDD.t1221 50.3539
R15383 VDD.t53 VDD.t2588 50.3539
R15384 VDD.t1809 VDD.t513 50.3539
R15385 VDD.t978 VDD.n2171 50.3539
R15386 VDD.t2305 VDD.t327 50.3539
R15387 VDD.n207 VDD.n198 48.9417
R15388 VDD.t1471 VDD.t2114 48.6754
R15389 VDD.t1793 VDD.t2183 48.6754
R15390 VDD.t539 VDD.t1079 48.6754
R15391 VDD.t972 VDD.t840 48.6754
R15392 VDD.t31 VDD.t680 48.6754
R15393 VDD.t240 VDD.t1670 48.6754
R15394 VDD.n333 VDD.n332 48.6258
R15395 VDD.n122 VDD.t935 48.6146
R15396 VDD.t3480 VDD.n122 48.6146
R15397 VDD.t3642 VDD.t1722 46.997
R15398 VDD.t2333 VDD.t1024 46.997
R15399 VDD.t1111 VDD.t852 46.997
R15400 VDD.n1597 VDD.t3261 46.997
R15401 VDD.t157 VDD.t3543 46.997
R15402 VDD.t1531 VDD.t2219 46.997
R15403 VDD.n1079 VDD.t3625 46.997
R15404 VDD.t1695 VDD.t3526 46.997
R15405 VDD.n318 VDD.n317 46.2505
R15406 VDD.n321 VDD.n320 46.2505
R15407 VDD.n322 VDD.n321 46.2505
R15408 VDD.n204 VDD.n203 46.2505
R15409 VDD.n201 VDD.n198 46.2505
R15410 VDD.n118 VDD.n112 46.2505
R15411 VDD.n118 VDD.n117 46.2505
R15412 VDD.n116 VDD.n115 46.2505
R15413 VDD.n117 VDD.n116 46.2505
R15414 VDD.t2608 VDD.t2799 45.3185
R15415 VDD.t2122 VDD.t3416 45.3185
R15416 VDD.t2974 VDD.t1565 45.3185
R15417 VDD.t377 VDD.n3865 45.3185
R15418 VDD.t564 VDD.t668 45.3185
R15419 VDD.t2678 VDD.t2519 45.3185
R15420 VDD.t3682 VDD.t1507 45.3185
R15421 VDD.t2140 VDD.t1269 45.3185
R15422 VDD.t2964 VDD.t1853 45.3185
R15423 VDD.t1465 VDD.t1811 45.3185
R15424 VDD.n3703 VDD.t424 45.3105
R15425 VDD.n3209 VDD.t1493 45.3105
R15426 VDD.n3578 VDD.t3317 45.3105
R15427 VDD.n2364 VDD.t388 45.3105
R15428 VDD.n2831 VDD.t957 45.3105
R15429 VDD.n3025 VDD.t695 45.3105
R15430 VDD.t63 VDD.n296 44.5891
R15431 VDD.n301 VDD.t70 44.5891
R15432 VDD.t62 VDD.n296 44.5891
R15433 VDD.t66 VDD.n301 44.5891
R15434 VDD.n3593 VDD.t1130 44.3255
R15435 VDD.n3583 VDD.t532 44.3255
R15436 VDD.n3583 VDD.t3030 44.3255
R15437 VDD.n3620 VDD.t2603 44.3255
R15438 VDD.n3570 VDD.t1280 44.3255
R15439 VDD.n3570 VDD.t3024 44.3255
R15440 VDD.n825 VDD.t1311 44.3255
R15441 VDD.n829 VDD.t2983 44.3255
R15442 VDD.n829 VDD.t3016 44.3255
R15443 VDD.t2934 VDD.t1851 43.6401
R15444 VDD.t2797 VDD.t2999 43.6401
R15445 VDD.t1252 VDD.t2208 43.6401
R15446 VDD.t2415 VDD.t2427 43.6401
R15447 VDD.t1255 VDD.t3349 43.6401
R15448 VDD.t3025 VDD.t1003 43.6401
R15449 VDD.t847 VDD.t3664 43.6401
R15450 VDD.t443 VDD.t328 43.6401
R15451 VDD.n2510 VDD.t1256 43.3874
R15452 VDD.n1785 VDD.t753 43.3874
R15453 VDD.n1641 VDD.t1689 43.3874
R15454 VDD.n1660 VDD.t3340 43.3874
R15455 VDD.n1963 VDD.t2756 42.3555
R15456 VDD.n1602 VDD.t823 42.3555
R15457 VDD.n1871 VDD.t2566 42.3555
R15458 VDD.t2620 VDD.t789 41.9616
R15459 VDD.t2019 VDD.t2467 41.9616
R15460 VDD.t2476 VDD.t1751 41.9616
R15461 VDD.t2344 VDD.t2464 41.9616
R15462 VDD.t1063 VDD.t2818 41.9616
R15463 VDD.t535 VDD.t1067 41.9616
R15464 VDD.t2417 VDD.t633 41.9616
R15465 VDD.t2939 VDD.t1539 41.9616
R15466 VDD.t3 VDD.t611 41.9616
R15467 VDD.t2690 VDD.t447 41.9616
R15468 VDD.t130 VDD.t723 41.9616
R15469 VDD.n4670 VDD.t2209 41.5552
R15470 VDD.n4670 VDD.t3738 41.5552
R15471 VDD.n3989 VDD.t2798 41.5552
R15472 VDD.n3989 VDD.t3740 41.5552
R15473 VDD.n4013 VDD.t2468 41.5552
R15474 VDD.n4013 VDD.t3132 41.5552
R15475 VDD.n4462 VDD.t1092 41.5552
R15476 VDD.n4462 VDD.t3127 41.5552
R15477 VDD.n4057 VDD.t3163 41.5552
R15478 VDD.n4057 VDD.t712 41.5552
R15479 VDD.n4062 VDD.t640 41.5552
R15480 VDD.n4062 VDD.t3160 41.5552
R15481 VDD.n4285 VDD.t1721 41.5552
R15482 VDD.n4285 VDD.t3161 41.5552
R15483 VDD.n4125 VDD.t1197 41.5552
R15484 VDD.n4125 VDD.t3152 41.5552
R15485 VDD.n3669 VDD.t3131 41.5552
R15486 VDD.n3669 VDD.t2752 41.5552
R15487 VDD.n3248 VDD.t1625 41.5552
R15488 VDD.n3248 VDD.t3158 41.5552
R15489 VDD.n3267 VDD.t537 41.5552
R15490 VDD.n3267 VDD.t3167 41.5552
R15491 VDD.n3407 VDD.t2342 41.5552
R15492 VDD.n3407 VDD.t3156 41.5552
R15493 VDD.n3403 VDD.t2462 41.5552
R15494 VDD.n3403 VDD.t3154 41.5552
R15495 VDD.n3386 VDD.t2474 41.5552
R15496 VDD.n3386 VDD.t3165 41.5552
R15497 VDD.n3122 VDD.t1587 41.5552
R15498 VDD.n3122 VDD.t3744 41.5552
R15499 VDD.n2501 VDD.t3141 41.5552
R15500 VDD.n2501 VDD.t1648 41.5552
R15501 VDD.n2610 VDD.t3143 41.5552
R15502 VDD.n2610 VDD.t2657 41.5552
R15503 VDD.n2305 VDD.t1319 41.5552
R15504 VDD.n2305 VDD.t3750 41.5552
R15505 VDD.n1547 VDD.t2437 41.5552
R15506 VDD.n1547 VDD.t3098 41.5552
R15507 VDD.n1826 VDD.t1698 41.5552
R15508 VDD.n1826 VDD.t3146 41.5552
R15509 VDD.n2188 VDD.t1601 41.5552
R15510 VDD.n2188 VDD.t3746 41.5552
R15511 VDD.n2191 VDD.t2689 41.5552
R15512 VDD.n2191 VDD.t3742 41.5552
R15513 VDD.n793 VDD.t1669 41.5552
R15514 VDD.n793 VDD.t3139 41.5552
R15515 VDD.n1065 VDD.t3148 41.5552
R15516 VDD.n1065 VDD.t2507 41.5552
R15517 VDD.n989 VDD.t1120 41.5552
R15518 VDD.n989 VDD.t3135 41.5552
R15519 VDD.n768 VDD.t1676 41.5552
R15520 VDD.n768 VDD.t3129 41.5552
R15521 VDD.n1130 VDD.t3144 41.5552
R15522 VDD.n1130 VDD.t2698 41.5552
R15523 VDD.n1423 VDD.t1323 41.5552
R15524 VDD.n1423 VDD.t3748 41.5552
R15525 VDD.n4195 VDD.t2402 41.0422
R15526 VDD.n4134 VDD.t1392 41.0422
R15527 VDD.n4131 VDD.t2662 41.0422
R15528 VDD.n3231 VDD.t41 41.0422
R15529 VDD.n3241 VDD.t644 41.0422
R15530 VDD.n3802 VDD.t1376 41.0422
R15531 VDD.n3790 VDD.t3338 41.0422
R15532 VDD.n3185 VDD.t2827 41.0422
R15533 VDD.n2804 VDD.t268 41.0422
R15534 VDD.n2421 VDD.t1651 41.0422
R15535 VDD.n2424 VDD.t2206 41.0422
R15536 VDD.n422 VDD.n421 40.6709
R15537 VDD.t2455 VDD.t2810 40.2832
R15538 VDD.t3696 VDD.t2205 40.2832
R15539 VDD.t2679 VDD.t1004 40.2832
R15540 VDD.t3620 VDD.t3294 40.2832
R15541 VDD.t2581 VDD.t914 40.2832
R15542 VDD.t1403 VDD.t1674 40.2832
R15543 VDD.t1979 VDD.t3466 40.2832
R15544 VDD.t812 VDD.t1451 40.2832
R15545 VDD.t1660 VDD.t3061 40.2832
R15546 VDD.t2409 VDD.t3057 40.2832
R15547 VDD.n410 VDD.n409 39.2805
R15548 VDD.t658 VDD.t3414 38.6047
R15549 VDD.t1931 VDD.t2443 38.6047
R15550 VDD.t1085 VDD.t3353 38.6047
R15551 VDD.t1997 VDD.t2941 38.6047
R15552 VDD.t3241 VDD.t429 38.6047
R15553 VDD.t2787 VDD.t3675 38.6047
R15554 VDD.t533 VDD.t3114 38.6047
R15555 VDD.t2177 VDD.t3420 38.6047
R15556 VDD.t572 VDD.t2479 38.6047
R15557 VDD.n3170 VDD.t1928 38.4155
R15558 VDD.n3815 VDD.t3436 38.4155
R15559 VDD.n2968 VDD.t2900 38.4155
R15560 VDD.n2614 VDD.t1536 38.4155
R15561 VDD.n2674 VDD.t3115 38.4155
R15562 VDD.n1990 VDD.t522 38.4155
R15563 VDD.n1578 VDD.t3321 38.4155
R15564 VDD.n134 VDD.t1246 38.4155
R15565 VDD.n4612 VDD.t2310 37.4305
R15566 VDD.n4600 VDD.t2115 37.4305
R15567 VDD.n4549 VDD.t2398 37.4305
R15568 VDD.n4029 VDD.t1339 37.4305
R15569 VDD.n4457 VDD.t739 37.4305
R15570 VDD.n4489 VDD.t1212 37.4305
R15571 VDD.n4058 VDD.t466 37.4305
R15572 VDD.n4081 VDD.t796 37.4305
R15573 VDD.n4081 VDD.t3199 37.4305
R15574 VDD.n4099 VDD.t2131 37.4305
R15575 VDD.n4107 VDD.t2176 37.4305
R15576 VDD.n3925 VDD.t422 37.4305
R15577 VDD.n3170 VDD.t726 37.4305
R15578 VDD.n3189 VDD.t2228 37.4305
R15579 VDD.n3815 VDD.t2589 37.4305
R15580 VDD.n2968 VDD.t1568 37.4305
R15581 VDD.n2374 VDD.t669 37.4305
R15582 VDD.n2674 VDD.t2718 37.4305
R15583 VDD.n1990 VDD.t2821 37.4305
R15584 VDD.n1578 VDD.t2936 37.4305
R15585 VDD.n851 VDD.t1241 37.4305
R15586 VDD.n304 VDD.n189 37.2235
R15587 VDD.n304 VDD.n299 37.2235
R15588 VDD.n313 VDD.n299 37.2235
R15589 VDD.n332 VDD.n189 37.1499
R15590 VDD.t2628 VDD.t2706 36.9263
R15591 VDD.t958 VDD.t3563 36.9263
R15592 VDD.t2471 VDD.t3435 36.9263
R15593 VDD.t2149 VDD.t1649 36.9263
R15594 VDD.t2658 VDD.t2369 36.9263
R15595 VDD.t1298 VDD.t3679 36.9263
R15596 VDD.t2433 VDD.t830 36.9263
R15597 VDD.t962 VDD.t2625 36.9263
R15598 VDD.t2413 VDD.t2699 36.9263
R15599 VDD.t2553 VDD.t3373 36.9263
R15600 VDD.n4305 VDD.t1186 36.4455
R15601 VDD.n3585 VDD.t953 36.4455
R15602 VDD.n3245 VDD.t837 36.4455
R15603 VDD.n3257 VDD.t2488 36.4455
R15604 VDD.n3419 VDD.t2184 36.4455
R15605 VDD.n3004 VDD.t681 36.4455
R15606 VDD.n2388 VDD.t1313 36.4455
R15607 VDD.n1412 VDD.t2497 36.4455
R15608 VDD.t1776 VDD.n57 36.2048
R15609 VDD.t3080 VDD.n20 36.2048
R15610 VDD.n3915 VDD.t2466 36.1587
R15611 VDD.n3915 VDD.t1934 36.1587
R15612 VDD.n4087 VDD.t410 36.1587
R15613 VDD.n4087 VDD.t1769 36.1587
R15614 VDD.n4121 VDD.t2874 36.1587
R15615 VDD.n4121 VDD.t2796 36.1587
R15616 VDD.n4141 VDD.t2872 36.1587
R15617 VDD.n4141 VDD.t1053 36.1587
R15618 VDD.n4149 VDD.t2870 36.1587
R15619 VDD.n4149 VDD.t1528 36.1587
R15620 VDD.n4156 VDD.t3573 36.1587
R15621 VDD.n4156 VDD.t675 36.1587
R15622 VDD.n2302 VDD.t3092 36.1587
R15623 VDD.n2302 VDD.t2635 36.1587
R15624 VDD.n2564 VDD.t2243 36.1587
R15625 VDD.n2564 VDD.t3575 36.1587
R15626 VDD.n1534 VDD.t3429 36.1587
R15627 VDD.n1534 VDD.t1224 36.1587
R15628 VDD.n1673 VDD.t3032 36.1587
R15629 VDD.n1673 VDD.t1138 36.1587
R15630 VDD.n719 VDD.t1696 36.1587
R15631 VDD.n719 VDD.t1980 36.1587
R15632 VDD.n752 VDD.t2053 36.1587
R15633 VDD.n752 VDD.t2297 36.1587
R15634 VDD.n775 VDD.t2234 36.1587
R15635 VDD.n775 VDD.t3688 36.1587
R15636 VDD.n814 VDD.t3232 36.1587
R15637 VDD.n814 VDD.t2572 36.1587
R15638 VDD.n1022 VDD.t2885 36.1587
R15639 VDD.n1022 VDD.t730 36.1587
R15640 VDD.n821 VDD.t2374 36.1587
R15641 VDD.n821 VDD.t2925 36.1587
R15642 VDD.n714 VDD.t3617 36.1587
R15643 VDD.n714 VDD.t2852 36.1587
R15644 VDD.n770 VDD.t1260 36.1587
R15645 VDD.n770 VDD.t3234 36.1587
R15646 VDD.n1136 VDD.t2108 36.1587
R15647 VDD.n1136 VDD.t2539 36.1587
R15648 VDD.n295 VDD.t3598 36.035
R15649 VDD.n2392 VDD.t2902 35.4605
R15650 VDD.n1548 VDD.t3571 35.4605
R15651 VDD.n2117 VDD.t3249 35.4605
R15652 VDD.n2129 VDD.t3007 35.4605
R15653 VDD.n658 VDD.t338 35.4605
R15654 VDD.n657 VDD.t2317 35.4605
R15655 VDD.n650 VDD.t1572 35.4605
R15656 VDD.n615 VDD.t3063 35.4605
R15657 VDD.n614 VDD.t2923 35.4605
R15658 VDD.n635 VDD.t2892 35.4605
R15659 VDD.n532 VDD.t2037 35.4605
R15660 VDD.n531 VDD.t3081 35.4605
R15661 VDD.n553 VDD.t2024 35.4605
R15662 VDD.n552 VDD.t3031 35.4605
R15663 VDD.n563 VDD.t2524 35.4605
R15664 VDD.n562 VDD.t370 35.4605
R15665 VDD.n573 VDD.t1552 35.4605
R15666 VDD.n572 VDD.t778 35.4605
R15667 VDD.n452 VDD.t2028 35.4605
R15668 VDD.n451 VDD.t3230 35.4605
R15669 VDD.n473 VDD.t3639 35.4605
R15670 VDD.n472 VDD.t2888 35.4605
R15671 VDD.n483 VDD.t2550 35.4605
R15672 VDD.n482 VDD.t1380 35.4605
R15673 VDD.n493 VDD.t1708 35.4605
R15674 VDD.n492 VDD.t2363 35.4605
R15675 VDD.t3754 VDD.t1829 35.2479
R15676 VDD.t1617 VDD.t3379 35.2479
R15677 VDD.t2800 VDD.t2606 35.2479
R15678 VDD.t3387 VDD.t2354 35.2479
R15679 VDD.t1247 VDD.t2063 35.2479
R15680 VDD.t1292 VDD.t2717 35.2479
R15681 VDD.t855 VDD.t521 35.2479
R15682 VDD.t1991 VDD.t2569 35.2479
R15683 VDD.t3657 VDD.t2505 35.2479
R15684 VDD.t47 VDD.t977 35.2479
R15685 VDD.n209 VDD.n207 34.7055
R15686 VDD.n3978 VDD.n3977 34.6358
R15687 VDD.n4291 VDD.n4094 34.6358
R15688 VDD.n3710 VDD.n3709 34.6358
R15689 VDD.n3561 VDD.n3559 34.6358
R15690 VDD.n3548 VDD.n3547 34.6358
R15691 VDD.n3529 VDD.n3526 34.6358
R15692 VDD.n3850 VDD.n3817 34.6358
R15693 VDD.n2337 VDD.n2336 34.6358
R15694 VDD.n1734 VDD.n1733 34.6358
R15695 VDD.n1085 VDD.n815 34.6358
R15696 VDD.n1034 VDD.n1023 34.6358
R15697 VDD.n1348 VDD.n1347 34.6358
R15698 VDD.n1280 VDD.n753 34.6358
R15699 VDD.n1225 VDD.n773 34.6358
R15700 VDD.n1161 VDD.n1151 34.6358
R15701 VDD.n1486 VDD.n1485 34.6358
R15702 VDD.n1467 VDD.n1466 34.6358
R15703 VDD.n4645 VDD.n4644 34.6358
R15704 VDD.n4588 VDD.n3987 34.6358
R15705 VDD.n4574 VDD.n3994 34.6358
R15706 VDD.n4575 VDD.n4574 34.6358
R15707 VDD.n4570 VDD.n4567 34.6358
R15708 VDD.n4564 VDD.n3998 34.6358
R15709 VDD.n4556 VDD.n4002 34.6358
R15710 VDD.n4542 VDD.n4541 34.6358
R15711 VDD.n4534 VDD.n4017 34.6358
R15712 VDD.n4537 VDD.n4536 34.6358
R15713 VDD.n4472 VDD.n4471 34.6358
R15714 VDD.n4429 VDD.n4428 34.6358
R15715 VDD.n4409 VDD.n4408 34.6358
R15716 VDD.n4401 VDD.n4055 34.6358
R15717 VDD.n4405 VDD.n4055 34.6358
R15718 VDD.n4367 VDD.n4366 34.6358
R15719 VDD.n4364 VDD.n4079 34.6358
R15720 VDD.n4321 VDD.n4276 34.6358
R15721 VDD.n4331 VDD.n4330 34.6358
R15722 VDD.n4327 VDD.n4274 34.6358
R15723 VDD.n4323 VDD.n4274 34.6358
R15724 VDD.n4266 VDD.n4265 34.6358
R15725 VDD.n4238 VDD.n4115 34.6358
R15726 VDD.n4242 VDD.n4115 34.6358
R15727 VDD.n4199 VDD.n4198 34.6358
R15728 VDD.n3710 VDD.n3700 34.6358
R15729 VDD.n3716 VDD.n3715 34.6358
R15730 VDD.n3720 VDD.n3719 34.6358
R15731 VDD.n3726 VDD.n3725 34.6358
R15732 VDD.n3740 VDD.n3739 34.6358
R15733 VDD.n3739 VDD.n3738 34.6358
R15734 VDD.n3749 VDD.n3200 34.6358
R15735 VDD.n3664 VDD.n3663 34.6358
R15736 VDD.n3668 VDD.n3667 34.6358
R15737 VDD.n3661 VDD.n3210 34.6358
R15738 VDD.n3650 VDD.n3219 34.6358
R15739 VDD.n3640 VDD.n3223 34.6358
R15740 VDD.n3589 VDD.n3588 34.6358
R15741 VDD.n3589 VDD.n3227 34.6358
R15742 VDD.n3623 VDD.n3622 34.6358
R15743 VDD.n3533 VDD.n3255 34.6358
R15744 VDD.n3534 VDD.n3533 34.6358
R15745 VDD.n3535 VDD.n3534 34.6358
R15746 VDD.n3447 VDD.n3446 34.6358
R15747 VDD.n3453 VDD.n3452 34.6358
R15748 VDD.n3452 VDD.n3398 34.6358
R15749 VDD.n3390 VDD.n3385 34.6358
R15750 VDD.n3374 VDD.n3373 34.6358
R15751 VDD.n3378 VDD.n3377 34.6358
R15752 VDD.n3371 VDD.n3300 34.6358
R15753 VDD.n3364 VDD.n3303 34.6358
R15754 VDD.n3173 VDD.n3172 34.6358
R15755 VDD.n3177 VDD.n3106 34.6358
R15756 VDD.n3770 VDD.n3769 34.6358
R15757 VDD.n3774 VDD.n3773 34.6358
R15758 VDD.n3798 VDD.n3797 34.6358
R15759 VDD.n3805 VDD.n3804 34.6358
R15760 VDD.n3805 VDD.n3179 34.6358
R15761 VDD.n3846 VDD.n3845 34.6358
R15762 VDD.n3843 VDD.n3822 34.6358
R15763 VDD.n3839 VDD.n3822 34.6358
R15764 VDD.n3875 VDD.n3874 34.6358
R15765 VDD.n2867 VDD.n2866 34.6358
R15766 VDD.n2531 VDD.n2530 34.6358
R15767 VDD.n2535 VDD.n2534 34.6358
R15768 VDD.n2543 VDD.n2542 34.6358
R15769 VDD.n2542 VDD.n2507 34.6358
R15770 VDD.n2538 VDD.n2507 34.6358
R15771 VDD.n2356 VDD.n2355 34.6358
R15772 VDD.n3066 VDD.n2359 34.6358
R15773 VDD.n2950 VDD.n2949 34.6358
R15774 VDD.n2971 VDD.n2966 34.6358
R15775 VDD.n2977 VDD.n2976 34.6358
R15776 VDD.n2986 VDD.n2984 34.6358
R15777 VDD.n3084 VDD.n3083 34.6358
R15778 VDD.n3083 VDD.n2282 34.6358
R15779 VDD.n3072 VDD.n3071 34.6358
R15780 VDD.n2787 VDD.n2786 34.6358
R15781 VDD.n2748 VDD.n2747 34.6358
R15782 VDD.n2748 VDD.n2456 34.6358
R15783 VDD.n2752 VDD.n2456 34.6358
R15784 VDD.n2741 VDD.n2740 34.6358
R15785 VDD.n2729 VDD.n2728 34.6358
R15786 VDD.n2602 VDD.n2601 34.6358
R15787 VDD.n2631 VDD.n2630 34.6358
R15788 VDD.n2637 VDD.n2636 34.6358
R15789 VDD.n2649 VDD.n2648 34.6358
R15790 VDD.n2724 VDD.n2474 34.6358
R15791 VDD.n2719 VDD.n2718 34.6358
R15792 VDD.n2718 VDD.n2653 34.6358
R15793 VDD.n2692 VDD.n2691 34.6358
R15794 VDD.n2686 VDD.n2685 34.6358
R15795 VDD.n2685 VDD.n2672 34.6358
R15796 VDD.n2681 VDD.n2672 34.6358
R15797 VDD.n2333 VDD.n2332 34.6358
R15798 VDD.n2332 VDD.n2331 34.6358
R15799 VDD.n2058 VDD.n2056 34.6358
R15800 VDD.n2041 VDD.n2040 34.6358
R15801 VDD.n2035 VDD.n2034 34.6358
R15802 VDD.n1987 VDD.n1971 34.6358
R15803 VDD.n2004 VDD.n2003 34.6358
R15804 VDD.n2007 VDD.n1960 34.6358
R15805 VDD.n1788 VDD.n1784 34.6358
R15806 VDD.n1792 VDD.n1638 34.6358
R15807 VDD.n1796 VDD.n1794 34.6358
R15808 VDD.n1782 VDD.n1642 34.6358
R15809 VDD.n1770 VDD.n1648 34.6358
R15810 VDD.n1753 VDD.n1657 34.6358
R15811 VDD.n1747 VDD.n1746 34.6358
R15812 VDD.n1747 VDD.n1661 34.6358
R15813 VDD.n1751 VDD.n1661 34.6358
R15814 VDD.n2090 VDD.n1528 34.6358
R15815 VDD.n2110 VDD.n2109 34.6358
R15816 VDD.n2013 VDD.n2012 34.6358
R15817 VDD.n2026 VDD.n2025 34.6358
R15818 VDD.n1931 VDD.n1567 34.6358
R15819 VDD.n1935 VDD.n1567 34.6358
R15820 VDD.n1936 VDD.n1935 34.6358
R15821 VDD.n1937 VDD.n1936 34.6358
R15822 VDD.n2165 VDD.n2164 34.6358
R15823 VDD.n2151 VDD.n2133 34.6358
R15824 VDD.n2147 VDD.n2146 34.6358
R15825 VDD.n2144 VDD.n2141 34.6358
R15826 VDD.n2240 VDD.n2176 34.6358
R15827 VDD.n2236 VDD.n2235 34.6358
R15828 VDD.n2229 VDD.n2228 34.6358
R15829 VDD.n2225 VDD.n2186 34.6358
R15830 VDD.n2219 VDD.n2189 34.6358
R15831 VDD.n2215 VDD.n2189 34.6358
R15832 VDD.n1116 VDD.n798 34.6358
R15833 VDD.n1120 VDD.n798 34.6358
R15834 VDD.n1113 VDD.n1112 34.6358
R15835 VDD.n1107 VDD.n1106 34.6358
R15836 VDD.n1108 VDD.n1107 34.6358
R15837 VDD.n1092 VDD.n1091 34.6358
R15838 VDD.n1081 VDD.n815 34.6358
R15839 VDD.n1030 VDD.n1029 34.6358
R15840 VDD.n1045 VDD.n1044 34.6358
R15841 VDD.n1050 VDD.n1049 34.6358
R15842 VDD.n1058 VDD.n1057 34.6358
R15843 VDD.n1064 VDD.n1063 34.6358
R15844 VDD.n1000 VDD.n999 34.6358
R15845 VDD.n995 VDD.n994 34.6358
R15846 VDD.n996 VDD.n995 34.6358
R15847 VDD.n991 VDD.n988 34.6358
R15848 VDD.n981 VDD.n831 34.6358
R15849 VDD.n985 VDD.n831 34.6358
R15850 VDD.n930 VDD.n885 34.6358
R15851 VDD.n940 VDD.n880 34.6358
R15852 VDD.n876 VDD.n849 34.6358
R15853 VDD.n1352 VDD.n1351 34.6358
R15854 VDD.n1340 VDD.n1339 34.6358
R15855 VDD.n1316 VDD.n1315 34.6358
R15856 VDD.n1319 VDD.n1316 34.6358
R15857 VDD.n1323 VDD.n729 34.6358
R15858 VDD.n1305 VDD.n735 34.6358
R15859 VDD.n1309 VDD.n735 34.6358
R15860 VDD.n1295 VDD.n1294 34.6358
R15861 VDD.n1296 VDD.n1295 34.6358
R15862 VDD.n1296 VDD.n742 34.6358
R15863 VDD.n1300 VDD.n742 34.6358
R15864 VDD.n1287 VDD.n748 34.6358
R15865 VDD.n1229 VDD.n773 34.6358
R15866 VDD.n1230 VDD.n1229 34.6358
R15867 VDD.n1223 VDD.n1222 34.6358
R15868 VDD.n1194 VDD.n791 34.6358
R15869 VDD.n1186 VDD.n1185 34.6358
R15870 VDD.n1180 VDD.n1179 34.6358
R15871 VDD.n1176 VDD.n1140 34.6358
R15872 VDD.n1157 VDD.n1156 34.6358
R15873 VDD.n1202 VDD.n787 34.6358
R15874 VDD.n1206 VDD.n785 34.6358
R15875 VDD.n1402 VDD.n1358 34.6358
R15876 VDD.n1390 VDD.n1389 34.6358
R15877 VDD.n1496 VDD.n703 34.6358
R15878 VDD.n1463 VDD.n1462 34.6358
R15879 VDD.n1460 VDD.n1418 34.6358
R15880 VDD.n624 VDD.n623 34.6358
R15881 VDD.n628 VDD.n627 34.6358
R15882 VDD.n629 VDD.n628 34.6358
R15883 VDD.n633 VDD.n632 34.6358
R15884 VDD.n690 VDD.n689 34.6358
R15885 VDD.n684 VDD.n683 34.6358
R15886 VDD.n683 VDD.n682 34.6358
R15887 VDD.n679 VDD.n678 34.6358
R15888 VDD.n673 VDD.n672 34.6358
R15889 VDD.n670 VDD.n652 34.6358
R15890 VDD.n666 VDD.n665 34.6358
R15891 VDD.n541 VDD.n540 34.6358
R15892 VDD.n545 VDD.n544 34.6358
R15893 VDD.n546 VDD.n545 34.6358
R15894 VDD.n550 VDD.n549 34.6358
R15895 VDD.n602 VDD.n601 34.6358
R15896 VDD.n599 VDD.n554 34.6358
R15897 VDD.n595 VDD.n554 34.6358
R15898 VDD.n595 VDD.n594 34.6358
R15899 VDD.n592 VDD.n557 34.6358
R15900 VDD.n586 VDD.n585 34.6358
R15901 VDD.n582 VDD.n581 34.6358
R15902 VDD.n579 VDD.n566 34.6358
R15903 VDD.n461 VDD.n460 34.6358
R15904 VDD.n465 VDD.n464 34.6358
R15905 VDD.n466 VDD.n465 34.6358
R15906 VDD.n470 VDD.n469 34.6358
R15907 VDD.n522 VDD.n521 34.6358
R15908 VDD.n519 VDD.n474 34.6358
R15909 VDD.n515 VDD.n474 34.6358
R15910 VDD.n515 VDD.n514 34.6358
R15911 VDD.n512 VDD.n477 34.6358
R15912 VDD.n506 VDD.n505 34.6358
R15913 VDD.n502 VDD.n501 34.6358
R15914 VDD.n499 VDD.n486 34.6358
R15915 VDD.n425 VDD.n424 34.6358
R15916 VDD.n140 VDD.n132 34.6358
R15917 VDD.n3214 VDD.t3299 34.4755
R15918 VDD.n3251 VDD.t3291 34.4755
R15919 VDD.n3413 VDD.t1794 34.4755
R15920 VDD.n3413 VDD.t1956 34.4755
R15921 VDD.n3409 VDD.t2379 34.4755
R15922 VDD.n3816 VDD.t54 34.4755
R15923 VDD.n3826 VDD.t728 34.4755
R15924 VDD.n2395 VDD.t3289 34.4755
R15925 VDD.n2395 VDD.t1100 34.4755
R15926 VDD.n2396 VDD.t1481 34.4755
R15927 VDD.n2369 VDD.t3469 34.4755
R15928 VDD.n2463 VDD.t3731 34.4755
R15929 VDD.n2472 VDD.t3293 34.4755
R15930 VDD.n2662 VDD.t3727 34.4755
R15931 VDD.n1605 VDD.t3301 34.4755
R15932 VDD.n1645 VDD.t3014 34.4755
R15933 VDD.n1591 VDD.t3295 34.4755
R15934 VDD.n1942 VDD.t3461 34.4755
R15935 VDD.n1559 VDD.t3285 34.4755
R15936 VDD.n2135 VDD.t3459 34.4755
R15937 VDD.n2135 VDD.t685 34.4755
R15938 VDD.n807 VDD.t3018 34.4755
R15939 VDD.n1005 VDD.t2099 34.4755
R15940 VDD.n734 VDD.t3479 34.4755
R15941 VDD.n738 VDD.t3473 34.4755
R15942 VDD.n747 VDD.t3475 34.4755
R15943 VDD.n1274 VDD.t2095 34.4755
R15944 VDD.n765 VDD.t2093 34.4755
R15945 VDD.n1129 VDD.t3012 34.4755
R15946 VDD.n1149 VDD.t3020 34.4755
R15947 VDD.n702 VDD.t2097 34.4755
R15948 VDD.n709 VDD.t2101 34.4755
R15949 VDD.n658 VDD.t3077 34.4755
R15950 VDD.n657 VDD.t2079 34.4755
R15951 VDD.n650 VDD.t3612 34.4755
R15952 VDD.n615 VDD.t1049 34.4755
R15953 VDD.n614 VDD.t1374 34.4755
R15954 VDD.n635 VDD.t720 34.4755
R15955 VDD.n532 VDD.t2650 34.4755
R15956 VDD.n531 VDD.t400 34.4755
R15957 VDD.n553 VDD.t885 34.4755
R15958 VDD.n552 VDD.t2161 34.4755
R15959 VDD.n563 VDD.t3229 34.4755
R15960 VDD.n562 VDD.t3605 34.4755
R15961 VDD.n573 VDD.t2920 34.4755
R15962 VDD.n572 VDD.t1971 34.4755
R15963 VDD.n452 VDD.t1152 34.4755
R15964 VDD.n451 VDD.t709 34.4755
R15965 VDD.n473 VDD.t286 34.4755
R15966 VDD.n472 VDD.t1615 34.4755
R15967 VDD.n483 VDD.t2957 34.4755
R15968 VDD.n482 VDD.t3765 34.4755
R15969 VDD.n493 VDD.t3760 34.4755
R15970 VDD.n492 VDD.t3095 34.4755
R15971 VDD.n3946 VDD.n3927 34.2593
R15972 VDD.n2104 VDD.n2102 34.2593
R15973 VDD.n1941 VDD.n1565 34.2593
R15974 VDD.n2152 VDD.n2151 34.2593
R15975 VDD.n2254 VDD.n1515 34.2593
R15976 VDD.n1059 VDD.n1058 34.2593
R15977 VDD.n627 VDD.n616 34.2593
R15978 VDD.n688 VDD.n687 34.2593
R15979 VDD.n663 VDD.n659 34.2593
R15980 VDD.n544 VDD.n533 34.2593
R15981 VDD.n600 VDD.n599 34.2593
R15982 VDD.n588 VDD.n587 34.2593
R15983 VDD.n575 VDD.n574 34.2593
R15984 VDD.n464 VDD.n453 34.2593
R15985 VDD.n520 VDD.n519 34.2593
R15986 VDD.n508 VDD.n507 34.2593
R15987 VDD.n495 VDD.n494 34.2593
R15988 VDD.n4290 VDD.t811 34.0906
R15989 VDD.n4112 VDD.t456 34.0906
R15990 VDD.n4144 VDD.t1266 34.0906
R15991 VDD.n4147 VDD.t2270 34.0906
R15992 VDD.n4155 VDD.t1683 34.0906
R15993 VDD.n4159 VDD.t2562 34.0906
R15994 VDD.n4160 VDD.t945 34.0906
R15995 VDD.n3959 VDD.t1172 34.0906
R15996 VDD.n3918 VDD.t3329 34.0906
R15997 VDD.n3921 VDD.t846 34.0906
R15998 VDD.n3922 VDD.t576 34.0906
R15999 VDD.n3929 VDD.t1132 34.0906
R16000 VDD.n3704 VDD.t1335 34.0906
R16001 VDD.n3315 VDD.t1331 34.0906
R16002 VDD.n3316 VDD.t1433 34.0906
R16003 VDD.n3762 VDD.t2695 34.0906
R16004 VDD.n3323 VDD.t2285 34.0906
R16005 VDD.n3325 VDD.t2211 34.0906
R16006 VDD.n3326 VDD.t476 34.0906
R16007 VDD.n3126 VDD.t1731 34.0906
R16008 VDD.n3128 VDD.t2526 34.0906
R16009 VDD.n3131 VDD.t1408 34.0906
R16010 VDD.n3132 VDD.t2568 34.0906
R16011 VDD.n2515 VDD.t2150 34.0906
R16012 VDD.n2562 VDD.t1229 34.0906
R16013 VDD.n2573 VDD.t594 34.0906
R16014 VDD.n2575 VDD.t577 34.0906
R16015 VDD.n2576 VDD.t396 34.0906
R16016 VDD.n2308 VDD.t1160 34.0906
R16017 VDD.n2310 VDD.t258 34.0906
R16018 VDD.n2311 VDD.t2168 34.0906
R16019 VDD.n1653 VDD.t745 34.0906
R16020 VDD.n1676 VDD.t949 34.0906
R16021 VDD.n1681 VDD.t2144 34.0906
R16022 VDD.n1683 VDD.t1277 34.0906
R16023 VDD.n1684 VDD.t1561 34.0906
R16024 VDD.n1687 VDD.t2535 34.0906
R16025 VDD.n1691 VDD.t1170 34.0906
R16026 VDD.n1692 VDD.t2431 34.0906
R16027 VDD.n1954 VDD.t895 34.0906
R16028 VDD.n2138 VDD.t1126 34.0906
R16029 VDD.n2192 VDD.t2216 34.0906
R16030 VDD.n2194 VDD.t460 34.0906
R16031 VDD.n2195 VDD.t290 34.0906
R16032 VDD.n795 VDD.t454 34.0906
R16033 VDD.n813 VDD.t2771 34.0906
R16034 VDD.n1007 VDD.t558 34.0906
R16035 VDD.n839 VDD.t2182 34.0906
R16036 VDD.n843 VDD.t264 34.0906
R16037 VDD.n900 VDD.t2220 34.0906
R16038 VDD.n896 VDD.t1727 34.0906
R16039 VDD.n889 VDD.t2790 34.0906
R16040 VDD.n931 VDD.t2809 34.0906
R16041 VDD.n881 VDD.t1440 34.0906
R16042 VDD.n855 VDD.t3333 34.0906
R16043 VDD.n723 VDD.t48 34.0906
R16044 VDD.n750 VDD.t2858 34.0906
R16045 VDD.n762 VDD.t911 34.0906
R16046 VDD.n779 VDD.t1402 34.0906
R16047 VDD.n1142 VDD.t2414 34.0906
R16048 VDD.n1360 VDD.t272 34.0906
R16049 VDD.n1368 VDD.t984 34.0906
R16050 VDD.n1371 VDD.t774 34.0906
R16051 VDD.n1409 VDD.t2556 34.0906
R16052 VDD.n1417 VDD.t901 34.0906
R16053 VDD.n1422 VDD.t314 34.0906
R16054 VDD.n1426 VDD.t2824 34.0906
R16055 VDD.n1427 VDD.t2448 34.0906
R16056 VDD.n1430 VDD.t1356 34.0906
R16057 VDD.n1431 VDD.t928 34.0906
R16058 VDD.n4620 VDD.n4619 33.8829
R16059 VDD.n4577 VDD.n4576 33.8829
R16060 VDD.n4496 VDD.n4495 33.8829
R16061 VDD.n3746 VDD.n3745 33.8829
R16062 VDD.n3667 VDD.n3206 33.8829
R16063 VDD.n3597 VDD.n3596 33.8829
R16064 VDD.n3427 VDD.n3426 33.8829
R16065 VDD.n3442 VDD.n3441 33.8829
R16066 VDD.n3377 VDD.n3297 33.8829
R16067 VDD.n3860 VDD.n3810 33.8829
R16068 VDD.n3869 VDD.n3104 33.8829
R16069 VDD.n2922 VDD.n2921 33.8829
R16070 VDD.n3068 VDD.n2286 33.8829
R16071 VDD.n2687 VDD.n2686 33.8829
R16072 VDD.n2678 VDD.n2677 33.8829
R16073 VDD.n2063 VDD.n2062 33.8829
R16074 VDD.n2040 VDD.n1553 33.8829
R16075 VDD.n1842 VDD.n1606 33.8829
R16076 VDD.n1708 VDD.n1707 33.8829
R16077 VDD.n2156 VDD.n2130 33.8829
R16078 VDD.n2257 VDD.n2256 33.8829
R16079 VDD.n981 VDD.n980 33.8829
R16080 VDD.n895 VDD.n892 33.8829
R16081 VDD.n919 VDD.n890 33.8829
R16082 VDD.n872 VDD.n853 33.8829
R16083 VDD.n1332 VDD.n1331 33.8829
R16084 VDD.n1395 VDD.n1362 33.8829
R16085 VDD.n3497 VDD.n3496 33.6462
R16086 VDD.n3479 VDD.n3478 33.6462
R16087 VDD.n2901 VDD.n2900 33.6462
R16088 VDD.n2897 VDD.n2413 33.6462
R16089 VDD.n3000 VDD.n2997 33.6462
R16090 VDD.n3063 VDD.n2360 33.6462
R16091 VDD.n3060 VDD.n3059 33.6462
R16092 VDD.n2893 VDD.n2418 33.6462
R16093 VDD.n2822 VDD.n2821 33.6462
R16094 VDD.n2820 VDD.n2422 33.6462
R16095 VDD.n1832 VDD.n1831 33.6462
R16096 VDD.n1828 VDD.n1825 33.6462
R16097 VDD.n1816 VDD.n1625 33.6462
R16098 VDD.t3184 VDD.t2171 33.5694
R16099 VDD.t1923 VDD.t942 33.5694
R16100 VDD.t874 VDD.t501 33.5694
R16101 VDD.t1026 VDD.t1882 33.5694
R16102 VDD.t3493 VDD.t1006 33.5694
R16103 VDD.t2041 VDD.t3190 33.5694
R16104 VDD.t2867 VDD.t3677 33.5694
R16105 VDD.t729 VDD.t1636 33.5694
R16106 VDD.t1652 VDD.t2600 33.5694
R16107 VDD.t1523 VDD.t1271 33.5694
R16108 VDD.t3531 VDD.t3437 33.5694
R16109 VDD.n4204 VDD.n4132 33.5064
R16110 VDD.n3645 VDD.n3219 33.5064
R16111 VDD.n3594 VDD.n3588 33.5064
R16112 VDD.n3621 VDD.n3575 33.5064
R16113 VDD.n3764 VDD.n3195 33.5064
R16114 VDD.n2951 VDD.n2950 33.5064
R16115 VDD.n2792 VDD.n2437 33.5064
R16116 VDD.n2788 VDD.n2787 33.5064
R16117 VDD.n1847 VDD.n1846 33.5064
R16118 VDD.n1738 VDD.n1737 33.5064
R16119 VDD.n677 VDD.n676 33.5064
R16120 VDD.n664 VDD.n663 33.5064
R16121 VDD.n588 VDD.n561 33.5064
R16122 VDD.n575 VDD.n571 33.5064
R16123 VDD.n508 VDD.n481 33.5064
R16124 VDD.n495 VDD.n491 33.5064
R16125 VDD.n3214 VDD.t2591 33.4905
R16126 VDD.n3251 VDD.t2300 33.4905
R16127 VDD.n3409 VDD.t3521 33.4905
R16128 VDD.n3816 VDD.t2472 33.4905
R16129 VDD.n3826 VDD.t3509 33.4905
R16130 VDD.n2369 VDD.t566 33.4905
R16131 VDD.n2463 VDD.t2850 33.4905
R16132 VDD.n2662 VDD.t1388 33.4905
R16133 VDD.n1559 VDD.t296 33.4905
R16134 VDD.n738 VDD.t1424 33.4905
R16135 VDD.n2906 VDD.n2905 33.2805
R16136 VDD.n3644 VDD.n3643 33.1299
R16137 VDD.n3510 VDD.n3509 33.1299
R16138 VDD.n3394 VDD.n3291 33.1299
R16139 VDD.n3379 VDD.n3378 33.1299
R16140 VDD.n3513 VDD.n3512 33.1299
R16141 VDD.n3406 VDD.n3404 33.1299
R16142 VDD.n2642 VDD.n2641 33.1299
R16143 VDD.n2697 VDD.n2665 33.1299
R16144 VDD.n1741 VDD.n1664 33.1299
R16145 VDD.n1711 VDD.n1710 33.1299
R16146 VDD.n1391 VDD.n1390 33.1299
R16147 VDD.n245 VDD.t2038 33.0605
R16148 VDD.n245 VDD.t3403 33.0605
R16149 VDD.n2889 VDD.n2888 32.9148
R16150 VDD.n1999 VDD.n1998 32.7534
R16151 VDD.n1335 VDD.n1334 32.7534
R16152 VDD.n433 VDD.n432 32.7534
R16153 VDD.n243 VDD.n242 32.6405
R16154 VDD.n3217 VDD.t959 32.5055
R16155 VDD.n3217 VDD.t517 32.5055
R16156 VDD.n3252 VDD.t3305 32.5055
R16157 VDD.n3252 VDD.t3623 32.5055
R16158 VDD.n3428 VDD.t1194 32.5055
R16159 VDD.n3428 VDD.t1694 32.5055
R16160 VDD.n3814 VDD.t1798 32.5055
R16161 VDD.n3814 VDD.t825 32.5055
R16162 VDD.n3824 VDD.t2091 32.5055
R16163 VDD.n3824 VDD.t2724 32.5055
R16164 VDD.n2373 VDD.t440 32.5055
R16165 VDD.n2373 VDD.t1930 32.5055
R16166 VDD.n2466 VDD.t1365 32.5055
R16167 VDD.n2466 VDD.t243 32.5055
R16168 VDD.n2657 VDD.t3644 32.5055
R16169 VDD.n2657 VDD.t3026 32.5055
R16170 VDD.n2660 VDD.t3665 32.5055
R16171 VDD.n2660 VDD.t3106 32.5055
R16172 VDD.n2083 VDD.t3050 32.5055
R16173 VDD.n1523 VDD.t3049 32.5055
R16174 VDD.n1949 VDD.t963 32.5055
R16175 VDD.n1949 VDD.t3271 32.5055
R16176 VDD.n739 VDD.t426 32.5055
R16177 VDD.n739 VDD.t2908 32.5055
R16178 VDD.n645 VDD.n643 32.4617
R16179 VDD.n4614 VDD.n4611 32.377
R16180 VDD.n4641 VDD.n4601 32.377
R16181 VDD.n4577 VDD.n3991 32.377
R16182 VDD.n4552 VDD.n4551 32.377
R16183 VDD.n4537 VDD.n4014 32.377
R16184 VDD.n4469 VDD.n4452 32.377
R16185 VDD.n4399 VDD.n4398 32.377
R16186 VDD.n2353 VDD.n2292 32.377
R16187 VDD.n2952 VDD.n2382 32.377
R16188 VDD.n1728 VDD.n1679 32.377
R16189 VDD.n2086 VDD.n2085 32.377
R16190 VDD.n986 VDD.n985 32.377
R16191 VDD.n946 VDD.n945 32.377
R16192 VDD.n876 VDD.n875 32.377
R16193 VDD.n873 VDD.n872 32.377
R16194 VDD.n1342 VDD.n721 32.377
R16195 VDD.n1231 VDD.n1230 32.377
R16196 VDD.n1186 VDD.n1133 32.377
R16197 VDD.n672 VDD.n671 32.377
R16198 VDD.n585 VDD.n564 32.377
R16199 VDD.n505 VDD.n484 32.377
R16200 VDD.n2919 VDD.n2402 32.377
R16201 VDD.n2704 VDD.n2703 32.377
R16202 VDD.n1842 VDD.n1841 32.377
R16203 VDD.n1951 VDD.n1560 32.377
R16204 VDD.n1304 VDD.n1303 32.377
R16205 VDD.n4294 VDD.n4293 32.0005
R16206 VDD.n4323 VDD.n4322 32.0005
R16207 VDD.n3942 VDD.n3941 32.0005
R16208 VDD.n3708 VDD.n3707 32.0005
R16209 VDD.n3740 VDD.n3685 32.0005
R16210 VDD.n3448 VDD.n3398 32.0005
R16211 VDD.n3367 VDD.n3366 32.0005
R16212 VDD.n3169 VDD.n3117 32.0005
R16213 VDD.n2328 VDD.n2309 32.0005
R16214 VDD.n1763 VDD.n1654 32.0005
R16215 VDD.n1724 VDD.n1723 32.0005
R16216 VDD.n2233 VDD.n2182 32.0005
R16217 VDD.n2213 VDD.n2212 32.0005
R16218 VDD.n1108 VDD.n802 32.0005
R16219 VDD.n1087 VDD.n1086 32.0005
R16220 VDD.n1072 VDD.n1071 32.0005
R16221 VDD.n912 VDD.n911 32.0005
R16222 VDD.n925 VDD.n924 32.0005
R16223 VDD.n868 VDD.n867 32.0005
R16224 VDD.n1218 VDD.n1217 32.0005
R16225 VDD.n430 VDD.n348 32.0005
R16226 VDD.t98 VDD.t2207 31.891
R16227 VDD.t94 VDD.t1909 31.891
R16228 VDD.t2473 VDD.t3424 31.891
R16229 VDD.t3322 VDD.t1413 31.891
R16230 VDD.t2785 VDD.t1399 31.891
R16231 VDD.t3629 VDD.t797 31.891
R16232 VDD.t1627 VDD.n3468 31.891
R16233 VDD.t1018 VDD.t1272 31.891
R16234 VDD.t303 VDD.t2380 31.891
R16235 VDD.n2029 VDD.t2438 31.891
R16236 VDD.t51 VDD.t1490 31.891
R16237 VDD.t832 VDD.t2480 31.891
R16238 VDD.t271 VDD.t696 31.891
R16239 VDD.n3057 VDD.n3006 31.8176
R16240 VDD.n2092 VDD.n1526 31.624
R16241 VDD.n3703 VDD.t3477 31.5205
R16242 VDD.n3209 VDD.t1349 31.5205
R16243 VDD.n3578 VDD.t3297 31.5205
R16244 VDD.n2364 VDD.t2776 31.5205
R16245 VDD.n2831 VDD.t3287 31.5205
R16246 VDD.n3025 VDD.t3465 31.5205
R16247 VDD.n244 VDD.n223 31.4672
R16248 VDD.n186 VDD.t3597 31.2992
R16249 VDD.n1018 VDD.n1015 31.2476
R16250 VDD.n623 VDD.n622 31.2476
R16251 VDD.n690 VDD.n634 31.2476
R16252 VDD.n540 VDD.n539 31.2476
R16253 VDD.n602 VDD.n551 31.2476
R16254 VDD.n460 VDD.n459 31.2476
R16255 VDD.n522 VDD.n471 31.2476
R16256 VDD.n185 VDD.t3593 31.2448
R16257 VDD.n186 VDD.t3596 30.9042
R16258 VDD.n3941 VDD.n3940 30.8711
R16259 VDD.n2986 VDD.n2985 30.8711
R16260 VDD.n1848 VDD.n1847 30.8711
R16261 VDD.n1772 VDD.n1646 30.8711
R16262 VDD.n1759 VDD.n1758 30.8711
R16263 VDD.n1094 VDD.n808 30.8711
R16264 VDD.n1006 VDD.n818 30.8711
R16265 VDD.n1276 VDD.n1275 30.8711
R16266 VDD.n1784 VDD.n1783 30.8711
R16267 VDD.n1753 VDD.n1752 30.8711
R16268 VDD.n185 VDD.t3594 30.8498
R16269 VDD.n420 VDD.n419 30.8338
R16270 VDD.n421 VDD.n420 30.8338
R16271 VDD.n358 VDD.n354 30.8338
R16272 VDD.n421 VDD.n354 30.8338
R16273 VDD.n374 VDD.n373 30.8338
R16274 VDD.n375 VDD.n374 30.8338
R16275 VDD.n382 VDD.n379 30.8338
R16276 VDD.n379 VDD.n375 30.8338
R16277 VDD.n3499 VDD.n3270 30.7205
R16278 VDD.n2083 VDD.t3001 30.5355
R16279 VDD.n1523 VDD.t3256 30.5355
R16280 VDD.n4357 VDD.n4356 30.4946
R16281 VDD.n867 VDD.n866 30.4946
R16282 VDD.t69 VDD.t58 30.2868
R16283 VDD.t58 VDD.t65 30.2868
R16284 VDD.t65 VDD.t62 30.2868
R16285 VDD.t59 VDD.t63 30.2868
R16286 VDD.t60 VDD.t59 30.2868
R16287 VDD.t71 VDD.t60 30.2868
R16288 VDD.t61 VDD.t67 30.2868
R16289 VDD.t57 VDD.t61 30.2868
R16290 VDD.t70 VDD.t57 30.2868
R16291 VDD.t66 VDD.t64 30.2868
R16292 VDD.t64 VDD.t68 30.2868
R16293 VDD.t68 VDD.t72 30.2868
R16294 VDD.t3192 VDD.t2175 30.2125
R16295 VDD.t3088 VDD.t2886 30.2125
R16296 VDD.t2841 VDD.t2111 30.2125
R16297 VDD.t1338 VDD.t3383 30.2125
R16298 VDD.t2783 VDD.t2509 30.2125
R16299 VDD.t2727 VDD.t3499 30.2125
R16300 VDD.t3764 VDD.t1346 30.2125
R16301 VDD.t2346 VDD.t1059 30.2125
R16302 VDD.t2723 VDD.t3640 30.2125
R16303 VDD.n2727 VDD.t238 30.2125
R16304 VDD.t605 VDD.t1699 30.2125
R16305 VDD.t3280 VDD.t277 30.2125
R16306 VDD.t518 VDD.t1258 30.2125
R16307 VDD.t1261 VDD.t3720 30.2125
R16308 VDD.t1307 VDD.t2861 30.2125
R16309 VDD.t2903 VDD.t212 30.2125
R16310 VDD.t898 VDD.t586 30.2125
R16311 VDD.n2247 VDD.n2174 30.1181
R16312 VDD.n1476 VDD.n1475 30.1181
R16313 VDD.n75 VDD.n72 30.1181
R16314 VDD.n32 VDD.n31 30.1181
R16315 VDD.n3517 VDD.n3516 30.1181
R16316 VDD.n2525 VDD.n2523 30.1181
R16317 VDD.n1980 VDD.n1979 30.1181
R16318 VDD.n1802 VDD.n1801 30.1181
R16319 VDD.n1038 VDD.n1020 30.1181
R16320 VDD.n1211 VDD.n782 30.1181
R16321 VDD.n1170 VDD.n1169 30.1181
R16322 VDD.n172 VDD.n171 29.8672
R16323 VDD.n3388 VDD.n3292 29.7417
R16324 VDD.n2349 VDD.n2348 29.7417
R16325 VDD.n2637 VDD.n2480 29.7417
R16326 VDD.n1101 VDD.n805 29.7417
R16327 VDD.n2816 VDD.n2813 29.6234
R16328 VDD.n897 VDD.t3022 29.5505
R16329 VDD.n897 VDD.t998 29.5505
R16330 VDD.n287 VDD.t3583 29.4286
R16331 VDD.n222 VDD.t3589 29.4286
R16332 VDD.n251 VDD.t3599 29.4286
R16333 VDD.n254 VDD.t3579 29.4286
R16334 VDD.n258 VDD.t3601 29.4286
R16335 VDD.n263 VDD.t3587 29.4286
R16336 VDD.n266 VDD.t3577 29.4286
R16337 VDD.n270 VDD.t3591 29.4286
R16338 VDD.n275 VDD.t3603 29.4286
R16339 VDD.n278 VDD.t3581 29.4286
R16340 VDD.n282 VDD.t3585 29.4286
R16341 VDD.n3535 VDD.n3253 29.3652
R16342 VDD.n2982 VDD.n2981 29.3652
R16343 VDD.n2707 VDD.n2706 29.3652
R16344 VDD.n2005 VDD.n2004 29.3652
R16345 VDD.n1852 VDD.n1603 29.3652
R16346 VDD.n3484 VDD.n3483 29.2576
R16347 VDD.n2848 VDD.n2844 29.2576
R16348 VDD.n1818 VDD.n1817 29.2576
R16349 VDD.n973 VDD.n967 29.1064
R16350 VDD.n4349 VDD.n4085 28.9887
R16351 VDD.n2928 VDD.n2927 28.9887
R16352 VDD.n1944 VDD.n1943 28.9887
R16353 VDD.n1311 VDD.n1310 28.9887
R16354 VDD.n666 VDD.n654 28.9887
R16355 VDD.n593 VDD.n592 28.9887
R16356 VDD.n580 VDD.n579 28.9887
R16357 VDD.n513 VDD.n512 28.9887
R16358 VDD.n500 VDD.n499 28.9887
R16359 VDD.n3482 VDD.n3284 28.8919
R16360 VDD.n2886 VDD.n2885 28.8919
R16361 VDD.n3904 VDD.t1548 28.752
R16362 VDD.n4590 VDD.t1714 28.752
R16363 VDD.n3993 VDD.t665 28.752
R16364 VDD.n4012 VDD.t1593 28.752
R16365 VDD.n4513 VDD.t2848 28.752
R16366 VDD.n4084 VDD.t1623 28.752
R16367 VDD.n4279 VDD.t1585 28.752
R16368 VDD.n3701 VDD.t589 28.752
R16369 VDD.n3684 VDD.t2383 28.752
R16370 VDD.n3205 VDD.t842 28.752
R16371 VDD.n3587 VDD.t766 28.752
R16372 VDD.n3573 VDD.t1200 28.752
R16373 VDD.n3296 VDD.t2490 28.752
R16374 VDD.n3809 VDD.t1386 28.752
R16375 VDD.n3825 VDD.t350 28.752
R16376 VDD.n3103 VDD.t2811 28.752
R16377 VDD.n2846 VDD.t3494 28.752
R16378 VDD.n2285 VDD.t1231 28.752
R16379 VDD.n2455 VDD.t2230 28.752
R16380 VDD.n2675 VDD.t534 28.752
R16381 VDD.n733 VDD.t2308 28.752
R16382 VDD.n4263 VDD.n4262 28.6123
R16383 VDD.t2253 VDD.t2126 28.5341
R16384 VDD.t906 VDD.t1211 28.5341
R16385 VDD.t1220 VDD.t3257 28.5341
R16386 VDD.t664 VDD.t1684 28.5341
R16387 VDD.t643 VDD.t1366 28.5341
R16388 VDD.t2830 VDD.t970 28.5341
R16389 VDD.t439 VDD.t670 28.5341
R16390 VDD.t694 VDD.t2103 28.5341
R16391 VDD.t3745 VDD.t582 28.5341
R16392 VDD.t3478 VDD.t3533 28.5341
R16393 VDD.n1613 VDD.t4 28.5169
R16394 VDD.n3910 VDD.t638 28.4453
R16395 VDD.n4449 VDD.t2542 28.4453
R16396 VDD.n4053 VDD.t2546 28.4453
R16397 VDD.n4358 VDD.t2528 28.4453
R16398 VDD.n2908 VDD.t1273 28.4453
R16399 VDD.n2288 VDD.t2263 28.4453
R16400 VDD.n2137 VDD.t3519 28.4453
R16401 VDD.n887 VDD.t2291 28.4453
R16402 VDD.n938 VDD.t1148 28.4453
R16403 VDD.n4042 VDD.t1233 28.4453
R16404 VDD.n3697 VDD.t1136 28.4453
R16405 VDD.n3192 VDD.t2726 28.4453
R16406 VDD.n2491 VDD.t2676 28.4453
R16407 VDD.n4560 VDD.n3998 28.2358
R16408 VDD.n4519 VDD.n4032 28.2358
R16409 VDD.n4506 VDD.n4035 28.2358
R16410 VDD.n4379 VDD.n4074 28.2358
R16411 VDD.n1999 VDD.n1965 28.2358
R16412 VDD.n1855 VDD.n1854 28.2358
R16413 VDD.n2963 VDD.n2380 28.2358
R16414 VDD.n4637 VDD.n4636 27.8593
R16415 VDD.n4526 VDD.n4525 27.8593
R16416 VDD.n4497 VDD.n4039 27.8593
R16417 VDD.n4258 VDD.n4257 27.8593
R16418 VDD.n3868 VDD.n3867 27.8593
R16419 VDD.n1983 VDD.n1973 27.8593
R16420 VDD.n2250 VDD.n2249 27.8593
R16421 VDD.n1099 VDD.n1098 27.8593
R16422 VDD.n1036 VDD.n1035 27.8593
R16423 VDD.n1044 VDD.n1043 27.8593
R16424 VDD.n906 VDD.n898 27.8593
R16425 VDD.n1166 VDD.n1165 27.8593
R16426 VDD.n1479 VDD.n710 27.8593
R16427 VDD.n432 VDD.n431 27.8593
R16428 VDD.n977 VDD.n835 27.724
R16429 VDD.n679 VDD.n639 27.7228
R16430 VDD.n4612 VDD.t3500 27.5805
R16431 VDD.n4610 VDD.t2316 27.5805
R16432 VDD.n4610 VDD.t2312 27.5805
R16433 VDD.n4600 VDD.t2359 27.5805
R16434 VDD.n4598 VDD.t2117 27.5805
R16435 VDD.n4598 VDD.t2119 27.5805
R16436 VDD.n4549 VDD.t1622 27.5805
R16437 VDD.n4004 VDD.t2400 27.5805
R16438 VDD.n4004 VDD.t2394 27.5805
R16439 VDD.n4025 VDD.t1341 27.5805
R16440 VDD.n4025 VDD.t1343 27.5805
R16441 VDD.n4029 VDD.t2977 27.5805
R16442 VDD.n4457 VDD.t2241 27.5805
R16443 VDD.n4455 VDD.t735 27.5805
R16444 VDD.n4455 VDD.t737 27.5805
R16445 VDD.n4489 VDD.t2192 27.5805
R16446 VDD.n4436 VDD.t1216 27.5805
R16447 VDD.n4436 VDD.t1218 27.5805
R16448 VDD.n4058 VDD.t2518 27.5805
R16449 VDD.n4059 VDD.t468 27.5805
R16450 VDD.n4059 VDD.t464 27.5805
R16451 VDD.n4298 VDD.t2764 27.5805
R16452 VDD.n4298 VDD.t2670 27.5805
R16453 VDD.n4305 VDD.t1996 27.5805
R16454 VDD.n4098 VDD.t2125 27.5805
R16455 VDD.n4098 VDD.t2129 27.5805
R16456 VDD.n4099 VDD.t1852 27.5805
R16457 VDD.n4103 VDD.t2172 27.5805
R16458 VDD.n4103 VDD.t2170 27.5805
R16459 VDD.n4107 VDD.t1597 27.5805
R16460 VDD.n4120 VDD.t2067 27.5805
R16461 VDD.n4120 VDD.t2664 27.5805
R16462 VDD.n3925 VDD.t2641 27.5805
R16463 VDD.n3926 VDD.t416 27.5805
R16464 VDD.n3926 VDD.t418 27.5805
R16465 VDD.n3585 VDD.t1864 27.5805
R16466 VDD.n3245 VDD.t1998 27.5805
R16467 VDD.n3257 VDD.t3087 27.5805
R16468 VDD.n3232 VDD.t3502 27.5805
R16469 VDD.n3232 VDD.t2367 27.5805
R16470 VDD.n3238 VDD.t1367 27.5805
R16471 VDD.n3238 VDD.t1369 27.5805
R16472 VDD.n3286 VDD.t1086 27.5805
R16473 VDD.n3286 VDD.t1084 27.5805
R16474 VDD.n3268 VDD.t3213 27.5805
R16475 VDD.n3268 VDD.t3217 27.5805
R16476 VDD.n3269 VDD.t1088 27.5805
R16477 VDD.n3269 VDD.t3169 27.5805
R16478 VDD.n3272 VDD.t1068 27.5805
R16479 VDD.n3272 VDD.t1076 27.5805
R16480 VDD.n3273 VDD.t1074 27.5805
R16481 VDD.n3273 VDD.t1090 27.5805
R16482 VDD.n3277 VDD.t1070 27.5805
R16483 VDD.n3277 VDD.t1072 27.5805
R16484 VDD.n3280 VDD.t1080 27.5805
R16485 VDD.n3281 VDD.t1062 27.5805
R16486 VDD.n3281 VDD.t1078 27.5805
R16487 VDD.n3287 VDD.t1082 27.5805
R16488 VDD.n3287 VDD.t1064 27.5805
R16489 VDD.n3419 VDD.t2272 27.5805
R16490 VDD.n3189 VDD.t3283 27.5805
R16491 VDD.n3782 VDD.t1570 27.5805
R16492 VDD.n3782 VDD.t2293 27.5805
R16493 VDD.n3781 VDD.t2224 27.5805
R16494 VDD.n3781 VDD.t2222 27.5805
R16495 VDD.n3004 VDD.t438 27.5805
R16496 VDD.n2388 VDD.t2744 27.5805
R16497 VDD.n2401 VDD.t3209 27.5805
R16498 VDD.n2401 VDD.t3219 27.5805
R16499 VDD.n2879 VDD.t496 27.5805
R16500 VDD.n2879 VDD.t502 27.5805
R16501 VDD.n2826 VDD.t500 27.5805
R16502 VDD.n2826 VDD.t488 27.5805
R16503 VDD.n2825 VDD.t498 27.5805
R16504 VDD.n2825 VDD.t482 27.5805
R16505 VDD.n2417 VDD.t478 27.5805
R16506 VDD.n2404 VDD.t1009 27.5805
R16507 VDD.n2404 VDD.t3221 27.5805
R16508 VDD.n2407 VDD.t1013 27.5805
R16509 VDD.n2407 VDD.t1019 27.5805
R16510 VDD.n2408 VDD.t1033 27.5805
R16511 VDD.n2408 VDD.t1015 27.5805
R16512 VDD.n2840 VDD.t1011 27.5805
R16513 VDD.n2840 VDD.t1005 27.5805
R16514 VDD.n2842 VDD.t1023 27.5805
R16515 VDD.n2842 VDD.t1029 27.5805
R16516 VDD.n2843 VDD.t1027 27.5805
R16517 VDD.n2843 VDD.t1031 27.5805
R16518 VDD.n2412 VDD.t1017 27.5805
R16519 VDD.n2411 VDD.t1021 27.5805
R16520 VDD.n2411 VDD.t1035 27.5805
R16521 VDD.n3015 VDD.t24 27.5805
R16522 VDD.n3015 VDD.t8 27.5805
R16523 VDD.n2374 VDD.t1968 27.5805
R16524 VDD.n2372 VDD.t671 27.5805
R16525 VDD.n2372 VDD.t673 27.5805
R16526 VDD.n2366 VDD.t3227 27.5805
R16527 VDD.n2366 VDD.t3173 27.5805
R16528 VDD.n2365 VDD.t3215 27.5805
R16529 VDD.n2365 VDD.t36 27.5805
R16530 VDD.n2998 VDD.t12 27.5805
R16531 VDD.n2998 VDD.t38 27.5805
R16532 VDD.n2361 VDD.t34 27.5805
R16533 VDD.n2361 VDD.t22 27.5805
R16534 VDD.n3005 VDD.t14 27.5805
R16535 VDD.n3005 VDD.t32 27.5805
R16536 VDD.n3008 VDD.t10 27.5805
R16537 VDD.n3011 VDD.t28 27.5805
R16538 VDD.n3011 VDD.t30 27.5805
R16539 VDD.n3014 VDD.t18 27.5805
R16540 VDD.n3014 VDD.t26 27.5805
R16541 VDD.n2415 VDD.t506 27.5805
R16542 VDD.n2415 VDD.t494 27.5805
R16543 VDD.n2420 VDD.t504 27.5805
R16544 VDD.n2420 VDD.t490 27.5805
R16545 VDD.n2814 VDD.t484 27.5805
R16546 VDD.n2814 VDD.t508 27.5805
R16547 VDD.n2425 VDD.t3697 27.5805
R16548 VDD.n2425 VDD.t480 27.5805
R16549 VDD.n2426 VDD.t3701 27.5805
R16550 VDD.n2426 VDD.t3699 27.5805
R16551 VDD.n2454 VDD.t250 27.5805
R16552 VDD.n2454 VDD.t1642 27.5805
R16553 VDD.n2462 VDD.t3117 27.5805
R16554 VDD.n2462 VDD.t651 27.5805
R16555 VDD.n1552 VDD.t3344 27.5805
R16556 VDD.n1552 VDD.t3567 27.5805
R16557 VDD.n1974 VDD.t2146 27.5805
R16558 VDD.n1974 VDD.t741 27.5805
R16559 VDD.n1624 VDD.t608 27.5805
R16560 VDD.n1624 VDD.t628 27.5805
R16561 VDD.n1608 VDD.t3175 27.5805
R16562 VDD.n1608 VDD.t3211 27.5805
R16563 VDD.n1610 VDD.t614 27.5805
R16564 VDD.n1610 VDD.t3207 27.5805
R16565 VDD.n1614 VDD.t624 27.5805
R16566 VDD.n1614 VDD.t612 27.5805
R16567 VDD.n1615 VDD.t626 27.5805
R16568 VDD.n1615 VDD.t598 27.5805
R16569 VDD.n1618 VDD.t604 27.5805
R16570 VDD.n1618 VDD.t616 27.5805
R16571 VDD.n1621 VDD.t602 27.5805
R16572 VDD.n1622 VDD.t606 27.5805
R16573 VDD.n1622 VDD.t610 27.5805
R16574 VDD.n1627 VDD.t620 27.5805
R16575 VDD.n1627 VDD.t600 27.5805
R16576 VDD.n1666 VDD.t636 27.5805
R16577 VDD.n1666 VDD.t2927 27.5805
R16578 VDD.n2082 VDD.t2915 27.5805
R16579 VDD.n2082 VDD.t325 27.5805
R16580 VDD.n1958 VDD.t3268 27.5805
R16581 VDD.n1958 VDD.t757 27.5805
R16582 VDD.n2126 VDD.t827 27.5805
R16583 VDD.n2126 VDD.t3251 27.5805
R16584 VDD.n1513 VDD.t1903 27.5805
R16585 VDD.n1513 VDD.t1914 27.5805
R16586 VDD.n1412 VDD.t1936 27.5805
R16587 VDD.n1012 VDD.t2985 27.5805
R16588 VDD.n1012 VDD.t1900 27.5805
R16589 VDD.n894 VDD.t3028 27.5805
R16590 VDD.n894 VDD.t3515 27.5805
R16591 VDD.n851 VDD.t2570 27.5805
R16592 VDD.n852 VDD.t1237 27.5805
R16593 VDD.n852 VDD.t1235 27.5805
R16594 VDD.n656 VDD.t336 27.5805
R16595 VDD.n656 VDD.t340 27.5805
R16596 VDD.n655 VDD.t2319 27.5805
R16597 VDD.n655 VDD.t2318 27.5805
R16598 VDD.n641 VDD.t1574 27.5805
R16599 VDD.n641 VDD.t1578 27.5805
R16600 VDD.n560 VDD.t2523 27.5805
R16601 VDD.n560 VDD.t2522 27.5805
R16602 VDD.n559 VDD.t366 27.5805
R16603 VDD.n559 VDD.t364 27.5805
R16604 VDD.n570 VDD.t1551 27.5805
R16605 VDD.n570 VDD.t1553 27.5805
R16606 VDD.n569 VDD.t782 27.5805
R16607 VDD.n569 VDD.t784 27.5805
R16608 VDD.n480 VDD.t2548 27.5805
R16609 VDD.n480 VDD.t2549 27.5805
R16610 VDD.n479 VDD.t1384 27.5805
R16611 VDD.n479 VDD.t1378 27.5805
R16612 VDD.n490 VDD.t1706 27.5805
R16613 VDD.n490 VDD.t1710 27.5805
R16614 VDD.n489 VDD.t2360 27.5805
R16615 VDD.n489 VDD.t2361 27.5805
R16616 VDD.n2996 VDD.n2995 27.5797
R16617 VDD.n2811 VDD.n2810 27.5797
R16618 VDD.n4356 VDD.n4355 27.4829
R16619 VDD.n3727 VDD.n3726 27.4829
R16620 VDD.n3655 VDD.n3654 27.4829
R16621 VDD.n3434 VDD.n3433 27.4829
R16622 VDD.n3854 VDD.n3853 27.4829
R16623 VDD.n3838 VDD.n3837 27.4829
R16624 VDD.n3833 VDD.n3827 27.4829
R16625 VDD.n2740 VDD.n2464 27.4829
R16626 VDD.n2736 VDD.n2735 27.4829
R16627 VDD.n1951 VDD.n1950 27.4829
R16628 VDD.n1303 VDD.n1302 27.4829
R16629 VDD.n3540 VDD.n3539 27.4829
R16630 VDD.n3435 VDD.n3434 27.4829
R16631 VDD.n3383 VDD.n3294 27.4829
R16632 VDD.n2548 VDD.n2504 27.4829
R16633 VDD.n2333 VDD.n2303 27.4829
R16634 VDD.n1063 VDD.n1010 27.4829
R16635 VDD.n1235 VDD.n771 27.4829
R16636 VDD.n1456 VDD.n1421 27.4829
R16637 VDD.n1593 VDD.t1361 27.3647
R16638 VDD.n1569 VDD.t3307 27.3647
R16639 VDD.n801 VDD.t3303 27.3647
R16640 VDD.n822 VDD.t3660 27.3647
R16641 VDD.n1325 VDD.t428 27.3647
R16642 VDD.n746 VDD.t1098 27.3647
R16643 VDD.n784 VDD.t969 27.3647
R16644 VDD.n3504 VDD.n3503 27.1064
R16645 VDD.n2544 VDD.n2543 27.1064
R16646 VDD.n2995 VDD.n2367 27.1064
R16647 VDD.n2810 VDD.n2427 27.1064
R16648 VDD.n2797 VDD.n2796 27.1064
R16649 VDD.n1777 VDD.n1776 27.1064
R16650 VDD.n1746 VDD.n1745 27.1064
R16651 VDD.n70 VDD.n69 27.1064
R16652 VDD.n41 VDD.n40 27.1064
R16653 VDD.n1884 VDD.n1883 27.0566
R16654 VDD.n2014 VDD.t2440 26.9729
R16655 VDD.t1880 VDD.t1135 26.8556
R16656 VDD.t3638 VDD.t2451 26.8556
R16657 VDD.t2671 VDD.t3733 26.8556
R16658 VDD.t315 VDD.t2896 26.8556
R16659 VDD.n3065 VDD.t1795 26.8556
R16660 VDD.t3718 VDD.t613 26.8556
R16661 VDD.t1302 VDD.t807 26.8556
R16662 VDD.t1515 VDD.t2435 26.8556
R16663 VDD.t2139 VDD.t1304 26.8556
R16664 VDD.t2138 VDD.t3246 26.8556
R16665 VDD.t2994 VDD.t2990 26.8556
R16666 VDD.n4589 VDD.n4588 26.7299
R16667 VDD.n3609 VDD.n3608 26.7299
R16668 VDD.n3441 VDD.n3440 26.7299
R16669 VDD.n2711 VDD.n2658 26.7299
R16670 VDD.n1733 VDD.n1732 26.7299
R16671 VDD.n4491 VDD.n4437 26.7299
R16672 VDD.n1823 VDD.n1619 26.6976
R16673 VDD.n3264 VDD.t581 26.5955
R16674 VDD.n2877 VDD.t875 26.5955
R16675 VDD.n3027 VDD.t2701 26.5955
R16676 VDD.n2478 VDD.t851 26.5955
R16677 VDD.n1962 VDD.t2278 26.5955
R16678 VDD.n726 VDD.t2503 26.5955
R16679 VDD.n1364 VDD.t787 26.5955
R16680 VDD.n1365 VDD.t592 26.5955
R16681 VDD.n4599 VDD.t1470 26.5955
R16682 VDD.n4599 VDD.t1478 26.5955
R16683 VDD.n4082 VDD.t792 26.5955
R16684 VDD.n4082 VDD.t794 26.5955
R16685 VDD.n4102 VDD.t3179 26.5955
R16686 VDD.n4102 VDD.t3189 26.5955
R16687 VDD.n4106 VDD.t3193 26.5955
R16688 VDD.n4106 VDD.t3185 26.5955
R16689 VDD.n4109 VDD.t2949 26.5955
R16690 VDD.n4109 VDD.t2938 26.5955
R16691 VDD.n3280 VDD.t1066 26.5955
R16692 VDD.n3102 VDD.t2460 26.5955
R16693 VDD.n3102 VDD.t2458 26.5955
R16694 VDD.n2392 VDD.t2148 26.5955
R16695 VDD.n2396 VDD.t1116 26.5955
R16696 VDD.n2417 VDD.t486 26.5955
R16697 VDD.n2412 VDD.t1007 26.5955
R16698 VDD.n2967 VDD.t436 26.5955
R16699 VDD.n2967 VDD.t3457 26.5955
R16700 VDD.n3008 VDD.t16 26.5955
R16701 VDD.n2613 VDD.t2748 26.5955
R16702 VDD.n2472 VDD.t1639 26.5955
R16703 VDD.n2661 VDD.t848 26.5955
R16704 VDD.n2661 VDD.t3549 26.5955
R16705 VDD.n1548 VDD.t2823 26.5955
R16706 VDD.n1970 VDD.t858 26.5955
R16707 VDD.n1970 VDD.t862 26.5955
R16708 VDD.n1605 VDD.t1734 26.5955
R16709 VDD.n1621 VDD.t618 26.5955
R16710 VDD.n1637 VDD.t306 26.5955
R16711 VDD.n1637 VDD.t302 26.5955
R16712 VDD.n1645 VDD.t2434 26.5955
R16713 VDD.n2117 VDD.t1162 26.5955
R16714 VDD.n1591 VDD.t278 26.5955
R16715 VDD.n1564 VDD.t1808 26.5955
R16716 VDD.n1564 VDD.t2722 26.5955
R16717 VDD.n1942 VDD.t1550 26.5955
R16718 VDD.n2129 VDD.t2495 26.5955
R16719 VDD.n1514 VDD.t552 26.5955
R16720 VDD.n1514 VDD.t554 26.5955
R16721 VDD.n807 VDD.t1653 26.5955
R16722 VDD.n810 VDD.t2595 26.5955
R16723 VDD.n810 VDD.t2593 26.5955
R16724 VDD.n1026 VDD.t1631 26.5955
R16725 VDD.n1026 VDD.t1635 26.5955
R16726 VDD.n1017 VDD.t3672 26.5955
R16727 VDD.n1017 VDD.t3658 26.5955
R16728 VDD.n1005 VDD.t2375 26.5955
R16729 VDD.n716 VDD.t3527 26.5955
R16730 VDD.n716 VDD.t3467 26.5955
R16731 VDD.n715 VDD.t3471 26.5955
R16732 VDD.n715 VDD.t3455 26.5955
R16733 VDD.n720 VDD.t3530 26.5955
R16734 VDD.n720 VDD.t3553 26.5955
R16735 VDD.n734 VDD.t1442 26.5955
R16736 VDD.n747 VDD.t1560 26.5955
R16737 VDD.n1274 VDD.t1416 26.5955
R16738 VDD.n765 VDD.t1517 26.5955
R16739 VDD.n1129 VDD.t866 26.5955
R16740 VDD.n1149 VDD.t2582 26.5955
R16741 VDD.n1150 VDD.t917 26.5955
R16742 VDD.n1150 VDD.t923 26.5955
R16743 VDD.n788 VDD.t1464 26.5955
R16744 VDD.n788 VDD.t1458 26.5955
R16745 VDD.n702 VDD.t585 26.5955
R16746 VDD.n707 VDD.t817 26.5955
R16747 VDD.n707 VDD.t815 26.5955
R16748 VDD.n709 VDD.t1452 26.5955
R16749 VDD.n619 VDD.t1045 26.5955
R16750 VDD.n619 VDD.t1051 26.5955
R16751 VDD.n618 VDD.t1372 26.5955
R16752 VDD.n618 VDD.t1373 26.5955
R16753 VDD.n608 VDD.t722 26.5955
R16754 VDD.n608 VDD.t718 26.5955
R16755 VDD.n536 VDD.t2648 26.5955
R16756 VDD.n536 VDD.t2651 26.5955
R16757 VDD.n535 VDD.t402 26.5955
R16758 VDD.n535 VDD.t398 26.5955
R16759 VDD.n528 VDD.t879 26.5955
R16760 VDD.n528 VDD.t881 26.5955
R16761 VDD.n527 VDD.t2159 26.5955
R16762 VDD.n527 VDD.t2162 26.5955
R16763 VDD.n456 VDD.t1153 26.5955
R16764 VDD.n456 VDD.t1154 26.5955
R16765 VDD.n455 VDD.t703 26.5955
R16766 VDD.n455 VDD.t707 26.5955
R16767 VDD.n448 VDD.t284 26.5955
R16768 VDD.n448 VDD.t280 26.5955
R16769 VDD.n447 VDD.t1613 26.5955
R16770 VDD.n447 VDD.t1614 26.5955
R16771 VDD.n346 VDD.t356 26.5955
R16772 VDD.n346 VDD.t352 26.5955
R16773 VDD.n345 VDD.t2687 26.5955
R16774 VDD.n345 VDD.t2637 26.5955
R16775 VDD.n347 VDD.t2685 26.5955
R16776 VDD.n347 VDD.t2681 26.5955
R16777 VDD.n351 VDD.t1210 26.5955
R16778 VDD.n351 VDD.t1204 26.5955
R16779 VDD.n134 VDD.t663 26.5955
R16780 VDD.n65 VDD.t1665 26.5955
R16781 VDD.n65 VDD.t1663 26.5955
R16782 VDD.n71 VDD.t3069 26.5955
R16783 VDD.n71 VDD.t3065 26.5955
R16784 VDD.n39 VDD.t2406 26.5955
R16785 VDD.n39 VDD.t2404 26.5955
R16786 VDD.n36 VDD.t3067 26.5955
R16787 VDD.n36 VDD.t3056 26.5955
R16788 VDD.n239 VDD.n238 26.4291
R16789 VDD.n240 VDD.n239 26.4291
R16790 VDD.n236 VDD.n235 26.4291
R16791 VDD.n235 VDD.n234 26.4291
R16792 VDD.n233 VDD.n223 26.4291
R16793 VDD.n234 VDD.n233 26.4291
R16794 VDD.n242 VDD.n241 26.4291
R16795 VDD.n241 VDD.n240 26.4291
R16796 VDD.n121 VDD.n101 26.4291
R16797 VDD.n122 VDD.n121 26.4291
R16798 VDD.n109 VDD.n102 26.4291
R16799 VDD.n122 VDD.n109 26.4291
R16800 VDD.n114 VDD.n110 26.4291
R16801 VDD.n122 VDD.n110 26.4291
R16802 VDD.n3108 VDD.t683 26.3637
R16803 VDD.n3819 VDD.t372 26.3637
R16804 VDD.n2379 VDD.t442 26.3637
R16805 VDD.n2470 VDD.t1371 26.3637
R16806 VDD.n1967 VDD.t1102 26.3637
R16807 VDD.n1581 VDD.t3279 26.3637
R16808 VDD.n4592 VDD.n4589 26.3534
R16809 VDD.n4243 VDD.n4242 26.3534
R16810 VDD.n2623 VDD.n2622 26.3534
R16811 VDD.n3629 VDD.n3628 25.977
R16812 VDD.n3519 VDD.n3518 25.977
R16813 VDD.n3425 VDD.n3411 25.977
R16814 VDD.n3859 VDD.n3858 25.977
R16815 VDD.n2975 VDD.n2377 25.977
R16816 VDD.n3073 VDD.n2282 25.977
R16817 VDD.n2733 VDD.n2468 25.977
R16818 VDD.n2627 VDD.n2485 25.977
R16819 VDD.n2056 VDD.n2055 25.977
R16820 VDD.n2054 VDD.n2053 25.977
R16821 VDD.n1861 VDD.n1860 25.977
R16822 VDD.n2111 VDD.n1519 25.977
R16823 VDD.n2165 VDD.n2123 25.977
R16824 VDD.n2153 VDD.n2152 25.977
R16825 VDD.n1385 VDD.n1384 25.977
R16826 VDD.n162 VDD.n161 25.977
R16827 VDD.n3984 VDD.t3034 25.6105
R16828 VDD.n4114 VDD.t3668 25.6105
R16829 VDD.n4117 VDD.t1595 25.6105
R16830 VDD.n3775 VDD.t761 25.6105
R16831 VDD.n2386 VDD.t2906 25.6105
R16832 VDD.n2834 VDD.t1 25.6105
R16833 VDD.n2621 VDD.t2746 25.6105
R16834 VDD.n2483 VDD.t2370 25.6105
R16835 VDD.n2655 VDD.t751 25.6105
R16836 VDD.n1540 VDD.t1150 25.6105
R16837 VDD.n1650 VDD.t2759 25.6105
R16838 VDD.n2103 VDD.t1270 25.6105
R16839 VDD.n1907 VDD.t524 25.6105
R16840 VDD.n2122 VDD.t2166 25.6105
R16841 VDD.n2132 VDD.t1039 25.6105
R16842 VDD.n4528 VDD.n4527 25.6005
R16843 VDD.n4294 VDD.n4288 25.6005
R16844 VDD.n4256 VDD.n4104 25.6005
R16845 VDD.n4250 VDD.n4249 25.6005
R16846 VDD.n4188 VDD.n4187 25.6005
R16847 VDD.n4171 VDD.n4170 25.6005
R16848 VDD.n3707 VDD.n3199 25.6005
R16849 VDD.n3347 VDD.n3317 25.6005
R16850 VDD.n3337 VDD.n3336 25.6005
R16851 VDD.n3149 VDD.n3129 25.6005
R16852 VDD.n3143 VDD.n3133 25.6005
R16853 VDD.n3032 VDD.n3029 25.6005
R16854 VDD.n2636 VDD.n2635 25.6005
R16855 VDD.n2587 VDD.n2586 25.6005
R16856 VDD.n2328 VDD.n2327 25.6005
R16857 VDD.n2322 VDD.n2321 25.6005
R16858 VDD.n1764 VDD.n1763 25.6005
R16859 VDD.n1723 VDD.n1722 25.6005
R16860 VDD.n1717 VDD.n1716 25.6005
R16861 VDD.n1703 VDD.n1702 25.6005
R16862 VDD.n2021 VDD.n2020 25.6005
R16863 VDD.n2268 VDD.n1509 25.6005
R16864 VDD.n2212 VDD.n2211 25.6005
R16865 VDD.n2206 VDD.n2205 25.6005
R16866 VDD.n1088 VDD.n1087 25.6005
R16867 VDD.n966 VDD.n965 25.6005
R16868 VDD.n905 VDD.n904 25.6005
R16869 VDD.n911 VDD.n910 25.6005
R16870 VDD.n1217 VDD.n1216 25.6005
R16871 VDD.n1389 VDD.n1366 25.6005
R16872 VDD.n1448 VDD.n1447 25.6005
R16873 VDD.n1442 VDD.n1441 25.6005
R16874 VDD.n3982 VDD.n3908 25.224
R16875 VDD.n4618 VDD.n4611 25.224
R16876 VDD.n4515 VDD.n4512 25.224
R16877 VDD.n4510 VDD.n4035 25.224
R16878 VDD.n4511 VDD.n4510 25.224
R16879 VDD.n4458 VDD.n4038 25.224
R16880 VDD.n4258 VDD.n4100 25.224
R16881 VDD.n3948 VDD.n3947 25.224
R16882 VDD.n3608 VDD.n3607 25.224
R16883 VDD.n3607 VDD.n3581 25.224
R16884 VDD.n3440 VDD.n3404 25.224
R16885 VDD.n3792 VDD.n3184 25.224
R16886 VDD.n2959 VDD.n2958 25.224
R16887 VDD.n2959 VDD.n2380 25.224
R16888 VDD.n2977 VDD.n2375 25.224
R16889 VDD.n2605 VDD.n2489 25.224
R16890 VDD.n2698 VDD.n2697 25.224
R16891 VDD.n2064 VDD.n2063 25.224
R16892 VDD.n2109 VDD.n1521 25.224
R16893 VDD.n632 VDD.n612 25.224
R16894 VDD.n549 VDD.n529 25.224
R16895 VDD.n469 VDD.n449 25.224
R16896 VDD.n76 VDD.n75 25.224
R16897 VDD.n37 VDD.n31 25.224
R16898 VDD.n4660 VDD.n3901 25.1912
R16899 VDD.n4479 VDD.n4478 25.1912
R16900 VDD.n4425 VDD.n4423 25.1912
R16901 VDD.n4380 VDD.n4379 25.1912
R16902 VDD.n4317 VDD.n4316 25.1912
R16903 VDD.n4210 VDD.n4209 25.1912
R16904 VDD.n3672 VDD.n3668 25.1912
R16905 VDD.n3833 VDD.n3832 25.1912
R16906 VDD.n3885 VDD.n3098 25.1912
R16907 VDD.n3152 VDD.n3151 25.1912
R16908 VDD.n2549 VDD.n2548 25.1912
R16909 VDD.n2561 VDD.n2497 25.1912
R16910 VDD.n2338 VDD.n2337 25.1912
R16911 VDD.n1276 VDD.n1273 25.1912
R16912 VDD.t1849 VDD.t2401 25.1772
R16913 VDD.t871 VDD.t1594 25.1772
R16914 VDD.t2251 VDD.t2128 25.1772
R16915 VDD.t2244 VDD.t180 25.1772
R16916 VDD.t1789 VDD.t2294 25.1772
R16917 VDD.t2210 VDD.t2309 25.1772
R16918 VDD.t2610 VDD.t2060 25.1772
R16919 VDD.t3408 VDD.t3666 25.1772
R16920 VDD.t2585 VDD.t2002 25.1772
R16921 VDD.t389 VDD.t2758 25.1772
R16922 VDD.t255 VDD.t1437 25.1772
R16923 VDD.t2652 VDD.t1831 25.1772
R16924 VDD.t519 VDD.t3326 25.1772
R16925 VDD.n2885 VDD.n2827 24.8691
R16926 VDD.n2853 VDD.n2852 24.8691
R16927 VDD.n3485 VDD.n3484 24.8691
R16928 VDD.n1819 VDD.n1818 24.8691
R16929 VDD.n4521 VDD.n4520 24.8476
R16930 VDD.n4371 VDD.n4077 24.8476
R16931 VDD.n4335 VDD.n4334 24.8476
R16932 VDD.n4191 VDD.n4190 24.8476
R16933 VDD.n4183 VDD.n4182 24.8476
R16934 VDD.n4183 VDD.n4145 24.8476
R16935 VDD.n4175 VDD.n4161 24.8476
R16936 VDD.n3958 VDD.n3919 24.8476
R16937 VDD.n3954 VDD.n3953 24.8476
R16938 VDD.n3952 VDD.n3923 24.8476
R16939 VDD.n3732 VDD.n3731 24.8476
R16940 VDD.n3349 VDD.n3348 24.8476
R16941 VDD.n3764 VDD.n3763 24.8476
R16942 VDD.n3341 VDD.n3327 24.8476
R16943 VDD.n3151 VDD.n3150 24.8476
R16944 VDD.n3145 VDD.n3144 24.8476
R16945 VDD.n2521 VDD.n2517 24.8476
R16946 VDD.n2529 VDD.n2514 24.8476
R16947 VDD.n2563 VDD.n2561 24.8476
R16948 VDD.n2644 VDD.n2476 24.8476
R16949 VDD.n2591 VDD.n2577 24.8476
R16950 VDD.n2326 VDD.n2312 24.8476
R16951 VDD.n1721 VDD.n1685 24.8476
R16952 VDD.n1707 VDD.n1693 24.8476
R16953 VDD.n2025 VDD.n1955 24.8476
R16954 VDD.n2243 VDD.n2242 24.8476
R16955 VDD.n2210 VDD.n2196 24.8476
R16956 VDD.n1124 VDD.n1123 24.8476
R16957 VDD.n961 VDD.n840 24.8476
R16958 VDD.n959 VDD.n958 24.8476
R16959 VDD.n932 VDD.n930 24.8476
R16960 VDD.n944 VDD.n880 24.8476
R16961 VDD.n1351 VDD.n717 24.8476
R16962 VDD.n1339 VDD.n724 24.8476
R16963 VDD.n1283 VDD.n748 24.8476
R16964 VDD.n1252 VDD.n1251 24.8476
R16965 VDD.n1172 VDD.n1171 24.8476
R16966 VDD.n1398 VDD.n1358 24.8476
R16967 VDD.n1383 VDD.n1369 24.8476
R16968 VDD.n1377 VDD.n1372 24.8476
R16969 VDD.n1474 VDD.n1473 24.8476
R16970 VDD.n1462 VDD.n1461 24.8476
R16971 VDD.n1456 VDD.n1455 24.8476
R16972 VDD.n1452 VDD.n1428 24.8476
R16973 VDD.n1446 VDD.n1432 24.8476
R16974 VDD.n409 VDD.n340 24.8005
R16975 VDD.n3475 VDD.n3288 24.6862
R16976 VDD.n2854 VDD.n2853 24.5034
R16977 VDD.n4203 VDD.n4202 24.4711
R16978 VDD.n4514 VDD.n4032 24.4711
R16979 VDD.n4398 VDD.n4397 24.4711
R16980 VDD.n3715 VDD.n3714 24.4711
R16981 VDD.n3643 VDD.n3642 24.4711
R16982 VDD.n3616 VDD.n3575 24.4711
R16983 VDD.n3628 VDD.n3627 24.4711
R16984 VDD.n3509 VDD.n3265 24.4711
R16985 VDD.n3421 VDD.n3411 24.4711
R16986 VDD.n3858 VDD.n3812 24.4711
R16987 VDD.n2921 VDD.n2920 24.4711
R16988 VDD.n2957 VDD.n2382 24.4711
R16989 VDD.n2990 VDD.n2989 24.4711
R16990 VDD.n2802 VDD.n2801 24.4711
R16991 VDD.n2793 VDD.n2792 24.4711
R16992 VDD.n2779 VDD.n2778 24.4711
R16993 VDD.n2734 VDD.n2733 24.4711
R16994 VDD.n2053 VDD.n1545 24.4711
R16995 VDD.n1865 VDD.n1594 24.4711
R16996 VDD.n1772 VDD.n1771 24.4711
R16997 VDD.n2019 VDD.n1957 24.4711
R16998 VDD.n917 VDD.n892 24.4711
R16999 VDD.n1327 VDD.n1324 24.4711
R17000 VDD.n162 VDD.n123 24.4711
R17001 VDD.n4301 VDD.n4300 24.0946
R17002 VDD.n4249 VDD.n4110 24.0946
R17003 VDD.n4236 VDD.n4118 24.0946
R17004 VDD.n4176 VDD.n4175 24.0946
R17005 VDD.n3641 VDD.n3640 24.0946
R17006 VDD.n3796 VDD.n3184 24.0946
R17007 VDD.n3145 VDD.n3129 24.0946
R17008 VDD.n2945 VDD.n2944 24.0946
R17009 VDD.n2327 VDD.n2326 24.0946
R17010 VDD.n1765 VDD.n1764 24.0946
R17011 VDD.n1729 VDD.n1728 24.0946
R17012 VDD.n1722 VDD.n1721 24.0946
R17013 VDD.n1883 VDD.n1588 24.0946
R17014 VDD.n1929 VDD.n1928 24.0946
R17015 VDD.n2268 VDD.n2267 24.0946
R17016 VDD.n2211 VDD.n2210 24.0946
R17017 VDD.n1121 VDD.n1120 24.0946
R17018 VDD.n967 VDD.n966 24.0946
R17019 VDD.n906 VDD.n905 24.0946
R17020 VDD.n937 VDD.n936 24.0946
R17021 VDD.n1216 VDD.n1215 24.0946
R17022 VDD.n1396 VDD.n1395 24.0946
R17023 VDD.n1378 VDD.n1377 24.0946
R17024 VDD.n1473 VDD.n1410 24.0946
R17025 VDD.n1453 VDD.n1452 24.0946
R17026 VDD.n1447 VDD.n1446 24.0946
R17027 VDD.n3049 VDD.n3048 23.7719
R17028 VDD.n1834 VDD.n1611 23.7719
R17029 VDD.n3523 VDD.n3258 23.7181
R17030 VDD.n3470 VDD.n3290 23.7181
R17031 VDD.n3173 VDD.n3111 23.7181
R17032 VDD.n2966 VDD.n2965 23.7181
R17033 VDD.n2677 VDD.n2471 23.7181
R17034 VDD.n1996 VDD.n1995 23.7181
R17035 VDD.n4649 VDD.n3983 23.7181
R17036 VDD.n4552 VDD.n4548 23.7181
R17037 VDD.n4547 VDD.n4009 23.7181
R17038 VDD.n4504 VDD.n4038 23.7181
R17039 VDD.n4501 VDD.n4039 23.7181
R17040 VDD.n4413 VDD.n4412 23.7181
R17041 VDD.n4347 VDD.n4092 23.7181
R17042 VDD.n4343 VDD.n4094 23.7181
R17043 VDD.n4229 VDD.n4123 23.7181
R17044 VDD.n3753 VDD.n3200 23.7181
R17045 VDD.n3651 VDD.n3650 23.7181
R17046 VDD.n3636 VDD.n3227 23.7181
R17047 VDD.n3633 VDD.n3228 23.7181
R17048 VDD.n3629 VDD.n3228 23.7181
R17049 VDD.n3466 VDD.n3291 23.7181
R17050 VDD.n3466 VDD.n3292 23.7181
R17051 VDD.n3349 VDD.n3313 23.7181
R17052 VDD.n3864 VDD.n3179 23.7181
R17053 VDD.n3864 VDD.n3863 23.7181
R17054 VDD.n3860 VDD.n3859 23.7181
R17055 VDD.n3342 VDD.n3341 23.7181
R17056 VDD.n2945 VDD.n2384 23.7181
R17057 VDD.n2866 VDD.n2865 23.7181
R17058 VDD.n2872 VDD.n2871 23.7181
R17059 VDD.n2348 VDD.n2347 23.7181
R17060 VDD.n2949 VDD.n2384 23.7181
R17061 VDD.n2976 VDD.n2975 23.7181
R17062 VDD.n3033 VDD.n3032 23.7181
R17063 VDD.n3073 VDD.n3072 23.7181
R17064 VDD.n2776 VDD.n2445 23.7181
R17065 VDD.n2729 VDD.n2468 23.7181
R17066 VDD.n2598 VDD.n2596 23.7181
R17067 VDD.n2623 VDD.n2485 23.7181
R17068 VDD.n2714 VDD.n2653 23.7181
R17069 VDD.n2712 VDD.n2711 23.7181
R17070 VDD.n2707 VDD.n2658 23.7181
R17071 VDD.n2592 VDD.n2591 23.7181
R17072 VDD.n2068 VDD.n1538 23.7181
R17073 VDD.n2030 VDD.n1558 23.7181
R17074 VDD.n2012 VDD.n1960 23.7181
R17075 VDD.n1860 VDD.n1859 23.7181
R17076 VDD.n1806 VDD.n1630 23.7181
R17077 VDD.n1758 VDD.n1757 23.7181
R17078 VDD.n1757 VDD.n1657 23.7181
R17079 VDD.n2111 VDD.n2110 23.7181
R17080 VDD.n2170 VDD.n1517 23.7181
R17081 VDD.n1902 VDD.n1576 23.7181
R17082 VDD.n2170 VDD.n2169 23.7181
R17083 VDD.n1198 VDD.n790 23.7181
R17084 VDD.n1081 VDD.n1080 23.7181
R17085 VDD.n1077 VDD.n818 23.7181
R17086 VDD.n1077 VDD.n819 23.7181
R17087 VDD.n957 VDD.n844 23.7181
R17088 VDD.n950 VDD.n849 23.7181
R17089 VDD.n1331 VDD.n727 23.7181
R17090 VDD.n1324 VDD.n1323 23.7181
R17091 VDD.n1252 VDD.n760 23.7181
R17092 VDD.n1198 VDD.n791 23.7181
R17093 VDD.n1403 VDD.n1402 23.7181
R17094 VDD.n1384 VDD.n1383 23.7181
R17095 VDD.n161 VDD.n160 23.7181
R17096 VDD.t890 VDD.t3202 23.4987
R17097 VDD.t3418 VDD.t2616 23.4987
R17098 VDD.t1193 VDD.t3155 23.4987
R17099 VDD.t3259 VDD.t3763 23.4987
R17100 VDD.t3142 VDD.t1543 23.4987
R17101 VDD.t2656 VDD.t1535 23.4987
R17102 VDD.t3548 VDD.t3105 23.4987
R17103 VDD.t804 VDD.t1448 23.4987
R17104 VDD.t2279 VDD.t499 23.4987
R17105 VDD.t3214 VDD.t2775 23.4987
R17106 VDD.t29 VDD.t379 23.4987
R17107 VDD.t621 VDD.t991 23.4987
R17108 VDD.t253 VDD.t1362 23.4987
R17109 VDD.t2328 VDD.t3389 23.4987
R17110 VDD.n146 VDD.t1760 23.3739
R17111 VDD.n150 VDD.t1756 23.3739
R17112 VDD.n88 VDD.t3434 23.3739
R17113 VDD.n130 VDD.t3432 23.3739
R17114 VDD.n4591 VDD.n3985 23.3417
R17115 VDD.n3526 VDD.n3525 23.3417
R17116 VDD.n3461 VDD.n3460 23.3417
R17117 VDD.n2534 VDD.n2511 23.3417
R17118 VDD.n2236 VDD.n2180 23.3417
R17119 VDD.n1122 VDD.n1121 23.3417
R17120 VDD.n1222 VDD.n777 23.3417
R17121 VDD.n1179 VDD.n1178 23.3417
R17122 VDD.n1468 VDD.n1467 23.3417
R17123 VDD.n230 VDD.n229 23.1255
R17124 VDD.n231 VDD.n224 23.1255
R17125 VDD.n232 VDD.n231 23.1255
R17126 VDD.n227 VDD.n225 23.1255
R17127 VDD.n3937 VDD.n3930 22.9652
R17128 VDD.n2781 VDD.n2439 22.9652
R17129 VDD.n950 VDD.n848 22.9652
R17130 VDD.n863 VDD.n856 22.9652
R17131 VDD.n4672 VDD.n4671 22.9652
R17132 VDD.n4584 VDD.n4583 22.9652
R17133 VDD.n4543 VDD.n4542 22.9652
R17134 VDD.n4464 VDD.n4463 22.9652
R17135 VDD.n4432 VDD.n4040 22.9652
R17136 VDD.n4300 VDD.n4299 22.9652
R17137 VDD.n4232 VDD.n4231 22.9652
R17138 VDD.n3727 VDD.n3692 22.9652
R17139 VDD.n3565 VDD.n3564 22.9652
R17140 VDD.n3559 VDD.n3558 22.9652
R17141 VDD.n3547 VDD.n3546 22.9652
R17142 VDD.n3541 VDD.n3540 22.9652
R17143 VDD.n3783 VDD.n3780 22.9652
R17144 VDD.n3837 VDD.n3827 22.9652
R17145 VDD.n2736 VDD.n2464 22.9652
R17146 VDD.n2703 VDD.n2663 22.9652
R17147 VDD.n1766 VDD.n1765 22.9652
R17148 VDD.n1741 VDD.n1740 22.9652
R17149 VDD.n2164 VDD.n2163 22.9652
R17150 VDD.n2221 VDD.n2186 22.9652
R17151 VDD.n1125 VDD.n1124 22.9652
R17152 VDD.n1053 VDD.n1013 22.9652
R17153 VDD.n1066 VDD.n1064 22.9652
R17154 VDD.n651 VDD.n648 22.9652
R17155 VDD.t62 VDD.n328 22.9315
R17156 VDD.n328 VDD.t63 22.9315
R17157 VDD.n324 VDD.t70 22.9315
R17158 VDD.n324 VDD.t66 22.9315
R17159 VDD.n3489 VDD.n3278 22.6748
R17160 VDD.n3776 VDD.n3774 22.5887
R17161 VDD.n3853 VDD.n3852 22.5887
R17162 VDD.n2936 VDD.n2935 22.5887
R17163 VDD.n2931 VDD.n2393 22.5887
R17164 VDD.n2920 VDD.n2919 22.5887
R17165 VDD.n3029 VDD.n3028 22.5887
R17166 VDD.n2681 VDD.n2680 22.5887
R17167 VDD.n2047 VDD.n2046 22.5887
R17168 VDD.n1839 VDD.n1838 22.5887
R17169 VDD.n2102 VDD.n1524 22.5887
R17170 VDD.n2116 VDD.n2115 22.5887
R17171 VDD.n2118 VDD.n1517 22.5887
R17172 VDD.n2157 VDD.n2156 22.5887
R17173 VDD.n990 VDD.n826 22.5887
R17174 VDD.n1385 VDD.n1366 22.5887
R17175 VDD.n4355 VDD.n4354 22.2123
R17176 VDD.n4349 VDD.n4348 22.2123
R17177 VDD.n4348 VDD.n4347 22.2123
R17178 VDD.n4307 VDD.n4306 22.2123
R17179 VDD.n4238 VDD.n4237 22.2123
R17180 VDD.n4231 VDD.n4230 22.2123
R17181 VDD.n4230 VDD.n4229 22.2123
R17182 VDD.n3663 VDD.n3662 22.2123
R17183 VDD.n3662 VDD.n3661 22.2123
R17184 VDD.n3602 VDD.n3601 22.2123
R17185 VDD.n3609 VDD.n3579 22.2123
R17186 VDD.n3613 VDD.n3579 22.2123
R17187 VDD.n3420 VDD.n3418 22.2123
R17188 VDD.n3421 VDD.n3420 22.2123
R17189 VDD.n2943 VDD.n2942 22.2123
R17190 VDD.n2867 VDD.n2832 22.2123
R17191 VDD.n2969 VDD.n2377 22.2123
R17192 VDD.n2747 VDD.n2746 22.2123
R17193 VDD.n2746 VDD.n2745 22.2123
R17194 VDD.n2069 VDD.n2068 22.2123
R17195 VDD.n2057 VDD.n1541 22.2123
R17196 VDD.n1975 VDD.n1558 22.2123
R17197 VDD.n2091 VDD.n2090 22.2123
R17198 VDD.n2092 VDD.n2091 22.2123
R17199 VDD.n2097 VDD.n2096 22.2123
R17200 VDD.n2015 VDD.n2013 22.2123
R17201 VDD.n2015 VDD.n1957 22.2123
R17202 VDD.n2169 VDD.n2123 22.2123
R17203 VDD.n1001 VDD.n819 22.2123
R17204 VDD.n1001 VDD.n1000 22.2123
R17205 VDD.n919 VDD.n918 22.2123
R17206 VDD.n1236 VDD.n1235 22.2123
R17207 VDD.n1185 VDD.n1184 22.2123
R17208 VDD.n1184 VDD.n1183 22.2123
R17209 VDD.n4642 VDD.n4641 21.8358
R17210 VDD.n3873 VDD.n3872 21.8358
R17211 VDD.n2935 VDD.n2393 21.8358
R17212 VDD.n1988 VDD.n1987 21.8358
R17213 VDD.n1794 VDD.n1793 21.8358
R17214 VDD.n2098 VDD.n1524 21.8358
R17215 VDD.n2118 VDD.n2116 21.8358
R17216 VDD.n1930 VDD.n1929 21.8358
R17217 VDD.n2255 VDD.n2254 21.8358
R17218 VDD.n1094 VDD.n1093 21.8358
R17219 VDD.n1027 VDD.n1023 21.8358
R17220 VDD.n789 VDD.n785 21.8358
R17221 VDD.n427 VDD.n426 21.8358
R17222 VDD.t769 VDD.t872 21.8203
R17223 VDD.n3467 VDD.t2301 21.8203
R17224 VDD.t3691 VDD.t2826 21.8203
R17225 VDD.t1589 VDD.t725 21.8203
R17226 VDD.t2197 VDD.t3186 21.8203
R17227 VDD.t2843 VDD.t1957 21.8203
R17228 VDD.t3091 VDD.t645 21.8203
R17229 VDD.t1598 VDD.t635 21.8203
R17230 VDD.t3244 VDD.t391 21.8203
R17231 VDD.t297 VDD.t1328 21.8203
R17232 VDD.t989 VDD.n1631 21.8203
R17233 VDD.t3250 VDD.t3523 21.8203
R17234 VDD.n2172 VDD.t543 21.8203
R17235 VDD.t3269 VDD.t2583 21.8203
R17236 VDD.t1155 VDD.t2235 21.8203
R17237 VDD.t3375 VDD.t3336 21.8203
R17238 VDD.t2963 VDD.t1679 21.8203
R17239 VDD.n4671 VDD.n3901 21.4593
R17240 VDD.n4584 VDD.n3987 21.4593
R17241 VDD.n4543 VDD.n4009 21.4593
R17242 VDD.n4524 VDD.n4030 21.4593
R17243 VDD.n4520 VDD.n4519 21.4593
R17244 VDD.n4463 VDD.n4454 21.4593
R17245 VDD.n4367 VDD.n4077 21.4593
R17246 VDD.n4353 VDD.n4085 21.4593
R17247 VDD.n4237 VDD.n4236 21.4593
R17248 VDD.n3731 VDD.n3692 21.4593
R17249 VDD.n3558 VDD.n3557 21.4593
R17250 VDD.n3545 VDD.n3249 21.4593
R17251 VDD.n3546 VDD.n3545 21.4593
R17252 VDD.n3178 VDD.n3177 21.4593
R17253 VDD.n3784 VDD.n3783 21.4593
R17254 VDD.n2938 VDD.n2937 21.4593
R17255 VDD.n2929 VDD.n2928 21.4593
R17256 VDD.n2927 VDD.n2398 21.4593
R17257 VDD.n2777 VDD.n2776 21.4593
R17258 VDD.n2622 VDD.n2620 21.4593
R17259 VDD.n2648 VDD.n2476 21.4593
R17260 VDD.n2720 VDD.n2474 21.4593
R17261 VDD.n2042 VDD.n2041 21.4593
R17262 VDD.n1981 VDD.n1980 21.4593
R17263 VDD.n1853 VDD.n1852 21.4593
R17264 VDD.n1801 VDD.n1800 21.4593
R17265 VDD.n1778 VDD.n1777 21.4593
R17266 VDD.n1766 VDD.n1648 21.4593
R17267 VDD.n2086 VDD.n2081 21.4593
R17268 VDD.n2098 VDD.n2097 21.4593
R17269 VDD.n1876 VDD.n1590 21.4593
R17270 VDD.n1943 VDD.n1941 21.4593
R17271 VDD.n1944 VDD.n1562 21.4593
R17272 VDD.n2163 VDD.n2162 21.4593
R17273 VDD.n2248 VDD.n2247 21.4593
R17274 VDD.n1125 VDD.n790 21.4593
R17275 VDD.n1102 VDD.n1100 21.4593
R17276 VDD.n1057 VDD.n1013 21.4593
R17277 VDD.n1066 VDD.n1008 21.4593
R17278 VDD.n1071 VDD.n1070 21.4593
R17279 VDD.n1311 VDD.n731 21.4593
R17280 VDD.n1310 VDD.n1309 21.4593
R17281 VDD.n1290 VDD.n744 21.4593
R17282 VDD.n1288 VDD.n1287 21.4593
R17283 VDD.n1281 VDD.n1280 21.4593
R17284 VDD.n1194 VDD.n1193 21.4593
R17285 VDD.n1169 VDD.n1145 21.4593
R17286 VDD.n1164 VDD.n1163 21.4593
R17287 VDD.n1497 VDD.n1496 21.4593
R17288 VDD.n1483 VDD.n1482 21.4593
R17289 VDD.n3359 VDD.n3303 21.1975
R17290 VDD.n3548 VDD.n3243 21.0829
R17291 VDD.n2923 VDD.n2398 21.0829
R17292 VDD.n2786 VDD.n2439 21.0829
R17293 VDD.n2720 VDD.n2719 21.0829
R17294 VDD.n2030 VDD.n1556 21.0829
R17295 VDD.n1778 VDD.n1642 21.0829
R17296 VDD.n1948 VDD.n1562 21.0829
R17297 VDD.n1070 VDD.n1008 21.0829
R17298 VDD.n1315 VDD.n731 21.0829
R17299 VDD.n1294 VDD.n744 21.0829
R17300 VDD.n1282 VDD.n1281 21.0829
R17301 VDD.n1250 VDD.n763 21.0829
R17302 VDD.n1191 VDD.n1190 21.0829
R17303 VDD.n3478 VDD.n3477 20.8462
R17304 VDD.n2616 VDD.n2611 20.7661
R17305 VDD.n3960 VDD.n3958 20.755
R17306 VDD.n4619 VDD.n4618 20.7064
R17307 VDD.n4634 VDD.n4604 20.7064
R17308 VDD.n4559 VDD.n4558 20.7064
R17309 VDD.n4458 VDD.n4454 20.7064
R17310 VDD.n4375 VDD.n4374 20.7064
R17311 VDD.n4262 VDD.n4100 20.7064
R17312 VDD.n4252 VDD.n4104 20.7064
R17313 VDD.n3947 VDD.n3946 20.7064
R17314 VDD.n3780 VDD.n3190 20.7064
R17315 VDD.n2981 VDD.n2375 20.7064
R17316 VDD.n1478 VDD.n1477 20.7064
R17317 VDD.n77 VDD.n76 20.7064
R17318 VDD.n38 VDD.n37 20.7064
R17319 VDD.n202 VDD.n199 20.5561
R17320 VDD.n202 VDD.n193 20.5561
R17321 VDD.n148 VDD.n147 20.5174
R17322 VDD.n149 VDD.n145 20.5174
R17323 VDD.n128 VDD.n127 20.5174
R17324 VDD.n129 VDD.n126 20.5174
R17325 VDD.n2855 VDD.n2854 20.4805
R17326 VDD.n3048 VDD.n3016 20.4805
R17327 VDD.n1812 VDD.n1809 20.4805
R17328 VDD.n4199 VDD.n4135 20.3837
R17329 VDD.n4198 VDD.n4197 20.3299
R17330 VDD.n3738 VDD.n3688 20.3299
R17331 VDD.n3518 VDD.n3517 20.3299
R17332 VDD.n3455 VDD.n3453 20.3299
R17333 VDD.n2873 VDD.n2829 20.3299
R17334 VDD.n2880 VDD.n2878 20.3299
R17335 VDD.n2525 VDD.n2514 20.3299
R17336 VDD.n1802 VDD.n1630 20.3299
R17337 VDD.n1795 VDD.n1635 20.3299
R17338 VDD.n2075 VDD.n2074 20.3299
R17339 VDD.n1106 VDD.n805 20.3299
R17340 VDD.n1042 VDD.n1020 20.3299
R17341 VDD.n1215 VDD.n782 20.3299
R17342 VDD.n1171 VDD.n1170 20.3299
R17343 VDD.t2340 VDD.t2302 20.1418
R17344 VDD.t2483 VDD.t1075 20.1418
R17345 VDD.t531 VDD.t1863 20.1418
R17346 VDD.t2622 VDD.t3562 20.1418
R17347 VDD.t509 VDD.t2423 20.1418
R17348 VDD.t27 VDD.t383 20.1418
R17349 VDD.t3097 VDD.t3524 20.1418
R17350 VDD.t3732 VDD.t2217 20.1418
R17351 VDD.t571 VDD.t1122 20.1418
R17352 VDD.t451 VDD.t2321 20.1418
R17353 VDD.t174 VDD.t1575 20.1418
R17354 VDD.n3483 VDD.n3482 20.1148
R17355 VDD.n2852 VDD.n2844 20.1148
R17356 VDD.n3052 VDD.n3051 20.1148
R17357 VDD.n1817 VDD.n1816 20.1148
R17358 VDD.n4625 VDD.n4606 19.9534
R17359 VDD.n4529 VDD.n4528 19.9534
R17360 VDD.n4465 VDD.n4464 19.9534
R17361 VDD.n4497 VDD.n4496 19.9534
R17362 VDD.n4257 VDD.n4256 19.9534
R17363 VDD.n3714 VDD.n3700 19.9534
R17364 VDD.n3657 VDD.n3210 19.9534
R17365 VDD.n3603 VDD.n3602 19.9534
R17366 VDD.n3616 VDD.n3615 19.9534
R17367 VDD.n3627 VDD.n3571 19.9534
R17368 VDD.n3552 VDD.n3551 19.9534
R17369 VDD.n3769 VDD.n3768 19.9534
R17370 VDD.n3784 VDD.n3187 19.9534
R17371 VDD.n2942 VDD.n2389 19.9534
R17372 VDD.n2937 VDD.n2936 19.9534
R17373 VDD.n2915 VDD.n2914 19.9534
R17374 VDD.n2873 VDD.n2872 19.9534
R17375 VDD.n2359 VDD.n2289 19.9534
R17376 VDD.n2742 VDD.n2741 19.9534
R17377 VDD.n2635 VDD.n2482 19.9534
R17378 VDD.n2650 VDD.n2649 19.9534
R17379 VDD.n2650 VDD.n2473 19.9534
R17380 VDD.n2042 VDD.n1550 19.9534
R17381 VDD.n1855 VDD.n1596 19.9534
R17382 VDD.n1771 VDD.n1770 19.9534
R17383 VDD.n2115 VDD.n1519 19.9534
R17384 VDD.n2162 VDD.n2127 19.9534
R17385 VDD.n924 VDD.n923 19.9534
R17386 VDD.n1301 VDD.n1300 19.9534
R17387 VDD.n1469 VDD.n1410 19.9534
R17388 VDD.n381 VDD.n380 19.828
R17389 VDD.n380 VDD.n372 19.828
R17390 VDD.n2898 VDD.n2897 19.7491
R17391 VDD.n2893 VDD.n2416 19.7491
R17392 VDD.n3058 VDD.n3057 19.7491
R17393 VDD.n4187 VDD.n4145 19.577
R17394 VDD.n4171 VDD.n4161 19.577
R17395 VDD.n3954 VDD.n3919 19.577
R17396 VDD.n3953 VDD.n3952 19.577
R17397 VDD.n3948 VDD.n3923 19.577
R17398 VDD.n3471 VDD.n3470 19.577
R17399 VDD.n3348 VDD.n3347 19.577
R17400 VDD.n3337 VDD.n3327 19.577
R17401 VDD.n3150 VDD.n3149 19.577
R17402 VDD.n3144 VDD.n3143 19.577
R17403 VDD.n2861 VDD.n2860 19.577
R17404 VDD.n2530 VDD.n2529 19.577
R17405 VDD.n2699 VDD.n2698 19.577
R17406 VDD.n2587 VDD.n2577 19.577
R17407 VDD.n2322 VDD.n2312 19.577
R17408 VDD.n1807 VDD.n1806 19.577
R17409 VDD.n1717 VDD.n1685 19.577
R17410 VDD.n1711 VDD.n1688 19.577
R17411 VDD.n1703 VDD.n1693 19.577
R17412 VDD.n2021 VDD.n1955 19.577
R17413 VDD.n2206 VDD.n2196 19.577
R17414 VDD.n965 VDD.n840 19.577
R17415 VDD.n958 VDD.n957 19.577
R17416 VDD.n904 VDD.n901 19.577
R17417 VDD.n933 VDD.n932 19.577
R17418 VDD.n945 VDD.n944 19.577
R17419 VDD.n1335 VDD.n724 19.577
R17420 VDD.n1283 VDD.n1282 19.577
R17421 VDD.n1251 VDD.n1250 19.577
R17422 VDD.n1172 VDD.n1140 19.577
R17423 VDD.n1461 VDD.n1460 19.577
R17424 VDD.n1448 VDD.n1428 19.577
R17425 VDD.n1442 VDD.n1432 19.577
R17426 VDD.n417 VDD.n359 19.4467
R17427 VDD.n418 VDD.n417 19.4467
R17428 VDD.n2754 VDD.n2753 19.2005
R17429 VDD.n1730 VDD.n1729 19.2005
R17430 VDD.n2105 VDD.n1521 19.2005
R17431 VDD.n2221 VDD.n2220 19.2005
R17432 VDD.n4512 VDD.n4511 18.824
R17433 VDD.n4359 VDD.n4079 18.824
R17434 VDD.n3653 VDD.n3652 18.824
R17435 VDD.n3101 VDD.n3098 18.824
R17436 VDD.n3067 VDD.n3066 18.824
R17437 VDD.n1995 VDD.n1968 18.824
R17438 VDD.n2267 VDD.n1510 18.824
R17439 VDD.n926 VDD.n888 18.824
R17440 VDD.n1347 VDD.n1346 18.824
R17441 VDD.n1157 VDD.n1154 18.824
R17442 VDD.n1156 VDD.n1155 18.824
R17443 VDD.n706 VDD.n703 18.824
R17444 VDD.n4308 VDD.n4307 18.7213
R17445 VDD.t2265 VDD.t892 18.4634
R17446 VDD.t808 VDD.t1822 18.4634
R17447 VDD.t2345 VDD.t1393 18.4634
R17448 VDD.t3312 VDD.t3501 18.4634
R17449 VDD.n2894 VDD.t493 18.4634
R17450 VDD.n2896 VDD.t1020 18.4634
R17451 VDD.t1480 VDD.t854 18.4634
R17452 VDD.t433 VDD.t441 18.4634
R17453 VDD.t435 VDD.t2899 18.4634
R17454 VDD.t869 VDD.t744 18.4634
R17455 VDD.t2757 VDD.t746 18.4634
R17456 VDD.t169 VDD.t3040 18.4634
R17457 VDD.t826 VDD.t654 18.4634
R17458 VDD.t910 VDD.t1898 18.4634
R17459 VDD.t2857 VDD.t1901 18.4634
R17460 VDD.t591 VDD.t785 18.4634
R17461 VDD.n4621 VDD.n4609 18.4476
R17462 VDD.n4317 VDD.n4281 18.4476
R17463 VDD.n4209 VDD.n4208 18.4476
R17464 VDD.n3601 VDD.n3584 18.4476
R17465 VDD.n3528 VDD.n3255 18.4476
R17466 VDD.n3443 VDD.n3401 18.4476
R17467 VDD.n2860 VDD.n2859 18.4476
R17468 VDD.n2538 VDD.n2537 18.4476
R17469 VDD.n2694 VDD.n2693 18.4476
R17470 VDD.n2037 VDD.n2036 18.4476
R17471 VDD.n1734 VDD.n1671 18.4476
R17472 VDD.n1116 VDD.n1115 18.4476
R17473 VDD.n979 VDD.n978 18.4476
R17474 VDD.n1354 VDD.n1353 18.4476
R17475 VDD.n1225 VDD.n1224 18.4476
R17476 VDD.n1497 VDD.n701 18.4476
R17477 VDD.n2904 VDD.n2409 18.2862
R17478 VDD.n3063 VDD.n2362 18.2862
R17479 VDD.n3053 VDD.n3052 18.2862
R17480 VDD.n1831 VDD.n1616 18.2862
R17481 VDD.n158 VDD.n125 18.2003
R17482 VDD.n4614 VDD.n4613 18.0711
R17483 VDD.n4581 VDD.n3991 18.0711
R17484 VDD.n4541 VDD.n4014 18.0711
R17485 VDD.n4406 VDD.n4405 18.0711
R17486 VDD.n3503 VDD.n3270 18.0711
R17487 VDD.n3415 VDD.n3414 18.0711
R17488 VDD.n2914 VDD.n2913 18.0711
R17489 VDD.n2801 VDD.n2431 18.0711
R17490 VDD.n2782 VDD.n2780 18.0711
R17491 VDD.n2046 VDD.n1550 18.0711
R17492 VDD.n1838 VDD.n1611 18.0711
R17493 VDD.n2080 VDD.n1530 18.0711
R17494 VDD.n2226 VDD.n2225 18.0711
R17495 VDD.n2220 VDD.n2219 18.0711
R17496 VDD.n953 VDD.n847 18.0711
R17497 VDD.n1190 VDD.n1133 18.0711
R17498 VDD.n687 VDD.n636 18.0711
R17499 VDD.n1811 VDD.n1625 17.9205
R17500 VDD.n4245 VDD.n4110 17.6946
R17501 VDD.n3603 VDD.n3581 17.6946
R17502 VDD.n3557 VDD.n3239 17.6946
R17503 VDD.n2597 VDD.n2492 17.6946
R17504 VDD.n648 VDD.n647 17.6181
R17505 VDD.n144 VDD.n143 17.5829
R17506 VDD.n300 VDD.n297 17.4665
R17507 VDD.n3912 VDD.n3911 17.3181
R17508 VDD.n4613 VDD.n3900 17.3181
R17509 VDD.n4672 VDD.n3900 17.3181
R17510 VDD.n4630 VDD.n4629 17.3181
R17511 VDD.n4582 VDD.n4581 17.3181
R17512 VDD.n4583 VDD.n4582 17.3181
R17513 VDD.n4565 VDD.n4564 17.3181
R17514 VDD.n4535 VDD.n4534 17.3181
R17515 VDD.n4536 VDD.n4535 17.3181
R17516 VDD.n4506 VDD.n4505 17.3181
R17517 VDD.n4328 VDD.n4327 17.3181
R17518 VDD.n3725 VDD.n3695 17.3181
R17519 VDD.n3722 VDD.n3695 17.3181
R17520 VDD.n3734 VDD.n3691 17.3181
R17521 VDD.n3656 VDD.n3655 17.3181
R17522 VDD.n3226 VDD.n3223 17.3181
R17523 VDD.n3615 VDD.n3614 17.3181
R17524 VDD.n3614 VDD.n3613 17.3181
R17525 VDD.n3365 VDD.n3364 17.3181
R17526 VDD.n3366 VDD.n3365 17.3181
R17527 VDD.n3798 VDD.n3182 17.3181
R17528 VDD.n3801 VDD.n3182 17.3181
R17529 VDD.n3845 VDD.n3844 17.3181
R17530 VDD.n3844 VDD.n3843 17.3181
R17531 VDD.n2859 VDD.n2838 17.3181
R17532 VDD.n3028 VDD.n2281 17.3181
R17533 VDD.n3084 VDD.n2281 17.3181
R17534 VDD.n2772 VDD.n2445 17.3181
R17535 VDD.n2745 VDD.n2460 17.3181
R17536 VDD.n2604 VDD.n2603 17.3181
R17537 VDD.n2691 VDD.n2669 17.3181
R17538 VDD.n2688 VDD.n2669 17.3181
R17539 VDD.n2064 VDD.n1538 17.3181
R17540 VDD.n2140 VDD.n2139 17.3181
R17541 VDD.n1319 VDD.n1318 17.3181
R17542 VDD.n1318 VDD.n729 17.3181
R17543 VDD.n2770 VDD.n2769 17.2853
R17544 VDD.n4529 VDD.n4023 16.9417
R17545 VDD.n4431 VDD.n4430 16.9417
R17546 VDD.n4395 VDD.n4394 16.9417
R17547 VDD.n3429 VDD.n3427 16.9417
R17548 VDD.n3761 VDD.n3197 16.9417
R17549 VDD.n3839 VDD.n3838 16.9417
R17550 VDD.n2861 VDD.n2835 16.9417
R17551 VDD.n1872 VDD.n1590 16.9417
R17552 VDD.n1950 VDD.n1948 16.9417
R17553 VDD.t2325 VDD.t1884 16.785
R17554 VDD.t417 VDD.t1131 16.785
R17555 VDD.t2489 VDD.t2475 16.785
R17556 VDD.t516 VDD.t960 16.785
R17557 VDD.t423 VDD.t1334 16.785
R17558 VDD.t1095 VDD.t1505 16.785
R17559 VDD.t3270 VDD.t758 16.785
R17560 VDD.t2909 VDD.t2712 16.785
R17561 VDD.t1236 VDD.t3332 16.785
R17562 VDD.t1726 VDD.t3514 16.785
R17563 VDD.t3634 VDD.t2697 16.785
R17564 VDD.t2107 VDD.t2696 16.785
R17565 VDD.t900 VDD.t2773 16.785
R17566 VDD.t353 VDD.t2684 16.785
R17567 VDD.t355 VDD.t2680 16.785
R17568 VDD.t351 VDD.t2686 16.785
R17569 VDD.t357 VDD.t2636 16.785
R17570 VDD.n316 VDD.t1770 16.7394
R17571 VDD.n3792 VDD.n3791 16.619
R17572 VDD.n4501 VDD.n4040 16.5652
R17573 VDD.n4340 VDD.n4095 16.5652
R17574 VDD.n2798 VDD.n2431 16.5652
R17575 VDD.n2780 VDD.n2779 16.5652
R17576 VDD.n2771 VDD.n2770 16.5652
R17577 VDD.n684 VDD.n636 16.5652
R17578 VDD.n4609 VDD.n4606 16.1887
R17579 VDD.n4208 VDD.n4207 16.1887
R17580 VDD.n3529 VDD.n3528 16.1887
R17581 VDD.n3446 VDD.n3401 16.1887
R17582 VDD.n3776 VDD.n3190 16.1887
R17583 VDD.n3797 VDD.n3796 16.1887
R17584 VDD.n2693 VDD.n2692 16.1887
R17585 VDD.n2036 VDD.n2035 16.1887
R17586 VDD.n2003 VDD.n1965 16.1887
R17587 VDD.n1737 VDD.n1671 16.1887
R17588 VDD.n978 VDD.n977 16.1887
R17589 VDD.n1224 VDD.n1223 16.1887
R17590 VDD.n1163 VDD.n1162 16.1887
R17591 VDD.n1484 VDD.n1483 16.1887
R17592 VDD.n3911 VDD.n3908 15.8123
R17593 VDD.n4652 VDD.n3982 15.8123
R17594 VDD.n4645 VDD.n4597 15.8123
R17595 VDD.n4432 VDD.n4431 15.8123
R17596 VDD.n4360 VDD.n4359 15.8123
R17597 VDD.n3560 VDD.n3234 15.8123
R17598 VDD.n3541 VDD.n3249 15.8123
R17599 VDD.n3875 VDD.n3101 15.8123
R17600 VDD.n2958 VDD.n2957 15.8123
R17601 VDD.n3068 VDD.n3067 15.8123
R17602 VDD.n2794 VDD.n2793 15.8123
R17603 VDD.n2605 VDD.n2604 15.8123
R17604 VDD.n2609 VDD.n2489 15.8123
R17605 VDD.n2699 VDD.n2663 15.8123
R17606 VDD.n2070 VDD.n2069 15.8123
R17607 VDD.n1992 VDD.n1968 15.8123
R17608 VDD.n1808 VDD.n1807 15.8123
R17609 VDD.n1786 VDD.n1638 15.8123
R17610 VDD.n1740 VDD.n1739 15.8123
R17611 VDD.n2258 VDD.n1510 15.8123
R17612 VDD.n1091 VDD.n811 15.8123
R17613 VDD.n1029 VDD.n1028 15.8123
R17614 VDD.n888 VDD.n885 15.8123
R17615 VDD.n1346 VDD.n1345 15.8123
R17616 VDD.n1193 VDD.n1192 15.8123
R17617 VDD.n1155 VDD.n787 15.8123
R17618 VDD.n1486 VDD.n706 15.8123
R17619 VDD.n2889 VDD.n2418 15.7262
R17620 VDD.n1812 VDD.n1811 15.7262
R17621 VDD.n4649 VDD.n3985 15.4358
R17622 VDD.n4281 VDD.n4280 15.4358
R17623 VDD.n4251 VDD.n4250 15.4358
R17624 VDD.n3553 VDD.n3239 15.4358
R17625 VDD.n2713 VDD.n2712 15.4358
R17626 VDD.n1732 VDD.n1731 15.4358
R17627 VDD.n1154 VDD.n1153 15.4358
R17628 VDD.n2901 VDD.n2409 15.3605
R17629 VDD.n3060 VDD.n2362 15.3605
R17630 VDD.n3050 VDD.n3049 15.3605
R17631 VDD.n3973 VDD.n3972 15.1657
R17632 VDD.t465 VDD.t3162 15.1065
R17633 VDD.t1215 VDD.t3235 15.1065
R17634 VDD.t2397 VDD.t1057 15.1065
R17635 VDD.t2299 VDD.t1624 15.1065
R17636 VDD.t1504 VDD.t929 15.1065
R17637 VDD.t727 VDD.t1419 15.1065
R17638 VDD.t948 VDD.t3082 15.1065
R17639 VDD.t49 VDD.t3174 15.1065
R17640 VDD.t3381 VDD.t445 15.1065
R17641 VDD.t1600 VDD.t2327 15.1065
R17642 VDD.t2984 VDD.t2508 15.1065
R17643 VDD.t3302 VDD.t1837 15.1065
R17644 VDD.t3274 VDD.t1525 15.1065
R17645 VDD.t45 VDD.t698 15.1065
R17646 VDD.t786 VDD.t3722 15.1065
R17647 VDD.n3642 VDD.n3641 15.0593
R17648 VDD.n3633 VDD.n3229 15.0593
R17649 VDD.n2076 VDD.n1530 15.0593
R17650 VDD.n1879 VDD.n1878 15.0593
R17651 VDD.n1208 VDD.n1207 15.0593
R17652 VDD.n1397 VDD.n1396 15.0593
R17653 VDD.n2847 VDD.n2413 14.9948
R17654 VDD.n47 VDD.n46 14.7184
R17655 VDD.n25 VDD.n11 14.7184
R17656 VDD.n4425 VDD.n4424 14.6829
R17657 VDD.n2598 VDD.n2597 14.6829
R17658 VDD.n2139 VDD.n1509 14.6829
R17659 VDD.n4597 VDD.n4596 14.6829
R17660 VDD.n4566 VDD.n4565 14.6829
R17661 VDD.n3418 VDD.n3415 14.6829
R17662 VDD.n3768 VDD.n3767 14.6829
R17663 VDD.n3788 VDD.n3187 14.6829
R17664 VDD.n2916 VDD.n2915 14.6829
R17665 VDD.n923 VDD.n922 14.6829
R17666 VDD.n1379 VDD.n1378 14.6829
R17667 VDD.n1827 VDD.n1616 14.6291
R17668 VDD.n3974 VDD.n3973 14.4912
R17669 VDD.n57 VDD.n56 14.4822
R17670 VDD.n20 VDD.n19 14.4822
R17671 VDD.n308 VDD.n296 14.4039
R17672 VDD.n310 VDD.n301 14.4039
R17673 VDD.n4244 VDD.n4243 14.3064
R17674 VDD.n3429 VDD.n3408 14.3064
R17675 VDD.n3820 VDD.n3817 14.3064
R17676 VDD.n2772 VDD.n2771 14.3064
R17677 VDD.n2070 VDD.n1532 14.3064
R17678 VDD.n2074 VDD.n1532 14.3064
R17679 VDD.n2076 VDD.n2075 14.3064
R17680 VDD.n987 VDD.n986 14.3064
R17681 VDD.n4653 VDD.n4652 14.2735
R17682 VDD.n4393 VDD.n4068 14.2735
R17683 VDD.n4225 VDD.n4123 14.2735
R17684 VDD.n3753 VDD.n3201 14.2735
R17685 VDD.n3165 VDD.n3117 14.2735
R17686 VDD.n3045 VDD.n3044 14.2735
R17687 VDD.n3036 VDD.n3035 14.2735
R17688 VDD.n1912 VDD.n1911 14.2735
R17689 VDD.n327 VDD.n189 14.2313
R17690 VDD.n328 VDD.n327 14.2313
R17691 VDD.n325 VDD.n299 14.2313
R17692 VDD.n325 VDD.n324 14.2313
R17693 VDD.n311 VDD.n310 14.2313
R17694 VDD.n308 VDD.n307 14.2313
R17695 VDD.n2757 VDD.n2450 14.2227
R17696 VDD.n2620 VDD.n2487 13.9478
R17697 VDD.n4488 VDD.n4441 13.9299
R17698 VDD.n4179 VDD.n4178 13.9299
R17699 VDD.n3757 VDD.n3197 13.9299
R17700 VDD.n2944 VDD.n2943 13.9299
R17701 VDD.n2714 VDD.n2713 13.9299
R17702 VDD.n1783 VDD.n1782 13.9299
R17703 VDD.n1752 VDD.n1751 13.9299
R17704 VDD.n1715 VDD.n1688 13.9299
R17705 VDD.n3059 VDD.n3058 13.8976
R17706 VDD.n2822 VDD.n2416 13.8976
R17707 VDD.n1256 VDD.n760 13.8432
R17708 VDD.n4374 VDD.n4373 13.5534
R17709 VDD.n4336 VDD.n4335 13.5534
R17710 VDD.n4336 VDD.n4095 13.5534
R17711 VDD.n3597 VDD.n3584 13.5534
R17712 VDD.n3564 VDD.n3234 13.5534
R17713 VDD.n3551 VDD.n3243 13.5534
R17714 VDD.n2938 VDD.n2389 13.5534
R17715 VDD.n2871 VDD.n2832 13.5534
R17716 VDD.n2596 VDD.n2494 13.5534
R17717 VDD.n3034 VDD.n3033 13.5534
R17718 VDD.n2803 VDD.n2802 13.5534
R17719 VDD.n2796 VDD.n2795 13.5534
R17720 VDD.n2757 VDD.n2756 13.5534
R17721 VDD.n2755 VDD.n2754 13.5534
R17722 VDD.n2081 VDD.n2080 13.5534
R17723 VDD.n1911 VDD.n1906 13.5534
R17724 VDD.n988 VDD.n987 13.5534
R17725 VDD.n1354 VDD.n712 13.5534
R17726 VDD.t419 VDD.t1133 13.4281
R17727 VDD.t760 VDD.t3282 13.4281
R17728 VDD.t682 VDD.t2453 13.4281
R17729 VDD.t1927 VDD.t1591 13.4281
R17730 VDD.t2504 VDD.t3111 13.4281
R17731 VDD.t2350 VDD.t3310 13.4281
R17732 VDD.t3700 VDD.t265 13.4281
R17733 VDD.t489 VDD.t1973 13.4281
R17734 VDD.t481 VDD.t3045 13.4281
R17735 VDD.t3044 VDD.t2445 13.4281
R17736 VDD.t1262 VDD.t1113 13.4281
R17737 VDD.t326 VDD.t3172 13.4281
R17738 VDD.t3439 VDD.t25 13.4281
R17739 VDD.t2986 VDD.t3490 13.4281
R17740 VDD.t1815 VDD.t2280 13.4281
R17741 VDD.t1107 VDD.t2794 13.4281
R17742 VDD.t324 VDD.t3000 13.4281
R17743 VDD.t1238 VDD.t3334 13.4281
R17744 VDD.n1201 VDD.t1463 13.4281
R17745 VDD.t3233 VDD.t1675 13.4281
R17746 VDD.t269 VDD.t976 13.4281
R17747 VDD.t2203 VDD.t1904 13.4281
R17748 VDD.t3064 VDD.t1654 13.4281
R17749 VDD.t3070 VDD.t1656 13.4281
R17750 VDD.t3059 VDD.t2195 13.4281
R17751 VDD.t3066 VDD.t2193 13.4281
R17752 VDD.n415 VDD.n359 13.2148
R17753 VDD.n415 VDD.n414 13.2148
R17754 VDD.n370 VDD.n365 13.2148
R17755 VDD.n370 VDD.n362 13.2148
R17756 VDD.n376 VDD.n372 13.2148
R17757 VDD.n376 VDD.n368 13.2148
R17758 VDD.n4521 VDD.n4030 13.177
R17759 VDD.n4428 VDD.n4043 13.177
R17760 VDD.n4266 VDD.n4096 13.177
R17761 VDD.n4232 VDD.n4118 13.177
R17762 VDD.n4181 VDD.n4180 13.177
R17763 VDD.n4180 VDD.n4179 13.177
R17764 VDD.n4177 VDD.n4176 13.177
R17765 VDD.n3756 VDD.n3199 13.177
R17766 VDD.n3343 VDD.n3317 13.177
R17767 VDD.n3867 VDD.n3178 13.177
R17768 VDD.n2565 VDD.n2495 13.177
R17769 VDD.n2593 VDD.n2495 13.177
R17770 VDD.n2291 VDD.n2289 13.177
R17771 VDD.n2806 VDD.n2803 13.177
R17772 VDD.n1859 VDD.n1596 13.177
R17773 VDD.n1800 VDD.n1799 13.177
R17774 VDD.n1716 VDD.n1715 13.177
R17775 VDD.n1937 VDD.n1565 13.177
R17776 VDD.n2249 VDD.n2248 13.177
R17777 VDD.n1100 VDD.n1099 13.177
R17778 VDD.n910 VDD.n898 13.177
R17779 VDD.n1403 VDD.n712 13.177
R17780 VDD.n1479 VDD.n1478 13.177
R17781 VDD.n3499 VDD.n3498 13.1662
R17782 VDD.n2910 VDD.n2907 13.1662
R17783 VDD.n3000 VDD.n2999 13.1662
R17784 VDD.n2816 VDD.n2815 13.1662
R17785 VDD.n4548 VDD.n4547 12.8005
R17786 VDD.n4394 VDD.n4393 12.8005
R17787 VDD.n4373 VDD.n4372 12.8005
R17788 VDD.n4343 VDD.n4092 12.8005
R17789 VDD.n4340 VDD.n4096 12.8005
R17790 VDD.n3691 VDD.n3688 12.8005
R17791 VDD.n3574 VDD.n3571 12.8005
R17792 VDD.n3519 VDD.n3258 12.8005
R17793 VDD.n3757 VDD.n3756 12.8005
R17794 VDD.n3789 VDD.n3788 12.8005
R17795 VDD.n3874 VDD.n3873 12.8005
R17796 VDD.n3343 VDD.n3342 12.8005
R17797 VDD.n2899 VDD.n2898 12.8005
R17798 VDD.n2593 VDD.n2592 12.8005
R17799 VDD.n2055 VDD.n2054 12.8005
R17800 VDD.n1989 VDD.n1988 12.8005
R17801 VDD.n1872 VDD.n1867 12.8005
R17802 VDD.n1861 VDD.n1594 12.8005
R17803 VDD.n1793 VDD.n1792 12.8005
R17804 VDD.n1931 VDD.n1930 12.8005
R17805 VDD.n2256 VDD.n2255 12.8005
R17806 VDD.n1114 VDD.n1113 12.8005
R17807 VDD.n1093 VDD.n1092 12.8005
R17808 VDD.n1030 VDD.n1027 12.8005
R17809 VDD.n1209 VDD.n1208 12.8005
R17810 VDD.n1162 VDD.n1161 12.8005
R17811 VDD.n1202 VDD.n789 12.8005
R17812 VDD.n1485 VDD.n1484 12.8005
R17813 VDD.n426 VDD.n425 12.8005
R17814 VDD.n4397 VDD.n4396 12.424
R17815 VDD.n4329 VDD.n4328 12.424
R17816 VDD.n3566 VDD.n3229 12.424
R17817 VDD.n2865 VDD.n2835 12.424
R17818 VDD.n2991 VDD.n2990 12.424
R17819 VDD.n1982 VDD.n1981 12.424
R17820 VDD.n953 VDD.n844 12.424
R17821 VDD.n1373 VDD.n701 12.424
R17822 VDD.n1454 VDD.n1453 12.424
R17823 VDD.n4643 VDD.n4642 12.0476
R17824 VDD.n4490 VDD.n4488 12.0476
R17825 VDD.n3654 VDD.n3653 12.0476
R17826 VDD.n3035 VDD.n3034 12.0476
R17827 VDD.n2795 VDD.n2794 12.0476
R17828 VDD.n2778 VDD.n2777 12.0476
R17829 VDD.n2756 VDD.n2755 12.0476
R17830 VDD.n2680 VDD.n2679 12.0476
R17831 VDD.n2061 VDD.n1541 12.0476
R17832 VDD.n1840 VDD.n1839 12.0476
R17833 VDD.n1246 VDD.n763 12.0147
R17834 VDD.n1239 VDD.n1237 12.0147
R17835 VDD.n315 VDD.n314 11.7586
R17836 VDD.t3159 VDD.t467 11.7496
R17837 VDD.t1213 VDD.t3237 11.7496
R17838 VDD.t1073 VDD.t2816 11.7496
R17839 VDD.t2604 VDD.t2429 11.7496
R17840 VDD.t293 VDD.t2745 11.7496
R17841 VDD.t529 VDD.t1959 11.7496
R17842 VDD.t1929 VDD.t672 11.7496
R17843 VDD.t33 VDD.n3064 11.7496
R17844 VDD.t2530 VDD.t3464 11.7496
R17845 VDD.t3749 VDD.t1159 11.7496
R17846 VDD.t2932 VDD.t3206 11.7496
R17847 VDD.t3741 VDD.t2215 11.7496
R17848 VDD.t263 VDD.t2134 11.7496
R17849 VDD.t2995 VDD.t559 11.7496
R17850 VDD.t2571 VDD.t2770 11.7496
R17851 VDD.t983 VDD.t3714 11.7496
R17852 VDD.n4189 VDD.n4188 11.6711
R17853 VDD.n3171 VDD.n3169 11.6711
R17854 VDD.n2856 VDD.n2838 11.6711
R17855 VDD.n1991 VDD.n1989 11.6711
R17856 VDD.n621 VDD.n620 11.4713
R17857 VDD.n538 VDD.n537 11.4713
R17858 VDD.n458 VDD.n457 11.4713
R17859 VDD.n209 VDD.n208 11.4643
R17860 VDD.n80 VDD.n62 11.4138
R17861 VDD.n44 VDD.n26 11.4138
R17862 VDD.n2881 VDD.n2827 11.3376
R17863 VDD.n4465 VDD.n4452 11.2946
R17864 VDD.n4245 VDD.n4244 11.2946
R17865 VDD.n3433 VDD.n3408 11.2946
R17866 VDD.n3462 VDD.n3461 11.2946
R17867 VDD.n994 VDD.n826 11.2946
R17868 VDD.n1219 VDD.n777 11.2946
R17869 VDD.n1469 VDD.n1468 11.2946
R17870 VDD.n676 VDD.n648 11.2946
R17871 VDD.n56 VDD.t1780 11.1031
R17872 VDD.n19 VDD.t3073 11.1031
R17873 VDD.n3486 VDD.n3278 10.9719
R17874 VDD.n3051 VDD.n3050 10.9719
R17875 VDD.n2805 VDD.n2427 10.9719
R17876 VDD.n4630 VDD.n4604 10.9181
R17877 VDD.n4560 VDD.n4559 10.9181
R17878 VDD.n4375 VDD.n4074 10.9181
R17879 VDD.n4299 VDD.n4288 10.9181
R17880 VDD.n3595 VDD.n3594 10.9181
R17881 VDD.n3622 VDD.n3621 10.9181
R17882 VDD.n3505 VDD.n3504 10.9181
R17883 VDD.n2728 VDD.n2471 10.9181
R17884 VDD.n1997 VDD.n1996 10.9181
R17885 VDD.n1147 VDD.n1145 10.9181
R17886 VDD.n1379 VDD.n1369 10.9181
R17887 VDD.n153 VDD.n152 10.9067
R17888 VDD.n3976 VDD.n3913 10.5744
R17889 VDD.n166 VDD.n165 10.5561
R17890 VDD.n4306 VDD.n4286 10.5417
R17891 VDD.n3553 VDD.n3552 10.5417
R17892 VDD.n2513 VDD.n2511 10.5417
R17893 VDD.n1878 VDD.n1876 10.5417
R17894 VDD.n1237 VDD.n1236 10.5417
R17895 VDD.n1178 VDD.n1177 10.5417
R17896 VDD.n142 VDD.n141 10.5417
R17897 VDD.n143 VDD.n142 10.5417
R17898 VDD.n622 VDD.n621 10.4058
R17899 VDD.n539 VDD.n538 10.4058
R17900 VDD.n459 VDD.n458 10.4058
R17901 VDD.n3490 VDD.n3489 10.2405
R17902 VDD.n2881 VDD.n2880 10.2405
R17903 VDD.n1824 VDD.n1823 10.2405
R17904 VDD.n74 VDD.n73 10.1732
R17905 VDD.n34 VDD.n33 10.1732
R17906 VDD.n4527 VDD.n4526 10.1652
R17907 VDD.n2048 VDD.n2047 10.1652
R17908 VDD.n1787 VDD.n1786 10.1652
R17909 VDD.n1731 VDD.n1730 10.1652
R17910 VDD.n2105 VDD.n2104 10.1652
R17911 VDD.n246 VDD.n244 10.1337
R17912 VDD.t2376 VDD.t455 10.0712
R17913 VDD.t2937 VDD.t1596 10.0712
R17914 VDD.t413 VDD.t2541 10.0712
R17915 VDD.t573 VDD.t2640 10.0712
R17916 VDD.t1522 VDD.t2271 10.0712
R17917 VDD.t3505 VDD.t1087 10.0712
R17918 VDD.n3635 VDD.t1747 10.0712
R17919 VDD.t2013 VDD.t931 10.0712
R17920 VDD.t2015 VDD.t933 10.0712
R17921 VDD.t1498 VDD.t3483 10.0712
R17922 VDD.t3486 VDD.t3337 10.0712
R17923 VDD.t2163 VDD.t2845 10.0712
R17924 VDD.t2849 VDD.t1296 10.0712
R17925 VDD.t1281 VDD.t3627 10.0712
R17926 VDD.t3226 VDD.t686 10.0712
R17927 VDD.t700 VDD.t23 10.0712
R17928 VDD.t307 VDD.t1146 10.0712
R17929 VDD.t3686 VDD.t896 10.0712
R17930 VDD.t1602 VDD.t2329 10.0712
R17931 VDD.t43 VDD.t1320 10.0712
R17932 VDD.t3481 VDD.t660 10.0712
R17933 VDD.n3852 VDD.n3851 9.78874
R17934 VDD.n1348 VDD.n717 9.78874
R17935 VDD.n1192 VDD.n1191 9.78874
R17936 VDD.n77 VDD.n70 9.78874
R17937 VDD.n41 VDD.n38 9.78874
R17938 VDD.n3803 VDD.n3801 9.73495
R17939 VDD.n1892 VDD.n1582 9.73273
R17940 VDD.n1895 VDD.n1894 9.73273
R17941 VDD.n2853 VDD.n2841 9.56172
R17942 VDD.n2850 VDD.n2844 9.56172
R17943 VDD.n2845 VDD.n2413 9.56172
R17944 VDD.n3051 VDD.n3010 9.56172
R17945 VDD.n3977 VDD.n3976 9.41227
R17946 VDD.n4567 VDD.n4566 9.41227
R17947 VDD.n4471 VDD.n4470 9.41227
R17948 VDD.n4409 VDD.n4051 9.41227
R17949 VDD.n4365 VDD.n4364 9.41227
R17950 VDD.n4322 VDD.n4321 9.41227
R17951 VDD.n4204 VDD.n4203 9.41227
R17952 VDD.n3721 VDD.n3720 9.41227
R17953 VDD.n3744 VDD.n3685 9.41227
R17954 VDD.n3505 VDD.n3265 9.41227
R17955 VDD.n3448 VDD.n3447 9.41227
R17956 VDD.n3367 VDD.n3300 9.41227
R17957 VDD.n2631 VDD.n2482 9.41227
R17958 VDD.n2049 VDD.n2048 9.41227
R17959 VDD.n2034 VDD.n1556 9.41227
R17960 VDD.n2020 VDD.n2019 9.41227
R17961 VDD.n2158 VDD.n2127 9.41227
R17962 VDD.n2158 VDD.n2157 9.41227
R17963 VDD.n2229 VDD.n2182 9.41227
R17964 VDD.n1112 VDD.n802 9.41227
R17965 VDD.n1049 VDD.n1015 9.41227
R17966 VDD.n996 VDD.n823 9.41227
R17967 VDD.n1341 VDD.n1340 9.41227
R17968 VDD.n629 VDD.n612 9.41227
R17969 VDD.n546 VDD.n529 9.41227
R17970 VDD.n466 VDD.n449 9.41227
R17971 VDD.n1928 VDD.n1570 9.3794
R17972 VDD.n4172 VDD.n4171 9.3005
R17973 VDD.n4173 VDD.n4161 9.3005
R17974 VDD.n4175 VDD.n4174 9.3005
R17975 VDD.n4176 VDD.n4158 9.3005
R17976 VDD.n4177 VDD.n4157 9.3005
R17977 VDD.n4178 VDD.n4154 9.3005
R17978 VDD.n4179 VDD.n4153 9.3005
R17979 VDD.n4180 VDD.n4150 9.3005
R17980 VDD.n4181 VDD.n4148 9.3005
R17981 VDD.n4182 VDD.n4146 9.3005
R17982 VDD.n4184 VDD.n4183 9.3005
R17983 VDD.n4185 VDD.n4145 9.3005
R17984 VDD.n4187 VDD.n4186 9.3005
R17985 VDD.n4188 VDD.n4143 9.3005
R17986 VDD.n4189 VDD.n4142 9.3005
R17987 VDD.n4190 VDD.n4140 9.3005
R17988 VDD.n4192 VDD.n4191 9.3005
R17989 VDD.n4194 VDD.n4193 9.3005
R17990 VDD.n4197 VDD.n4137 9.3005
R17991 VDD.n4198 VDD.n4136 9.3005
R17992 VDD.n4200 VDD.n4199 9.3005
R17993 VDD.n4202 VDD.n4201 9.3005
R17994 VDD.n4203 VDD.n4133 9.3005
R17995 VDD.n4205 VDD.n4204 9.3005
R17996 VDD.n4207 VDD.n4206 9.3005
R17997 VDD.n4209 VDD.n4129 9.3005
R17998 VDD.n4211 VDD.n4210 9.3005
R17999 VDD.n4213 VDD.n4212 9.3005
R18000 VDD.n4215 VDD.n4127 9.3005
R18001 VDD.n4218 VDD.n4217 9.3005
R18002 VDD.n4219 VDD.n4126 9.3005
R18003 VDD.n4221 VDD.n4220 9.3005
R18004 VDD.n4222 VDD.n4124 9.3005
R18005 VDD.n4226 VDD.n4225 9.3005
R18006 VDD.n4227 VDD.n4123 9.3005
R18007 VDD.n4229 VDD.n4228 9.3005
R18008 VDD.n4230 VDD.n4122 9.3005
R18009 VDD.n4231 VDD.n4119 9.3005
R18010 VDD.n4233 VDD.n4232 9.3005
R18011 VDD.n4234 VDD.n4118 9.3005
R18012 VDD.n4236 VDD.n4235 9.3005
R18013 VDD.n4237 VDD.n4116 9.3005
R18014 VDD.n4239 VDD.n4238 9.3005
R18015 VDD.n4240 VDD.n4115 9.3005
R18016 VDD.n4242 VDD.n4241 9.3005
R18017 VDD.n4243 VDD.n4113 9.3005
R18018 VDD.n4244 VDD.n4111 9.3005
R18019 VDD.n4246 VDD.n4245 9.3005
R18020 VDD.n4247 VDD.n4110 9.3005
R18021 VDD.n4249 VDD.n4248 9.3005
R18022 VDD.n4250 VDD.n4108 9.3005
R18023 VDD.n4251 VDD.n4105 9.3005
R18024 VDD.n4253 VDD.n4252 9.3005
R18025 VDD.n4254 VDD.n4104 9.3005
R18026 VDD.n4256 VDD.n4255 9.3005
R18027 VDD.n4257 VDD.n4101 9.3005
R18028 VDD.n4259 VDD.n4258 9.3005
R18029 VDD.n4260 VDD.n4100 9.3005
R18030 VDD.n4262 VDD.n4261 9.3005
R18031 VDD.n4265 VDD.n4097 9.3005
R18032 VDD.n4267 VDD.n4266 9.3005
R18033 VDD.n4268 VDD.n4096 9.3005
R18034 VDD.n4340 VDD.n4339 9.3005
R18035 VDD.n4338 VDD.n4095 9.3005
R18036 VDD.n4337 VDD.n4336 9.3005
R18037 VDD.n4335 VDD.n4269 9.3005
R18038 VDD.n4334 VDD.n4333 9.3005
R18039 VDD.n4332 VDD.n4331 9.3005
R18040 VDD.n4330 VDD.n4271 9.3005
R18041 VDD.n4327 VDD.n4326 9.3005
R18042 VDD.n4325 VDD.n4274 9.3005
R18043 VDD.n4324 VDD.n4323 9.3005
R18044 VDD.n4322 VDD.n4275 9.3005
R18045 VDD.n4321 VDD.n4320 9.3005
R18046 VDD.n4319 VDD.n4276 9.3005
R18047 VDD.n4318 VDD.n4317 9.3005
R18048 VDD.n4316 VDD.n4277 9.3005
R18049 VDD.n4313 VDD.n4312 9.3005
R18050 VDD.n4311 VDD.n4282 9.3005
R18051 VDD.n4310 VDD.n4309 9.3005
R18052 VDD.n4307 VDD.n4283 9.3005
R18053 VDD.n4306 VDD.n4304 9.3005
R18054 VDD.n4303 VDD.n4286 9.3005
R18055 VDD.n4302 VDD.n4301 9.3005
R18056 VDD.n4300 VDD.n4287 9.3005
R18057 VDD.n4299 VDD.n4297 9.3005
R18058 VDD.n4296 VDD.n4288 9.3005
R18059 VDD.n4295 VDD.n4294 9.3005
R18060 VDD.n4291 VDD.n4289 9.3005
R18061 VDD.n4094 VDD.n4093 9.3005
R18062 VDD.n4344 VDD.n4343 9.3005
R18063 VDD.n4347 VDD.n4346 9.3005
R18064 VDD.n4348 VDD.n4086 9.3005
R18065 VDD.n4350 VDD.n4349 9.3005
R18066 VDD.n4351 VDD.n4085 9.3005
R18067 VDD.n4353 VDD.n4352 9.3005
R18068 VDD.n4355 VDD.n4083 9.3005
R18069 VDD.n4356 VDD.n4080 9.3005
R18070 VDD.n4361 VDD.n4360 9.3005
R18071 VDD.n4362 VDD.n4079 9.3005
R18072 VDD.n4364 VDD.n4363 9.3005
R18073 VDD.n4366 VDD.n4078 9.3005
R18074 VDD.n4368 VDD.n4367 9.3005
R18075 VDD.n4369 VDD.n4077 9.3005
R18076 VDD.n4371 VDD.n4370 9.3005
R18077 VDD.n4374 VDD.n4075 9.3005
R18078 VDD.n4376 VDD.n4375 9.3005
R18079 VDD.n4377 VDD.n4074 9.3005
R18080 VDD.n4379 VDD.n4378 9.3005
R18081 VDD.n4380 VDD.n4073 9.3005
R18082 VDD.n4383 VDD.n4382 9.3005
R18083 VDD.n4385 VDD.n4384 9.3005
R18084 VDD.n4386 VDD.n4070 9.3005
R18085 VDD.n4390 VDD.n4389 9.3005
R18086 VDD.n4391 VDD.n4068 9.3005
R18087 VDD.n4393 VDD.n4392 9.3005
R18088 VDD.n4395 VDD.n4063 9.3005
R18089 VDD.n4396 VDD.n4061 9.3005
R18090 VDD.n4397 VDD.n4060 9.3005
R18091 VDD.n4398 VDD.n4056 9.3005
R18092 VDD.n4402 VDD.n4401 9.3005
R18093 VDD.n4403 VDD.n4055 9.3005
R18094 VDD.n4405 VDD.n4404 9.3005
R18095 VDD.n4406 VDD.n4054 9.3005
R18096 VDD.n4408 VDD.n4052 9.3005
R18097 VDD.n4410 VDD.n4409 9.3005
R18098 VDD.n4412 VDD.n4411 9.3005
R18099 VDD.n4417 VDD.n4416 9.3005
R18100 VDD.n4418 VDD.n4046 9.3005
R18101 VDD.n4420 VDD.n4419 9.3005
R18102 VDD.n4423 VDD.n4044 9.3005
R18103 VDD.n4426 VDD.n4425 9.3005
R18104 VDD.n4428 VDD.n4427 9.3005
R18105 VDD.n4429 VDD.n4041 9.3005
R18106 VDD.n4433 VDD.n4432 9.3005
R18107 VDD.n4434 VDD.n4040 9.3005
R18108 VDD.n4501 VDD.n4500 9.3005
R18109 VDD.n4499 VDD.n4039 9.3005
R18110 VDD.n4498 VDD.n4497 9.3005
R18111 VDD.n4496 VDD.n4435 9.3005
R18112 VDD.n4494 VDD.n4493 9.3005
R18113 VDD.n4492 VDD.n4491 9.3005
R18114 VDD.n4490 VDD.n4438 9.3005
R18115 VDD.n4488 VDD.n4487 9.3005
R18116 VDD.n4485 VDD.n4484 9.3005
R18117 VDD.n4483 VDD.n4442 9.3005
R18118 VDD.n4482 VDD.n4481 9.3005
R18119 VDD.n4480 VDD.n4479 9.3005
R18120 VDD.n4478 VDD.n4447 9.3005
R18121 VDD.n4475 VDD.n4474 9.3005
R18122 VDD.n4473 VDD.n4472 9.3005
R18123 VDD.n4471 VDD.n4451 9.3005
R18124 VDD.n4469 VDD.n4468 9.3005
R18125 VDD.n4467 VDD.n4452 9.3005
R18126 VDD.n4466 VDD.n4465 9.3005
R18127 VDD.n4464 VDD.n4453 9.3005
R18128 VDD.n4463 VDD.n4461 9.3005
R18129 VDD.n4460 VDD.n4454 9.3005
R18130 VDD.n4459 VDD.n4458 9.3005
R18131 VDD.n4456 VDD.n4038 9.3005
R18132 VDD.n4504 VDD.n4036 9.3005
R18133 VDD.n4507 VDD.n4506 9.3005
R18134 VDD.n4508 VDD.n4035 9.3005
R18135 VDD.n4510 VDD.n4509 9.3005
R18136 VDD.n4511 VDD.n4034 9.3005
R18137 VDD.n4512 VDD.n4033 9.3005
R18138 VDD.n4516 VDD.n4515 9.3005
R18139 VDD.n4517 VDD.n4032 9.3005
R18140 VDD.n4519 VDD.n4518 9.3005
R18141 VDD.n4520 VDD.n4031 9.3005
R18142 VDD.n4522 VDD.n4521 9.3005
R18143 VDD.n4524 VDD.n4523 9.3005
R18144 VDD.n4526 VDD.n4027 9.3005
R18145 VDD.n4527 VDD.n4026 9.3005
R18146 VDD.n4528 VDD.n4024 9.3005
R18147 VDD.n4530 VDD.n4529 9.3005
R18148 VDD.n4532 VDD.n4017 9.3005
R18149 VDD.n4534 VDD.n4533 9.3005
R18150 VDD.n4536 VDD.n4015 9.3005
R18151 VDD.n4538 VDD.n4537 9.3005
R18152 VDD.n4539 VDD.n4014 9.3005
R18153 VDD.n4541 VDD.n4540 9.3005
R18154 VDD.n4542 VDD.n4011 9.3005
R18155 VDD.n4544 VDD.n4543 9.3005
R18156 VDD.n4545 VDD.n4009 9.3005
R18157 VDD.n4547 VDD.n4546 9.3005
R18158 VDD.n4553 VDD.n4552 9.3005
R18159 VDD.n4554 VDD.n4002 9.3005
R18160 VDD.n4556 VDD.n4555 9.3005
R18161 VDD.n4558 VDD.n4001 9.3005
R18162 VDD.n4559 VDD.n3999 9.3005
R18163 VDD.n4561 VDD.n4560 9.3005
R18164 VDD.n4562 VDD.n3998 9.3005
R18165 VDD.n4564 VDD.n4563 9.3005
R18166 VDD.n4566 VDD.n3996 9.3005
R18167 VDD.n4567 VDD.n3995 9.3005
R18168 VDD.n4571 VDD.n4570 9.3005
R18169 VDD.n4572 VDD.n3994 9.3005
R18170 VDD.n4574 VDD.n4573 9.3005
R18171 VDD.n4575 VDD.n3992 9.3005
R18172 VDD.n4578 VDD.n4577 9.3005
R18173 VDD.n4579 VDD.n3991 9.3005
R18174 VDD.n4581 VDD.n4580 9.3005
R18175 VDD.n4583 VDD.n3988 9.3005
R18176 VDD.n4585 VDD.n4584 9.3005
R18177 VDD.n4586 VDD.n3987 9.3005
R18178 VDD.n4588 VDD.n4587 9.3005
R18179 VDD.n4589 VDD.n3986 9.3005
R18180 VDD.n4593 VDD.n4592 9.3005
R18181 VDD.n4594 VDD.n3985 9.3005
R18182 VDD.n4649 VDD.n4648 9.3005
R18183 VDD.n4647 VDD.n3983 9.3005
R18184 VDD.n4646 VDD.n4645 9.3005
R18185 VDD.n4644 VDD.n4595 9.3005
R18186 VDD.n4641 VDD.n4640 9.3005
R18187 VDD.n4639 VDD.n4638 9.3005
R18188 VDD.n4636 VDD.n4602 9.3005
R18189 VDD.n4634 VDD.n4633 9.3005
R18190 VDD.n4632 VDD.n4604 9.3005
R18191 VDD.n4631 VDD.n4630 9.3005
R18192 VDD.n4625 VDD.n4624 9.3005
R18193 VDD.n4623 VDD.n4606 9.3005
R18194 VDD.n4622 VDD.n4621 9.3005
R18195 VDD.n4619 VDD.n4607 9.3005
R18196 VDD.n4618 VDD.n4617 9.3005
R18197 VDD.n4616 VDD.n4611 9.3005
R18198 VDD.n4615 VDD.n4614 9.3005
R18199 VDD.n4613 VDD.n3897 9.3005
R18200 VDD.n4673 VDD.n4672 9.3005
R18201 VDD.n4671 VDD.n4669 9.3005
R18202 VDD.n4662 VDD.n3901 9.3005
R18203 VDD.n4661 VDD.n4660 9.3005
R18204 VDD.n4657 VDD.n3903 9.3005
R18205 VDD.n4656 VDD.n4655 9.3005
R18206 VDD.n4654 VDD.n4653 9.3005
R18207 VDD.n4652 VDD.n3906 9.3005
R18208 VDD.n3982 VDD.n3981 9.3005
R18209 VDD.n3980 VDD.n3908 9.3005
R18210 VDD.n3979 VDD.n3978 9.3005
R18211 VDD.n3977 VDD.n3909 9.3005
R18212 VDD.n3967 VDD.n3966 9.3005
R18213 VDD.n3965 VDD.n3916 9.3005
R18214 VDD.n3964 VDD.n3963 9.3005
R18215 VDD.n3961 VDD.n3917 9.3005
R18216 VDD.n3958 VDD.n3957 9.3005
R18217 VDD.n3956 VDD.n3919 9.3005
R18218 VDD.n3955 VDD.n3954 9.3005
R18219 VDD.n3953 VDD.n3920 9.3005
R18220 VDD.n3952 VDD.n3951 9.3005
R18221 VDD.n3950 VDD.n3923 9.3005
R18222 VDD.n3949 VDD.n3948 9.3005
R18223 VDD.n3947 VDD.n3924 9.3005
R18224 VDD.n3946 VDD.n3945 9.3005
R18225 VDD.n3944 VDD.n3943 9.3005
R18226 VDD.n3941 VDD.n3928 9.3005
R18227 VDD.n3939 VDD.n3938 9.3005
R18228 VDD.n3338 VDD.n3337 9.3005
R18229 VDD.n3339 VDD.n3327 9.3005
R18230 VDD.n3341 VDD.n3340 9.3005
R18231 VDD.n3344 VDD.n3343 9.3005
R18232 VDD.n3345 VDD.n3317 9.3005
R18233 VDD.n3347 VDD.n3346 9.3005
R18234 VDD.n3348 VDD.n3314 9.3005
R18235 VDD.n3350 VDD.n3349 9.3005
R18236 VDD.n3352 VDD.n3305 9.3005
R18237 VDD.n3354 VDD.n3353 9.3005
R18238 VDD.n3356 VDD.n3304 9.3005
R18239 VDD.n3361 VDD.n3360 9.3005
R18240 VDD.n3362 VDD.n3303 9.3005
R18241 VDD.n3364 VDD.n3363 9.3005
R18242 VDD.n3366 VDD.n3301 9.3005
R18243 VDD.n3368 VDD.n3367 9.3005
R18244 VDD.n3369 VDD.n3300 9.3005
R18245 VDD.n3371 VDD.n3370 9.3005
R18246 VDD.n3373 VDD.n3298 9.3005
R18247 VDD.n3375 VDD.n3374 9.3005
R18248 VDD.n3377 VDD.n3376 9.3005
R18249 VDD.n3378 VDD.n3295 9.3005
R18250 VDD.n3381 VDD.n3380 9.3005
R18251 VDD.n3383 VDD.n3382 9.3005
R18252 VDD.n3385 VDD.n3293 9.3005
R18253 VDD.n3391 VDD.n3390 9.3005
R18254 VDD.n3392 VDD.n3292 9.3005
R18255 VDD.n3466 VDD.n3465 9.3005
R18256 VDD.n3464 VDD.n3291 9.3005
R18257 VDD.n3463 VDD.n3462 9.3005
R18258 VDD.n3460 VDD.n3393 9.3005
R18259 VDD.n3458 VDD.n3457 9.3005
R18260 VDD.n3456 VDD.n3455 9.3005
R18261 VDD.n3453 VDD.n3397 9.3005
R18262 VDD.n3452 VDD.n3451 9.3005
R18263 VDD.n3450 VDD.n3398 9.3005
R18264 VDD.n3449 VDD.n3448 9.3005
R18265 VDD.n3447 VDD.n3399 9.3005
R18266 VDD.n3446 VDD.n3445 9.3005
R18267 VDD.n3444 VDD.n3443 9.3005
R18268 VDD.n3441 VDD.n3402 9.3005
R18269 VDD.n3440 VDD.n3439 9.3005
R18270 VDD.n3438 VDD.n3404 9.3005
R18271 VDD.n3437 VDD.n3436 9.3005
R18272 VDD.n3434 VDD.n3405 9.3005
R18273 VDD.n3433 VDD.n3432 9.3005
R18274 VDD.n3431 VDD.n3408 9.3005
R18275 VDD.n3430 VDD.n3429 9.3005
R18276 VDD.n3427 VDD.n3410 9.3005
R18277 VDD.n3425 VDD.n3424 9.3005
R18278 VDD.n3423 VDD.n3411 9.3005
R18279 VDD.n3422 VDD.n3421 9.3005
R18280 VDD.n3420 VDD.n3412 9.3005
R18281 VDD.n3418 VDD.n3417 9.3005
R18282 VDD.n3416 VDD.n3290 9.3005
R18283 VDD.n3470 VDD.n3289 9.3005
R18284 VDD.n3472 VDD.n3471 9.3005
R18285 VDD.n3473 VDD.n3288 9.3005
R18286 VDD.n3475 VDD.n3474 9.3005
R18287 VDD.n3478 VDD.n3285 9.3005
R18288 VDD.n3480 VDD.n3479 9.3005
R18289 VDD.n3482 VDD.n3481 9.3005
R18290 VDD.n3483 VDD.n3282 9.3005
R18291 VDD.n3484 VDD.n3279 9.3005
R18292 VDD.n3487 VDD.n3486 9.3005
R18293 VDD.n3489 VDD.n3488 9.3005
R18294 VDD.n3491 VDD.n3275 9.3005
R18295 VDD.n3494 VDD.n3493 9.3005
R18296 VDD.n3496 VDD.n3495 9.3005
R18297 VDD.n3497 VDD.n3271 9.3005
R18298 VDD.n3500 VDD.n3499 9.3005
R18299 VDD.n3501 VDD.n3270 9.3005
R18300 VDD.n3503 VDD.n3502 9.3005
R18301 VDD.n3504 VDD.n3266 9.3005
R18302 VDD.n3506 VDD.n3505 9.3005
R18303 VDD.n3507 VDD.n3265 9.3005
R18304 VDD.n3509 VDD.n3508 9.3005
R18305 VDD.n3511 VDD.n3263 9.3005
R18306 VDD.n3514 VDD.n3513 9.3005
R18307 VDD.n3516 VDD.n3515 9.3005
R18308 VDD.n3517 VDD.n3261 9.3005
R18309 VDD.n3518 VDD.n3259 9.3005
R18310 VDD.n3520 VDD.n3519 9.3005
R18311 VDD.n3521 VDD.n3258 9.3005
R18312 VDD.n3523 VDD.n3522 9.3005
R18313 VDD.n3526 VDD.n3256 9.3005
R18314 VDD.n3530 VDD.n3529 9.3005
R18315 VDD.n3531 VDD.n3255 9.3005
R18316 VDD.n3533 VDD.n3532 9.3005
R18317 VDD.n3534 VDD.n3254 9.3005
R18318 VDD.n3536 VDD.n3535 9.3005
R18319 VDD.n3538 VDD.n3537 9.3005
R18320 VDD.n3540 VDD.n3250 9.3005
R18321 VDD.n3542 VDD.n3541 9.3005
R18322 VDD.n3543 VDD.n3249 9.3005
R18323 VDD.n3545 VDD.n3544 9.3005
R18324 VDD.n3546 VDD.n3246 9.3005
R18325 VDD.n3547 VDD.n3244 9.3005
R18326 VDD.n3549 VDD.n3548 9.3005
R18327 VDD.n3551 VDD.n3550 9.3005
R18328 VDD.n3552 VDD.n3240 9.3005
R18329 VDD.n3554 VDD.n3553 9.3005
R18330 VDD.n3555 VDD.n3239 9.3005
R18331 VDD.n3557 VDD.n3556 9.3005
R18332 VDD.n3558 VDD.n3236 9.3005
R18333 VDD.n3559 VDD.n3235 9.3005
R18334 VDD.n3562 VDD.n3561 9.3005
R18335 VDD.n3564 VDD.n3563 9.3005
R18336 VDD.n3565 VDD.n3230 9.3005
R18337 VDD.n3567 VDD.n3566 9.3005
R18338 VDD.n3568 VDD.n3229 9.3005
R18339 VDD.n3633 VDD.n3632 9.3005
R18340 VDD.n3631 VDD.n3228 9.3005
R18341 VDD.n3630 VDD.n3629 9.3005
R18342 VDD.n3628 VDD.n3569 9.3005
R18343 VDD.n3627 VDD.n3626 9.3005
R18344 VDD.n3625 VDD.n3571 9.3005
R18345 VDD.n3624 VDD.n3623 9.3005
R18346 VDD.n3622 VDD.n3572 9.3005
R18347 VDD.n3621 VDD.n3619 9.3005
R18348 VDD.n3618 VDD.n3575 9.3005
R18349 VDD.n3617 VDD.n3616 9.3005
R18350 VDD.n3615 VDD.n3576 9.3005
R18351 VDD.n3613 VDD.n3612 9.3005
R18352 VDD.n3611 VDD.n3579 9.3005
R18353 VDD.n3610 VDD.n3609 9.3005
R18354 VDD.n3608 VDD.n3580 9.3005
R18355 VDD.n3607 VDD.n3606 9.3005
R18356 VDD.n3605 VDD.n3581 9.3005
R18357 VDD.n3604 VDD.n3603 9.3005
R18358 VDD.n3602 VDD.n3582 9.3005
R18359 VDD.n3601 VDD.n3600 9.3005
R18360 VDD.n3599 VDD.n3584 9.3005
R18361 VDD.n3598 VDD.n3597 9.3005
R18362 VDD.n3595 VDD.n3586 9.3005
R18363 VDD.n3594 VDD.n3592 9.3005
R18364 VDD.n3591 VDD.n3588 9.3005
R18365 VDD.n3590 VDD.n3589 9.3005
R18366 VDD.n3227 VDD.n3224 9.3005
R18367 VDD.n3637 VDD.n3636 9.3005
R18368 VDD.n3638 VDD.n3223 9.3005
R18369 VDD.n3640 VDD.n3639 9.3005
R18370 VDD.n3641 VDD.n3222 9.3005
R18371 VDD.n3642 VDD.n3221 9.3005
R18372 VDD.n3643 VDD.n3220 9.3005
R18373 VDD.n3647 VDD.n3646 9.3005
R18374 VDD.n3648 VDD.n3219 9.3005
R18375 VDD.n3650 VDD.n3649 9.3005
R18376 VDD.n3651 VDD.n3218 9.3005
R18377 VDD.n3652 VDD.n3216 9.3005
R18378 VDD.n3653 VDD.n3215 9.3005
R18379 VDD.n3654 VDD.n3213 9.3005
R18380 VDD.n3655 VDD.n3211 9.3005
R18381 VDD.n3658 VDD.n3657 9.3005
R18382 VDD.n3659 VDD.n3210 9.3005
R18383 VDD.n3661 VDD.n3660 9.3005
R18384 VDD.n3662 VDD.n3208 9.3005
R18385 VDD.n3663 VDD.n3207 9.3005
R18386 VDD.n3665 VDD.n3664 9.3005
R18387 VDD.n3667 VDD.n3666 9.3005
R18388 VDD.n3668 VDD.n3204 9.3005
R18389 VDD.n3673 VDD.n3672 9.3005
R18390 VDD.n3674 VDD.n3203 9.3005
R18391 VDD.n3676 VDD.n3675 9.3005
R18392 VDD.n3677 VDD.n3202 9.3005
R18393 VDD.n3681 VDD.n3680 9.3005
R18394 VDD.n3682 VDD.n3201 9.3005
R18395 VDD.n3753 VDD.n3752 9.3005
R18396 VDD.n3751 VDD.n3200 9.3005
R18397 VDD.n3750 VDD.n3749 9.3005
R18398 VDD.n3746 VDD.n3683 9.3005
R18399 VDD.n3744 VDD.n3743 9.3005
R18400 VDD.n3742 VDD.n3685 9.3005
R18401 VDD.n3741 VDD.n3740 9.3005
R18402 VDD.n3739 VDD.n3686 9.3005
R18403 VDD.n3738 VDD.n3737 9.3005
R18404 VDD.n3736 VDD.n3688 9.3005
R18405 VDD.n3735 VDD.n3734 9.3005
R18406 VDD.n3732 VDD.n3689 9.3005
R18407 VDD.n3731 VDD.n3730 9.3005
R18408 VDD.n3729 VDD.n3692 9.3005
R18409 VDD.n3728 VDD.n3727 9.3005
R18410 VDD.n3726 VDD.n3693 9.3005
R18411 VDD.n3725 VDD.n3724 9.3005
R18412 VDD.n3723 VDD.n3722 9.3005
R18413 VDD.n3720 VDD.n3696 9.3005
R18414 VDD.n3719 VDD.n3718 9.3005
R18415 VDD.n3717 VDD.n3716 9.3005
R18416 VDD.n3715 VDD.n3699 9.3005
R18417 VDD.n3714 VDD.n3713 9.3005
R18418 VDD.n3712 VDD.n3700 9.3005
R18419 VDD.n3711 VDD.n3710 9.3005
R18420 VDD.n3709 VDD.n3702 9.3005
R18421 VDD.n3707 VDD.n3706 9.3005
R18422 VDD.n3705 VDD.n3199 9.3005
R18423 VDD.n3756 VDD.n3198 9.3005
R18424 VDD.n3758 VDD.n3757 9.3005
R18425 VDD.n3759 VDD.n3197 9.3005
R18426 VDD.n3761 VDD.n3760 9.3005
R18427 VDD.n3763 VDD.n3196 9.3005
R18428 VDD.n3765 VDD.n3764 9.3005
R18429 VDD.n3767 VDD.n3766 9.3005
R18430 VDD.n3769 VDD.n3194 9.3005
R18431 VDD.n3771 VDD.n3770 9.3005
R18432 VDD.n3773 VDD.n3772 9.3005
R18433 VDD.n3774 VDD.n3191 9.3005
R18434 VDD.n3777 VDD.n3776 9.3005
R18435 VDD.n3778 VDD.n3190 9.3005
R18436 VDD.n3780 VDD.n3779 9.3005
R18437 VDD.n3783 VDD.n3188 9.3005
R18438 VDD.n3785 VDD.n3784 9.3005
R18439 VDD.n3786 VDD.n3187 9.3005
R18440 VDD.n3788 VDD.n3787 9.3005
R18441 VDD.n3789 VDD.n3186 9.3005
R18442 VDD.n3793 VDD.n3792 9.3005
R18443 VDD.n3794 VDD.n3184 9.3005
R18444 VDD.n3796 VDD.n3795 9.3005
R18445 VDD.n3797 VDD.n3183 9.3005
R18446 VDD.n3799 VDD.n3798 9.3005
R18447 VDD.n3801 VDD.n3800 9.3005
R18448 VDD.n3804 VDD.n3180 9.3005
R18449 VDD.n3806 VDD.n3805 9.3005
R18450 VDD.n3807 VDD.n3179 9.3005
R18451 VDD.n3864 VDD.n3808 9.3005
R18452 VDD.n3863 VDD.n3862 9.3005
R18453 VDD.n3861 VDD.n3860 9.3005
R18454 VDD.n3859 VDD.n3811 9.3005
R18455 VDD.n3858 VDD.n3857 9.3005
R18456 VDD.n3856 VDD.n3812 9.3005
R18457 VDD.n3855 VDD.n3854 9.3005
R18458 VDD.n3853 VDD.n3813 9.3005
R18459 VDD.n3850 VDD.n3849 9.3005
R18460 VDD.n3848 VDD.n3817 9.3005
R18461 VDD.n3847 VDD.n3846 9.3005
R18462 VDD.n3845 VDD.n3818 9.3005
R18463 VDD.n3843 VDD.n3842 9.3005
R18464 VDD.n3841 VDD.n3822 9.3005
R18465 VDD.n3840 VDD.n3839 9.3005
R18466 VDD.n3838 VDD.n3823 9.3005
R18467 VDD.n3837 VDD.n3836 9.3005
R18468 VDD.n3835 VDD.n3827 9.3005
R18469 VDD.n3834 VDD.n3833 9.3005
R18470 VDD.n3832 VDD.n3828 9.3005
R18471 VDD.n3829 VDD.n3094 9.3005
R18472 VDD.n3888 VDD.n3887 9.3005
R18473 VDD.n3885 VDD.n3884 9.3005
R18474 VDD.n3877 VDD.n3098 9.3005
R18475 VDD.n3876 VDD.n3875 9.3005
R18476 VDD.n3874 VDD.n3100 9.3005
R18477 VDD.n3872 VDD.n3871 9.3005
R18478 VDD.n3870 VDD.n3869 9.3005
R18479 VDD.n3867 VDD.n3105 9.3005
R18480 VDD.n3177 VDD.n3176 9.3005
R18481 VDD.n3175 VDD.n3106 9.3005
R18482 VDD.n3174 VDD.n3173 9.3005
R18483 VDD.n3172 VDD.n3107 9.3005
R18484 VDD.n3169 VDD.n3168 9.3005
R18485 VDD.n3166 VDD.n3165 9.3005
R18486 VDD.n3163 VDD.n3118 9.3005
R18487 VDD.n3161 VDD.n3160 9.3005
R18488 VDD.n3159 VDD.n3119 9.3005
R18489 VDD.n3158 VDD.n3157 9.3005
R18490 VDD.n3156 VDD.n3120 9.3005
R18491 VDD.n3155 VDD.n3154 9.3005
R18492 VDD.n3153 VDD.n3152 9.3005
R18493 VDD.n3151 VDD.n3124 9.3005
R18494 VDD.n3150 VDD.n3127 9.3005
R18495 VDD.n3149 VDD.n3148 9.3005
R18496 VDD.n3147 VDD.n3129 9.3005
R18497 VDD.n3146 VDD.n3145 9.3005
R18498 VDD.n3144 VDD.n3130 9.3005
R18499 VDD.n3143 VDD.n3142 9.3005
R18500 VDD.n2588 VDD.n2587 9.3005
R18501 VDD.n2589 VDD.n2577 9.3005
R18502 VDD.n2591 VDD.n2590 9.3005
R18503 VDD.n2593 VDD.n2568 9.3005
R18504 VDD.n2567 VDD.n2495 9.3005
R18505 VDD.n2566 VDD.n2565 9.3005
R18506 VDD.n2563 VDD.n2496 9.3005
R18507 VDD.n2561 VDD.n2560 9.3005
R18508 VDD.n2559 VDD.n2497 9.3005
R18509 VDD.n2558 VDD.n2557 9.3005
R18510 VDD.n2555 VDD.n2498 9.3005
R18511 VDD.n2554 VDD.n2553 9.3005
R18512 VDD.n2552 VDD.n2551 9.3005
R18513 VDD.n2549 VDD.n2503 9.3005
R18514 VDD.n2548 VDD.n2547 9.3005
R18515 VDD.n2546 VDD.n2545 9.3005
R18516 VDD.n2543 VDD.n2505 9.3005
R18517 VDD.n2542 VDD.n2541 9.3005
R18518 VDD.n2540 VDD.n2507 9.3005
R18519 VDD.n2539 VDD.n2538 9.3005
R18520 VDD.n2535 VDD.n2508 9.3005
R18521 VDD.n2534 VDD.n2533 9.3005
R18522 VDD.n2532 VDD.n2531 9.3005
R18523 VDD.n2530 VDD.n2512 9.3005
R18524 VDD.n2529 VDD.n2528 9.3005
R18525 VDD.n2527 VDD.n2514 9.3005
R18526 VDD.n2526 VDD.n2525 9.3005
R18527 VDD.n2523 VDD.n2516 9.3005
R18528 VDD.n2521 VDD.n2520 9.3005
R18529 VDD.n2519 VDD.n2517 9.3005
R18530 VDD.n2518 VDD.n2494 9.3005
R18531 VDD.n2596 VDD.n2493 9.3005
R18532 VDD.n2599 VDD.n2598 9.3005
R18533 VDD.n2601 VDD.n2600 9.3005
R18534 VDD.n2602 VDD.n2490 9.3005
R18535 VDD.n2606 VDD.n2605 9.3005
R18536 VDD.n2607 VDD.n2489 9.3005
R18537 VDD.n2609 VDD.n2608 9.3005
R18538 VDD.n2611 VDD.n2488 9.3005
R18539 VDD.n2617 VDD.n2616 9.3005
R18540 VDD.n2618 VDD.n2487 9.3005
R18541 VDD.n2620 VDD.n2619 9.3005
R18542 VDD.n2622 VDD.n2486 9.3005
R18543 VDD.n2624 VDD.n2623 9.3005
R18544 VDD.n2625 VDD.n2485 9.3005
R18545 VDD.n2627 VDD.n2626 9.3005
R18546 VDD.n2630 VDD.n2484 9.3005
R18547 VDD.n2632 VDD.n2631 9.3005
R18548 VDD.n2633 VDD.n2482 9.3005
R18549 VDD.n2635 VDD.n2634 9.3005
R18550 VDD.n2636 VDD.n2481 9.3005
R18551 VDD.n2638 VDD.n2637 9.3005
R18552 VDD.n2640 VDD.n2639 9.3005
R18553 VDD.n2642 VDD.n2477 9.3005
R18554 VDD.n2645 VDD.n2644 9.3005
R18555 VDD.n2646 VDD.n2476 9.3005
R18556 VDD.n2648 VDD.n2647 9.3005
R18557 VDD.n2649 VDD.n2475 9.3005
R18558 VDD.n2651 VDD.n2650 9.3005
R18559 VDD.n2724 VDD.n2723 9.3005
R18560 VDD.n2722 VDD.n2474 9.3005
R18561 VDD.n2721 VDD.n2720 9.3005
R18562 VDD.n2719 VDD.n2652 9.3005
R18563 VDD.n2718 VDD.n2717 9.3005
R18564 VDD.n2716 VDD.n2653 9.3005
R18565 VDD.n2715 VDD.n2714 9.3005
R18566 VDD.n2713 VDD.n2654 9.3005
R18567 VDD.n2712 VDD.n2656 9.3005
R18568 VDD.n2711 VDD.n2710 9.3005
R18569 VDD.n2709 VDD.n2658 9.3005
R18570 VDD.n2708 VDD.n2707 9.3005
R18571 VDD.n2705 VDD.n2659 9.3005
R18572 VDD.n2703 VDD.n2702 9.3005
R18573 VDD.n2701 VDD.n2663 9.3005
R18574 VDD.n2700 VDD.n2699 9.3005
R18575 VDD.n2698 VDD.n2664 9.3005
R18576 VDD.n2697 VDD.n2696 9.3005
R18577 VDD.n2695 VDD.n2694 9.3005
R18578 VDD.n2692 VDD.n2666 9.3005
R18579 VDD.n2691 VDD.n2690 9.3005
R18580 VDD.n2689 VDD.n2688 9.3005
R18581 VDD.n2686 VDD.n2670 9.3005
R18582 VDD.n2685 VDD.n2684 9.3005
R18583 VDD.n2683 VDD.n2672 9.3005
R18584 VDD.n2682 VDD.n2681 9.3005
R18585 VDD.n2679 VDD.n2673 9.3005
R18586 VDD.n2677 VDD.n2676 9.3005
R18587 VDD.n2728 VDD.n2469 9.3005
R18588 VDD.n2730 VDD.n2729 9.3005
R18589 VDD.n2731 VDD.n2468 9.3005
R18590 VDD.n2733 VDD.n2732 9.3005
R18591 VDD.n2734 VDD.n2467 9.3005
R18592 VDD.n2735 VDD.n2465 9.3005
R18593 VDD.n2737 VDD.n2736 9.3005
R18594 VDD.n2738 VDD.n2464 9.3005
R18595 VDD.n2740 VDD.n2739 9.3005
R18596 VDD.n2741 VDD.n2461 9.3005
R18597 VDD.n2743 VDD.n2742 9.3005
R18598 VDD.n2745 VDD.n2744 9.3005
R18599 VDD.n2746 VDD.n2458 9.3005
R18600 VDD.n2747 VDD.n2457 9.3005
R18601 VDD.n2749 VDD.n2748 9.3005
R18602 VDD.n2750 VDD.n2456 9.3005
R18603 VDD.n2752 VDD.n2751 9.3005
R18604 VDD.n2754 VDD.n2453 9.3005
R18605 VDD.n2755 VDD.n2452 9.3005
R18606 VDD.n2756 VDD.n2451 9.3005
R18607 VDD.n2758 VDD.n2757 9.3005
R18608 VDD.n2760 VDD.n2759 9.3005
R18609 VDD.n2763 VDD.n2449 9.3005
R18610 VDD.n2767 VDD.n2766 9.3005
R18611 VDD.n2769 VDD.n2768 9.3005
R18612 VDD.n2770 VDD.n2447 9.3005
R18613 VDD.n2771 VDD.n2446 9.3005
R18614 VDD.n2773 VDD.n2772 9.3005
R18615 VDD.n2774 VDD.n2445 9.3005
R18616 VDD.n2776 VDD.n2775 9.3005
R18617 VDD.n2777 VDD.n2444 9.3005
R18618 VDD.n2778 VDD.n2442 9.3005
R18619 VDD.n2779 VDD.n2440 9.3005
R18620 VDD.n2783 VDD.n2782 9.3005
R18621 VDD.n2784 VDD.n2439 9.3005
R18622 VDD.n2786 VDD.n2785 9.3005
R18623 VDD.n2787 VDD.n2438 9.3005
R18624 VDD.n2790 VDD.n2789 9.3005
R18625 VDD.n2792 VDD.n2791 9.3005
R18626 VDD.n2793 VDD.n2436 9.3005
R18627 VDD.n2794 VDD.n2435 9.3005
R18628 VDD.n2795 VDD.n2434 9.3005
R18629 VDD.n2796 VDD.n2432 9.3005
R18630 VDD.n2799 VDD.n2798 9.3005
R18631 VDD.n2801 VDD.n2800 9.3005
R18632 VDD.n2802 VDD.n2429 9.3005
R18633 VDD.n2803 VDD.n2428 9.3005
R18634 VDD.n2807 VDD.n2806 9.3005
R18635 VDD.n2808 VDD.n2427 9.3005
R18636 VDD.n2810 VDD.n2809 9.3005
R18637 VDD.n2812 VDD.n2423 9.3005
R18638 VDD.n2817 VDD.n2816 9.3005
R18639 VDD.n2818 VDD.n2422 9.3005
R18640 VDD.n2820 VDD.n2819 9.3005
R18641 VDD.n2821 VDD.n2419 9.3005
R18642 VDD.n2823 VDD.n2822 9.3005
R18643 VDD.n2893 VDD.n2892 9.3005
R18644 VDD.n2891 VDD.n2418 9.3005
R18645 VDD.n2890 VDD.n2889 9.3005
R18646 VDD.n2887 VDD.n2824 9.3005
R18647 VDD.n2885 VDD.n2884 9.3005
R18648 VDD.n2883 VDD.n2827 9.3005
R18649 VDD.n2882 VDD.n2881 9.3005
R18650 VDD.n2880 VDD.n2828 9.3005
R18651 VDD.n2878 VDD.n2876 9.3005
R18652 VDD.n2875 VDD.n2829 9.3005
R18653 VDD.n2874 VDD.n2873 9.3005
R18654 VDD.n2872 VDD.n2830 9.3005
R18655 VDD.n2871 VDD.n2870 9.3005
R18656 VDD.n2869 VDD.n2832 9.3005
R18657 VDD.n2868 VDD.n2867 9.3005
R18658 VDD.n2866 VDD.n2833 9.3005
R18659 VDD.n2865 VDD.n2864 9.3005
R18660 VDD.n2863 VDD.n2835 9.3005
R18661 VDD.n2862 VDD.n2861 9.3005
R18662 VDD.n2860 VDD.n2836 9.3005
R18663 VDD.n2859 VDD.n2858 9.3005
R18664 VDD.n2857 VDD.n2856 9.3005
R18665 VDD.n2854 VDD.n2839 9.3005
R18666 VDD.n2852 VDD.n2851 9.3005
R18667 VDD.n2849 VDD.n2848 9.3005
R18668 VDD.n2897 VDD.n2414 9.3005
R18669 VDD.n2900 VDD.n2410 9.3005
R18670 VDD.n2902 VDD.n2901 9.3005
R18671 VDD.n2904 VDD.n2903 9.3005
R18672 VDD.n2906 VDD.n2406 9.3005
R18673 VDD.n2911 VDD.n2910 9.3005
R18674 VDD.n2913 VDD.n2912 9.3005
R18675 VDD.n2914 VDD.n2403 9.3005
R18676 VDD.n2917 VDD.n2916 9.3005
R18677 VDD.n2919 VDD.n2918 9.3005
R18678 VDD.n2920 VDD.n2400 9.3005
R18679 VDD.n2921 VDD.n2399 9.3005
R18680 VDD.n2924 VDD.n2923 9.3005
R18681 VDD.n2925 VDD.n2398 9.3005
R18682 VDD.n2927 VDD.n2926 9.3005
R18683 VDD.n2928 VDD.n2397 9.3005
R18684 VDD.n2929 VDD.n2394 9.3005
R18685 VDD.n2932 VDD.n2931 9.3005
R18686 VDD.n2933 VDD.n2393 9.3005
R18687 VDD.n2935 VDD.n2934 9.3005
R18688 VDD.n2936 VDD.n2391 9.3005
R18689 VDD.n2937 VDD.n2390 9.3005
R18690 VDD.n2939 VDD.n2938 9.3005
R18691 VDD.n2940 VDD.n2389 9.3005
R18692 VDD.n2942 VDD.n2941 9.3005
R18693 VDD.n2943 VDD.n2387 9.3005
R18694 VDD.n2944 VDD.n2385 9.3005
R18695 VDD.n2946 VDD.n2945 9.3005
R18696 VDD.n2947 VDD.n2384 9.3005
R18697 VDD.n2949 VDD.n2948 9.3005
R18698 VDD.n2950 VDD.n2383 9.3005
R18699 VDD.n2954 VDD.n2953 9.3005
R18700 VDD.n2955 VDD.n2382 9.3005
R18701 VDD.n2957 VDD.n2956 9.3005
R18702 VDD.n2958 VDD.n2381 9.3005
R18703 VDD.n2960 VDD.n2959 9.3005
R18704 VDD.n2961 VDD.n2380 9.3005
R18705 VDD.n2963 VDD.n2962 9.3005
R18706 VDD.n2966 VDD.n2378 9.3005
R18707 VDD.n2972 VDD.n2971 9.3005
R18708 VDD.n2973 VDD.n2377 9.3005
R18709 VDD.n2975 VDD.n2974 9.3005
R18710 VDD.n2976 VDD.n2376 9.3005
R18711 VDD.n2978 VDD.n2977 9.3005
R18712 VDD.n2979 VDD.n2375 9.3005
R18713 VDD.n2981 VDD.n2980 9.3005
R18714 VDD.n2984 VDD.n2371 9.3005
R18715 VDD.n2987 VDD.n2986 9.3005
R18716 VDD.n2989 VDD.n2988 9.3005
R18717 VDD.n2990 VDD.n2368 9.3005
R18718 VDD.n2992 VDD.n2991 9.3005
R18719 VDD.n2993 VDD.n2367 9.3005
R18720 VDD.n2995 VDD.n2994 9.3005
R18721 VDD.n2997 VDD.n2363 9.3005
R18722 VDD.n3001 VDD.n3000 9.3005
R18723 VDD.n3002 VDD.n2360 9.3005
R18724 VDD.n3063 VDD.n3062 9.3005
R18725 VDD.n3061 VDD.n3060 9.3005
R18726 VDD.n3059 VDD.n3003 9.3005
R18727 VDD.n3057 VDD.n3056 9.3005
R18728 VDD.n3055 VDD.n3054 9.3005
R18729 VDD.n3009 VDD.n3007 9.3005
R18730 VDD.n3017 VDD.n3012 9.3005
R18731 VDD.n3018 VDD.n3013 9.3005
R18732 VDD.n3048 VDD.n3047 9.3005
R18733 VDD.n3046 VDD.n3045 9.3005
R18734 VDD.n3044 VDD.n3019 9.3005
R18735 VDD.n3040 VDD.n3039 9.3005
R18736 VDD.n3038 VDD.n3020 9.3005
R18737 VDD.n3037 VDD.n3036 9.3005
R18738 VDD.n3035 VDD.n3021 9.3005
R18739 VDD.n3034 VDD.n3024 9.3005
R18740 VDD.n3033 VDD.n3026 9.3005
R18741 VDD.n3032 VDD.n3031 9.3005
R18742 VDD.n3030 VDD.n3029 9.3005
R18743 VDD.n3028 VDD.n2278 9.3005
R18744 VDD.n3085 VDD.n3084 9.3005
R18745 VDD.n3083 VDD.n3082 9.3005
R18746 VDD.n3075 VDD.n2282 9.3005
R18747 VDD.n3074 VDD.n3073 9.3005
R18748 VDD.n3072 VDD.n2284 9.3005
R18749 VDD.n3071 VDD.n3070 9.3005
R18750 VDD.n3069 VDD.n3068 9.3005
R18751 VDD.n3066 VDD.n2287 9.3005
R18752 VDD.n2359 VDD.n2358 9.3005
R18753 VDD.n2357 VDD.n2356 9.3005
R18754 VDD.n2355 VDD.n2290 9.3005
R18755 VDD.n2353 VDD.n2352 9.3005
R18756 VDD.n2351 VDD.n2350 9.3005
R18757 VDD.n2348 VDD.n2293 9.3005
R18758 VDD.n2345 VDD.n2344 9.3005
R18759 VDD.n2342 VDD.n2296 9.3005
R18760 VDD.n2341 VDD.n2340 9.3005
R18761 VDD.n2339 VDD.n2338 9.3005
R18762 VDD.n2337 VDD.n2301 9.3005
R18763 VDD.n2336 VDD.n2335 9.3005
R18764 VDD.n2334 VDD.n2333 9.3005
R18765 VDD.n2332 VDD.n2304 9.3005
R18766 VDD.n2331 VDD.n2330 9.3005
R18767 VDD.n2329 VDD.n2328 9.3005
R18768 VDD.n2327 VDD.n2307 9.3005
R18769 VDD.n2326 VDD.n2325 9.3005
R18770 VDD.n2324 VDD.n2312 9.3005
R18771 VDD.n2323 VDD.n2322 9.3005
R18772 VDD.n1704 VDD.n1703 9.3005
R18773 VDD.n1705 VDD.n1693 9.3005
R18774 VDD.n1707 VDD.n1706 9.3005
R18775 VDD.n1709 VDD.n1690 9.3005
R18776 VDD.n1712 VDD.n1711 9.3005
R18777 VDD.n1713 VDD.n1688 9.3005
R18778 VDD.n1715 VDD.n1714 9.3005
R18779 VDD.n1716 VDD.n1686 9.3005
R18780 VDD.n1718 VDD.n1717 9.3005
R18781 VDD.n1719 VDD.n1685 9.3005
R18782 VDD.n1721 VDD.n1720 9.3005
R18783 VDD.n1722 VDD.n1682 9.3005
R18784 VDD.n1723 VDD.n1680 9.3005
R18785 VDD.n1726 VDD.n1725 9.3005
R18786 VDD.n1728 VDD.n1727 9.3005
R18787 VDD.n1729 VDD.n1678 9.3005
R18788 VDD.n1730 VDD.n1677 9.3005
R18789 VDD.n1731 VDD.n1675 9.3005
R18790 VDD.n1732 VDD.n1674 9.3005
R18791 VDD.n1733 VDD.n1672 9.3005
R18792 VDD.n1735 VDD.n1734 9.3005
R18793 VDD.n1737 VDD.n1736 9.3005
R18794 VDD.n1738 VDD.n1669 9.3005
R18795 VDD.n1739 VDD.n1668 9.3005
R18796 VDD.n1740 VDD.n1665 9.3005
R18797 VDD.n1742 VDD.n1741 9.3005
R18798 VDD.n1744 VDD.n1743 9.3005
R18799 VDD.n1746 VDD.n1662 9.3005
R18800 VDD.n1748 VDD.n1747 9.3005
R18801 VDD.n1749 VDD.n1661 9.3005
R18802 VDD.n1751 VDD.n1750 9.3005
R18803 VDD.n1752 VDD.n1659 9.3005
R18804 VDD.n1754 VDD.n1753 9.3005
R18805 VDD.n1755 VDD.n1657 9.3005
R18806 VDD.n1757 VDD.n1756 9.3005
R18807 VDD.n1758 VDD.n1655 9.3005
R18808 VDD.n1761 VDD.n1760 9.3005
R18809 VDD.n1763 VDD.n1762 9.3005
R18810 VDD.n1764 VDD.n1652 9.3005
R18811 VDD.n1765 VDD.n1649 9.3005
R18812 VDD.n1768 VDD.n1648 9.3005
R18813 VDD.n1770 VDD.n1769 9.3005
R18814 VDD.n1771 VDD.n1647 9.3005
R18815 VDD.n1773 VDD.n1772 9.3005
R18816 VDD.n1775 VDD.n1774 9.3005
R18817 VDD.n1777 VDD.n1643 9.3005
R18818 VDD.n1779 VDD.n1778 9.3005
R18819 VDD.n1780 VDD.n1642 9.3005
R18820 VDD.n1782 VDD.n1781 9.3005
R18821 VDD.n1783 VDD.n1640 9.3005
R18822 VDD.n1784 VDD.n1639 9.3005
R18823 VDD.n1789 VDD.n1788 9.3005
R18824 VDD.n1790 VDD.n1638 9.3005
R18825 VDD.n1792 VDD.n1791 9.3005
R18826 VDD.n1794 VDD.n1636 9.3005
R18827 VDD.n1797 VDD.n1796 9.3005
R18828 VDD.n1799 VDD.n1798 9.3005
R18829 VDD.n1801 VDD.n1632 9.3005
R18830 VDD.n1803 VDD.n1802 9.3005
R18831 VDD.n1804 VDD.n1630 9.3005
R18832 VDD.n1806 VDD.n1805 9.3005
R18833 VDD.n1807 VDD.n1629 9.3005
R18834 VDD.n1808 VDD.n1628 9.3005
R18835 VDD.n1809 VDD.n1626 9.3005
R18836 VDD.n1813 VDD.n1812 9.3005
R18837 VDD.n1814 VDD.n1625 9.3005
R18838 VDD.n1816 VDD.n1815 9.3005
R18839 VDD.n1817 VDD.n1623 9.3005
R18840 VDD.n1818 VDD.n1620 9.3005
R18841 VDD.n1821 VDD.n1820 9.3005
R18842 VDD.n1823 VDD.n1822 9.3005
R18843 VDD.n1825 VDD.n1617 9.3005
R18844 VDD.n1829 VDD.n1828 9.3005
R18845 VDD.n1831 VDD.n1830 9.3005
R18846 VDD.n1832 VDD.n1612 9.3005
R18847 VDD.n1835 VDD.n1834 9.3005
R18848 VDD.n1836 VDD.n1611 9.3005
R18849 VDD.n1838 VDD.n1837 9.3005
R18850 VDD.n1840 VDD.n1607 9.3005
R18851 VDD.n1843 VDD.n1842 9.3005
R18852 VDD.n1845 VDD.n1844 9.3005
R18853 VDD.n1847 VDD.n1604 9.3005
R18854 VDD.n1850 VDD.n1849 9.3005
R18855 VDD.n1852 VDD.n1851 9.3005
R18856 VDD.n1853 VDD.n1601 9.3005
R18857 VDD.n1854 VDD.n1599 9.3005
R18858 VDD.n1856 VDD.n1855 9.3005
R18859 VDD.n1857 VDD.n1596 9.3005
R18860 VDD.n1859 VDD.n1858 9.3005
R18861 VDD.n1860 VDD.n1595 9.3005
R18862 VDD.n1862 VDD.n1861 9.3005
R18863 VDD.n1863 VDD.n1594 9.3005
R18864 VDD.n1865 VDD.n1864 9.3005
R18865 VDD.n1867 VDD.n1592 9.3005
R18866 VDD.n1874 VDD.n1590 9.3005
R18867 VDD.n1876 VDD.n1875 9.3005
R18868 VDD.n1878 VDD.n1589 9.3005
R18869 VDD.n1880 VDD.n1879 9.3005
R18870 VDD.n1881 VDD.n1588 9.3005
R18871 VDD.n1883 VDD.n1882 9.3005
R18872 VDD.n1884 VDD.n1587 9.3005
R18873 VDD.n1888 VDD.n1887 9.3005
R18874 VDD.n1890 VDD.n1582 9.3005
R18875 VDD.n1892 VDD.n1891 9.3005
R18876 VDD.n1894 VDD.n1580 9.3005
R18877 VDD.n1896 VDD.n1895 9.3005
R18878 VDD.n1898 VDD.n1897 9.3005
R18879 VDD.n1900 VDD.n1577 9.3005
R18880 VDD.n1903 VDD.n1902 9.3005
R18881 VDD.n1904 VDD.n1576 9.3005
R18882 VDD.n1906 VDD.n1905 9.3005
R18883 VDD.n1913 VDD.n1912 9.3005
R18884 VDD.n1915 VDD.n1914 9.3005
R18885 VDD.n1917 VDD.n1573 9.3005
R18886 VDD.n1919 VDD.n1918 9.3005
R18887 VDD.n1921 VDD.n1920 9.3005
R18888 VDD.n1922 VDD.n1571 9.3005
R18889 VDD.n1925 VDD.n1924 9.3005
R18890 VDD.n1926 VDD.n1570 9.3005
R18891 VDD.n1928 VDD.n1927 9.3005
R18892 VDD.n1929 VDD.n1568 9.3005
R18893 VDD.n1932 VDD.n1931 9.3005
R18894 VDD.n1933 VDD.n1567 9.3005
R18895 VDD.n1935 VDD.n1934 9.3005
R18896 VDD.n1936 VDD.n1566 9.3005
R18897 VDD.n1938 VDD.n1937 9.3005
R18898 VDD.n1939 VDD.n1565 9.3005
R18899 VDD.n1941 VDD.n1940 9.3005
R18900 VDD.n1943 VDD.n1563 9.3005
R18901 VDD.n1945 VDD.n1944 9.3005
R18902 VDD.n1946 VDD.n1562 9.3005
R18903 VDD.n1948 VDD.n1947 9.3005
R18904 VDD.n1950 VDD.n1561 9.3005
R18905 VDD.n1952 VDD.n1951 9.3005
R18906 VDD.n2026 VDD.n1953 9.3005
R18907 VDD.n2025 VDD.n2024 9.3005
R18908 VDD.n2023 VDD.n1955 9.3005
R18909 VDD.n2022 VDD.n2021 9.3005
R18910 VDD.n2020 VDD.n1956 9.3005
R18911 VDD.n2019 VDD.n2018 9.3005
R18912 VDD.n2017 VDD.n1957 9.3005
R18913 VDD.n2016 VDD.n2015 9.3005
R18914 VDD.n2013 VDD.n1959 9.3005
R18915 VDD.n2009 VDD.n1960 9.3005
R18916 VDD.n2008 VDD.n2007 9.3005
R18917 VDD.n2004 VDD.n1961 9.3005
R18918 VDD.n2003 VDD.n2002 9.3005
R18919 VDD.n2001 VDD.n1965 9.3005
R18920 VDD.n2000 VDD.n1999 9.3005
R18921 VDD.n1997 VDD.n1966 9.3005
R18922 VDD.n1995 VDD.n1994 9.3005
R18923 VDD.n1993 VDD.n1992 9.3005
R18924 VDD.n1989 VDD.n1969 9.3005
R18925 VDD.n1987 VDD.n1986 9.3005
R18926 VDD.n1985 VDD.n1971 9.3005
R18927 VDD.n1984 VDD.n1983 9.3005
R18928 VDD.n1980 VDD.n1972 9.3005
R18929 VDD.n1979 VDD.n1977 9.3005
R18930 VDD.n1976 VDD.n1975 9.3005
R18931 VDD.n1558 VDD.n1557 9.3005
R18932 VDD.n2031 VDD.n2030 9.3005
R18933 VDD.n2032 VDD.n1556 9.3005
R18934 VDD.n2034 VDD.n2033 9.3005
R18935 VDD.n2035 VDD.n1554 9.3005
R18936 VDD.n2038 VDD.n2037 9.3005
R18937 VDD.n2040 VDD.n2039 9.3005
R18938 VDD.n2041 VDD.n1551 9.3005
R18939 VDD.n2043 VDD.n2042 9.3005
R18940 VDD.n2044 VDD.n1550 9.3005
R18941 VDD.n2046 VDD.n2045 9.3005
R18942 VDD.n2047 VDD.n1549 9.3005
R18943 VDD.n2048 VDD.n1546 9.3005
R18944 VDD.n2050 VDD.n2049 9.3005
R18945 VDD.n2051 VDD.n1545 9.3005
R18946 VDD.n2053 VDD.n2052 9.3005
R18947 VDD.n2054 VDD.n1544 9.3005
R18948 VDD.n2055 VDD.n1543 9.3005
R18949 VDD.n2056 VDD.n1542 9.3005
R18950 VDD.n2059 VDD.n2058 9.3005
R18951 VDD.n2061 VDD.n2060 9.3005
R18952 VDD.n2063 VDD.n1539 9.3005
R18953 VDD.n2065 VDD.n2064 9.3005
R18954 VDD.n2068 VDD.n2067 9.3005
R18955 VDD.n2069 VDD.n1533 9.3005
R18956 VDD.n2071 VDD.n2070 9.3005
R18957 VDD.n2072 VDD.n1532 9.3005
R18958 VDD.n2074 VDD.n2073 9.3005
R18959 VDD.n2075 VDD.n1531 9.3005
R18960 VDD.n2077 VDD.n2076 9.3005
R18961 VDD.n2078 VDD.n1530 9.3005
R18962 VDD.n2080 VDD.n2079 9.3005
R18963 VDD.n2081 VDD.n1529 9.3005
R18964 VDD.n2087 VDD.n2086 9.3005
R18965 VDD.n2088 VDD.n1528 9.3005
R18966 VDD.n2090 VDD.n2089 9.3005
R18967 VDD.n2091 VDD.n1527 9.3005
R18968 VDD.n2093 VDD.n2092 9.3005
R18969 VDD.n2095 VDD.n2094 9.3005
R18970 VDD.n2097 VDD.n1525 9.3005
R18971 VDD.n2099 VDD.n2098 9.3005
R18972 VDD.n2100 VDD.n1524 9.3005
R18973 VDD.n2102 VDD.n2101 9.3005
R18974 VDD.n2104 VDD.n1522 9.3005
R18975 VDD.n2106 VDD.n2105 9.3005
R18976 VDD.n2107 VDD.n1521 9.3005
R18977 VDD.n2109 VDD.n2108 9.3005
R18978 VDD.n2110 VDD.n1520 9.3005
R18979 VDD.n2112 VDD.n2111 9.3005
R18980 VDD.n2113 VDD.n1519 9.3005
R18981 VDD.n2115 VDD.n2114 9.3005
R18982 VDD.n2116 VDD.n1518 9.3005
R18983 VDD.n2119 VDD.n2118 9.3005
R18984 VDD.n2120 VDD.n1517 9.3005
R18985 VDD.n2170 VDD.n2121 9.3005
R18986 VDD.n2169 VDD.n2168 9.3005
R18987 VDD.n2167 VDD.n2123 9.3005
R18988 VDD.n2166 VDD.n2165 9.3005
R18989 VDD.n2164 VDD.n2124 9.3005
R18990 VDD.n2163 VDD.n2125 9.3005
R18991 VDD.n2162 VDD.n2161 9.3005
R18992 VDD.n2160 VDD.n2127 9.3005
R18993 VDD.n2159 VDD.n2158 9.3005
R18994 VDD.n2157 VDD.n2128 9.3005
R18995 VDD.n2156 VDD.n2155 9.3005
R18996 VDD.n2154 VDD.n2153 9.3005
R18997 VDD.n2151 VDD.n2150 9.3005
R18998 VDD.n2149 VDD.n2133 9.3005
R18999 VDD.n2148 VDD.n2147 9.3005
R19000 VDD.n2146 VDD.n2134 9.3005
R19001 VDD.n2144 VDD.n2143 9.3005
R19002 VDD.n2142 VDD.n2141 9.3005
R19003 VDD.n1509 VDD.n1507 9.3005
R19004 VDD.n2269 VDD.n2268 9.3005
R19005 VDD.n2267 VDD.n2266 9.3005
R19006 VDD.n2259 VDD.n2258 9.3005
R19007 VDD.n2256 VDD.n1512 9.3005
R19008 VDD.n2254 VDD.n2253 9.3005
R19009 VDD.n2252 VDD.n2251 9.3005
R19010 VDD.n2249 VDD.n1516 9.3005
R19011 VDD.n2247 VDD.n2246 9.3005
R19012 VDD.n2245 VDD.n2174 9.3005
R19013 VDD.n2244 VDD.n2243 9.3005
R19014 VDD.n2242 VDD.n2175 9.3005
R19015 VDD.n2240 VDD.n2239 9.3005
R19016 VDD.n2238 VDD.n2176 9.3005
R19017 VDD.n2237 VDD.n2236 9.3005
R19018 VDD.n2235 VDD.n2177 9.3005
R19019 VDD.n2233 VDD.n2232 9.3005
R19020 VDD.n2231 VDD.n2182 9.3005
R19021 VDD.n2230 VDD.n2229 9.3005
R19022 VDD.n2228 VDD.n2183 9.3005
R19023 VDD.n2226 VDD.n2185 9.3005
R19024 VDD.n2225 VDD.n2224 9.3005
R19025 VDD.n2223 VDD.n2186 9.3005
R19026 VDD.n2222 VDD.n2221 9.3005
R19027 VDD.n2220 VDD.n2187 9.3005
R19028 VDD.n2219 VDD.n2218 9.3005
R19029 VDD.n2217 VDD.n2189 9.3005
R19030 VDD.n2216 VDD.n2215 9.3005
R19031 VDD.n2212 VDD.n2190 9.3005
R19032 VDD.n2211 VDD.n2193 9.3005
R19033 VDD.n2210 VDD.n2209 9.3005
R19034 VDD.n2208 VDD.n2196 9.3005
R19035 VDD.n2207 VDD.n2206 9.3005
R19036 VDD.n865 VDD.n864 9.3005
R19037 VDD.n867 VDD.n854 9.3005
R19038 VDD.n870 VDD.n869 9.3005
R19039 VDD.n872 VDD.n871 9.3005
R19040 VDD.n874 VDD.n850 9.3005
R19041 VDD.n877 VDD.n876 9.3005
R19042 VDD.n878 VDD.n849 9.3005
R19043 VDD.n950 VDD.n949 9.3005
R19044 VDD.n948 VDD.n947 9.3005
R19045 VDD.n945 VDD.n879 9.3005
R19046 VDD.n944 VDD.n943 9.3005
R19047 VDD.n942 VDD.n880 9.3005
R19048 VDD.n941 VDD.n940 9.3005
R19049 VDD.n937 VDD.n882 9.3005
R19050 VDD.n936 VDD.n935 9.3005
R19051 VDD.n934 VDD.n933 9.3005
R19052 VDD.n932 VDD.n884 9.3005
R19053 VDD.n930 VDD.n929 9.3005
R19054 VDD.n928 VDD.n885 9.3005
R19055 VDD.n927 VDD.n926 9.3005
R19056 VDD.n924 VDD.n886 9.3005
R19057 VDD.n922 VDD.n921 9.3005
R19058 VDD.n920 VDD.n919 9.3005
R19059 VDD.n918 VDD.n891 9.3005
R19060 VDD.n917 VDD.n916 9.3005
R19061 VDD.n915 VDD.n892 9.3005
R19062 VDD.n914 VDD.n913 9.3005
R19063 VDD.n911 VDD.n893 9.3005
R19064 VDD.n910 VDD.n909 9.3005
R19065 VDD.n908 VDD.n898 9.3005
R19066 VDD.n907 VDD.n906 9.3005
R19067 VDD.n905 VDD.n899 9.3005
R19068 VDD.n904 VDD.n903 9.3005
R19069 VDD.n902 VDD.n901 9.3005
R19070 VDD.n847 VDD.n845 9.3005
R19071 VDD.n954 VDD.n953 9.3005
R19072 VDD.n955 VDD.n844 9.3005
R19073 VDD.n957 VDD.n956 9.3005
R19074 VDD.n958 VDD.n842 9.3005
R19075 VDD.n959 VDD.n841 9.3005
R19076 VDD.n962 VDD.n961 9.3005
R19077 VDD.n963 VDD.n840 9.3005
R19078 VDD.n965 VDD.n964 9.3005
R19079 VDD.n966 VDD.n837 9.3005
R19080 VDD.n967 VDD.n836 9.3005
R19081 VDD.n974 VDD.n973 9.3005
R19082 VDD.n975 VDD.n835 9.3005
R19083 VDD.n977 VDD.n976 9.3005
R19084 VDD.n979 VDD.n832 9.3005
R19085 VDD.n982 VDD.n981 9.3005
R19086 VDD.n983 VDD.n831 9.3005
R19087 VDD.n985 VDD.n984 9.3005
R19088 VDD.n986 VDD.n830 9.3005
R19089 VDD.n987 VDD.n828 9.3005
R19090 VDD.n988 VDD.n827 9.3005
R19091 VDD.n992 VDD.n991 9.3005
R19092 VDD.n994 VDD.n993 9.3005
R19093 VDD.n995 VDD.n824 9.3005
R19094 VDD.n997 VDD.n996 9.3005
R19095 VDD.n999 VDD.n998 9.3005
R19096 VDD.n1000 VDD.n820 9.3005
R19097 VDD.n1002 VDD.n1001 9.3005
R19098 VDD.n1003 VDD.n819 9.3005
R19099 VDD.n1077 VDD.n1076 9.3005
R19100 VDD.n1075 VDD.n818 9.3005
R19101 VDD.n1074 VDD.n1073 9.3005
R19102 VDD.n1071 VDD.n1004 9.3005
R19103 VDD.n1070 VDD.n1069 9.3005
R19104 VDD.n1068 VDD.n1008 9.3005
R19105 VDD.n1067 VDD.n1066 9.3005
R19106 VDD.n1064 VDD.n1009 9.3005
R19107 VDD.n1063 VDD.n1062 9.3005
R19108 VDD.n1061 VDD.n1060 9.3005
R19109 VDD.n1058 VDD.n1011 9.3005
R19110 VDD.n1057 VDD.n1056 9.3005
R19111 VDD.n1055 VDD.n1013 9.3005
R19112 VDD.n1054 VDD.n1053 9.3005
R19113 VDD.n1050 VDD.n1014 9.3005
R19114 VDD.n1049 VDD.n1048 9.3005
R19115 VDD.n1047 VDD.n1015 9.3005
R19116 VDD.n1046 VDD.n1045 9.3005
R19117 VDD.n1044 VDD.n1016 9.3005
R19118 VDD.n1042 VDD.n1041 9.3005
R19119 VDD.n1040 VDD.n1020 9.3005
R19120 VDD.n1039 VDD.n1038 9.3005
R19121 VDD.n1036 VDD.n1021 9.3005
R19122 VDD.n1034 VDD.n1033 9.3005
R19123 VDD.n1032 VDD.n1023 9.3005
R19124 VDD.n1031 VDD.n1030 9.3005
R19125 VDD.n1029 VDD.n1025 9.3005
R19126 VDD.n1024 VDD.n817 9.3005
R19127 VDD.n1080 VDD.n816 9.3005
R19128 VDD.n1082 VDD.n1081 9.3005
R19129 VDD.n1083 VDD.n815 9.3005
R19130 VDD.n1085 VDD.n1084 9.3005
R19131 VDD.n1087 VDD.n812 9.3005
R19132 VDD.n1089 VDD.n1088 9.3005
R19133 VDD.n1091 VDD.n1090 9.3005
R19134 VDD.n1092 VDD.n809 9.3005
R19135 VDD.n1095 VDD.n1094 9.3005
R19136 VDD.n1097 VDD.n1096 9.3005
R19137 VDD.n1099 VDD.n806 9.3005
R19138 VDD.n1103 VDD.n1102 9.3005
R19139 VDD.n1104 VDD.n805 9.3005
R19140 VDD.n1106 VDD.n1105 9.3005
R19141 VDD.n1107 VDD.n803 9.3005
R19142 VDD.n1109 VDD.n1108 9.3005
R19143 VDD.n1110 VDD.n802 9.3005
R19144 VDD.n1112 VDD.n1111 9.3005
R19145 VDD.n1113 VDD.n799 9.3005
R19146 VDD.n1117 VDD.n1116 9.3005
R19147 VDD.n1118 VDD.n798 9.3005
R19148 VDD.n1120 VDD.n1119 9.3005
R19149 VDD.n1121 VDD.n797 9.3005
R19150 VDD.n1122 VDD.n796 9.3005
R19151 VDD.n1123 VDD.n794 9.3005
R19152 VDD.n1124 VDD.n792 9.3005
R19153 VDD.n1126 VDD.n1125 9.3005
R19154 VDD.n1127 VDD.n790 9.3005
R19155 VDD.n1198 VDD.n1197 9.3005
R19156 VDD.n1196 VDD.n791 9.3005
R19157 VDD.n1195 VDD.n1194 9.3005
R19158 VDD.n1193 VDD.n1128 9.3005
R19159 VDD.n1192 VDD.n1131 9.3005
R19160 VDD.n1191 VDD.n1132 9.3005
R19161 VDD.n1190 VDD.n1189 9.3005
R19162 VDD.n1188 VDD.n1133 9.3005
R19163 VDD.n1187 VDD.n1186 9.3005
R19164 VDD.n1185 VDD.n1134 9.3005
R19165 VDD.n1184 VDD.n1135 9.3005
R19166 VDD.n1183 VDD.n1182 9.3005
R19167 VDD.n1181 VDD.n1180 9.3005
R19168 VDD.n1179 VDD.n1139 9.3005
R19169 VDD.n1176 VDD.n1175 9.3005
R19170 VDD.n1174 VDD.n1140 9.3005
R19171 VDD.n1173 VDD.n1172 9.3005
R19172 VDD.n1171 VDD.n1141 9.3005
R19173 VDD.n1170 VDD.n1144 9.3005
R19174 VDD.n1169 VDD.n1168 9.3005
R19175 VDD.n1167 VDD.n1166 9.3005
R19176 VDD.n1164 VDD.n1146 9.3005
R19177 VDD.n1163 VDD.n1148 9.3005
R19178 VDD.n1161 VDD.n1160 9.3005
R19179 VDD.n1159 VDD.n1151 9.3005
R19180 VDD.n1158 VDD.n1157 9.3005
R19181 VDD.n1156 VDD.n1152 9.3005
R19182 VDD.n787 VDD.n786 9.3005
R19183 VDD.n1203 VDD.n1202 9.3005
R19184 VDD.n1204 VDD.n785 9.3005
R19185 VDD.n1206 VDD.n1205 9.3005
R19186 VDD.n1209 VDD.n783 9.3005
R19187 VDD.n1212 VDD.n1211 9.3005
R19188 VDD.n1213 VDD.n782 9.3005
R19189 VDD.n1215 VDD.n1214 9.3005
R19190 VDD.n1216 VDD.n780 9.3005
R19191 VDD.n1217 VDD.n778 9.3005
R19192 VDD.n1220 VDD.n1219 9.3005
R19193 VDD.n1222 VDD.n1221 9.3005
R19194 VDD.n1223 VDD.n774 9.3005
R19195 VDD.n1226 VDD.n1225 9.3005
R19196 VDD.n1227 VDD.n773 9.3005
R19197 VDD.n1229 VDD.n1228 9.3005
R19198 VDD.n1230 VDD.n772 9.3005
R19199 VDD.n1233 VDD.n1232 9.3005
R19200 VDD.n1235 VDD.n1234 9.3005
R19201 VDD.n1236 VDD.n769 9.3005
R19202 VDD.n1237 VDD.n767 9.3005
R19203 VDD.n1240 VDD.n1239 9.3005
R19204 VDD.n1242 VDD.n1241 9.3005
R19205 VDD.n1244 VDD.n764 9.3005
R19206 VDD.n1247 VDD.n1246 9.3005
R19207 VDD.n1248 VDD.n763 9.3005
R19208 VDD.n1250 VDD.n1249 9.3005
R19209 VDD.n1251 VDD.n761 9.3005
R19210 VDD.n1253 VDD.n1252 9.3005
R19211 VDD.n1254 VDD.n760 9.3005
R19212 VDD.n1256 VDD.n1255 9.3005
R19213 VDD.n759 VDD.n758 9.3005
R19214 VDD.n1263 VDD.n1262 9.3005
R19215 VDD.n1265 VDD.n1264 9.3005
R19216 VDD.n1267 VDD.n756 9.3005
R19217 VDD.n1269 VDD.n1268 9.3005
R19218 VDD.n1271 VDD.n1270 9.3005
R19219 VDD.n1273 VDD.n754 9.3005
R19220 VDD.n1277 VDD.n1276 9.3005
R19221 VDD.n1278 VDD.n753 9.3005
R19222 VDD.n1280 VDD.n1279 9.3005
R19223 VDD.n1281 VDD.n751 9.3005
R19224 VDD.n1282 VDD.n749 9.3005
R19225 VDD.n1284 VDD.n1283 9.3005
R19226 VDD.n1285 VDD.n748 9.3005
R19227 VDD.n1287 VDD.n1286 9.3005
R19228 VDD.n1288 VDD.n745 9.3005
R19229 VDD.n1291 VDD.n1290 9.3005
R19230 VDD.n1292 VDD.n744 9.3005
R19231 VDD.n1294 VDD.n1293 9.3005
R19232 VDD.n1295 VDD.n743 9.3005
R19233 VDD.n1297 VDD.n1296 9.3005
R19234 VDD.n1298 VDD.n742 9.3005
R19235 VDD.n1300 VDD.n1299 9.3005
R19236 VDD.n1301 VDD.n741 9.3005
R19237 VDD.n1302 VDD.n740 9.3005
R19238 VDD.n1303 VDD.n736 9.3005
R19239 VDD.n1306 VDD.n1305 9.3005
R19240 VDD.n1307 VDD.n735 9.3005
R19241 VDD.n1309 VDD.n1308 9.3005
R19242 VDD.n1310 VDD.n732 9.3005
R19243 VDD.n1312 VDD.n1311 9.3005
R19244 VDD.n1313 VDD.n731 9.3005
R19245 VDD.n1315 VDD.n1314 9.3005
R19246 VDD.n1316 VDD.n730 9.3005
R19247 VDD.n1320 VDD.n1319 9.3005
R19248 VDD.n1321 VDD.n729 9.3005
R19249 VDD.n1323 VDD.n1322 9.3005
R19250 VDD.n1324 VDD.n728 9.3005
R19251 VDD.n1328 VDD.n1327 9.3005
R19252 VDD.n1329 VDD.n727 9.3005
R19253 VDD.n1331 VDD.n1330 9.3005
R19254 VDD.n1333 VDD.n725 9.3005
R19255 VDD.n1336 VDD.n1335 9.3005
R19256 VDD.n1337 VDD.n724 9.3005
R19257 VDD.n1339 VDD.n1338 9.3005
R19258 VDD.n1340 VDD.n722 9.3005
R19259 VDD.n1343 VDD.n1342 9.3005
R19260 VDD.n1345 VDD.n1344 9.3005
R19261 VDD.n1347 VDD.n718 9.3005
R19262 VDD.n1349 VDD.n1348 9.3005
R19263 VDD.n1351 VDD.n1350 9.3005
R19264 VDD.n1352 VDD.n713 9.3005
R19265 VDD.n1355 VDD.n1354 9.3005
R19266 VDD.n1356 VDD.n712 9.3005
R19267 VDD.n1403 VDD.n1357 9.3005
R19268 VDD.n1402 VDD.n1401 9.3005
R19269 VDD.n1400 VDD.n1358 9.3005
R19270 VDD.n1399 VDD.n1398 9.3005
R19271 VDD.n1397 VDD.n1359 9.3005
R19272 VDD.n1396 VDD.n1361 9.3005
R19273 VDD.n1395 VDD.n1394 9.3005
R19274 VDD.n1393 VDD.n1392 9.3005
R19275 VDD.n1390 VDD.n1363 9.3005
R19276 VDD.n1389 VDD.n1388 9.3005
R19277 VDD.n1387 VDD.n1366 9.3005
R19278 VDD.n1386 VDD.n1385 9.3005
R19279 VDD.n1384 VDD.n1367 9.3005
R19280 VDD.n1383 VDD.n1382 9.3005
R19281 VDD.n1381 VDD.n1369 9.3005
R19282 VDD.n1380 VDD.n1379 9.3005
R19283 VDD.n1378 VDD.n1370 9.3005
R19284 VDD.n1377 VDD.n1376 9.3005
R19285 VDD.n1375 VDD.n1372 9.3005
R19286 VDD.n1374 VDD.n1373 9.3005
R19287 VDD.n701 VDD.n699 9.3005
R19288 VDD.n1498 VDD.n1497 9.3005
R19289 VDD.n1496 VDD.n1495 9.3005
R19290 VDD.n1488 VDD.n703 9.3005
R19291 VDD.n1487 VDD.n1486 9.3005
R19292 VDD.n1485 VDD.n705 9.3005
R19293 VDD.n1483 VDD.n708 9.3005
R19294 VDD.n1482 VDD.n1481 9.3005
R19295 VDD.n1480 VDD.n1479 9.3005
R19296 VDD.n1476 VDD.n711 9.3005
R19297 VDD.n1475 VDD.n1407 9.3005
R19298 VDD.n1474 VDD.n1408 9.3005
R19299 VDD.n1473 VDD.n1472 9.3005
R19300 VDD.n1471 VDD.n1410 9.3005
R19301 VDD.n1470 VDD.n1469 9.3005
R19302 VDD.n1467 VDD.n1411 9.3005
R19303 VDD.n1466 VDD.n1465 9.3005
R19304 VDD.n1464 VDD.n1463 9.3005
R19305 VDD.n1462 VDD.n1415 9.3005
R19306 VDD.n1461 VDD.n1416 9.3005
R19307 VDD.n1460 VDD.n1459 9.3005
R19308 VDD.n1458 VDD.n1418 9.3005
R19309 VDD.n1457 VDD.n1456 9.3005
R19310 VDD.n1455 VDD.n1419 9.3005
R19311 VDD.n1454 VDD.n1424 9.3005
R19312 VDD.n1453 VDD.n1425 9.3005
R19313 VDD.n1452 VDD.n1451 9.3005
R19314 VDD.n1450 VDD.n1428 9.3005
R19315 VDD.n1449 VDD.n1448 9.3005
R19316 VDD.n1447 VDD.n1429 9.3005
R19317 VDD.n1446 VDD.n1445 9.3005
R19318 VDD.n1444 VDD.n1432 9.3005
R19319 VDD.n1443 VDD.n1442 9.3005
R19320 VDD.n668 VDD.n652 9.3005
R19321 VDD.n665 VDD.n653 9.3005
R19322 VDD.n663 VDD.n662 9.3005
R19323 VDD.n667 VDD.n666 9.3005
R19324 VDD.n670 VDD.n669 9.3005
R19325 VDD.n672 VDD.n649 9.3005
R19326 VDD.n674 VDD.n673 9.3005
R19327 VDD.n676 VDD.n675 9.3005
R19328 VDD.n678 VDD.n640 9.3005
R19329 VDD.n680 VDD.n679 9.3005
R19330 VDD.n682 VDD.n681 9.3005
R19331 VDD.n683 VDD.n637 9.3005
R19332 VDD.n685 VDD.n684 9.3005
R19333 VDD.n687 VDD.n686 9.3005
R19334 VDD.n689 VDD.n607 9.3005
R19335 VDD.n691 VDD.n690 9.3005
R19336 VDD.n623 VDD.n617 9.3005
R19337 VDD.n625 VDD.n624 9.3005
R19338 VDD.n627 VDD.n626 9.3005
R19339 VDD.n628 VDD.n613 9.3005
R19340 VDD.n630 VDD.n629 9.3005
R19341 VDD.n632 VDD.n631 9.3005
R19342 VDD.n633 VDD.n606 9.3005
R19343 VDD.n594 VDD.n555 9.3005
R19344 VDD.n590 VDD.n557 9.3005
R19345 VDD.n586 VDD.n558 9.3005
R19346 VDD.n583 VDD.n582 9.3005
R19347 VDD.n581 VDD.n565 9.3005
R19348 VDD.n577 VDD.n566 9.3005
R19349 VDD.n576 VDD.n575 9.3005
R19350 VDD.n579 VDD.n578 9.3005
R19351 VDD.n585 VDD.n584 9.3005
R19352 VDD.n589 VDD.n588 9.3005
R19353 VDD.n592 VDD.n591 9.3005
R19354 VDD.n596 VDD.n595 9.3005
R19355 VDD.n540 VDD.n534 9.3005
R19356 VDD.n542 VDD.n541 9.3005
R19357 VDD.n544 VDD.n543 9.3005
R19358 VDD.n545 VDD.n530 9.3005
R19359 VDD.n547 VDD.n546 9.3005
R19360 VDD.n549 VDD.n548 9.3005
R19361 VDD.n550 VDD.n525 9.3005
R19362 VDD.n603 VDD.n602 9.3005
R19363 VDD.n601 VDD.n526 9.3005
R19364 VDD.n599 VDD.n598 9.3005
R19365 VDD.n597 VDD.n554 9.3005
R19366 VDD.n514 VDD.n475 9.3005
R19367 VDD.n510 VDD.n477 9.3005
R19368 VDD.n506 VDD.n478 9.3005
R19369 VDD.n503 VDD.n502 9.3005
R19370 VDD.n501 VDD.n485 9.3005
R19371 VDD.n497 VDD.n486 9.3005
R19372 VDD.n496 VDD.n495 9.3005
R19373 VDD.n499 VDD.n498 9.3005
R19374 VDD.n505 VDD.n504 9.3005
R19375 VDD.n509 VDD.n508 9.3005
R19376 VDD.n512 VDD.n511 9.3005
R19377 VDD.n516 VDD.n515 9.3005
R19378 VDD.n460 VDD.n454 9.3005
R19379 VDD.n462 VDD.n461 9.3005
R19380 VDD.n464 VDD.n463 9.3005
R19381 VDD.n465 VDD.n450 9.3005
R19382 VDD.n467 VDD.n466 9.3005
R19383 VDD.n469 VDD.n468 9.3005
R19384 VDD.n470 VDD.n445 9.3005
R19385 VDD.n523 VDD.n522 9.3005
R19386 VDD.n521 VDD.n446 9.3005
R19387 VDD.n519 VDD.n518 9.3005
R19388 VDD.n517 VDD.n474 9.3005
R19389 VDD.n432 VDD.n344 9.3005
R19390 VDD.n430 VDD.n429 9.3005
R19391 VDD.n428 VDD.n427 9.3005
R19392 VDD.n425 VDD.n349 9.3005
R19393 VDD.n439 VDD.n438 9.3005
R19394 VDD.n440 VDD.n339 9.3005
R19395 VDD.n442 VDD.n441 9.3005
R19396 VDD.n340 VDD.n338 9.3005
R19397 VDD.n210 VDD.n196 9.3005
R19398 VDD.n142 VDD.n131 9.3005
R19399 VDD.n138 VDD.n132 9.3005
R19400 VDD.n140 VDD.n139 9.3005
R19401 VDD.n163 VDD.n162 9.3005
R19402 VDD.n161 VDD.n124 9.3005
R19403 VDD.n160 VDD.n159 9.3005
R19404 VDD.n70 VDD.n63 9.3005
R19405 VDD.n78 VDD.n77 9.3005
R19406 VDD.n76 VDD.n64 9.3005
R19407 VDD.n75 VDD.n74 9.3005
R19408 VDD.n42 VDD.n41 9.3005
R19409 VDD.n38 VDD.n27 9.3005
R19410 VDD.n34 VDD.n31 9.3005
R19411 VDD.n37 VDD.n35 9.3005
R19412 VDD.n3054 VDD.n3053 9.14336
R19413 VDD.n1887 VDD.n1885 9.09802
R19414 VDD.n1899 VDD.n1898 9.09802
R19415 VDD.n4491 VDD.n4490 9.03579
R19416 VDD.n4331 VDD.n4270 9.03579
R19417 VDD.n4194 VDD.n4139 9.03579
R19418 VDD.n4190 VDD.n4189 9.03579
R19419 VDD.n3734 VDD.n3733 9.03579
R19420 VDD.n3525 VDD.n3524 9.03579
R19421 VDD.n3516 VDD.n3262 9.03579
R19422 VDD.n3459 VDD.n3458 9.03579
R19423 VDD.n3385 VDD.n3384 9.03579
R19424 VDD.n2523 VDD.n2522 9.03579
R19425 VDD.n2354 VDD.n2353 9.03579
R19426 VDD.n2643 VDD.n2642 9.03579
R19427 VDD.n2049 VDD.n1545 9.03579
R19428 VDD.n1906 VDD.n1576 9.03579
R19429 VDD.n2241 VDD.n2240 9.03579
R19430 VDD.n1080 VDD.n817 9.03579
R19431 VDD.n1038 VDD.n1037 9.03579
R19432 VDD.n961 VDD.n960 9.03579
R19433 VDD.n1211 VDD.n1210 9.03579
R19434 VDD.n3496 VDD.n3274 8.77764
R19435 VDD.n3486 VDD.n3485 8.77764
R19436 VDD.n3477 VDD.n3476 8.77764
R19437 VDD.n1820 VDD.n1819 8.77764
R19438 VDD.n661 VDD.n660 8.76674
R19439 VDD.n568 VDD.n567 8.76674
R19440 VDD.n488 VDD.n487 8.76674
R19441 VDD.n3763 VDD.n3761 8.65932
R19442 VDD.n2970 VDD.n2969 8.65932
R19443 VDD.n1788 VDD.n1787 8.65932
R19444 VDD.n1028 VDD.n817 8.65932
R19445 VDD.t1395 VDD.t3667 8.39273
R19446 VDD.t639 VDD.t461 8.39273
R19447 VDD.t908 VDD.t2191 8.39273
R19448 VDD.t3033 VDD.t1713 8.39273
R19449 VDD.t1173 VDD.t1987 8.39273
R19450 VDD.t3330 VDD.t3650 8.39273
R19451 VDD.t843 VDD.t2878 8.39273
R19452 VDD.t2364 VDD.t40 8.39273
R19453 VDD.t341 VDD.t588 8.39273
R19454 VDD.t1893 VDD.t2692 8.39273
R19455 VDD.t2743 VDD.t2017 8.39273
R19456 VDD.t1306 VDD.t3036 8.39273
R19457 VDD.n4396 VDD.n4395 8.28285
R19458 VDD.n2536 VDD.n2535 8.28285
R19459 VDD.n1088 VDD.n811 8.28285
R19460 VDD.n135 VDD.n132 8.28285
R19461 VDD.n141 VDD.n140 8.28285
R19462 VDD.n160 VDD.n125 8.28285
R19463 VDD.n314 VDD.n313 8.27619
R19464 VDD.n52 VDD.n48 8.22907
R19465 VDD.n24 VDD.n12 8.22907
R19466 VDD.n3566 VDD.n3565 7.90638
R19467 VDD.n2537 VDD.n2536 7.90638
R19468 VDD.n2991 VDD.n2367 7.90638
R19469 VDD.n1455 VDD.n1454 7.90638
R19470 VDD.n661 VDD.n659 7.61813
R19471 VDD.n574 VDD.n568 7.61813
R19472 VDD.n494 VDD.n488 7.61813
R19473 VDD.n2931 VDD.n2930 7.52991
R19474 VDD.n2545 VDD.n2544 7.52991
R19475 VDD.n2611 VDD.n2609 7.52991
R19476 VDD.n1799 VDD.n1635 7.52991
R19477 VDD.n1776 VDD.n1775 7.52991
R19478 VDD.n1745 VDD.n1744 7.52991
R19479 VDD.n2147 VDD.n2136 7.52991
R19480 VDD.n55 VDD.n54 7.4005
R19481 VDD.n59 VDD.n58 7.4005
R19482 VDD.n22 VDD.n21 7.4005
R19483 VDD.n18 VDD.n17 7.4005
R19484 VDD.n441 VDD.n340 7.3605
R19485 VDD.n441 VDD.n440 7.3605
R19486 VDD.n440 VDD.n439 7.3605
R19487 VDD.n439 VDD.n342 7.3605
R19488 VDD.n3972 VDD.n3971 7.23528
R19489 VDD.n4182 VDD.n4181 7.15344
R19490 VDD.n4178 VDD.n4177 7.15344
R19491 VDD.n3657 VDD.n3656 7.15344
R19492 VDD.n3539 VDD.n3538 7.15344
R19493 VDD.n3436 VDD.n3435 7.15344
R19494 VDD.n3380 VDD.n3294 7.15344
R19495 VDD.n2545 VDD.n2504 7.15344
R19496 VDD.n2565 VDD.n2563 7.15344
R19497 VDD.n2742 VDD.n2460 7.15344
R19498 VDD.n2336 VDD.n2303 7.15344
R19499 VDD.n1979 VDD.n1975 7.15344
R19500 VDD.n2243 VDD.n2174 7.15344
R19501 VDD.n1060 VDD.n1010 7.15344
R19502 VDD.n1232 VDD.n771 7.15344
R19503 VDD.n434 VDD.n433 7.13298
R19504 VDD.n1260 VDD.n1259 7.11866
R19505 VDD.n293 VDD.n292 7.11588
R19506 VDD.n331 VDD.n330 7.11588
R19507 VDD.n330 VDD.n329 7.11588
R19508 VDD.n3971 VDD.n3913 6.95702
R19509 VDD.n1820 VDD.n1619 6.94907
R19510 VDD.n2615 VDD.n2612 6.90844
R19511 VDD.n105 VDD.n89 6.9065
R19512 VDD.n137 VDD.n133 6.84103
R19513 VDD.n4638 VDD.n4637 6.77697
R19514 VDD.n4424 VDD.n4043 6.77697
R19515 VDD.n4301 VDD.n4286 6.77697
R19516 VDD.n3652 VDD.n3651 6.77697
R19517 VDD.n3869 VDD.n3868 6.77697
R19518 VDD.n2517 VDD.n2494 6.77697
R19519 VDD.n2964 VDD.n2963 6.77697
R19520 VDD.n1973 VDD.n1971 6.77697
R19521 VDD.n1796 VDD.n1795 6.77697
R19522 VDD.n1739 VDD.n1738 6.77697
R19523 VDD.n2251 VDD.n2250 6.77697
R19524 VDD.n1098 VDD.n1097 6.77697
R19525 VDD.n1035 VDD.n1034 6.77697
R19526 VDD.n1043 VDD.n1042 6.77697
R19527 VDD.n918 VDD.n917 6.77697
R19528 VDD.n1302 VDD.n1301 6.77697
R19529 VDD.n1165 VDD.n1164 6.77697
R19530 VDD.n1207 VDD.n1206 6.77697
R19531 VDD.n1482 VDD.n710 6.77697
R19532 VDD.n431 VDD.n430 6.77697
R19533 VDD.t1052 VDD.t1509 6.71428
R19534 VDD.t1352 VDD.t1861 6.71428
R19535 VDD.t2173 VDD.t3178 6.71428
R19536 VDD.t2378 VDD.t2341 6.71428
R19537 VDD.t3412 VDD.t1071 6.71428
R19538 VDD.t3318 VDD.t838 6.71428
R19539 VDD.t3632 VDD.t2366 6.71428
R19540 VDD.t2223 VDD.t1569 6.71428
R19541 VDD.t2221 VDD.t2292 6.71428
R19542 VDD.t3522 VDD.t985 6.71428
R19543 VDD.t42 VDD.t3726 6.71428
R19544 VDD.t309 VDD.t2425 6.71428
R19545 VDD.t1819 VDD.t1314 6.71428
R19546 VDD.t562 VDD.t1826 6.71428
R19547 VDD.t3488 VDD.t1318 6.71428
R19548 VDD.t2277 VDD.t2755 6.71428
R19549 VDD.t2371 VDD.t652 6.71428
R19550 VDD.t3051 VDD.t2688 6.71428
R19551 VDD.t1906 VDD.t3147 6.71428
R19552 VDD.t1690 VDD.t2506 6.71428
R19553 VDD.t2296 VDD.t2094 6.71428
R19554 VDD.t3616 VDD.t3454 6.71428
R19555 VDD.t3450 VDD.t584 6.71428
R19556 VDD.n137 VDD.n136 6.70566
R19557 VDD.n1887 VDD.n1886 6.66496
R19558 VDD.n1886 VDD.n1582 6.66496
R19559 VDD.n1894 VDD.n1893 6.66496
R19560 VDD.n2997 VDD.n2996 6.58336
R19561 VDD.n2812 VDD.n2811 6.58336
R19562 VDD.n61 VDD.n47 6.49269
R19563 VDD.n11 VDD.n10 6.49269
R19564 VDD.n4505 VDD.n4504 6.4005
R19565 VDD.n4472 VDD.n4450 6.4005
R19566 VDD.n4408 VDD.n4407 6.4005
R19567 VDD.n3719 VDD.n3698 6.4005
R19568 VDD.n3636 VDD.n3226 6.4005
R19569 VDD.n3770 VDD.n3193 6.4005
R19570 VDD.n1879 VDD.n1588 6.4005
R19571 VDD.n2145 VDD.n2144 6.4005
R19572 VDD.n2180 VDD.n2179 6.4005
R19573 VDD.n939 VDD.n937 6.4005
R19574 VDD.n1342 VDD.n1341 6.4005
R19575 VDD.n1398 VDD.n1397 6.4005
R19576 VDD.n1421 VDD.n1420 6.4005
R19577 VDD.n107 VDD.n106 6.39021
R19578 VDD.n252 VDD.n222 6.28433
R19579 VDD.n1898 VDD.n1579 6.24182
R19580 VDD.n4569 VDD.n3994 6.02403
R19581 VDD.n4023 VDD.n4017 6.02403
R19582 VDD.n4477 VDD.n4475 6.02403
R19583 VDD.n3749 VDD.n3748 6.02403
R19584 VDD.n3373 VDD.n3372 6.02403
R19585 VDD.n3111 VDD.n3110 6.02403
R19586 VDD.n3854 VDD.n3812 6.02403
R19587 VDD.n2878 VDD.n2829 6.02403
R19588 VDD.n2735 VDD.n2734 6.02403
R19589 VDD.n2629 VDD.n2627 6.02403
R19590 VDD.n2234 VDD.n2233 6.02403
R19591 VDD.n1053 VDD.n1052 6.02403
R19592 VDD.n1183 VDD.n1138 6.02403
R19593 VDD.n1373 VDD.n1372 6.02403
R19594 VDD.n1463 VDD.n1414 6.02403
R19595 VDD.n252 VDD.n251 5.94683
R19596 VDD.n254 VDD.n253 5.94683
R19597 VDD.n258 VDD.n219 5.94683
R19598 VDD.n264 VDD.n263 5.94683
R19599 VDD.n266 VDD.n265 5.94683
R19600 VDD.n270 VDD.n216 5.94683
R19601 VDD.n276 VDD.n275 5.94683
R19602 VDD.n278 VDD.n277 5.94683
R19603 VDD.n282 VDD.n211 5.94683
R19604 VDD.n288 VDD.n287 5.94683
R19605 VDD.n3493 VDD.n3492 5.85193
R19606 VDD.n3493 VDD.n3274 5.85193
R19607 VDD.n62 VDD.n46 5.80439
R19608 VDD.n26 VDD.n25 5.80403
R19609 VDD.n248 VDD.n247 5.78447
R19610 VDD.n250 VDD.n221 5.78447
R19611 VDD.n256 VDD.n255 5.78447
R19612 VDD.n259 VDD.n257 5.78447
R19613 VDD.n262 VDD.n218 5.78447
R19614 VDD.n268 VDD.n267 5.78447
R19615 VDD.n271 VDD.n269 5.78447
R19616 VDD.n274 VDD.n215 5.78447
R19617 VDD.n280 VDD.n279 5.78447
R19618 VDD.n283 VDD.n281 5.78447
R19619 VDD.n286 VDD.n213 5.78447
R19620 VDD.n99 VDD.n90 5.78175
R19621 VDD.n99 VDD.n98 5.78175
R19622 VDD.n97 VDD.n91 5.78175
R19623 VDD.n98 VDD.n97 5.78175
R19624 VDD.n168 VDD.n167 5.78175
R19625 VDD.n167 VDD.n166 5.78175
R19626 VDD.n172 VDD.n96 5.78175
R19627 VDD.n166 VDD.n96 5.78175
R19628 VDD.n157 VDD.n87 5.73998
R19629 VDD.n4264 VDD.n4263 5.64756
R19630 VDD.n4252 VDD.n4251 5.64756
R19631 VDD.n654 VDD.n652 5.64756
R19632 VDD.n594 VDD.n593 5.64756
R19633 VDD.n581 VDD.n580 5.64756
R19634 VDD.n514 VDD.n513 5.64756
R19635 VDD.n501 VDD.n500 5.64756
R19636 VDD.n2821 VDD.n2820 5.48621
R19637 VDD.n437 VDD.n342 5.37145
R19638 VDD.n400 VDD.n399 5.34555
R19639 VDD.n1901 VDD.n1900 5.32709
R19640 VDD.n3561 VDD.n3560 5.27109
R19641 VDD.n3538 VDD.n3253 5.27109
R19642 VDD.n3471 VDD.n3288 5.27109
R19643 VDD.n2706 VDD.n2705 5.27109
R19644 VDD.n1849 VDD.n1603 5.27109
R19645 VDD.n1902 VDD.n1901 5.27109
R19646 VDD.n1475 VDD.n1474 5.27109
R19647 VDD.n4197 VDD.n4196 5.21731
R19648 VDD.n969 VDD.n968 5.2005
R19649 VDD.n407 VDD.n406 5.14633
R19650 VDD.n647 VDD.n642 5.0887
R19651 VDD.n682 VDD.n639 5.06396
R19652 VDD.n213 VDD.n212 5.063
R19653 VDD.n285 VDD.n197 5.058
R19654 VDD.n289 VDD.n288 5.05712
R19655 VDD.t674 VDD.t1682 5.03584
R19656 VDD.t2269 VDD.t1527 5.03584
R19657 VDD.t2663 VDD.t1537 5.03584
R19658 VDD.t711 VDD.t2517 5.03584
R19659 VDD.t3216 VDD.t536 5.03584
R19660 VDD.t801 VDD.t580 5.03584
R19661 VDD.t1724 VDD.t1644 5.03584
R19662 VDD.t1225 VDD.t1869 5.03584
R19663 VDD.t39 VDD.t952 5.03584
R19664 VDD.t1857 VDD.t3476 5.03584
R19665 VDD.t2225 VDD.t1817 5.03584
R19666 VDD.t3395 VDD.t3446 5.03584
R19667 VDD.t3574 VDD.t1228 5.03584
R19668 VDD.t1878 VDD.t3286 5.03584
R19669 VDD.t3101 VDD.t0 5.03584
R19670 VDD.t1030 VDD.t2335 5.03584
R19671 VDD.t2962 VDD.t1439 5.03584
R19672 VDD.t557 VDD.t2098 5.03584
R19673 VDD.n423 VDD.t2946 5.03584
R19674 VDD.n4330 VDD.n4329 4.89462
R19675 VDD.n3110 VDD.n3106 4.89462
R19676 VDD.n2350 VDD.n2349 4.89462
R19677 VDD.n2983 VDD.n2982 4.89462
R19678 VDD.n2640 VDD.n2480 4.89462
R19679 VDD.n2179 VDD.n2176 4.89462
R19680 VDD.n249 VDD.n248 4.838
R19681 VDD.n247 VDD.n246 4.813
R19682 VDD.n4170 VDD.n4169 4.75748
R19683 VDD.n3336 VDD.n3335 4.75748
R19684 VDD.n3141 VDD.n3133 4.75748
R19685 VDD.n2586 VDD.n2585 4.75748
R19686 VDD.n2321 VDD.n2320 4.75748
R19687 VDD.n1702 VDD.n1701 4.75748
R19688 VDD.n2205 VDD.n2204 4.75748
R19689 VDD.n1441 VDD.n1440 4.75748
R19690 VDD.n3479 VDD.n3284 4.75479
R19691 VDD.n2887 VDD.n2886 4.75479
R19692 VDD.n208 VDD.n196 4.70477
R19693 VDD.n4657 VDD.n4656 4.67352
R19694 VDD.n4484 VDD.n4483 4.67352
R19695 VDD.n4483 VDD.n4482 4.67352
R19696 VDD.n4416 VDD.n4046 4.67352
R19697 VDD.n4420 VDD.n4046 4.67352
R19698 VDD.n4386 VDD.n4385 4.67352
R19699 VDD.n4313 VDD.n4282 4.67352
R19700 VDD.n4217 VDD.n4215 4.67352
R19701 VDD.n4221 VDD.n4126 4.67352
R19702 VDD.n4222 VDD.n4221 4.67352
R19703 VDD.n3967 VDD.n3916 4.67352
R19704 VDD.n3963 VDD.n3916 4.67352
R19705 VDD.n3676 VDD.n3203 4.67352
R19706 VDD.n3677 VDD.n3676 4.67352
R19707 VDD.n3354 VDD.n3305 4.67352
R19708 VDD.n3161 VDD.n3119 4.67352
R19709 VDD.n3157 VDD.n3156 4.67352
R19710 VDD.n3156 VDD.n3155 4.67352
R19711 VDD.n2555 VDD.n2554 4.67352
R19712 VDD.n3040 VDD.n3020 4.67352
R19713 VDD.n2766 VDD.n2763 4.67352
R19714 VDD.n2342 VDD.n2341 4.67352
R19715 VDD.n1918 VDD.n1917 4.67352
R19716 VDD.n1922 VDD.n1921 4.67352
R19717 VDD.n1924 VDD.n1922 4.67352
R19718 VDD.n1268 VDD.n1267 4.67352
R19719 VDD.n1767 VDD.n1766 4.62124
R19720 VDD.n2012 VDD.n2010 4.62124
R19721 VDD.n2152 VDD.n2131 4.62124
R19722 VDD.n400 VDD.n398 4.60988
R19723 VDD.n405 VDD.n404 4.60206
R19724 VDD.n350 VDD.n349 4.58437
R19725 VDD.n2557 VDD.n2556 4.57193
R19726 VDD.n2554 VDD.n2502 4.57193
R19727 VDD.n4676 VDD.n3895 4.51401
R19728 VDD.n4668 VDD.n4667 4.51401
R19729 VDD.n3891 VDD.n3092 4.51401
R19730 VDD.n3883 VDD.n3882 4.51401
R19731 VDD.n3088 VDD.n2276 4.51401
R19732 VDD.n3081 VDD.n3080 4.51401
R19733 VDD.n2272 VDD.n1505 4.51401
R19734 VDD.n2265 VDD.n2264 4.51401
R19735 VDD.n1501 VDD.n697 4.51401
R19736 VDD.n1494 VDD.n1493 4.51401
R19737 VDD.n305 VDD.n297 4.5127
R19738 VDD.n312 VDD.n298 4.5127
R19739 VDD.n323 VDD.n298 4.5127
R19740 VDD.n4675 VDD.n4674 4.5005
R19741 VDD.n4663 VDD.n3898 4.5005
R19742 VDD.n4666 VDD.n3902 4.5005
R19743 VDD.n3890 VDD.n3889 4.5005
R19744 VDD.n3878 VDD.n3095 4.5005
R19745 VDD.n3881 VDD.n3099 4.5005
R19746 VDD.n3087 VDD.n3086 4.5005
R19747 VDD.n3076 VDD.n2279 4.5005
R19748 VDD.n3079 VDD.n2283 4.5005
R19749 VDD.n2271 VDD.n2270 4.5005
R19750 VDD.n2260 VDD.n1508 4.5005
R19751 VDD.n2263 VDD.n1511 4.5005
R19752 VDD.n1500 VDD.n1499 4.5005
R19753 VDD.n1489 VDD.n700 4.5005
R19754 VDD.n1492 VDD.n704 4.5005
R19755 VDD.n436 VDD.n435 4.5005
R19756 VDD.n436 VDD.n343 4.5005
R19757 VDD.n402 VDD.n401 4.5005
R19758 VDD.n403 VDD.n397 4.5005
R19759 VDD.n279 VDD.n214 4.5005
R19760 VDD.n274 VDD.n273 4.5005
R19761 VDD.n272 VDD.n271 4.5005
R19762 VDD.n267 VDD.n217 4.5005
R19763 VDD.n262 VDD.n261 4.5005
R19764 VDD.n260 VDD.n259 4.5005
R19765 VDD.n255 VDD.n220 4.5005
R19766 VDD.n250 VDD.n249 4.5005
R19767 VDD.n284 VDD.n283 4.5005
R19768 VDD.n286 VDD.n285 4.5005
R19769 VDD.n83 VDD.n82 4.5005
R19770 VDD.n85 VDD.n84 4.5005
R19771 VDD.n8 VDD.n7 4.5005
R19772 VDD.n6 VDD.n5 4.5005
R19773 VDD.n3491 VDD.n3490 4.38907
R19774 VDD.n1834 VDD.n1833 4.38907
R19775 VDD.n1825 VDD.n1824 4.38907
R19776 VDD.n4382 VDD.n4381 4.36875
R19777 VDD.n4389 VDD.n4388 4.36875
R19778 VDD.n4284 VDD.n4282 4.36875
R19779 VDD.n4213 VDD.n4128 4.36875
R19780 VDD.n3963 VDD.n3962 4.36875
R19781 VDD.n3680 VDD.n3679 4.36875
R19782 VDD.n3357 VDD.n3356 4.36875
R19783 VDD.n3887 VDD.n3886 4.36875
R19784 VDD.n3164 VDD.n3163 4.36875
R19785 VDD.n2557 VDD.n2500 4.36875
R19786 VDD.n2551 VDD.n2550 4.36875
R19787 VDD.n2341 VDD.n2300 4.36875
R19788 VDD.n1915 VDD.n1574 4.36875
R19789 VDD.n1921 VDD.n1572 4.36875
R19790 VDD.n1924 VDD.n1923 4.36875
R19791 VDD.n1271 VDD.n755 4.36875
R19792 VDD.n1272 VDD.n1271 4.36875
R19793 VDD.n1245 VDD.n1244 4.36875
R19794 VDD.n3907 VDD.n3905 4.26717
R19795 VDD.n4224 VDD.n4223 4.26717
R19796 VDD.n3671 VDD.n3670 4.26717
R19797 VDD.n3125 VDD.n3123 4.26717
R19798 VDD.n605 VDD.n524 4.25409
R19799 VDD.n2765 VDD.n2764 4.21637
R19800 VDD.n4196 VDD.n4194 4.19546
R19801 VDD.n3804 VDD.n3803 4.19546
R19802 VDD.n1243 VDD.n1242 4.16558
R19803 VDD.n4596 VDD.n3983 4.14168
R19804 VDD.n4470 VDD.n4469 4.14168
R19805 VDD.n4412 VDD.n4051 4.14168
R19806 VDD.n4366 VDD.n4365 4.14168
R19807 VDD.n4360 VDD.n4357 4.14168
R19808 VDD.n3722 VDD.n3721 4.14168
R19809 VDD.n3389 VDD.n3388 4.14168
R19810 VDD.n2965 VDD.n2964 4.14168
R19811 VDD.n933 VDD.n883 4.14168
R19812 VDD.n866 VDD.n865 4.14168
R19813 VDD.n3023 VDD.n3022 4.06399
R19814 VDD.n3476 VDD.n3475 4.02336
R19815 VDD.n2813 VDD.n2812 4.02336
R19816 VDD.n4629 VDD.n4628 4.02033
R19817 VDD.n4548 VDD.n4008 4.02033
R19818 VDD.n4023 VDD.n4020 4.02033
R19819 VDD.n4394 VDD.n4066 4.02033
R19820 VDD.n4092 VDD.n4090 4.02033
R19821 VDD.n4168 VDD.n4164 4.02033
R19822 VDD.n4168 VDD.n4167 4.02033
R19823 VDD.n3937 VDD.n3933 4.02033
R19824 VDD.n3937 VDD.n3936 4.02033
R19825 VDD.n3342 VDD.n3322 4.02033
R19826 VDD.n3334 VDD.n3330 4.02033
R19827 VDD.n3334 VDD.n3333 4.02033
R19828 VDD.n3117 VDD.n3114 4.02033
R19829 VDD.n3140 VDD.n3136 4.02033
R19830 VDD.n3140 VDD.n3139 4.02033
R19831 VDD.n2592 VDD.n2571 4.02033
R19832 VDD.n2584 VDD.n2580 4.02033
R19833 VDD.n2584 VDD.n2583 4.02033
R19834 VDD.n2319 VDD.n2315 4.02033
R19835 VDD.n2319 VDD.n2318 4.02033
R19836 VDD.n1538 VDD.n1537 4.02033
R19837 VDD.n1700 VDD.n1696 4.02033
R19838 VDD.n1700 VDD.n1699 4.02033
R19839 VDD.n1872 VDD.n1870 4.02033
R19840 VDD.n1911 VDD.n1910 4.02033
R19841 VDD.n2203 VDD.n2199 4.02033
R19842 VDD.n2203 VDD.n2202 4.02033
R19843 VDD.n863 VDD.n859 4.02033
R19844 VDD.n863 VDD.n862 4.02033
R19845 VDD.n1439 VDD.n1435 4.02033
R19846 VDD.n1439 VDD.n1438 4.02033
R19847 VDD.n4421 VDD.n4420 4.0132
R19848 VDD.n693 VDD.n692 3.9555
R19849 VDD.n605 VDD.n604 3.9555
R19850 VDD.n1266 VDD.n1265 3.87908
R19851 VDD.n164 VDD.n123 3.77767
R19852 VDD.n4570 VDD.n4569 3.76521
R19853 VDD.n4478 VDD.n4477 3.76521
R19854 VDD.n3940 VDD.n3939 3.76521
R19855 VDD.n3748 VDD.n3746 3.76521
R19856 VDD.n3458 VDD.n3396 3.76521
R19857 VDD.n3372 VDD.n3371 3.76521
R19858 VDD.n2971 VDD.n2970 3.76521
R19859 VDD.n2630 VDD.n2629 3.76521
R19860 VDD.n2724 VDD.n2473 3.76521
R19861 VDD.n1849 VDD.n1848 3.76521
R19862 VDD.n1809 VDD.n1808 3.76521
R19863 VDD.n1775 VDD.n1646 3.76521
R19864 VDD.n1760 VDD.n1759 3.76521
R19865 VDD.n2235 VDD.n2234 3.76521
R19866 VDD.n2228 VDD.n2227 3.76521
R19867 VDD.n2227 VDD.n2226 3.76521
R19868 VDD.n1097 VDD.n808 3.76521
R19869 VDD.n1052 VDD.n1050 3.76521
R19870 VDD.n1073 VDD.n1006 3.76521
R19871 VDD.n1353 VDD.n1352 3.76521
R19872 VDD.n1289 VDD.n1288 3.76521
R19873 VDD.n1275 VDD.n753 3.76521
R19874 VDD.n1180 VDD.n1138 3.76521
R19875 VDD.n1466 VDD.n1414 3.76521
R19876 VDD.n73 VDD.n72 3.76521
R19877 VDD.n33 VDD.n32 3.76521
R19878 VDD.n3976 VDD.n3975 3.76495
R19879 VDD.n3313 VDD.n3312 3.76495
R19880 VDD.n642 VDD.n636 3.73715
R19881 VDD.n4216 VDD.n4126 3.70844
R19882 VDD.n3678 VDD.n3677 3.70844
R19883 VDD.n3157 VDD.n3121 3.70844
R19884 VDD.n3492 VDD.n3491 3.65764
R19885 VDD.n69 VDD.n68 3.63311
R19886 VDD.n40 VDD.n30 3.63295
R19887 VDD.n294 VDD.n188 3.62795
R19888 VDD.t3576 VDD.n294 3.62795
R19889 VDD.n206 VDD.n194 3.62795
R19890 VDD.t3576 VDD.n194 3.62795
R19891 VDD.n1895 VDD.n1579 3.49141
R19892 VDD.n4667 VDD.n0 3.43925
R19893 VDD.n4677 VDD.n4676 3.43925
R19894 VDD.n3882 VDD.n1 3.43925
R19895 VDD.n3892 VDD.n3891 3.43925
R19896 VDD.n3080 VDD.n2 3.43925
R19897 VDD.n3089 VDD.n3088 3.43925
R19898 VDD.n2264 VDD.n3 3.43925
R19899 VDD.n2273 VDD.n2272 3.43925
R19900 VDD.n1493 VDD.n4 3.43925
R19901 VDD.n1502 VDD.n1501 3.43925
R19902 VDD.n644 VDD.n636 3.43136
R19903 VDD.n3896 VDD.n3894 3.4105
R19904 VDD.n4665 VDD.n4664 3.4105
R19905 VDD.n3093 VDD.n3091 3.4105
R19906 VDD.n3880 VDD.n3879 3.4105
R19907 VDD.n2277 VDD.n2275 3.4105
R19908 VDD.n3078 VDD.n3077 3.4105
R19909 VDD.n1506 VDD.n1504 3.4105
R19910 VDD.n2262 VDD.n2261 3.4105
R19911 VDD.n698 VDD.n696 3.4105
R19912 VDD.n1491 VDD.n1490 3.4105
R19913 VDD.n4475 VDD.n4450 3.38874
R19914 VDD.n3716 VDD.n3698 3.38874
R19915 VDD.n3773 VDD.n3193 3.38874
R19916 VDD.n2006 VDD.n2005 3.38874
R19917 VDD.n2146 VDD.n2145 3.38874
R19918 VDD.n1115 VDD.n1114 3.38874
R19919 VDD.n940 VDD.n939 3.38874
R19920 VDD.n634 VDD.n633 3.38874
R19921 VDD.n551 VDD.n550 3.38874
R19922 VDD.n471 VDD.n470 3.38874
R19923 VDD.n136 VDD.n135 3.38874
R19924 VDD.t2972 VDD.t2575 3.35739
R19925 VDD.t82 VDD.t2618 3.35739
R19926 VDD.n4503 VDD.t1907 3.35739
R19927 VDD.t2441 VDD.t2847 3.35739
R19928 VDD.t203 VDD.t2465 3.35739
R19929 VDD.t225 VDD.t1739 3.35739
R19930 VDD.t1054 VDD.t2477 3.35739
R19931 VDD.t1975 VDD.t163 3.35739
R19932 VDD.t3618 VDD.t3607 3.35739
R19933 VDD.t966 VDD.t511 3.35739
R19934 VDD.t3084 VDD.t2031 3.35739
R19935 VDD.t894 VDD.t1297 3.35739
R19936 VDD.t2820 VDD.t857 3.35739
R19937 VDD.t5 VDD.t3006 3.35739
R19938 VDD.t2557 VDD.t2968 3.35739
R19939 VDD.t221 VDD.t1516 3.35739
R19940 VDD.t1555 VDD.t2011 3.35739
R19941 VDD.t2501 VDD.t1354 3.35739
R19942 VDD.n2909 VDD.n2405 3.29193
R19943 VDD.n2910 VDD.n2909 3.29193
R19944 VDD.n3938 VDD.n3937 3.28705
R19945 VDD.n864 VDD.n863 3.28705
R19946 VDD.n424 VDD.n350 3.21639
R19947 VDD.n437 VDD.n436 3.18654
R19948 VDD.n1262 VDD.n757 3.16454
R19949 VDD.n4385 VDD.n4072 3.14971
R19950 VDD.n632 VDD.n611 3.12116
R19951 VDD.n1893 VDD.n1892 3.06827
R19952 VDD.n4345 VDD.n4092 3.04861
R19953 VDD.n4394 VDD.n4067 3.04861
R19954 VDD.n4531 VDD.n4023 3.04861
R19955 VDD.n4548 VDD.n4003 3.04861
R19956 VDD.n4629 VDD.n4605 3.04861
R19957 VDD.n3342 VDD.n3318 3.04861
R19958 VDD.n2592 VDD.n2572 3.04861
R19959 VDD.n1911 VDD.n1575 3.04861
R19960 VDD.n2066 VDD.n1538 3.04861
R19961 VDD.n1873 VDD.n1872 3.04861
R19962 VDD.n183 VDD.n182 3.03833
R19963 VDD.n2095 VDD.n1526 3.01226
R19964 VDD.n1123 VDD.n1122 3.01226
R19965 VDD.n4484 VDD.n4445 2.99733
R19966 VDD.n4416 VDD.n4415 2.99733
R19967 VDD.n3968 VDD.n3967 2.99733
R19968 VDD.n2344 VDD.n2298 2.99733
R19969 VDD.n1586 VDD.n1585 2.91308
R19970 VDD.n164 VDD.n163 2.90013
R19971 VDD.n3356 VDD.n3355 2.89574
R19972 VDD.n4444 VDD.n4441 2.87861
R19973 VDD.n4414 VDD.n4413 2.87861
R19974 VDD.n3976 VDD.n3970 2.87861
R19975 VDD.n3313 VDD.n3309 2.87861
R19976 VDD.n2347 VDD.n2295 2.87861
R19977 VDD.t1754 VDD.n148 2.857
R19978 VDD.n148 VDD.t1759 2.857
R19979 VDD.t1756 VDD.n149 2.857
R19980 VDD.n149 VDD.t1754 2.857
R19981 VDD.t3430 VDD.n128 2.857
R19982 VDD.n128 VDD.t3433 2.857
R19983 VDD.t3432 VDD.n129 2.857
R19984 VDD.n129 VDD.t3430 2.857
R19985 VDD.n4448 VDD.n4446 2.84494
R19986 VDD.n3307 VDD.n3306 2.79415
R19987 VDD.n1261 VDD.n759 2.76904
R19988 VDD.n334 VDD.n187 2.76312
R19989 VDD.n3974 VDD.n3971 2.75091
R19990 VDD.n53 VDD.n49 2.66717
R19991 VDD.n16 VDD.n13 2.66717
R19992 VDD.n3975 VDD.n3971 2.64513
R19993 VDD.n4629 VDD.n4625 2.63579
R19994 VDD.n3943 VDD.n3942 2.63579
R19995 VDD.n3709 VDD.n3708 2.63579
R19996 VDD.n1854 VDD.n1853 2.63579
R19997 VDD.n1760 VDD.n1654 2.63579
R19998 VDD.n1725 VDD.n1724 2.63579
R19999 VDD.n2141 VDD.n2140 2.63579
R20000 VDD.n1086 VDD.n1085 2.63579
R20001 VDD.n1073 VDD.n1072 2.63579
R20002 VDD.n913 VDD.n912 2.63579
R20003 VDD.n926 VDD.n925 2.63579
R20004 VDD.n869 VDD.n868 2.63579
R20005 VDD.n1219 VDD.n1218 2.63579
R20006 VDD.n427 VDD.n348 2.63579
R20007 VDD.n4628 VDD.n4626 2.63539
R20008 VDD.n4008 VDD.n4006 2.63539
R20009 VDD.n4020 VDD.n4018 2.63539
R20010 VDD.n4066 VDD.n4064 2.63539
R20011 VDD.n4090 VDD.n4088 2.63539
R20012 VDD.n4164 VDD.n4162 2.63539
R20013 VDD.n4167 VDD.n4165 2.63539
R20014 VDD.n3933 VDD.n3931 2.63539
R20015 VDD.n3936 VDD.n3934 2.63539
R20016 VDD.n3312 VDD.n3310 2.63539
R20017 VDD.n3322 VDD.n3320 2.63539
R20018 VDD.n3330 VDD.n3328 2.63539
R20019 VDD.n3333 VDD.n3331 2.63539
R20020 VDD.n3114 VDD.n3112 2.63539
R20021 VDD.n3136 VDD.n3134 2.63539
R20022 VDD.n3139 VDD.n3137 2.63539
R20023 VDD.n2571 VDD.n2569 2.63539
R20024 VDD.n2580 VDD.n2578 2.63539
R20025 VDD.n2583 VDD.n2581 2.63539
R20026 VDD.n2315 VDD.n2313 2.63539
R20027 VDD.n2318 VDD.n2316 2.63539
R20028 VDD.n1537 VDD.n1535 2.63539
R20029 VDD.n1696 VDD.n1694 2.63539
R20030 VDD.n1699 VDD.n1697 2.63539
R20031 VDD.n1870 VDD.n1868 2.63539
R20032 VDD.n1910 VDD.n1908 2.63539
R20033 VDD.n2199 VDD.n2197 2.63539
R20034 VDD.n2202 VDD.n2200 2.63539
R20035 VDD.n859 VDD.n857 2.63539
R20036 VDD.n862 VDD.n860 2.63539
R20037 VDD.n1435 VDD.n1433 2.63539
R20038 VDD.n1438 VDD.n1436 2.63539
R20039 VDD.n611 VDD.n609 2.63539
R20040 VDD.n4445 VDD.n4443 2.61352
R20041 VDD.n4415 VDD.n4048 2.61352
R20042 VDD.n3969 VDD.n3968 2.61352
R20043 VDD.n3308 VDD.n3307 2.61352
R20044 VDD.n2298 VDD.n2297 2.61352
R20045 VDD.n183 VDD.n87 2.59875
R20046 VDD.n4389 VDD.n4387 2.48939
R20047 VDD.n2343 VDD.n2342 2.48939
R20048 VDD.n435 VDD.n434 2.48504
R20049 VDD.n4214 VDD.n4213 2.4386
R20050 VDD.n3163 VDD.n3162 2.4386
R20051 VDD.n1916 VDD.n1915 2.4386
R20052 VDD.n4627 VDD.n4626 2.37495
R20053 VDD.n4007 VDD.n4006 2.37495
R20054 VDD.n4019 VDD.n4018 2.37495
R20055 VDD.n4065 VDD.n4064 2.37495
R20056 VDD.n4089 VDD.n4088 2.37495
R20057 VDD.n4166 VDD.n4165 2.37495
R20058 VDD.n4163 VDD.n4162 2.37495
R20059 VDD.n3935 VDD.n3934 2.37495
R20060 VDD.n3932 VDD.n3931 2.37495
R20061 VDD.n3311 VDD.n3310 2.37495
R20062 VDD.n3321 VDD.n3320 2.37495
R20063 VDD.n3332 VDD.n3331 2.37495
R20064 VDD.n3329 VDD.n3328 2.37495
R20065 VDD.n3113 VDD.n3112 2.37495
R20066 VDD.n3138 VDD.n3137 2.37495
R20067 VDD.n3135 VDD.n3134 2.37495
R20068 VDD.n2570 VDD.n2569 2.37495
R20069 VDD.n2582 VDD.n2581 2.37495
R20070 VDD.n2579 VDD.n2578 2.37495
R20071 VDD.n2317 VDD.n2316 2.37495
R20072 VDD.n2314 VDD.n2313 2.37495
R20073 VDD.n1536 VDD.n1535 2.37495
R20074 VDD.n1698 VDD.n1697 2.37495
R20075 VDD.n1695 VDD.n1694 2.37495
R20076 VDD.n1869 VDD.n1868 2.37495
R20077 VDD.n1909 VDD.n1908 2.37495
R20078 VDD.n2201 VDD.n2200 2.37495
R20079 VDD.n2198 VDD.n2197 2.37495
R20080 VDD.n861 VDD.n860 2.37495
R20081 VDD.n858 VDD.n857 2.37495
R20082 VDD.n1437 VDD.n1436 2.37495
R20083 VDD.n1434 VDD.n1433 2.37495
R20084 VDD.n610 VDD.n609 2.37495
R20085 VDD.n4658 VDD.n4657 2.33701
R20086 VDD.n4314 VDD.n4313 2.33701
R20087 VDD.n3830 VDD.n3829 2.33701
R20088 VDD.n3829 VDD.n3097 2.33701
R20089 VDD.n3887 VDD.n3097 2.33701
R20090 VDD.n2763 VDD.n2762 2.33701
R20091 VDD.n1242 VDD.n766 2.33701
R20092 VDD.n51 VDD.n49 2.313
R20093 VDD.n57 VDD.n51 2.313
R20094 VDD.n15 VDD.n13 2.313
R20095 VDD.n20 VDD.n15 2.313
R20096 VDD.n52 VDD.n50 2.28445
R20097 VDD.n56 VDD.n50 2.28445
R20098 VDD.n14 VDD.n12 2.28445
R20099 VDD.n19 VDD.n14 2.28445
R20100 VDD.n155 VDD.n154 2.28415
R20101 VDD.n4638 VDD.n4601 2.25932
R20102 VDD.n4525 VDD.n4524 2.25932
R20103 VDD.n4293 VDD.n4292 2.25932
R20104 VDD.n3524 VDD.n3523 2.25932
R20105 VDD.n3851 VDD.n3850 2.25932
R20106 VDD.n2930 VDD.n2929 2.25932
R20107 VDD.n2916 VDD.n2402 2.25932
R20108 VDD.n2350 VDD.n2292 2.25932
R20109 VDD.n2953 VDD.n2952 2.25932
R20110 VDD.n2989 VDD.n2370 2.25932
R20111 VDD.n2601 VDD.n2492 2.25932
R20112 VDD.n2705 VDD.n2704 2.25932
R20113 VDD.n1841 VDD.n1840 2.25932
R20114 VDD.n1725 VDD.n1679 2.25932
R20115 VDD.n2096 VDD.n2095 2.25932
R20116 VDD.n2026 VDD.n1560 2.25932
R20117 VDD.n2136 VDD.n2133 2.25932
R20118 VDD.n947 VDD.n946 2.25932
R20119 VDD.n874 VDD.n873 2.25932
R20120 VDD.n875 VDD.n874 2.25932
R20121 VDD.n1345 VDD.n721 2.25932
R20122 VDD.n1305 VDD.n1304 2.25932
R20123 VDD.n1232 VDD.n1231 2.25932
R20124 VDD.n1166 VDD.n1147 2.25932
R20125 VDD.n671 VDD.n670 2.25932
R20126 VDD.n582 VDD.n564 2.25932
R20127 VDD.n502 VDD.n484 2.25932
R20128 VDD.n2347 VDD.n2346 2.25312
R20129 VDD.n1889 VDD.n1586 2.25312
R20130 VDD.n4413 VDD.n4047 2.25293
R20131 VDD.n4486 VDD.n4441 2.25293
R20132 VDD.n3351 VDD.n3313 2.25293
R20133 VDD.n3167 VDD.n3117 2.25293
R20134 VDD.n4215 VDD.n4214 2.23542
R20135 VDD.n3162 VDD.n3161 2.23542
R20136 VDD.n1917 VDD.n1916 2.23542
R20137 VDD.n4387 VDD.n4386 2.18463
R20138 VDD.n2344 VDD.n2343 2.18463
R20139 VDD.n1258 VDD.n1257 2.1578
R20140 VDD.n42 VDD.n30 2.05049
R20141 VDD.n68 VDD.n63 2.05017
R20142 VDD.n4659 VDD.n4658 2.03225
R20143 VDD.n4315 VDD.n4314 2.03225
R20144 VDD.n3831 VDD.n3830 2.03225
R20145 VDD.n3043 VDD.n3042 2.03225
R20146 VDD.n2762 VDD.n2761 2.03225
R20147 VDD.n1238 VDD.n766 2.03225
R20148 VDD.n1585 VDD.n1583 2.01703
R20149 VDD.n178 VDD.n177 2.01137
R20150 VDD.n177 VDD.t1753 2.01137
R20151 VDD.n104 VDD.n95 2.01137
R20152 VDD.t1753 VDD.n95 2.01137
R20153 VDD.n176 VDD.n175 2.01137
R20154 VDD.t1753 VDD.n176 2.01137
R20155 VDD.n180 VDD.n179 1.9205
R20156 VDD.n1584 VDD.n1583 1.88416
R20157 VDD.n4430 VDD.n4429 1.88285
R20158 VDD.n3414 VDD.n3290 1.88285
R20159 VDD.n2309 VDD.n2306 1.88285
R20160 VDD.n1998 VDD.n1997 1.88285
R20161 VDD.n2007 VDD.n2006 1.88285
R20162 VDD.n2085 VDD.n2084 1.88285
R20163 VDD.n2214 VDD.n2213 1.88285
R20164 VDD.n1334 VDD.n1333 1.88285
R20165 VDD.n30 VDD.n29 1.87577
R20166 VDD.n68 VDD.n67 1.87546
R20167 VDD.n3054 VDD.n3006 1.82907
R20168 VDD.n81 VDD.n80 1.79129
R20169 VDD.n3355 VDD.n3354 1.77828
R20170 VDD.n3976 VDD.n3914 1.76869
R20171 VDD.n1503 VDD.n4 1.69188
R20172 VDD.n1503 VDD.n1502 1.69188
R20173 VDD.n2274 VDD.n3 1.69188
R20174 VDD.n2274 VDD.n2273 1.69188
R20175 VDD.n3090 VDD.n2 1.69188
R20176 VDD.n3090 VDD.n3089 1.69188
R20177 VDD.n3893 VDD.n1 1.69188
R20178 VDD.n3893 VDD.n3892 1.69188
R20179 VDD.n4678 VDD.n0 1.69188
R20180 VDD.n4678 VDD.n4677 1.69188
R20181 VDD.n1886 VDD.n1586 1.68673
R20182 VDD.n4169 VDD.n4168 1.6819
R20183 VDD.n3335 VDD.n3334 1.6819
R20184 VDD.n3141 VDD.n3140 1.6819
R20185 VDD.n2585 VDD.n2584 1.6819
R20186 VDD.n2320 VDD.n2319 1.6819
R20187 VDD.n1701 VDD.n1700 1.6819
R20188 VDD.n2204 VDD.n2203 1.6819
R20189 VDD.n1440 VDD.n1439 1.6819
R20190 VDD.t1680 VDD.t3572 1.67895
R20191 VDD.t2869 VDD.t2267 1.67895
R20192 VDD.t2245 VDD.t1486 1.67895
R20193 VDD.t1091 VDD.t734 1.67895
R20194 VDD.t736 VDD.t3126 1.67895
R20195 VDD.t415 VDD.t2039 1.67895
R20196 VDD.t3170 VDD.t3166 1.67895
R20197 VDD.t3194 VDD.t1645 1.67895
R20198 VDD.t1579 VDD.t3314 1.67895
R20199 VDD.t1278 VDD.t954 1.67895
R20200 VDD.t349 VDD.t3508 1.67895
R20201 VDD.t160 VDD.t3371 1.67895
R20202 VDD.t1226 VDD.t2242 1.67895
R20203 VDD.t750 VDD.t805 1.67895
R20204 VDD.t249 VDD.t2229 1.67895
R20205 VDD.t236 VDD.t2189 1.67895
R20206 VDD.t267 VDD.t3694 1.67895
R20207 VDD.t1650 VDD.t503 1.67895
R20208 VDD.t666 VDD.t3468 1.67895
R20209 VDD.t629 VDD.t2532 1.67895
R20210 VDD.t631 VDD.t2534 1.67895
R20211 VDD.t3222 VDD.t3176 1.67895
R20212 VDD.t1234 VDD.t2034 1.67895
R20213 VDD.t2088 VDD.t3027 1.67895
R20214 VDD.t771 VDD.t3441 1.67895
R20215 VDD.t313 VDD.t1322 1.67895
R20216 VDD.t311 VDD.t3747 1.67895
R20217 VDD.n184 VDD.n86 1.65485
R20218 VDD.n2616 VDD.n2615 1.6259
R20219 VDD.n972 VDD.n968 1.6005
R20220 VDD.n45 VDD.n44 1.54166
R20221 VDD.n4482 VDD.n4446 1.52431
R20222 VDD.n4382 VDD.n4072 1.52431
R20223 VDD.n3042 VDD.n3041 1.52431
R20224 VDD.n3978 VDD.n3912 1.50638
R20225 VDD.n4550 VDD.n4002 1.50638
R20226 VDD.n4400 VDD.n4399 1.50638
R20227 VDD.n3646 VDD.n3644 1.50638
R20228 VDD.n3511 VDD.n3510 1.50638
R20229 VDD.n3512 VDD.n3511 1.50638
R20230 VDD.n3436 VDD.n3406 1.50638
R20231 VDD.n3455 VDD.n3396 1.50638
R20232 VDD.n3462 VDD.n3394 1.50638
R20233 VDD.n3380 VDD.n3379 1.50638
R20234 VDD.n3172 VDD.n3171 1.50638
R20235 VDD.n3846 VDD.n3820 1.50638
R20236 VDD.n2356 VDD.n2291 1.50638
R20237 VDD.n2985 VDD.n2370 1.50638
R20238 VDD.n2603 VDD.n2602 1.50638
R20239 VDD.n2641 VDD.n2640 1.50638
R20240 VDD.n2694 VDD.n2665 1.50638
R20241 VDD.n1992 VDD.n1991 1.50638
R20242 VDD.n1744 VDD.n1664 1.50638
R20243 VDD.n1710 VDD.n1709 1.50638
R20244 VDD.n1392 VDD.n1391 1.50638
R20245 VDD.n3498 VDD.n3497 1.46336
R20246 VDD.n2907 VDD.n2906 1.46336
R20247 VDD.n2999 VDD.n2360 1.46336
R20248 VDD.n2815 VDD.n2422 1.46336
R20249 VDD.n1833 VDD.n1832 1.46336
R20250 VDD.n335 VDD.n185 1.41175
R20251 VDD.n175 VDD.n174 1.4085
R20252 VDD.n973 VDD.n972 1.4005
R20253 VDD.n80 VDD.n79 1.3989
R20254 VDD.n44 VDD.n43 1.3989
R20255 VDD.n181 VDD.n89 1.3755
R20256 VDD.n184 VDD.n183 1.34504
R20257 VDD.n4172 VDD.n4169 1.30718
R20258 VDD.n3338 VDD.n3335 1.30718
R20259 VDD.n3142 VDD.n3141 1.30718
R20260 VDD.n2588 VDD.n2585 1.30718
R20261 VDD.n2323 VDD.n2320 1.30718
R20262 VDD.n1704 VDD.n1701 1.30718
R20263 VDD.n2207 VDD.n2204 1.30718
R20264 VDD.n1443 VDD.n1440 1.30718
R20265 VDD.n182 VDD.n181 1.2505
R20266 VDD.n4445 VDD.n4444 1.2502
R20267 VDD.n4415 VDD.n4414 1.2502
R20268 VDD.n3970 VDD.n3968 1.2502
R20269 VDD.n3309 VDD.n3307 1.2502
R20270 VDD.n2298 VDD.n2295 1.2502
R20271 VDD.n695 VDD.n45 1.22824
R20272 VDD.n444 VDD.n443 1.2116
R20273 VDD.n244 VDD.n243 1.17383
R20274 VDD.n4635 VDD.n4634 1.12991
R20275 VDD.n4558 VDD.n4557 1.12991
R20276 VDD.n4407 VDD.n4406 1.12991
R20277 VDD.n4207 VDD.n4132 1.12991
R20278 VDD.n3646 VDD.n3645 1.12991
R20279 VDD.n3767 VDD.n3195 1.12991
R20280 VDD.n2953 VDD.n2951 1.12991
R20281 VDD.n2798 VDD.n2797 1.12991
R20282 VDD.n2789 VDD.n2788 1.12991
R20283 VDD.n2789 VDD.n2437 1.12991
R20284 VDD.n2782 VDD.n2781 1.12991
R20285 VDD.n1846 VDD.n1845 1.12991
R20286 VDD.n678 VDD.n677 1.12991
R20287 VDD.n665 VDD.n664 1.12991
R20288 VDD.n561 VDD.n557 1.12991
R20289 VDD.n571 VDD.n566 1.12991
R20290 VDD.n481 VDD.n477 1.12991
R20291 VDD.n491 VDD.n486 1.12991
R20292 VDD.n2900 VDD.n2899 1.09764
R20293 VDD.n105 VDD.n104 1.09764
R20294 VDD.n337 VDD.n184 1.07996
R20295 VDD.n4202 VDD.n4135 1.07613
R20296 VDD.n444 VDD.n337 1.06614
R20297 VDD.n336 VDD.n335 1.03946
R20298 VDD.n969 VDD.n835 1.0005
R20299 VDD.n4217 VDD.n4216 0.965579
R20300 VDD.n3680 VDD.n3678 0.965579
R20301 VDD.n3121 VDD.n3119 0.965579
R20302 VDD.n1258 VDD.n759 0.935332
R20303 VDD.n4548 VDD.n4005 0.899674
R20304 VDD.n3342 VDD.n3324 0.899674
R20305 VDD.n2592 VDD.n2574 0.899674
R20306 VDD.n157 VDD.n156 0.841846
R20307 VDD.n4309 VDD.n4308 0.813843
R20308 VDD.n3041 VDD.n3040 0.813198
R20309 VDD.n2612 VDD.n2487 0.813198
R20310 VDD.n130 VDD.n126 0.757118
R20311 VDD.n127 VDD.n126 0.757118
R20312 VDD.n127 VDD.n88 0.757118
R20313 VDD.n150 VDD.n145 0.757118
R20314 VDD.n147 VDD.n145 0.757118
R20315 VDD.n147 VDD.n146 0.757118
R20316 VDD.n4621 VDD.n4620 0.753441
R20317 VDD.n4636 VDD.n4635 0.753441
R20318 VDD.n4644 VDD.n4643 0.753441
R20319 VDD.n4592 VDD.n4591 0.753441
R20320 VDD.n4576 VDD.n4575 0.753441
R20321 VDD.n4557 VDD.n4556 0.753441
R20322 VDD.n4551 VDD.n4550 0.753441
R20323 VDD.n4515 VDD.n4514 0.753441
R20324 VDD.n4495 VDD.n4494 0.753441
R20325 VDD.n4494 VDD.n4437 0.753441
R20326 VDD.n4401 VDD.n4400 0.753441
R20327 VDD.n4354 VDD.n4353 0.753441
R20328 VDD.n4280 VDD.n4276 0.753441
R20329 VDD.n4334 VDD.n4270 0.753441
R20330 VDD.n4191 VDD.n4139 0.753441
R20331 VDD.n3939 VDD.n3930 0.753441
R20332 VDD.n3733 VDD.n3732 0.753441
R20333 VDD.n3745 VDD.n3744 0.753441
R20334 VDD.n3664 VDD.n3206 0.753441
R20335 VDD.n3596 VDD.n3595 0.753441
R20336 VDD.n3623 VDD.n3574 0.753441
R20337 VDD.n3513 VDD.n3262 0.753441
R20338 VDD.n3426 VDD.n3425 0.753441
R20339 VDD.n3443 VDD.n3442 0.753441
R20340 VDD.n3460 VDD.n3459 0.753441
R20341 VDD.n3390 VDD.n3389 0.753441
R20342 VDD.n3384 VDD.n3383 0.753441
R20343 VDD.n3374 VDD.n3297 0.753441
R20344 VDD.n3863 VDD.n3810 0.753441
R20345 VDD.n3872 VDD.n3104 0.753441
R20346 VDD.n2923 VDD.n2922 0.753441
R20347 VDD.n2522 VDD.n2521 0.753441
R20348 VDD.n2531 VDD.n2513 0.753441
R20349 VDD.n2355 VDD.n2354 0.753441
R20350 VDD.n3071 VDD.n2286 0.753441
R20351 VDD.n2753 VDD.n2752 0.753441
R20352 VDD.n2644 VDD.n2643 0.753441
R20353 VDD.n2688 VDD.n2687 0.753441
R20354 VDD.n2679 VDD.n2678 0.753441
R20355 VDD.n2331 VDD.n2306 0.753441
R20356 VDD.n2062 VDD.n2061 0.753441
R20357 VDD.n2037 VDD.n1553 0.753441
R20358 VDD.n1983 VDD.n1982 0.753441
R20359 VDD.n1867 VDD.n1866 0.753441
R20360 VDD.n1845 VDD.n1606 0.753441
R20361 VDD.n1709 VDD.n1708 0.753441
R20362 VDD.n2153 VDD.n2130 0.753441
R20363 VDD.n2258 VDD.n2257 0.753441
R20364 VDD.n2242 VDD.n2241 0.753441
R20365 VDD.n2215 VDD.n2214 0.753441
R20366 VDD.n1037 VDD.n1036 0.753441
R20367 VDD.n1045 VDD.n1018 0.753441
R20368 VDD.n991 VDD.n990 0.753441
R20369 VDD.n980 VDD.n979 0.753441
R20370 VDD.n960 VDD.n959 0.753441
R20371 VDD.n901 VDD.n847 0.753441
R20372 VDD.n913 VDD.n895 0.753441
R20373 VDD.n922 VDD.n890 0.753441
R20374 VDD.n947 VDD.n848 0.753441
R20375 VDD.n869 VDD.n853 0.753441
R20376 VDD.n865 VDD.n856 0.753441
R20377 VDD.n1333 VDD.n1332 0.753441
R20378 VDD.n1326 VDD.n727 0.753441
R20379 VDD.n1210 VDD.n1209 0.753441
R20380 VDD.n1177 VDD.n1176 0.753441
R20381 VDD.n1392 VDD.n1362 0.753441
R20382 VDD.n1477 VDD.n1476 0.753441
R20383 VDD.n1420 VDD.n1418 0.753441
R20384 VDD.n156 VDD.n155 0.745692
R20385 VDD.n621 VDD.n617 0.732469
R20386 VDD.n538 VDD.n534 0.732469
R20387 VDD.n458 VDD.n454 0.732469
R20388 VDD.n2888 VDD.n2887 0.731929
R20389 VDD.n2848 VDD.n2847 0.731929
R20390 VDD.n1828 VDD.n1827 0.731929
R20391 VDD.n4441 VDD.n4440 0.644287
R20392 VDD.n4413 VDD.n4050 0.644287
R20393 VDD.n60 VDD.n59 0.6405
R20394 VDD.n23 VDD.n22 0.6405
R20395 VDD.n1885 VDD.n1884 0.635211
R20396 VDD.n1900 VDD.n1899 0.635211
R20397 VDD.n292 VDD.n291 0.622722
R20398 VDD.n138 VDD.n137 0.614477
R20399 VDD.n26 VDD.n10 0.600153
R20400 VDD.n62 VDD.n61 0.599785
R20401 VDD.n3360 VDD.n3359 0.597116
R20402 VDD.n151 VDD.n150 0.590759
R20403 VDD.n1262 VDD.n1261 0.539826
R20404 VDD.n290 VDD.n289 0.519731
R20405 VDD.n1244 VDD.n1243 0.508436
R20406 VDD.n662 VDD.n661 0.508344
R20407 VDD.n576 VDD.n568 0.508344
R20408 VDD.n496 VDD.n488 0.508344
R20409 VDD.n289 VDD.n210 0.491846
R20410 VDD.n335 VDD.n334 0.488781
R20411 VDD.n212 VDD.n197 0.481269
R20412 VDD.n9 VDD.n8 0.442135
R20413 VDD.n403 VDD.n402 0.438
R20414 VDD.n694 VDD.n693 0.430246
R20415 VDD.n337 VDD.n336 0.393625
R20416 VDD.n61 VDD.n60 0.388
R20417 VDD.n23 VDD.n10 0.388
R20418 VDD.n153 VDD.n151 0.383913
R20419 VDD.n4372 VDD.n4371 0.376971
R20420 VDD.n4292 VDD.n4291 0.376971
R20421 VDD.n4265 VDD.n4264 0.376971
R20422 VDD.n3943 VDD.n3927 0.376971
R20423 VDD.n2984 VDD.n2983 0.376971
R20424 VDD.n2058 VDD.n2057 0.376971
R20425 VDD.n1866 VDD.n1865 0.376971
R20426 VDD.n2084 VDD.n1528 0.376971
R20427 VDD.n2251 VDD.n1515 0.376971
R20428 VDD.n1102 VDD.n1101 0.376971
R20429 VDD.n1060 VDD.n1059 0.376971
R20430 VDD.n999 VDD.n823 0.376971
R20431 VDD.n936 VDD.n883 0.376971
R20432 VDD.n1327 VDD.n1326 0.376971
R20433 VDD.n1290 VDD.n1289 0.376971
R20434 VDD.n1153 VDD.n1151 0.376971
R20435 VDD.n624 VDD.n616 0.376971
R20436 VDD.n689 VDD.n688 0.376971
R20437 VDD.n673 VDD.n651 0.376971
R20438 VDD.n541 VDD.n533 0.376971
R20439 VDD.n601 VDD.n600 0.376971
R20440 VDD.n587 VDD.n586 0.376971
R20441 VDD.n461 VDD.n453 0.376971
R20442 VDD.n521 VDD.n520 0.376971
R20443 VDD.n507 VDD.n506 0.376971
R20444 VDD.n2905 VDD.n2904 0.366214
R20445 VDD.n154 VDD.n153 0.359875
R20446 VDD.n4422 VDD.n4421 0.356056
R20447 VDD.n3914 VDD.n3909 0.35457
R20448 VDD.n3966 VDD.n3914 0.354142
R20449 VDD.n284 VDD.n214 0.3505
R20450 VDD.n261 VDD.n260 0.3505
R20451 VDD.n281 VDD.n280 0.3505
R20452 VDD.n257 VDD.n218 0.3505
R20453 VDD.n277 VDD.n211 0.3505
R20454 VDD.n264 VDD.n219 0.3505
R20455 VDD.n158 VDD.n157 0.342872
R20456 VDD.n285 VDD.n284 0.338
R20457 VDD.n273 VDD.n214 0.338
R20458 VDD.n273 VDD.n272 0.338
R20459 VDD.n272 VDD.n217 0.338
R20460 VDD.n261 VDD.n217 0.338
R20461 VDD.n260 VDD.n220 0.338
R20462 VDD.n249 VDD.n220 0.338
R20463 VDD.n281 VDD.n213 0.338
R20464 VDD.n280 VDD.n215 0.338
R20465 VDD.n269 VDD.n215 0.338
R20466 VDD.n269 VDD.n268 0.338
R20467 VDD.n268 VDD.n218 0.338
R20468 VDD.n257 VDD.n256 0.338
R20469 VDD.n256 VDD.n221 0.338
R20470 VDD.n247 VDD.n221 0.338
R20471 VDD.n288 VDD.n211 0.338
R20472 VDD.n277 VDD.n276 0.338
R20473 VDD.n276 VDD.n216 0.338
R20474 VDD.n265 VDD.n216 0.338
R20475 VDD.n265 VDD.n264 0.338
R20476 VDD.n253 VDD.n219 0.338
R20477 VDD.n253 VDD.n252 0.338
R20478 VDD.n291 VDD.n290 0.332643
R20479 VDD.n3791 VDD.n3789 0.323189
R20480 VDD.n2806 VDD.n2805 0.323189
R20481 VDD.n4023 VDD.n4022 0.318972
R20482 VDD.n1503 VDD.n695 0.316225
R20483 VDD.n4660 VDD.n4659 0.305262
R20484 VDD.n4653 VDD.n3907 0.305262
R20485 VDD.n4479 VDD.n4448 0.305262
R20486 VDD.n4423 VDD.n4422 0.305262
R20487 VDD.n4381 VDD.n4380 0.305262
R20488 VDD.n4388 VDD.n4068 0.305262
R20489 VDD.n4316 VDD.n4315 0.305262
R20490 VDD.n4309 VDD.n4284 0.305262
R20491 VDD.n4210 VDD.n4128 0.305262
R20492 VDD.n4225 VDD.n4224 0.305262
R20493 VDD.n3962 VDD.n3961 0.305262
R20494 VDD.n3672 VDD.n3671 0.305262
R20495 VDD.n3679 VDD.n3201 0.305262
R20496 VDD.n3360 VDD.n3357 0.305262
R20497 VDD.n3832 VDD.n3831 0.305262
R20498 VDD.n3886 VDD.n3885 0.305262
R20499 VDD.n3165 VDD.n3164 0.305262
R20500 VDD.n3152 VDD.n3125 0.305262
R20501 VDD.n2550 VDD.n2549 0.305262
R20502 VDD.n3052 VDD.n3009 0.305262
R20503 VDD.n3044 VDD.n3043 0.305262
R20504 VDD.n3022 VDD.n3020 0.305262
R20505 VDD.n3036 VDD.n3023 0.305262
R20506 VDD.n2761 VDD.n2760 0.305262
R20507 VDD.n2338 VDD.n2300 0.305262
R20508 VDD.n1912 VDD.n1574 0.305262
R20509 VDD.n1918 VDD.n1572 0.305262
R20510 VDD.n1923 VDD.n1570 0.305262
R20511 VDD.n1267 VDD.n1266 0.305262
R20512 VDD.n1268 VDD.n755 0.305262
R20513 VDD.n1273 VDD.n1272 0.305262
R20514 VDD.n1239 VDD.n1238 0.305262
R20515 VDD.n1246 VDD.n1245 0.305262
R20516 VDD.n693 VDD.n605 0.301853
R20517 VDD.n409 VDD.n408 0.3005
R20518 VDD.n2346 VDD.n2293 0.298074
R20519 VDD.n1889 VDD.n1888 0.298074
R20520 VDD.n4411 VDD.n4047 0.29768
R20521 VDD.n4417 VDD.n4047 0.29768
R20522 VDD.n4487 VDD.n4486 0.29768
R20523 VDD.n4486 VDD.n4485 0.29768
R20524 VDD.n3351 VDD.n3350 0.29768
R20525 VDD.n3352 VDD.n3351 0.29768
R20526 VDD.n3167 VDD.n3166 0.29768
R20527 VDD.n3168 VDD.n3167 0.29768
R20528 VDD.n2346 VDD.n2345 0.297291
R20529 VDD.n1890 VDD.n1889 0.297291
R20530 VDD.n3961 VDD.n3960 0.281745
R20531 VDD.n3050 VDD.n3012 0.278761
R20532 VDD.n187 VDD.n186 0.278
R20533 VDD.n2764 VDD.n2448 0.254468
R20534 VDD.n2856 VDD.n2855 0.25148
R20535 VDD.n3045 VDD.n3016 0.25148
R20536 VDD.n2913 VDD.n2405 0.246654
R20537 VDD.n155 VDD.n144 0.243729
R20538 VDD.n4346 VDD.n4345 0.239726
R20539 VDD.n4067 VDD.n4063 0.239726
R20540 VDD.n4532 VDD.n4531 0.239726
R20541 VDD.n4553 VDD.n4003 0.239726
R20542 VDD.n4624 VDD.n4605 0.239726
R20543 VDD.n3344 VDD.n3318 0.239726
R20544 VDD.n2572 VDD.n2568 0.239726
R20545 VDD.n1913 VDD.n1575 0.239726
R20546 VDD.n2067 VDD.n2066 0.239726
R20547 VDD.n1873 VDD.n1592 0.239726
R20548 VDD.n4345 VDD.n4344 0.239381
R20549 VDD.n4392 VDD.n4067 0.239381
R20550 VDD.n4531 VDD.n4530 0.239381
R20551 VDD.n4546 VDD.n4003 0.239381
R20552 VDD.n4631 VDD.n4605 0.239381
R20553 VDD.n3340 VDD.n3318 0.239381
R20554 VDD.n2590 VDD.n2572 0.239381
R20555 VDD.n1874 VDD.n1873 0.239381
R20556 VDD.n1905 VDD.n1575 0.239381
R20557 VDD.n2066 VDD.n2065 0.239381
R20558 VDD.n3049 VDD.n3013 0.229071
R20559 VDD.n694 VDD.n444 0.227798
R20560 VDD.n401 VDD.n397 0.21925
R20561 VDD.n1257 VDD.n1256 0.21623
R20562 VDD.n695 VDD.n694 0.213625
R20563 VDD.n86 VDD.n85 0.209465
R20564 VDD.n3306 VDD.n3305 0.203675
R20565 VDD.n2499 VDD.n2497 0.203675
R20566 VDD.n407 VDD.n338 0.203144
R20567 VDD.n155 VDD.n100 0.202674
R20568 VDD.n210 VDD.n209 0.184982
R20569 VDD.n1767 VDD.n1649 0.180304
R20570 VDD.n1768 VDD.n1767 0.180304
R20571 VDD.n2010 VDD.n1959 0.180304
R20572 VDD.n2010 VDD.n2009 0.180304
R20573 VDD.n2154 VDD.n2131 0.180304
R20574 VDD.n2150 VDD.n2131 0.180304
R20575 VDD.n408 VDD.n405 0.168469
R20576 VDD.n2766 VDD.n2765 0.152881
R20577 VDD.n4678 VDD.n3893 0.15002
R20578 VDD.n3893 VDD.n3090 0.15002
R20579 VDD.n3090 VDD.n2274 0.15002
R20580 VDD.n2274 VDD.n1503 0.15002
R20581 VDD.n181 VDD.n180 0.148119
R20582 VDD.n1265 VDD.n757 0.14432
R20583 VDD.n248 VDD.n222 0.142484
R20584 VDD.n251 VDD.n250 0.142484
R20585 VDD.n255 VDD.n254 0.142484
R20586 VDD.n259 VDD.n258 0.142484
R20587 VDD.n263 VDD.n262 0.142484
R20588 VDD.n267 VDD.n266 0.142484
R20589 VDD.n271 VDD.n270 0.142484
R20590 VDD.n275 VDD.n274 0.142484
R20591 VDD.n279 VDD.n278 0.142484
R20592 VDD.n283 VDD.n282 0.142484
R20593 VDD.n287 VDD.n286 0.142484
R20594 VDD.n159 VDD.n158 0.141672
R20595 VDD.n45 VDD.n9 0.127382
R20596 VDD.n53 VDD.n47 0.122868
R20597 VDD.n16 VDD.n11 0.122868
R20598 VDD.n7 VDD.n6 0.120751
R20599 VDD.n84 VDD.n83 0.120751
R20600 VDD.n4173 VDD.n4172 0.120292
R20601 VDD.n4174 VDD.n4173 0.120292
R20602 VDD.n4174 VDD.n4158 0.120292
R20603 VDD.n4158 VDD.n4157 0.120292
R20604 VDD.n4157 VDD.n4154 0.120292
R20605 VDD.n4154 VDD.n4153 0.120292
R20606 VDD.n4153 VDD.n4150 0.120292
R20607 VDD.n4150 VDD.n4148 0.120292
R20608 VDD.n4148 VDD.n4146 0.120292
R20609 VDD.n4184 VDD.n4146 0.120292
R20610 VDD.n4185 VDD.n4184 0.120292
R20611 VDD.n4186 VDD.n4185 0.120292
R20612 VDD.n4186 VDD.n4143 0.120292
R20613 VDD.n4143 VDD.n4142 0.120292
R20614 VDD.n4142 VDD.n4140 0.120292
R20615 VDD.n4192 VDD.n4140 0.120292
R20616 VDD.n4193 VDD.n4192 0.120292
R20617 VDD.n4193 VDD.n4137 0.120292
R20618 VDD.n4137 VDD.n4136 0.120292
R20619 VDD.n4200 VDD.n4136 0.120292
R20620 VDD.n4201 VDD.n4200 0.120292
R20621 VDD.n4201 VDD.n4133 0.120292
R20622 VDD.n4205 VDD.n4133 0.120292
R20623 VDD.n4206 VDD.n4205 0.120292
R20624 VDD.n4206 VDD.n4129 0.120292
R20625 VDD.n4211 VDD.n4129 0.120292
R20626 VDD.n4212 VDD.n4211 0.120292
R20627 VDD.n4212 VDD.n4127 0.120292
R20628 VDD.n4218 VDD.n4127 0.120292
R20629 VDD.n4219 VDD.n4218 0.120292
R20630 VDD.n4220 VDD.n4219 0.120292
R20631 VDD.n4220 VDD.n4124 0.120292
R20632 VDD.n4226 VDD.n4124 0.120292
R20633 VDD.n4227 VDD.n4226 0.120292
R20634 VDD.n4228 VDD.n4227 0.120292
R20635 VDD.n4228 VDD.n4122 0.120292
R20636 VDD.n4122 VDD.n4119 0.120292
R20637 VDD.n4233 VDD.n4119 0.120292
R20638 VDD.n4234 VDD.n4233 0.120292
R20639 VDD.n4235 VDD.n4234 0.120292
R20640 VDD.n4235 VDD.n4116 0.120292
R20641 VDD.n4239 VDD.n4116 0.120292
R20642 VDD.n4240 VDD.n4239 0.120292
R20643 VDD.n4241 VDD.n4240 0.120292
R20644 VDD.n4241 VDD.n4113 0.120292
R20645 VDD.n4113 VDD.n4111 0.120292
R20646 VDD.n4246 VDD.n4111 0.120292
R20647 VDD.n4247 VDD.n4246 0.120292
R20648 VDD.n4248 VDD.n4247 0.120292
R20649 VDD.n4248 VDD.n4108 0.120292
R20650 VDD.n4108 VDD.n4105 0.120292
R20651 VDD.n4253 VDD.n4105 0.120292
R20652 VDD.n4254 VDD.n4253 0.120292
R20653 VDD.n4255 VDD.n4254 0.120292
R20654 VDD.n4255 VDD.n4101 0.120292
R20655 VDD.n4259 VDD.n4101 0.120292
R20656 VDD.n4260 VDD.n4259 0.120292
R20657 VDD.n4261 VDD.n4260 0.120292
R20658 VDD.n4261 VDD.n4097 0.120292
R20659 VDD.n4267 VDD.n4097 0.120292
R20660 VDD.n4268 VDD.n4267 0.120292
R20661 VDD.n4339 VDD.n4268 0.120292
R20662 VDD.n4339 VDD.n4338 0.120292
R20663 VDD.n4338 VDD.n4337 0.120292
R20664 VDD.n4337 VDD.n4269 0.120292
R20665 VDD.n4333 VDD.n4269 0.120292
R20666 VDD.n4333 VDD.n4332 0.120292
R20667 VDD.n4332 VDD.n4271 0.120292
R20668 VDD.n4326 VDD.n4271 0.120292
R20669 VDD.n4326 VDD.n4325 0.120292
R20670 VDD.n4325 VDD.n4324 0.120292
R20671 VDD.n4324 VDD.n4275 0.120292
R20672 VDD.n4320 VDD.n4275 0.120292
R20673 VDD.n4320 VDD.n4319 0.120292
R20674 VDD.n4319 VDD.n4318 0.120292
R20675 VDD.n4318 VDD.n4277 0.120292
R20676 VDD.n4312 VDD.n4277 0.120292
R20677 VDD.n4312 VDD.n4311 0.120292
R20678 VDD.n4311 VDD.n4310 0.120292
R20679 VDD.n4310 VDD.n4283 0.120292
R20680 VDD.n4304 VDD.n4283 0.120292
R20681 VDD.n4304 VDD.n4303 0.120292
R20682 VDD.n4303 VDD.n4302 0.120292
R20683 VDD.n4302 VDD.n4287 0.120292
R20684 VDD.n4297 VDD.n4287 0.120292
R20685 VDD.n4297 VDD.n4296 0.120292
R20686 VDD.n4296 VDD.n4295 0.120292
R20687 VDD.n4295 VDD.n4289 0.120292
R20688 VDD.n4289 VDD.n4093 0.120292
R20689 VDD.n4344 VDD.n4093 0.120292
R20690 VDD.n4346 VDD.n4086 0.120292
R20691 VDD.n4350 VDD.n4086 0.120292
R20692 VDD.n4351 VDD.n4350 0.120292
R20693 VDD.n4352 VDD.n4351 0.120292
R20694 VDD.n4352 VDD.n4083 0.120292
R20695 VDD.n4083 VDD.n4080 0.120292
R20696 VDD.n4361 VDD.n4080 0.120292
R20697 VDD.n4362 VDD.n4361 0.120292
R20698 VDD.n4363 VDD.n4362 0.120292
R20699 VDD.n4363 VDD.n4078 0.120292
R20700 VDD.n4368 VDD.n4078 0.120292
R20701 VDD.n4369 VDD.n4368 0.120292
R20702 VDD.n4370 VDD.n4369 0.120292
R20703 VDD.n4370 VDD.n4075 0.120292
R20704 VDD.n4376 VDD.n4075 0.120292
R20705 VDD.n4377 VDD.n4376 0.120292
R20706 VDD.n4378 VDD.n4377 0.120292
R20707 VDD.n4378 VDD.n4073 0.120292
R20708 VDD.n4383 VDD.n4073 0.120292
R20709 VDD.n4384 VDD.n4383 0.120292
R20710 VDD.n4384 VDD.n4070 0.120292
R20711 VDD.n4390 VDD.n4070 0.120292
R20712 VDD.n4391 VDD.n4390 0.120292
R20713 VDD.n4392 VDD.n4391 0.120292
R20714 VDD.n4063 VDD.n4061 0.120292
R20715 VDD.n4061 VDD.n4060 0.120292
R20716 VDD.n4060 VDD.n4056 0.120292
R20717 VDD.n4402 VDD.n4056 0.120292
R20718 VDD.n4403 VDD.n4402 0.120292
R20719 VDD.n4404 VDD.n4403 0.120292
R20720 VDD.n4404 VDD.n4054 0.120292
R20721 VDD.n4054 VDD.n4052 0.120292
R20722 VDD.n4410 VDD.n4052 0.120292
R20723 VDD.n4411 VDD.n4410 0.120292
R20724 VDD.n4418 VDD.n4417 0.120292
R20725 VDD.n4419 VDD.n4418 0.120292
R20726 VDD.n4419 VDD.n4044 0.120292
R20727 VDD.n4426 VDD.n4044 0.120292
R20728 VDD.n4427 VDD.n4426 0.120292
R20729 VDD.n4427 VDD.n4041 0.120292
R20730 VDD.n4433 VDD.n4041 0.120292
R20731 VDD.n4434 VDD.n4433 0.120292
R20732 VDD.n4500 VDD.n4434 0.120292
R20733 VDD.n4500 VDD.n4499 0.120292
R20734 VDD.n4499 VDD.n4498 0.120292
R20735 VDD.n4498 VDD.n4435 0.120292
R20736 VDD.n4493 VDD.n4435 0.120292
R20737 VDD.n4493 VDD.n4492 0.120292
R20738 VDD.n4492 VDD.n4438 0.120292
R20739 VDD.n4487 VDD.n4438 0.120292
R20740 VDD.n4485 VDD.n4442 0.120292
R20741 VDD.n4481 VDD.n4442 0.120292
R20742 VDD.n4481 VDD.n4480 0.120292
R20743 VDD.n4480 VDD.n4447 0.120292
R20744 VDD.n4474 VDD.n4447 0.120292
R20745 VDD.n4474 VDD.n4473 0.120292
R20746 VDD.n4473 VDD.n4451 0.120292
R20747 VDD.n4468 VDD.n4451 0.120292
R20748 VDD.n4468 VDD.n4467 0.120292
R20749 VDD.n4467 VDD.n4466 0.120292
R20750 VDD.n4466 VDD.n4453 0.120292
R20751 VDD.n4461 VDD.n4453 0.120292
R20752 VDD.n4461 VDD.n4460 0.120292
R20753 VDD.n4460 VDD.n4459 0.120292
R20754 VDD.n4459 VDD.n4456 0.120292
R20755 VDD.n4456 VDD.n4036 0.120292
R20756 VDD.n4507 VDD.n4036 0.120292
R20757 VDD.n4508 VDD.n4507 0.120292
R20758 VDD.n4509 VDD.n4508 0.120292
R20759 VDD.n4509 VDD.n4034 0.120292
R20760 VDD.n4034 VDD.n4033 0.120292
R20761 VDD.n4516 VDD.n4033 0.120292
R20762 VDD.n4517 VDD.n4516 0.120292
R20763 VDD.n4518 VDD.n4517 0.120292
R20764 VDD.n4518 VDD.n4031 0.120292
R20765 VDD.n4522 VDD.n4031 0.120292
R20766 VDD.n4523 VDD.n4522 0.120292
R20767 VDD.n4523 VDD.n4027 0.120292
R20768 VDD.n4027 VDD.n4026 0.120292
R20769 VDD.n4026 VDD.n4024 0.120292
R20770 VDD.n4530 VDD.n4024 0.120292
R20771 VDD.n4533 VDD.n4532 0.120292
R20772 VDD.n4533 VDD.n4015 0.120292
R20773 VDD.n4538 VDD.n4015 0.120292
R20774 VDD.n4539 VDD.n4538 0.120292
R20775 VDD.n4540 VDD.n4539 0.120292
R20776 VDD.n4540 VDD.n4011 0.120292
R20777 VDD.n4544 VDD.n4011 0.120292
R20778 VDD.n4545 VDD.n4544 0.120292
R20779 VDD.n4546 VDD.n4545 0.120292
R20780 VDD.n4554 VDD.n4553 0.120292
R20781 VDD.n4555 VDD.n4554 0.120292
R20782 VDD.n4555 VDD.n4001 0.120292
R20783 VDD.n4001 VDD.n3999 0.120292
R20784 VDD.n4561 VDD.n3999 0.120292
R20785 VDD.n4562 VDD.n4561 0.120292
R20786 VDD.n4563 VDD.n4562 0.120292
R20787 VDD.n4563 VDD.n3996 0.120292
R20788 VDD.n3996 VDD.n3995 0.120292
R20789 VDD.n4571 VDD.n3995 0.120292
R20790 VDD.n4572 VDD.n4571 0.120292
R20791 VDD.n4573 VDD.n4572 0.120292
R20792 VDD.n4573 VDD.n3992 0.120292
R20793 VDD.n4578 VDD.n3992 0.120292
R20794 VDD.n4579 VDD.n4578 0.120292
R20795 VDD.n4580 VDD.n4579 0.120292
R20796 VDD.n4580 VDD.n3988 0.120292
R20797 VDD.n4585 VDD.n3988 0.120292
R20798 VDD.n4586 VDD.n4585 0.120292
R20799 VDD.n4587 VDD.n4586 0.120292
R20800 VDD.n4587 VDD.n3986 0.120292
R20801 VDD.n4593 VDD.n3986 0.120292
R20802 VDD.n4594 VDD.n4593 0.120292
R20803 VDD.n4648 VDD.n4594 0.120292
R20804 VDD.n4648 VDD.n4647 0.120292
R20805 VDD.n4647 VDD.n4646 0.120292
R20806 VDD.n4646 VDD.n4595 0.120292
R20807 VDD.n4640 VDD.n4595 0.120292
R20808 VDD.n4640 VDD.n4639 0.120292
R20809 VDD.n4639 VDD.n4602 0.120292
R20810 VDD.n4633 VDD.n4602 0.120292
R20811 VDD.n4633 VDD.n4632 0.120292
R20812 VDD.n4632 VDD.n4631 0.120292
R20813 VDD.n4624 VDD.n4623 0.120292
R20814 VDD.n4623 VDD.n4622 0.120292
R20815 VDD.n4622 VDD.n4607 0.120292
R20816 VDD.n4617 VDD.n4607 0.120292
R20817 VDD.n4617 VDD.n4616 0.120292
R20818 VDD.n4616 VDD.n4615 0.120292
R20819 VDD.n4662 VDD.n4661 0.120292
R20820 VDD.n4661 VDD.n3903 0.120292
R20821 VDD.n4655 VDD.n3903 0.120292
R20822 VDD.n4655 VDD.n4654 0.120292
R20823 VDD.n4654 VDD.n3906 0.120292
R20824 VDD.n3981 VDD.n3906 0.120292
R20825 VDD.n3981 VDD.n3980 0.120292
R20826 VDD.n3980 VDD.n3979 0.120292
R20827 VDD.n3979 VDD.n3909 0.120292
R20828 VDD.n3966 VDD.n3965 0.120292
R20829 VDD.n3965 VDD.n3964 0.120292
R20830 VDD.n3964 VDD.n3917 0.120292
R20831 VDD.n3957 VDD.n3917 0.120292
R20832 VDD.n3957 VDD.n3956 0.120292
R20833 VDD.n3956 VDD.n3955 0.120292
R20834 VDD.n3955 VDD.n3920 0.120292
R20835 VDD.n3951 VDD.n3920 0.120292
R20836 VDD.n3951 VDD.n3950 0.120292
R20837 VDD.n3950 VDD.n3949 0.120292
R20838 VDD.n3949 VDD.n3924 0.120292
R20839 VDD.n3945 VDD.n3924 0.120292
R20840 VDD.n3945 VDD.n3944 0.120292
R20841 VDD.n3944 VDD.n3928 0.120292
R20842 VDD.n3938 VDD.n3928 0.120292
R20843 VDD.n3339 VDD.n3338 0.120292
R20844 VDD.n3340 VDD.n3339 0.120292
R20845 VDD.n3345 VDD.n3344 0.120292
R20846 VDD.n3346 VDD.n3345 0.120292
R20847 VDD.n3346 VDD.n3314 0.120292
R20848 VDD.n3350 VDD.n3314 0.120292
R20849 VDD.n3353 VDD.n3352 0.120292
R20850 VDD.n3353 VDD.n3304 0.120292
R20851 VDD.n3361 VDD.n3304 0.120292
R20852 VDD.n3362 VDD.n3361 0.120292
R20853 VDD.n3363 VDD.n3362 0.120292
R20854 VDD.n3363 VDD.n3301 0.120292
R20855 VDD.n3368 VDD.n3301 0.120292
R20856 VDD.n3369 VDD.n3368 0.120292
R20857 VDD.n3370 VDD.n3369 0.120292
R20858 VDD.n3370 VDD.n3298 0.120292
R20859 VDD.n3375 VDD.n3298 0.120292
R20860 VDD.n3376 VDD.n3375 0.120292
R20861 VDD.n3376 VDD.n3295 0.120292
R20862 VDD.n3381 VDD.n3295 0.120292
R20863 VDD.n3382 VDD.n3381 0.120292
R20864 VDD.n3382 VDD.n3293 0.120292
R20865 VDD.n3391 VDD.n3293 0.120292
R20866 VDD.n3392 VDD.n3391 0.120292
R20867 VDD.n3465 VDD.n3392 0.120292
R20868 VDD.n3465 VDD.n3464 0.120292
R20869 VDD.n3464 VDD.n3463 0.120292
R20870 VDD.n3463 VDD.n3393 0.120292
R20871 VDD.n3457 VDD.n3393 0.120292
R20872 VDD.n3457 VDD.n3456 0.120292
R20873 VDD.n3456 VDD.n3397 0.120292
R20874 VDD.n3451 VDD.n3397 0.120292
R20875 VDD.n3451 VDD.n3450 0.120292
R20876 VDD.n3450 VDD.n3449 0.120292
R20877 VDD.n3449 VDD.n3399 0.120292
R20878 VDD.n3445 VDD.n3399 0.120292
R20879 VDD.n3445 VDD.n3444 0.120292
R20880 VDD.n3444 VDD.n3402 0.120292
R20881 VDD.n3439 VDD.n3402 0.120292
R20882 VDD.n3439 VDD.n3438 0.120292
R20883 VDD.n3438 VDD.n3437 0.120292
R20884 VDD.n3437 VDD.n3405 0.120292
R20885 VDD.n3432 VDD.n3405 0.120292
R20886 VDD.n3432 VDD.n3431 0.120292
R20887 VDD.n3431 VDD.n3430 0.120292
R20888 VDD.n3430 VDD.n3410 0.120292
R20889 VDD.n3424 VDD.n3410 0.120292
R20890 VDD.n3424 VDD.n3423 0.120292
R20891 VDD.n3423 VDD.n3422 0.120292
R20892 VDD.n3422 VDD.n3412 0.120292
R20893 VDD.n3417 VDD.n3412 0.120292
R20894 VDD.n3417 VDD.n3416 0.120292
R20895 VDD.n3416 VDD.n3289 0.120292
R20896 VDD.n3472 VDD.n3289 0.120292
R20897 VDD.n3473 VDD.n3472 0.120292
R20898 VDD.n3474 VDD.n3473 0.120292
R20899 VDD.n3474 VDD.n3285 0.120292
R20900 VDD.n3480 VDD.n3285 0.120292
R20901 VDD.n3481 VDD.n3480 0.120292
R20902 VDD.n3481 VDD.n3282 0.120292
R20903 VDD.n3282 VDD.n3279 0.120292
R20904 VDD.n3487 VDD.n3279 0.120292
R20905 VDD.n3488 VDD.n3487 0.120292
R20906 VDD.n3488 VDD.n3275 0.120292
R20907 VDD.n3494 VDD.n3275 0.120292
R20908 VDD.n3495 VDD.n3494 0.120292
R20909 VDD.n3495 VDD.n3271 0.120292
R20910 VDD.n3500 VDD.n3271 0.120292
R20911 VDD.n3501 VDD.n3500 0.120292
R20912 VDD.n3502 VDD.n3501 0.120292
R20913 VDD.n3502 VDD.n3266 0.120292
R20914 VDD.n3506 VDD.n3266 0.120292
R20915 VDD.n3507 VDD.n3506 0.120292
R20916 VDD.n3508 VDD.n3507 0.120292
R20917 VDD.n3508 VDD.n3263 0.120292
R20918 VDD.n3514 VDD.n3263 0.120292
R20919 VDD.n3515 VDD.n3514 0.120292
R20920 VDD.n3515 VDD.n3261 0.120292
R20921 VDD.n3261 VDD.n3259 0.120292
R20922 VDD.n3520 VDD.n3259 0.120292
R20923 VDD.n3521 VDD.n3520 0.120292
R20924 VDD.n3522 VDD.n3521 0.120292
R20925 VDD.n3522 VDD.n3256 0.120292
R20926 VDD.n3530 VDD.n3256 0.120292
R20927 VDD.n3531 VDD.n3530 0.120292
R20928 VDD.n3532 VDD.n3531 0.120292
R20929 VDD.n3532 VDD.n3254 0.120292
R20930 VDD.n3536 VDD.n3254 0.120292
R20931 VDD.n3537 VDD.n3536 0.120292
R20932 VDD.n3537 VDD.n3250 0.120292
R20933 VDD.n3542 VDD.n3250 0.120292
R20934 VDD.n3543 VDD.n3542 0.120292
R20935 VDD.n3544 VDD.n3543 0.120292
R20936 VDD.n3544 VDD.n3246 0.120292
R20937 VDD.n3246 VDD.n3244 0.120292
R20938 VDD.n3549 VDD.n3244 0.120292
R20939 VDD.n3550 VDD.n3549 0.120292
R20940 VDD.n3550 VDD.n3240 0.120292
R20941 VDD.n3554 VDD.n3240 0.120292
R20942 VDD.n3555 VDD.n3554 0.120292
R20943 VDD.n3556 VDD.n3555 0.120292
R20944 VDD.n3556 VDD.n3236 0.120292
R20945 VDD.n3236 VDD.n3235 0.120292
R20946 VDD.n3562 VDD.n3235 0.120292
R20947 VDD.n3563 VDD.n3562 0.120292
R20948 VDD.n3563 VDD.n3230 0.120292
R20949 VDD.n3567 VDD.n3230 0.120292
R20950 VDD.n3568 VDD.n3567 0.120292
R20951 VDD.n3632 VDD.n3568 0.120292
R20952 VDD.n3632 VDD.n3631 0.120292
R20953 VDD.n3631 VDD.n3630 0.120292
R20954 VDD.n3630 VDD.n3569 0.120292
R20955 VDD.n3626 VDD.n3569 0.120292
R20956 VDD.n3626 VDD.n3625 0.120292
R20957 VDD.n3625 VDD.n3624 0.120292
R20958 VDD.n3624 VDD.n3572 0.120292
R20959 VDD.n3619 VDD.n3572 0.120292
R20960 VDD.n3619 VDD.n3618 0.120292
R20961 VDD.n3618 VDD.n3617 0.120292
R20962 VDD.n3617 VDD.n3576 0.120292
R20963 VDD.n3612 VDD.n3576 0.120292
R20964 VDD.n3612 VDD.n3611 0.120292
R20965 VDD.n3611 VDD.n3610 0.120292
R20966 VDD.n3610 VDD.n3580 0.120292
R20967 VDD.n3606 VDD.n3580 0.120292
R20968 VDD.n3606 VDD.n3605 0.120292
R20969 VDD.n3605 VDD.n3604 0.120292
R20970 VDD.n3604 VDD.n3582 0.120292
R20971 VDD.n3600 VDD.n3582 0.120292
R20972 VDD.n3600 VDD.n3599 0.120292
R20973 VDD.n3599 VDD.n3598 0.120292
R20974 VDD.n3598 VDD.n3586 0.120292
R20975 VDD.n3592 VDD.n3586 0.120292
R20976 VDD.n3592 VDD.n3591 0.120292
R20977 VDD.n3591 VDD.n3590 0.120292
R20978 VDD.n3590 VDD.n3224 0.120292
R20979 VDD.n3637 VDD.n3224 0.120292
R20980 VDD.n3638 VDD.n3637 0.120292
R20981 VDD.n3639 VDD.n3638 0.120292
R20982 VDD.n3639 VDD.n3222 0.120292
R20983 VDD.n3222 VDD.n3221 0.120292
R20984 VDD.n3221 VDD.n3220 0.120292
R20985 VDD.n3647 VDD.n3220 0.120292
R20986 VDD.n3648 VDD.n3647 0.120292
R20987 VDD.n3649 VDD.n3648 0.120292
R20988 VDD.n3649 VDD.n3218 0.120292
R20989 VDD.n3218 VDD.n3216 0.120292
R20990 VDD.n3216 VDD.n3215 0.120292
R20991 VDD.n3215 VDD.n3213 0.120292
R20992 VDD.n3213 VDD.n3211 0.120292
R20993 VDD.n3658 VDD.n3211 0.120292
R20994 VDD.n3659 VDD.n3658 0.120292
R20995 VDD.n3660 VDD.n3659 0.120292
R20996 VDD.n3660 VDD.n3208 0.120292
R20997 VDD.n3208 VDD.n3207 0.120292
R20998 VDD.n3665 VDD.n3207 0.120292
R20999 VDD.n3666 VDD.n3665 0.120292
R21000 VDD.n3666 VDD.n3204 0.120292
R21001 VDD.n3673 VDD.n3204 0.120292
R21002 VDD.n3674 VDD.n3673 0.120292
R21003 VDD.n3675 VDD.n3674 0.120292
R21004 VDD.n3675 VDD.n3202 0.120292
R21005 VDD.n3681 VDD.n3202 0.120292
R21006 VDD.n3682 VDD.n3681 0.120292
R21007 VDD.n3752 VDD.n3682 0.120292
R21008 VDD.n3752 VDD.n3751 0.120292
R21009 VDD.n3751 VDD.n3750 0.120292
R21010 VDD.n3750 VDD.n3683 0.120292
R21011 VDD.n3743 VDD.n3683 0.120292
R21012 VDD.n3743 VDD.n3742 0.120292
R21013 VDD.n3742 VDD.n3741 0.120292
R21014 VDD.n3741 VDD.n3686 0.120292
R21015 VDD.n3737 VDD.n3686 0.120292
R21016 VDD.n3737 VDD.n3736 0.120292
R21017 VDD.n3736 VDD.n3735 0.120292
R21018 VDD.n3735 VDD.n3689 0.120292
R21019 VDD.n3730 VDD.n3689 0.120292
R21020 VDD.n3730 VDD.n3729 0.120292
R21021 VDD.n3729 VDD.n3728 0.120292
R21022 VDD.n3728 VDD.n3693 0.120292
R21023 VDD.n3724 VDD.n3693 0.120292
R21024 VDD.n3724 VDD.n3723 0.120292
R21025 VDD.n3723 VDD.n3696 0.120292
R21026 VDD.n3718 VDD.n3696 0.120292
R21027 VDD.n3718 VDD.n3717 0.120292
R21028 VDD.n3717 VDD.n3699 0.120292
R21029 VDD.n3713 VDD.n3699 0.120292
R21030 VDD.n3713 VDD.n3712 0.120292
R21031 VDD.n3712 VDD.n3711 0.120292
R21032 VDD.n3711 VDD.n3702 0.120292
R21033 VDD.n3706 VDD.n3702 0.120292
R21034 VDD.n3706 VDD.n3705 0.120292
R21035 VDD.n3705 VDD.n3198 0.120292
R21036 VDD.n3758 VDD.n3198 0.120292
R21037 VDD.n3759 VDD.n3758 0.120292
R21038 VDD.n3760 VDD.n3759 0.120292
R21039 VDD.n3760 VDD.n3196 0.120292
R21040 VDD.n3765 VDD.n3196 0.120292
R21041 VDD.n3766 VDD.n3765 0.120292
R21042 VDD.n3766 VDD.n3194 0.120292
R21043 VDD.n3771 VDD.n3194 0.120292
R21044 VDD.n3772 VDD.n3771 0.120292
R21045 VDD.n3772 VDD.n3191 0.120292
R21046 VDD.n3777 VDD.n3191 0.120292
R21047 VDD.n3778 VDD.n3777 0.120292
R21048 VDD.n3779 VDD.n3778 0.120292
R21049 VDD.n3779 VDD.n3188 0.120292
R21050 VDD.n3785 VDD.n3188 0.120292
R21051 VDD.n3786 VDD.n3785 0.120292
R21052 VDD.n3787 VDD.n3786 0.120292
R21053 VDD.n3787 VDD.n3186 0.120292
R21054 VDD.n3793 VDD.n3186 0.120292
R21055 VDD.n3794 VDD.n3793 0.120292
R21056 VDD.n3795 VDD.n3794 0.120292
R21057 VDD.n3795 VDD.n3183 0.120292
R21058 VDD.n3799 VDD.n3183 0.120292
R21059 VDD.n3800 VDD.n3799 0.120292
R21060 VDD.n3800 VDD.n3180 0.120292
R21061 VDD.n3806 VDD.n3180 0.120292
R21062 VDD.n3807 VDD.n3806 0.120292
R21063 VDD.n3808 VDD.n3807 0.120292
R21064 VDD.n3862 VDD.n3808 0.120292
R21065 VDD.n3862 VDD.n3861 0.120292
R21066 VDD.n3861 VDD.n3811 0.120292
R21067 VDD.n3857 VDD.n3811 0.120292
R21068 VDD.n3857 VDD.n3856 0.120292
R21069 VDD.n3856 VDD.n3855 0.120292
R21070 VDD.n3855 VDD.n3813 0.120292
R21071 VDD.n3849 VDD.n3813 0.120292
R21072 VDD.n3849 VDD.n3848 0.120292
R21073 VDD.n3848 VDD.n3847 0.120292
R21074 VDD.n3847 VDD.n3818 0.120292
R21075 VDD.n3842 VDD.n3818 0.120292
R21076 VDD.n3842 VDD.n3841 0.120292
R21077 VDD.n3841 VDD.n3840 0.120292
R21078 VDD.n3840 VDD.n3823 0.120292
R21079 VDD.n3836 VDD.n3823 0.120292
R21080 VDD.n3836 VDD.n3835 0.120292
R21081 VDD.n3835 VDD.n3834 0.120292
R21082 VDD.n3834 VDD.n3828 0.120292
R21083 VDD.n3877 VDD.n3876 0.120292
R21084 VDD.n3876 VDD.n3100 0.120292
R21085 VDD.n3871 VDD.n3100 0.120292
R21086 VDD.n3871 VDD.n3870 0.120292
R21087 VDD.n3870 VDD.n3105 0.120292
R21088 VDD.n3176 VDD.n3105 0.120292
R21089 VDD.n3176 VDD.n3175 0.120292
R21090 VDD.n3175 VDD.n3174 0.120292
R21091 VDD.n3174 VDD.n3107 0.120292
R21092 VDD.n3168 VDD.n3107 0.120292
R21093 VDD.n3166 VDD.n3118 0.120292
R21094 VDD.n3160 VDD.n3118 0.120292
R21095 VDD.n3160 VDD.n3159 0.120292
R21096 VDD.n3159 VDD.n3158 0.120292
R21097 VDD.n3158 VDD.n3120 0.120292
R21098 VDD.n3154 VDD.n3120 0.120292
R21099 VDD.n3154 VDD.n3153 0.120292
R21100 VDD.n3153 VDD.n3124 0.120292
R21101 VDD.n3127 VDD.n3124 0.120292
R21102 VDD.n3148 VDD.n3127 0.120292
R21103 VDD.n3148 VDD.n3147 0.120292
R21104 VDD.n3147 VDD.n3146 0.120292
R21105 VDD.n3146 VDD.n3130 0.120292
R21106 VDD.n3142 VDD.n3130 0.120292
R21107 VDD.n2589 VDD.n2588 0.120292
R21108 VDD.n2590 VDD.n2589 0.120292
R21109 VDD.n2568 VDD.n2567 0.120292
R21110 VDD.n2567 VDD.n2566 0.120292
R21111 VDD.n2566 VDD.n2496 0.120292
R21112 VDD.n2560 VDD.n2496 0.120292
R21113 VDD.n2560 VDD.n2559 0.120292
R21114 VDD.n2559 VDD.n2558 0.120292
R21115 VDD.n2558 VDD.n2498 0.120292
R21116 VDD.n2553 VDD.n2498 0.120292
R21117 VDD.n2553 VDD.n2552 0.120292
R21118 VDD.n2552 VDD.n2503 0.120292
R21119 VDD.n2547 VDD.n2503 0.120292
R21120 VDD.n2547 VDD.n2546 0.120292
R21121 VDD.n2546 VDD.n2505 0.120292
R21122 VDD.n2541 VDD.n2505 0.120292
R21123 VDD.n2541 VDD.n2540 0.120292
R21124 VDD.n2540 VDD.n2539 0.120292
R21125 VDD.n2539 VDD.n2508 0.120292
R21126 VDD.n2533 VDD.n2508 0.120292
R21127 VDD.n2533 VDD.n2532 0.120292
R21128 VDD.n2532 VDD.n2512 0.120292
R21129 VDD.n2528 VDD.n2512 0.120292
R21130 VDD.n2528 VDD.n2527 0.120292
R21131 VDD.n2527 VDD.n2526 0.120292
R21132 VDD.n2526 VDD.n2516 0.120292
R21133 VDD.n2520 VDD.n2516 0.120292
R21134 VDD.n2520 VDD.n2519 0.120292
R21135 VDD.n2519 VDD.n2518 0.120292
R21136 VDD.n2518 VDD.n2493 0.120292
R21137 VDD.n2599 VDD.n2493 0.120292
R21138 VDD.n2600 VDD.n2599 0.120292
R21139 VDD.n2600 VDD.n2490 0.120292
R21140 VDD.n2606 VDD.n2490 0.120292
R21141 VDD.n2607 VDD.n2606 0.120292
R21142 VDD.n2608 VDD.n2607 0.120292
R21143 VDD.n2608 VDD.n2488 0.120292
R21144 VDD.n2617 VDD.n2488 0.120292
R21145 VDD.n2618 VDD.n2617 0.120292
R21146 VDD.n2619 VDD.n2618 0.120292
R21147 VDD.n2619 VDD.n2486 0.120292
R21148 VDD.n2624 VDD.n2486 0.120292
R21149 VDD.n2625 VDD.n2624 0.120292
R21150 VDD.n2626 VDD.n2625 0.120292
R21151 VDD.n2626 VDD.n2484 0.120292
R21152 VDD.n2632 VDD.n2484 0.120292
R21153 VDD.n2633 VDD.n2632 0.120292
R21154 VDD.n2634 VDD.n2633 0.120292
R21155 VDD.n2634 VDD.n2481 0.120292
R21156 VDD.n2638 VDD.n2481 0.120292
R21157 VDD.n2639 VDD.n2638 0.120292
R21158 VDD.n2639 VDD.n2477 0.120292
R21159 VDD.n2645 VDD.n2477 0.120292
R21160 VDD.n2646 VDD.n2645 0.120292
R21161 VDD.n2647 VDD.n2646 0.120292
R21162 VDD.n2647 VDD.n2475 0.120292
R21163 VDD.n2651 VDD.n2475 0.120292
R21164 VDD.n2723 VDD.n2651 0.120292
R21165 VDD.n2723 VDD.n2722 0.120292
R21166 VDD.n2722 VDD.n2721 0.120292
R21167 VDD.n2721 VDD.n2652 0.120292
R21168 VDD.n2717 VDD.n2652 0.120292
R21169 VDD.n2717 VDD.n2716 0.120292
R21170 VDD.n2716 VDD.n2715 0.120292
R21171 VDD.n2715 VDD.n2654 0.120292
R21172 VDD.n2656 VDD.n2654 0.120292
R21173 VDD.n2710 VDD.n2656 0.120292
R21174 VDD.n2710 VDD.n2709 0.120292
R21175 VDD.n2709 VDD.n2708 0.120292
R21176 VDD.n2708 VDD.n2659 0.120292
R21177 VDD.n2702 VDD.n2659 0.120292
R21178 VDD.n2702 VDD.n2701 0.120292
R21179 VDD.n2701 VDD.n2700 0.120292
R21180 VDD.n2700 VDD.n2664 0.120292
R21181 VDD.n2696 VDD.n2664 0.120292
R21182 VDD.n2696 VDD.n2695 0.120292
R21183 VDD.n2695 VDD.n2666 0.120292
R21184 VDD.n2690 VDD.n2666 0.120292
R21185 VDD.n2690 VDD.n2689 0.120292
R21186 VDD.n2689 VDD.n2670 0.120292
R21187 VDD.n2684 VDD.n2670 0.120292
R21188 VDD.n2684 VDD.n2683 0.120292
R21189 VDD.n2683 VDD.n2682 0.120292
R21190 VDD.n2682 VDD.n2673 0.120292
R21191 VDD.n2676 VDD.n2673 0.120292
R21192 VDD.n2676 VDD.n2469 0.120292
R21193 VDD.n2730 VDD.n2469 0.120292
R21194 VDD.n2731 VDD.n2730 0.120292
R21195 VDD.n2732 VDD.n2731 0.120292
R21196 VDD.n2732 VDD.n2467 0.120292
R21197 VDD.n2467 VDD.n2465 0.120292
R21198 VDD.n2737 VDD.n2465 0.120292
R21199 VDD.n2738 VDD.n2737 0.120292
R21200 VDD.n2739 VDD.n2738 0.120292
R21201 VDD.n2739 VDD.n2461 0.120292
R21202 VDD.n2743 VDD.n2461 0.120292
R21203 VDD.n2744 VDD.n2743 0.120292
R21204 VDD.n2744 VDD.n2458 0.120292
R21205 VDD.n2458 VDD.n2457 0.120292
R21206 VDD.n2749 VDD.n2457 0.120292
R21207 VDD.n2750 VDD.n2749 0.120292
R21208 VDD.n2751 VDD.n2750 0.120292
R21209 VDD.n2751 VDD.n2453 0.120292
R21210 VDD.n2453 VDD.n2452 0.120292
R21211 VDD.n2452 VDD.n2451 0.120292
R21212 VDD.n2758 VDD.n2451 0.120292
R21213 VDD.n2759 VDD.n2758 0.120292
R21214 VDD.n2759 VDD.n2449 0.120292
R21215 VDD.n2767 VDD.n2449 0.120292
R21216 VDD.n2768 VDD.n2767 0.120292
R21217 VDD.n2768 VDD.n2447 0.120292
R21218 VDD.n2447 VDD.n2446 0.120292
R21219 VDD.n2773 VDD.n2446 0.120292
R21220 VDD.n2774 VDD.n2773 0.120292
R21221 VDD.n2775 VDD.n2774 0.120292
R21222 VDD.n2775 VDD.n2444 0.120292
R21223 VDD.n2444 VDD.n2442 0.120292
R21224 VDD.n2442 VDD.n2440 0.120292
R21225 VDD.n2783 VDD.n2440 0.120292
R21226 VDD.n2784 VDD.n2783 0.120292
R21227 VDD.n2785 VDD.n2784 0.120292
R21228 VDD.n2785 VDD.n2438 0.120292
R21229 VDD.n2790 VDD.n2438 0.120292
R21230 VDD.n2791 VDD.n2790 0.120292
R21231 VDD.n2791 VDD.n2436 0.120292
R21232 VDD.n2436 VDD.n2435 0.120292
R21233 VDD.n2435 VDD.n2434 0.120292
R21234 VDD.n2434 VDD.n2432 0.120292
R21235 VDD.n2799 VDD.n2432 0.120292
R21236 VDD.n2800 VDD.n2799 0.120292
R21237 VDD.n2800 VDD.n2429 0.120292
R21238 VDD.n2429 VDD.n2428 0.120292
R21239 VDD.n2807 VDD.n2428 0.120292
R21240 VDD.n2808 VDD.n2807 0.120292
R21241 VDD.n2809 VDD.n2808 0.120292
R21242 VDD.n2809 VDD.n2423 0.120292
R21243 VDD.n2817 VDD.n2423 0.120292
R21244 VDD.n2818 VDD.n2817 0.120292
R21245 VDD.n2819 VDD.n2818 0.120292
R21246 VDD.n2819 VDD.n2419 0.120292
R21247 VDD.n2823 VDD.n2419 0.120292
R21248 VDD.n2892 VDD.n2823 0.120292
R21249 VDD.n2892 VDD.n2891 0.120292
R21250 VDD.n2891 VDD.n2890 0.120292
R21251 VDD.n2890 VDD.n2824 0.120292
R21252 VDD.n2884 VDD.n2824 0.120292
R21253 VDD.n2884 VDD.n2883 0.120292
R21254 VDD.n2883 VDD.n2882 0.120292
R21255 VDD.n2882 VDD.n2828 0.120292
R21256 VDD.n2876 VDD.n2828 0.120292
R21257 VDD.n2876 VDD.n2875 0.120292
R21258 VDD.n2875 VDD.n2874 0.120292
R21259 VDD.n2874 VDD.n2830 0.120292
R21260 VDD.n2870 VDD.n2830 0.120292
R21261 VDD.n2870 VDD.n2869 0.120292
R21262 VDD.n2869 VDD.n2868 0.120292
R21263 VDD.n2868 VDD.n2833 0.120292
R21264 VDD.n2864 VDD.n2833 0.120292
R21265 VDD.n2864 VDD.n2863 0.120292
R21266 VDD.n2863 VDD.n2862 0.120292
R21267 VDD.n2862 VDD.n2836 0.120292
R21268 VDD.n2858 VDD.n2836 0.120292
R21269 VDD.n2858 VDD.n2857 0.120292
R21270 VDD.n2857 VDD.n2839 0.120292
R21271 VDD.n2841 VDD.n2839 0.120292
R21272 VDD.n2851 VDD.n2841 0.120292
R21273 VDD.n2851 VDD.n2850 0.120292
R21274 VDD.n2850 VDD.n2849 0.120292
R21275 VDD.n2849 VDD.n2845 0.120292
R21276 VDD.n2845 VDD.n2414 0.120292
R21277 VDD.n2414 VDD.n2410 0.120292
R21278 VDD.n2902 VDD.n2410 0.120292
R21279 VDD.n2903 VDD.n2902 0.120292
R21280 VDD.n2903 VDD.n2406 0.120292
R21281 VDD.n2911 VDD.n2406 0.120292
R21282 VDD.n2912 VDD.n2911 0.120292
R21283 VDD.n2912 VDD.n2403 0.120292
R21284 VDD.n2917 VDD.n2403 0.120292
R21285 VDD.n2918 VDD.n2917 0.120292
R21286 VDD.n2918 VDD.n2400 0.120292
R21287 VDD.n2400 VDD.n2399 0.120292
R21288 VDD.n2924 VDD.n2399 0.120292
R21289 VDD.n2925 VDD.n2924 0.120292
R21290 VDD.n2926 VDD.n2925 0.120292
R21291 VDD.n2926 VDD.n2397 0.120292
R21292 VDD.n2397 VDD.n2394 0.120292
R21293 VDD.n2932 VDD.n2394 0.120292
R21294 VDD.n2933 VDD.n2932 0.120292
R21295 VDD.n2934 VDD.n2933 0.120292
R21296 VDD.n2934 VDD.n2391 0.120292
R21297 VDD.n2391 VDD.n2390 0.120292
R21298 VDD.n2939 VDD.n2390 0.120292
R21299 VDD.n2940 VDD.n2939 0.120292
R21300 VDD.n2941 VDD.n2940 0.120292
R21301 VDD.n2941 VDD.n2387 0.120292
R21302 VDD.n2387 VDD.n2385 0.120292
R21303 VDD.n2946 VDD.n2385 0.120292
R21304 VDD.n2947 VDD.n2946 0.120292
R21305 VDD.n2948 VDD.n2947 0.120292
R21306 VDD.n2948 VDD.n2383 0.120292
R21307 VDD.n2954 VDD.n2383 0.120292
R21308 VDD.n2955 VDD.n2954 0.120292
R21309 VDD.n2956 VDD.n2955 0.120292
R21310 VDD.n2956 VDD.n2381 0.120292
R21311 VDD.n2960 VDD.n2381 0.120292
R21312 VDD.n2961 VDD.n2960 0.120292
R21313 VDD.n2962 VDD.n2961 0.120292
R21314 VDD.n2962 VDD.n2378 0.120292
R21315 VDD.n2972 VDD.n2378 0.120292
R21316 VDD.n2973 VDD.n2972 0.120292
R21317 VDD.n2974 VDD.n2973 0.120292
R21318 VDD.n2974 VDD.n2376 0.120292
R21319 VDD.n2978 VDD.n2376 0.120292
R21320 VDD.n2979 VDD.n2978 0.120292
R21321 VDD.n2980 VDD.n2979 0.120292
R21322 VDD.n2980 VDD.n2371 0.120292
R21323 VDD.n2987 VDD.n2371 0.120292
R21324 VDD.n2988 VDD.n2987 0.120292
R21325 VDD.n2988 VDD.n2368 0.120292
R21326 VDD.n2992 VDD.n2368 0.120292
R21327 VDD.n2993 VDD.n2992 0.120292
R21328 VDD.n2994 VDD.n2993 0.120292
R21329 VDD.n2994 VDD.n2363 0.120292
R21330 VDD.n3001 VDD.n2363 0.120292
R21331 VDD.n3002 VDD.n3001 0.120292
R21332 VDD.n3062 VDD.n3002 0.120292
R21333 VDD.n3062 VDD.n3061 0.120292
R21334 VDD.n3061 VDD.n3003 0.120292
R21335 VDD.n3056 VDD.n3003 0.120292
R21336 VDD.n3056 VDD.n3055 0.120292
R21337 VDD.n3055 VDD.n3007 0.120292
R21338 VDD.n3010 VDD.n3007 0.120292
R21339 VDD.n3017 VDD.n3010 0.120292
R21340 VDD.n3018 VDD.n3017 0.120292
R21341 VDD.n3047 VDD.n3018 0.120292
R21342 VDD.n3047 VDD.n3046 0.120292
R21343 VDD.n3046 VDD.n3019 0.120292
R21344 VDD.n3039 VDD.n3019 0.120292
R21345 VDD.n3039 VDD.n3038 0.120292
R21346 VDD.n3038 VDD.n3037 0.120292
R21347 VDD.n3037 VDD.n3021 0.120292
R21348 VDD.n3024 VDD.n3021 0.120292
R21349 VDD.n3026 VDD.n3024 0.120292
R21350 VDD.n3031 VDD.n3026 0.120292
R21351 VDD.n3031 VDD.n3030 0.120292
R21352 VDD.n3075 VDD.n3074 0.120292
R21353 VDD.n3074 VDD.n2284 0.120292
R21354 VDD.n3070 VDD.n2284 0.120292
R21355 VDD.n3070 VDD.n3069 0.120292
R21356 VDD.n3069 VDD.n2287 0.120292
R21357 VDD.n2358 VDD.n2287 0.120292
R21358 VDD.n2358 VDD.n2357 0.120292
R21359 VDD.n2357 VDD.n2290 0.120292
R21360 VDD.n2352 VDD.n2290 0.120292
R21361 VDD.n2352 VDD.n2351 0.120292
R21362 VDD.n2351 VDD.n2293 0.120292
R21363 VDD.n2345 VDD.n2296 0.120292
R21364 VDD.n2340 VDD.n2296 0.120292
R21365 VDD.n2340 VDD.n2339 0.120292
R21366 VDD.n2339 VDD.n2301 0.120292
R21367 VDD.n2335 VDD.n2301 0.120292
R21368 VDD.n2335 VDD.n2334 0.120292
R21369 VDD.n2334 VDD.n2304 0.120292
R21370 VDD.n2330 VDD.n2304 0.120292
R21371 VDD.n2330 VDD.n2329 0.120292
R21372 VDD.n2329 VDD.n2307 0.120292
R21373 VDD.n2325 VDD.n2307 0.120292
R21374 VDD.n2325 VDD.n2324 0.120292
R21375 VDD.n2324 VDD.n2323 0.120292
R21376 VDD.n1705 VDD.n1704 0.120292
R21377 VDD.n1706 VDD.n1705 0.120292
R21378 VDD.n1706 VDD.n1690 0.120292
R21379 VDD.n1712 VDD.n1690 0.120292
R21380 VDD.n1713 VDD.n1712 0.120292
R21381 VDD.n1714 VDD.n1713 0.120292
R21382 VDD.n1714 VDD.n1686 0.120292
R21383 VDD.n1718 VDD.n1686 0.120292
R21384 VDD.n1719 VDD.n1718 0.120292
R21385 VDD.n1720 VDD.n1719 0.120292
R21386 VDD.n1720 VDD.n1682 0.120292
R21387 VDD.n1682 VDD.n1680 0.120292
R21388 VDD.n1726 VDD.n1680 0.120292
R21389 VDD.n1727 VDD.n1726 0.120292
R21390 VDD.n1727 VDD.n1678 0.120292
R21391 VDD.n1678 VDD.n1677 0.120292
R21392 VDD.n1677 VDD.n1675 0.120292
R21393 VDD.n1675 VDD.n1674 0.120292
R21394 VDD.n1674 VDD.n1672 0.120292
R21395 VDD.n1735 VDD.n1672 0.120292
R21396 VDD.n1736 VDD.n1735 0.120292
R21397 VDD.n1736 VDD.n1669 0.120292
R21398 VDD.n1669 VDD.n1668 0.120292
R21399 VDD.n1668 VDD.n1665 0.120292
R21400 VDD.n1742 VDD.n1665 0.120292
R21401 VDD.n1743 VDD.n1742 0.120292
R21402 VDD.n1743 VDD.n1662 0.120292
R21403 VDD.n1748 VDD.n1662 0.120292
R21404 VDD.n1749 VDD.n1748 0.120292
R21405 VDD.n1750 VDD.n1749 0.120292
R21406 VDD.n1750 VDD.n1659 0.120292
R21407 VDD.n1754 VDD.n1659 0.120292
R21408 VDD.n1755 VDD.n1754 0.120292
R21409 VDD.n1756 VDD.n1755 0.120292
R21410 VDD.n1756 VDD.n1655 0.120292
R21411 VDD.n1761 VDD.n1655 0.120292
R21412 VDD.n1762 VDD.n1761 0.120292
R21413 VDD.n1762 VDD.n1652 0.120292
R21414 VDD.n1652 VDD.n1649 0.120292
R21415 VDD.n1769 VDD.n1768 0.120292
R21416 VDD.n1769 VDD.n1647 0.120292
R21417 VDD.n1773 VDD.n1647 0.120292
R21418 VDD.n1774 VDD.n1773 0.120292
R21419 VDD.n1774 VDD.n1643 0.120292
R21420 VDD.n1779 VDD.n1643 0.120292
R21421 VDD.n1780 VDD.n1779 0.120292
R21422 VDD.n1781 VDD.n1780 0.120292
R21423 VDD.n1781 VDD.n1640 0.120292
R21424 VDD.n1640 VDD.n1639 0.120292
R21425 VDD.n1789 VDD.n1639 0.120292
R21426 VDD.n1790 VDD.n1789 0.120292
R21427 VDD.n1791 VDD.n1790 0.120292
R21428 VDD.n1791 VDD.n1636 0.120292
R21429 VDD.n1797 VDD.n1636 0.120292
R21430 VDD.n1798 VDD.n1797 0.120292
R21431 VDD.n1798 VDD.n1632 0.120292
R21432 VDD.n1803 VDD.n1632 0.120292
R21433 VDD.n1804 VDD.n1803 0.120292
R21434 VDD.n1805 VDD.n1804 0.120292
R21435 VDD.n1805 VDD.n1629 0.120292
R21436 VDD.n1629 VDD.n1628 0.120292
R21437 VDD.n1628 VDD.n1626 0.120292
R21438 VDD.n1813 VDD.n1626 0.120292
R21439 VDD.n1814 VDD.n1813 0.120292
R21440 VDD.n1815 VDD.n1814 0.120292
R21441 VDD.n1815 VDD.n1623 0.120292
R21442 VDD.n1623 VDD.n1620 0.120292
R21443 VDD.n1821 VDD.n1620 0.120292
R21444 VDD.n1822 VDD.n1821 0.120292
R21445 VDD.n1822 VDD.n1617 0.120292
R21446 VDD.n1829 VDD.n1617 0.120292
R21447 VDD.n1830 VDD.n1829 0.120292
R21448 VDD.n1830 VDD.n1612 0.120292
R21449 VDD.n1835 VDD.n1612 0.120292
R21450 VDD.n1836 VDD.n1835 0.120292
R21451 VDD.n1837 VDD.n1836 0.120292
R21452 VDD.n1837 VDD.n1607 0.120292
R21453 VDD.n1843 VDD.n1607 0.120292
R21454 VDD.n1844 VDD.n1843 0.120292
R21455 VDD.n1844 VDD.n1604 0.120292
R21456 VDD.n1850 VDD.n1604 0.120292
R21457 VDD.n1851 VDD.n1850 0.120292
R21458 VDD.n1851 VDD.n1601 0.120292
R21459 VDD.n1601 VDD.n1599 0.120292
R21460 VDD.n1856 VDD.n1599 0.120292
R21461 VDD.n1857 VDD.n1856 0.120292
R21462 VDD.n1858 VDD.n1857 0.120292
R21463 VDD.n1858 VDD.n1595 0.120292
R21464 VDD.n1862 VDD.n1595 0.120292
R21465 VDD.n1863 VDD.n1862 0.120292
R21466 VDD.n1864 VDD.n1863 0.120292
R21467 VDD.n1864 VDD.n1592 0.120292
R21468 VDD.n1875 VDD.n1874 0.120292
R21469 VDD.n1875 VDD.n1589 0.120292
R21470 VDD.n1880 VDD.n1589 0.120292
R21471 VDD.n1881 VDD.n1880 0.120292
R21472 VDD.n1882 VDD.n1881 0.120292
R21473 VDD.n1882 VDD.n1587 0.120292
R21474 VDD.n1888 VDD.n1587 0.120292
R21475 VDD.n1891 VDD.n1890 0.120292
R21476 VDD.n1891 VDD.n1580 0.120292
R21477 VDD.n1896 VDD.n1580 0.120292
R21478 VDD.n1897 VDD.n1896 0.120292
R21479 VDD.n1897 VDD.n1577 0.120292
R21480 VDD.n1903 VDD.n1577 0.120292
R21481 VDD.n1904 VDD.n1903 0.120292
R21482 VDD.n1905 VDD.n1904 0.120292
R21483 VDD.n1914 VDD.n1913 0.120292
R21484 VDD.n1914 VDD.n1573 0.120292
R21485 VDD.n1919 VDD.n1573 0.120292
R21486 VDD.n1920 VDD.n1919 0.120292
R21487 VDD.n1920 VDD.n1571 0.120292
R21488 VDD.n1925 VDD.n1571 0.120292
R21489 VDD.n1926 VDD.n1925 0.120292
R21490 VDD.n1927 VDD.n1926 0.120292
R21491 VDD.n1927 VDD.n1568 0.120292
R21492 VDD.n1932 VDD.n1568 0.120292
R21493 VDD.n1933 VDD.n1932 0.120292
R21494 VDD.n1934 VDD.n1933 0.120292
R21495 VDD.n1934 VDD.n1566 0.120292
R21496 VDD.n1938 VDD.n1566 0.120292
R21497 VDD.n1939 VDD.n1938 0.120292
R21498 VDD.n1940 VDD.n1939 0.120292
R21499 VDD.n1940 VDD.n1563 0.120292
R21500 VDD.n1945 VDD.n1563 0.120292
R21501 VDD.n1946 VDD.n1945 0.120292
R21502 VDD.n1947 VDD.n1946 0.120292
R21503 VDD.n1947 VDD.n1561 0.120292
R21504 VDD.n1952 VDD.n1561 0.120292
R21505 VDD.n1953 VDD.n1952 0.120292
R21506 VDD.n2024 VDD.n1953 0.120292
R21507 VDD.n2024 VDD.n2023 0.120292
R21508 VDD.n2023 VDD.n2022 0.120292
R21509 VDD.n2022 VDD.n1956 0.120292
R21510 VDD.n2018 VDD.n1956 0.120292
R21511 VDD.n2018 VDD.n2017 0.120292
R21512 VDD.n2017 VDD.n2016 0.120292
R21513 VDD.n2016 VDD.n1959 0.120292
R21514 VDD.n2009 VDD.n2008 0.120292
R21515 VDD.n2008 VDD.n1961 0.120292
R21516 VDD.n2002 VDD.n1961 0.120292
R21517 VDD.n2002 VDD.n2001 0.120292
R21518 VDD.n2001 VDD.n2000 0.120292
R21519 VDD.n2000 VDD.n1966 0.120292
R21520 VDD.n1994 VDD.n1966 0.120292
R21521 VDD.n1994 VDD.n1993 0.120292
R21522 VDD.n1993 VDD.n1969 0.120292
R21523 VDD.n1986 VDD.n1969 0.120292
R21524 VDD.n1986 VDD.n1985 0.120292
R21525 VDD.n1985 VDD.n1984 0.120292
R21526 VDD.n1984 VDD.n1972 0.120292
R21527 VDD.n1977 VDD.n1972 0.120292
R21528 VDD.n1977 VDD.n1976 0.120292
R21529 VDD.n1976 VDD.n1557 0.120292
R21530 VDD.n2031 VDD.n1557 0.120292
R21531 VDD.n2032 VDD.n2031 0.120292
R21532 VDD.n2033 VDD.n2032 0.120292
R21533 VDD.n2033 VDD.n1554 0.120292
R21534 VDD.n2038 VDD.n1554 0.120292
R21535 VDD.n2039 VDD.n2038 0.120292
R21536 VDD.n2039 VDD.n1551 0.120292
R21537 VDD.n2043 VDD.n1551 0.120292
R21538 VDD.n2044 VDD.n2043 0.120292
R21539 VDD.n2045 VDD.n2044 0.120292
R21540 VDD.n2045 VDD.n1549 0.120292
R21541 VDD.n1549 VDD.n1546 0.120292
R21542 VDD.n2050 VDD.n1546 0.120292
R21543 VDD.n2051 VDD.n2050 0.120292
R21544 VDD.n2052 VDD.n2051 0.120292
R21545 VDD.n2052 VDD.n1544 0.120292
R21546 VDD.n1544 VDD.n1543 0.120292
R21547 VDD.n1543 VDD.n1542 0.120292
R21548 VDD.n2059 VDD.n1542 0.120292
R21549 VDD.n2060 VDD.n2059 0.120292
R21550 VDD.n2060 VDD.n1539 0.120292
R21551 VDD.n2065 VDD.n1539 0.120292
R21552 VDD.n2067 VDD.n1533 0.120292
R21553 VDD.n2071 VDD.n1533 0.120292
R21554 VDD.n2072 VDD.n2071 0.120292
R21555 VDD.n2073 VDD.n2072 0.120292
R21556 VDD.n2073 VDD.n1531 0.120292
R21557 VDD.n2077 VDD.n1531 0.120292
R21558 VDD.n2078 VDD.n2077 0.120292
R21559 VDD.n2079 VDD.n2078 0.120292
R21560 VDD.n2079 VDD.n1529 0.120292
R21561 VDD.n2087 VDD.n1529 0.120292
R21562 VDD.n2088 VDD.n2087 0.120292
R21563 VDD.n2089 VDD.n2088 0.120292
R21564 VDD.n2089 VDD.n1527 0.120292
R21565 VDD.n2093 VDD.n1527 0.120292
R21566 VDD.n2094 VDD.n2093 0.120292
R21567 VDD.n2094 VDD.n1525 0.120292
R21568 VDD.n2099 VDD.n1525 0.120292
R21569 VDD.n2100 VDD.n2099 0.120292
R21570 VDD.n2101 VDD.n2100 0.120292
R21571 VDD.n2101 VDD.n1522 0.120292
R21572 VDD.n2106 VDD.n1522 0.120292
R21573 VDD.n2107 VDD.n2106 0.120292
R21574 VDD.n2108 VDD.n2107 0.120292
R21575 VDD.n2108 VDD.n1520 0.120292
R21576 VDD.n2112 VDD.n1520 0.120292
R21577 VDD.n2113 VDD.n2112 0.120292
R21578 VDD.n2114 VDD.n2113 0.120292
R21579 VDD.n2114 VDD.n1518 0.120292
R21580 VDD.n2119 VDD.n1518 0.120292
R21581 VDD.n2120 VDD.n2119 0.120292
R21582 VDD.n2121 VDD.n2120 0.120292
R21583 VDD.n2168 VDD.n2121 0.120292
R21584 VDD.n2168 VDD.n2167 0.120292
R21585 VDD.n2167 VDD.n2166 0.120292
R21586 VDD.n2166 VDD.n2124 0.120292
R21587 VDD.n2125 VDD.n2124 0.120292
R21588 VDD.n2161 VDD.n2125 0.120292
R21589 VDD.n2161 VDD.n2160 0.120292
R21590 VDD.n2160 VDD.n2159 0.120292
R21591 VDD.n2159 VDD.n2128 0.120292
R21592 VDD.n2155 VDD.n2128 0.120292
R21593 VDD.n2155 VDD.n2154 0.120292
R21594 VDD.n2150 VDD.n2149 0.120292
R21595 VDD.n2149 VDD.n2148 0.120292
R21596 VDD.n2148 VDD.n2134 0.120292
R21597 VDD.n2143 VDD.n2134 0.120292
R21598 VDD.n2143 VDD.n2142 0.120292
R21599 VDD.n2259 VDD.n1512 0.120292
R21600 VDD.n2253 VDD.n1512 0.120292
R21601 VDD.n2253 VDD.n2252 0.120292
R21602 VDD.n2252 VDD.n1516 0.120292
R21603 VDD.n2246 VDD.n1516 0.120292
R21604 VDD.n2246 VDD.n2245 0.120292
R21605 VDD.n2245 VDD.n2244 0.120292
R21606 VDD.n2244 VDD.n2175 0.120292
R21607 VDD.n2239 VDD.n2175 0.120292
R21608 VDD.n2239 VDD.n2238 0.120292
R21609 VDD.n2238 VDD.n2237 0.120292
R21610 VDD.n2237 VDD.n2177 0.120292
R21611 VDD.n2232 VDD.n2177 0.120292
R21612 VDD.n2232 VDD.n2231 0.120292
R21613 VDD.n2231 VDD.n2230 0.120292
R21614 VDD.n2230 VDD.n2183 0.120292
R21615 VDD.n2185 VDD.n2183 0.120292
R21616 VDD.n2224 VDD.n2185 0.120292
R21617 VDD.n2224 VDD.n2223 0.120292
R21618 VDD.n2223 VDD.n2222 0.120292
R21619 VDD.n2222 VDD.n2187 0.120292
R21620 VDD.n2218 VDD.n2187 0.120292
R21621 VDD.n2218 VDD.n2217 0.120292
R21622 VDD.n2217 VDD.n2216 0.120292
R21623 VDD.n2216 VDD.n2190 0.120292
R21624 VDD.n2193 VDD.n2190 0.120292
R21625 VDD.n2209 VDD.n2193 0.120292
R21626 VDD.n2209 VDD.n2208 0.120292
R21627 VDD.n2208 VDD.n2207 0.120292
R21628 VDD.n864 VDD.n854 0.120292
R21629 VDD.n870 VDD.n854 0.120292
R21630 VDD.n871 VDD.n870 0.120292
R21631 VDD.n871 VDD.n850 0.120292
R21632 VDD.n877 VDD.n850 0.120292
R21633 VDD.n878 VDD.n877 0.120292
R21634 VDD.n949 VDD.n878 0.120292
R21635 VDD.n949 VDD.n948 0.120292
R21636 VDD.n948 VDD.n879 0.120292
R21637 VDD.n943 VDD.n879 0.120292
R21638 VDD.n943 VDD.n942 0.120292
R21639 VDD.n942 VDD.n941 0.120292
R21640 VDD.n941 VDD.n882 0.120292
R21641 VDD.n935 VDD.n882 0.120292
R21642 VDD.n935 VDD.n934 0.120292
R21643 VDD.n934 VDD.n884 0.120292
R21644 VDD.n929 VDD.n884 0.120292
R21645 VDD.n929 VDD.n928 0.120292
R21646 VDD.n928 VDD.n927 0.120292
R21647 VDD.n927 VDD.n886 0.120292
R21648 VDD.n921 VDD.n886 0.120292
R21649 VDD.n921 VDD.n920 0.120292
R21650 VDD.n920 VDD.n891 0.120292
R21651 VDD.n916 VDD.n891 0.120292
R21652 VDD.n916 VDD.n915 0.120292
R21653 VDD.n915 VDD.n914 0.120292
R21654 VDD.n914 VDD.n893 0.120292
R21655 VDD.n909 VDD.n893 0.120292
R21656 VDD.n909 VDD.n908 0.120292
R21657 VDD.n908 VDD.n907 0.120292
R21658 VDD.n907 VDD.n899 0.120292
R21659 VDD.n903 VDD.n899 0.120292
R21660 VDD.n903 VDD.n902 0.120292
R21661 VDD.n902 VDD.n845 0.120292
R21662 VDD.n954 VDD.n845 0.120292
R21663 VDD.n955 VDD.n954 0.120292
R21664 VDD.n956 VDD.n955 0.120292
R21665 VDD.n956 VDD.n842 0.120292
R21666 VDD.n842 VDD.n841 0.120292
R21667 VDD.n962 VDD.n841 0.120292
R21668 VDD.n963 VDD.n962 0.120292
R21669 VDD.n964 VDD.n963 0.120292
R21670 VDD.n964 VDD.n837 0.120292
R21671 VDD.n837 VDD.n836 0.120292
R21672 VDD.n974 VDD.n836 0.120292
R21673 VDD.n975 VDD.n974 0.120292
R21674 VDD.n976 VDD.n975 0.120292
R21675 VDD.n976 VDD.n832 0.120292
R21676 VDD.n982 VDD.n832 0.120292
R21677 VDD.n983 VDD.n982 0.120292
R21678 VDD.n984 VDD.n983 0.120292
R21679 VDD.n984 VDD.n830 0.120292
R21680 VDD.n830 VDD.n828 0.120292
R21681 VDD.n828 VDD.n827 0.120292
R21682 VDD.n992 VDD.n827 0.120292
R21683 VDD.n993 VDD.n992 0.120292
R21684 VDD.n993 VDD.n824 0.120292
R21685 VDD.n997 VDD.n824 0.120292
R21686 VDD.n998 VDD.n997 0.120292
R21687 VDD.n998 VDD.n820 0.120292
R21688 VDD.n1002 VDD.n820 0.120292
R21689 VDD.n1003 VDD.n1002 0.120292
R21690 VDD.n1076 VDD.n1003 0.120292
R21691 VDD.n1076 VDD.n1075 0.120292
R21692 VDD.n1075 VDD.n1074 0.120292
R21693 VDD.n1074 VDD.n1004 0.120292
R21694 VDD.n1069 VDD.n1004 0.120292
R21695 VDD.n1069 VDD.n1068 0.120292
R21696 VDD.n1068 VDD.n1067 0.120292
R21697 VDD.n1067 VDD.n1009 0.120292
R21698 VDD.n1062 VDD.n1009 0.120292
R21699 VDD.n1062 VDD.n1061 0.120292
R21700 VDD.n1061 VDD.n1011 0.120292
R21701 VDD.n1056 VDD.n1011 0.120292
R21702 VDD.n1056 VDD.n1055 0.120292
R21703 VDD.n1055 VDD.n1054 0.120292
R21704 VDD.n1054 VDD.n1014 0.120292
R21705 VDD.n1048 VDD.n1014 0.120292
R21706 VDD.n1048 VDD.n1047 0.120292
R21707 VDD.n1047 VDD.n1046 0.120292
R21708 VDD.n1046 VDD.n1016 0.120292
R21709 VDD.n1041 VDD.n1016 0.120292
R21710 VDD.n1041 VDD.n1040 0.120292
R21711 VDD.n1040 VDD.n1039 0.120292
R21712 VDD.n1039 VDD.n1021 0.120292
R21713 VDD.n1033 VDD.n1021 0.120292
R21714 VDD.n1033 VDD.n1032 0.120292
R21715 VDD.n1032 VDD.n1031 0.120292
R21716 VDD.n1031 VDD.n1025 0.120292
R21717 VDD.n1025 VDD.n1024 0.120292
R21718 VDD.n1024 VDD.n816 0.120292
R21719 VDD.n1082 VDD.n816 0.120292
R21720 VDD.n1083 VDD.n1082 0.120292
R21721 VDD.n1084 VDD.n1083 0.120292
R21722 VDD.n1084 VDD.n812 0.120292
R21723 VDD.n1089 VDD.n812 0.120292
R21724 VDD.n1090 VDD.n1089 0.120292
R21725 VDD.n1090 VDD.n809 0.120292
R21726 VDD.n1095 VDD.n809 0.120292
R21727 VDD.n1096 VDD.n1095 0.120292
R21728 VDD.n1096 VDD.n806 0.120292
R21729 VDD.n1103 VDD.n806 0.120292
R21730 VDD.n1104 VDD.n1103 0.120292
R21731 VDD.n1105 VDD.n1104 0.120292
R21732 VDD.n1105 VDD.n803 0.120292
R21733 VDD.n1109 VDD.n803 0.120292
R21734 VDD.n1110 VDD.n1109 0.120292
R21735 VDD.n1111 VDD.n1110 0.120292
R21736 VDD.n1111 VDD.n799 0.120292
R21737 VDD.n1117 VDD.n799 0.120292
R21738 VDD.n1118 VDD.n1117 0.120292
R21739 VDD.n1119 VDD.n1118 0.120292
R21740 VDD.n1119 VDD.n797 0.120292
R21741 VDD.n797 VDD.n796 0.120292
R21742 VDD.n796 VDD.n794 0.120292
R21743 VDD.n794 VDD.n792 0.120292
R21744 VDD.n1126 VDD.n792 0.120292
R21745 VDD.n1127 VDD.n1126 0.120292
R21746 VDD.n1197 VDD.n1127 0.120292
R21747 VDD.n1197 VDD.n1196 0.120292
R21748 VDD.n1196 VDD.n1195 0.120292
R21749 VDD.n1195 VDD.n1128 0.120292
R21750 VDD.n1131 VDD.n1128 0.120292
R21751 VDD.n1132 VDD.n1131 0.120292
R21752 VDD.n1189 VDD.n1132 0.120292
R21753 VDD.n1189 VDD.n1188 0.120292
R21754 VDD.n1188 VDD.n1187 0.120292
R21755 VDD.n1187 VDD.n1134 0.120292
R21756 VDD.n1135 VDD.n1134 0.120292
R21757 VDD.n1182 VDD.n1135 0.120292
R21758 VDD.n1182 VDD.n1181 0.120292
R21759 VDD.n1181 VDD.n1139 0.120292
R21760 VDD.n1175 VDD.n1139 0.120292
R21761 VDD.n1175 VDD.n1174 0.120292
R21762 VDD.n1174 VDD.n1173 0.120292
R21763 VDD.n1173 VDD.n1141 0.120292
R21764 VDD.n1144 VDD.n1141 0.120292
R21765 VDD.n1168 VDD.n1144 0.120292
R21766 VDD.n1168 VDD.n1167 0.120292
R21767 VDD.n1167 VDD.n1146 0.120292
R21768 VDD.n1148 VDD.n1146 0.120292
R21769 VDD.n1160 VDD.n1148 0.120292
R21770 VDD.n1160 VDD.n1159 0.120292
R21771 VDD.n1159 VDD.n1158 0.120292
R21772 VDD.n1158 VDD.n1152 0.120292
R21773 VDD.n1152 VDD.n786 0.120292
R21774 VDD.n1203 VDD.n786 0.120292
R21775 VDD.n1204 VDD.n1203 0.120292
R21776 VDD.n1205 VDD.n1204 0.120292
R21777 VDD.n1205 VDD.n783 0.120292
R21778 VDD.n1212 VDD.n783 0.120292
R21779 VDD.n1213 VDD.n1212 0.120292
R21780 VDD.n1214 VDD.n1213 0.120292
R21781 VDD.n1214 VDD.n780 0.120292
R21782 VDD.n780 VDD.n778 0.120292
R21783 VDD.n1220 VDD.n778 0.120292
R21784 VDD.n1221 VDD.n1220 0.120292
R21785 VDD.n1221 VDD.n774 0.120292
R21786 VDD.n1226 VDD.n774 0.120292
R21787 VDD.n1227 VDD.n1226 0.120292
R21788 VDD.n1228 VDD.n1227 0.120292
R21789 VDD.n1228 VDD.n772 0.120292
R21790 VDD.n1233 VDD.n772 0.120292
R21791 VDD.n1234 VDD.n1233 0.120292
R21792 VDD.n1234 VDD.n769 0.120292
R21793 VDD.n769 VDD.n767 0.120292
R21794 VDD.n1240 VDD.n767 0.120292
R21795 VDD.n1241 VDD.n1240 0.120292
R21796 VDD.n1241 VDD.n764 0.120292
R21797 VDD.n1247 VDD.n764 0.120292
R21798 VDD.n1248 VDD.n1247 0.120292
R21799 VDD.n1249 VDD.n1248 0.120292
R21800 VDD.n1249 VDD.n761 0.120292
R21801 VDD.n1253 VDD.n761 0.120292
R21802 VDD.n1254 VDD.n1253 0.120292
R21803 VDD.n1255 VDD.n1254 0.120292
R21804 VDD.n1255 VDD.n758 0.120292
R21805 VDD.n1263 VDD.n758 0.120292
R21806 VDD.n1264 VDD.n1263 0.120292
R21807 VDD.n1264 VDD.n756 0.120292
R21808 VDD.n1269 VDD.n756 0.120292
R21809 VDD.n1270 VDD.n1269 0.120292
R21810 VDD.n1270 VDD.n754 0.120292
R21811 VDD.n1277 VDD.n754 0.120292
R21812 VDD.n1278 VDD.n1277 0.120292
R21813 VDD.n1279 VDD.n1278 0.120292
R21814 VDD.n1279 VDD.n751 0.120292
R21815 VDD.n751 VDD.n749 0.120292
R21816 VDD.n1284 VDD.n749 0.120292
R21817 VDD.n1285 VDD.n1284 0.120292
R21818 VDD.n1286 VDD.n1285 0.120292
R21819 VDD.n1286 VDD.n745 0.120292
R21820 VDD.n1291 VDD.n745 0.120292
R21821 VDD.n1292 VDD.n1291 0.120292
R21822 VDD.n1293 VDD.n1292 0.120292
R21823 VDD.n1293 VDD.n743 0.120292
R21824 VDD.n1297 VDD.n743 0.120292
R21825 VDD.n1298 VDD.n1297 0.120292
R21826 VDD.n1299 VDD.n1298 0.120292
R21827 VDD.n1299 VDD.n741 0.120292
R21828 VDD.n741 VDD.n740 0.120292
R21829 VDD.n740 VDD.n736 0.120292
R21830 VDD.n1306 VDD.n736 0.120292
R21831 VDD.n1307 VDD.n1306 0.120292
R21832 VDD.n1308 VDD.n1307 0.120292
R21833 VDD.n1308 VDD.n732 0.120292
R21834 VDD.n1312 VDD.n732 0.120292
R21835 VDD.n1313 VDD.n1312 0.120292
R21836 VDD.n1314 VDD.n1313 0.120292
R21837 VDD.n1314 VDD.n730 0.120292
R21838 VDD.n1320 VDD.n730 0.120292
R21839 VDD.n1321 VDD.n1320 0.120292
R21840 VDD.n1322 VDD.n1321 0.120292
R21841 VDD.n1322 VDD.n728 0.120292
R21842 VDD.n1328 VDD.n728 0.120292
R21843 VDD.n1329 VDD.n1328 0.120292
R21844 VDD.n1330 VDD.n1329 0.120292
R21845 VDD.n1330 VDD.n725 0.120292
R21846 VDD.n1336 VDD.n725 0.120292
R21847 VDD.n1337 VDD.n1336 0.120292
R21848 VDD.n1338 VDD.n1337 0.120292
R21849 VDD.n1338 VDD.n722 0.120292
R21850 VDD.n1343 VDD.n722 0.120292
R21851 VDD.n1344 VDD.n1343 0.120292
R21852 VDD.n1344 VDD.n718 0.120292
R21853 VDD.n1349 VDD.n718 0.120292
R21854 VDD.n1350 VDD.n1349 0.120292
R21855 VDD.n1350 VDD.n713 0.120292
R21856 VDD.n1355 VDD.n713 0.120292
R21857 VDD.n1356 VDD.n1355 0.120292
R21858 VDD.n1357 VDD.n1356 0.120292
R21859 VDD.n1401 VDD.n1357 0.120292
R21860 VDD.n1401 VDD.n1400 0.120292
R21861 VDD.n1400 VDD.n1399 0.120292
R21862 VDD.n1399 VDD.n1359 0.120292
R21863 VDD.n1361 VDD.n1359 0.120292
R21864 VDD.n1394 VDD.n1361 0.120292
R21865 VDD.n1394 VDD.n1393 0.120292
R21866 VDD.n1393 VDD.n1363 0.120292
R21867 VDD.n1388 VDD.n1363 0.120292
R21868 VDD.n1388 VDD.n1387 0.120292
R21869 VDD.n1387 VDD.n1386 0.120292
R21870 VDD.n1386 VDD.n1367 0.120292
R21871 VDD.n1382 VDD.n1367 0.120292
R21872 VDD.n1382 VDD.n1381 0.120292
R21873 VDD.n1381 VDD.n1380 0.120292
R21874 VDD.n1380 VDD.n1370 0.120292
R21875 VDD.n1376 VDD.n1370 0.120292
R21876 VDD.n1376 VDD.n1375 0.120292
R21877 VDD.n1375 VDD.n1374 0.120292
R21878 VDD.n1488 VDD.n1487 0.120292
R21879 VDD.n1487 VDD.n705 0.120292
R21880 VDD.n708 VDD.n705 0.120292
R21881 VDD.n1481 VDD.n708 0.120292
R21882 VDD.n1481 VDD.n1480 0.120292
R21883 VDD.n1480 VDD.n711 0.120292
R21884 VDD.n1407 VDD.n711 0.120292
R21885 VDD.n1408 VDD.n1407 0.120292
R21886 VDD.n1472 VDD.n1408 0.120292
R21887 VDD.n1472 VDD.n1471 0.120292
R21888 VDD.n1471 VDD.n1470 0.120292
R21889 VDD.n1470 VDD.n1411 0.120292
R21890 VDD.n1465 VDD.n1411 0.120292
R21891 VDD.n1465 VDD.n1464 0.120292
R21892 VDD.n1464 VDD.n1415 0.120292
R21893 VDD.n1416 VDD.n1415 0.120292
R21894 VDD.n1459 VDD.n1416 0.120292
R21895 VDD.n1459 VDD.n1458 0.120292
R21896 VDD.n1458 VDD.n1457 0.120292
R21897 VDD.n1457 VDD.n1419 0.120292
R21898 VDD.n1424 VDD.n1419 0.120292
R21899 VDD.n1425 VDD.n1424 0.120292
R21900 VDD.n1451 VDD.n1425 0.120292
R21901 VDD.n1451 VDD.n1450 0.120292
R21902 VDD.n1450 VDD.n1449 0.120292
R21903 VDD.n1449 VDD.n1429 0.120292
R21904 VDD.n1445 VDD.n1429 0.120292
R21905 VDD.n1445 VDD.n1444 0.120292
R21906 VDD.n1444 VDD.n1443 0.120292
R21907 VDD.n625 VDD.n617 0.120292
R21908 VDD.n626 VDD.n625 0.120292
R21909 VDD.n626 VDD.n613 0.120292
R21910 VDD.n630 VDD.n613 0.120292
R21911 VDD.n631 VDD.n630 0.120292
R21912 VDD.n631 VDD.n606 0.120292
R21913 VDD.n691 VDD.n607 0.120292
R21914 VDD.n686 VDD.n607 0.120292
R21915 VDD.n686 VDD.n685 0.120292
R21916 VDD.n685 VDD.n637 0.120292
R21917 VDD.n681 VDD.n637 0.120292
R21918 VDD.n681 VDD.n680 0.120292
R21919 VDD.n680 VDD.n640 0.120292
R21920 VDD.n675 VDD.n640 0.120292
R21921 VDD.n675 VDD.n674 0.120292
R21922 VDD.n674 VDD.n649 0.120292
R21923 VDD.n669 VDD.n649 0.120292
R21924 VDD.n669 VDD.n668 0.120292
R21925 VDD.n668 VDD.n667 0.120292
R21926 VDD.n667 VDD.n653 0.120292
R21927 VDD.n662 VDD.n653 0.120292
R21928 VDD.n542 VDD.n534 0.120292
R21929 VDD.n543 VDD.n542 0.120292
R21930 VDD.n543 VDD.n530 0.120292
R21931 VDD.n547 VDD.n530 0.120292
R21932 VDD.n548 VDD.n547 0.120292
R21933 VDD.n548 VDD.n525 0.120292
R21934 VDD.n603 VDD.n526 0.120292
R21935 VDD.n598 VDD.n526 0.120292
R21936 VDD.n598 VDD.n597 0.120292
R21937 VDD.n597 VDD.n596 0.120292
R21938 VDD.n596 VDD.n555 0.120292
R21939 VDD.n591 VDD.n555 0.120292
R21940 VDD.n591 VDD.n590 0.120292
R21941 VDD.n590 VDD.n589 0.120292
R21942 VDD.n589 VDD.n558 0.120292
R21943 VDD.n584 VDD.n558 0.120292
R21944 VDD.n584 VDD.n583 0.120292
R21945 VDD.n583 VDD.n565 0.120292
R21946 VDD.n578 VDD.n565 0.120292
R21947 VDD.n578 VDD.n577 0.120292
R21948 VDD.n577 VDD.n576 0.120292
R21949 VDD.n462 VDD.n454 0.120292
R21950 VDD.n463 VDD.n462 0.120292
R21951 VDD.n463 VDD.n450 0.120292
R21952 VDD.n467 VDD.n450 0.120292
R21953 VDD.n468 VDD.n467 0.120292
R21954 VDD.n468 VDD.n445 0.120292
R21955 VDD.n523 VDD.n446 0.120292
R21956 VDD.n518 VDD.n446 0.120292
R21957 VDD.n518 VDD.n517 0.120292
R21958 VDD.n517 VDD.n516 0.120292
R21959 VDD.n516 VDD.n475 0.120292
R21960 VDD.n511 VDD.n475 0.120292
R21961 VDD.n511 VDD.n510 0.120292
R21962 VDD.n510 VDD.n509 0.120292
R21963 VDD.n509 VDD.n478 0.120292
R21964 VDD.n504 VDD.n478 0.120292
R21965 VDD.n504 VDD.n503 0.120292
R21966 VDD.n503 VDD.n485 0.120292
R21967 VDD.n498 VDD.n485 0.120292
R21968 VDD.n498 VDD.n497 0.120292
R21969 VDD.n497 VDD.n496 0.120292
R21970 VDD.n428 VDD.n349 0.120292
R21971 VDD.n429 VDD.n428 0.120292
R21972 VDD.n139 VDD.n138 0.120292
R21973 VDD.n139 VDD.n131 0.120292
R21974 VDD.n144 VDD.n131 0.120292
R21975 VDD.n163 VDD.n124 0.120292
R21976 VDD.n159 VDD.n124 0.120292
R21977 VDD.n78 VDD.n64 0.120292
R21978 VDD.n74 VDD.n64 0.120292
R21979 VDD.n35 VDD.n34 0.120292
R21980 VDD.n35 VDD.n27 0.120292
R21981 VDD.n48 VDD.n46 0.119731
R21982 VDD.n25 VDD.n24 0.119731
R21983 VDD.n334 VDD.n333 0.111214
R21984 VDD.n402 VDD.n398 0.109875
R21985 VDD.n401 VDD.n400 0.109875
R21986 VDD.n174 VDD.n87 0.107397
R21987 VDD.n4656 VDD.n3905 0.102087
R21988 VDD.n4223 VDD.n4222 0.102087
R21989 VDD.n3670 VDD.n3203 0.102087
R21990 VDD.n3155 VDD.n3123 0.102087
R21991 VDD.n2500 VDD.n2499 0.102087
R21992 VDD.n2556 VDD.n2555 0.102087
R21993 VDD.n2551 VDD.n2502 0.102087
R21994 VDD.n404 VDD.n403 0.102062
R21995 VDD.n405 VDD.n397 0.102062
R21996 VDD.n692 VDD.n691 0.0968542
R21997 VDD.n604 VDD.n603 0.0968542
R21998 VDD.n524 VDD.n523 0.0968542
R21999 VDD.n4676 VDD.n4675 0.0950946
R22000 VDD.n4667 VDD.n4666 0.0950946
R22001 VDD.n3891 VDD.n3890 0.0950946
R22002 VDD.n3882 VDD.n3881 0.0950946
R22003 VDD.n3088 VDD.n3087 0.0950946
R22004 VDD.n3080 VDD.n3079 0.0950946
R22005 VDD.n2272 VDD.n2271 0.0950946
R22006 VDD.n2264 VDD.n2263 0.0950946
R22007 VDD.n1501 VDD.n1500 0.0950946
R22008 VDD.n1493 VDD.n1492 0.0950946
R22009 VDD.n79 VDD.n63 0.0890417
R22010 VDD.n43 VDD.n42 0.0877396
R22011 VDD.n86 VDD.n81 0.0867212
R22012 VDD.n3902 VDD.n3898 0.0838333
R22013 VDD.n3099 VDD.n3095 0.0838333
R22014 VDD.n2283 VDD.n2279 0.0838333
R22015 VDD.n1511 VDD.n1508 0.0838333
R22016 VDD.n704 VDD.n700 0.0838333
R22017 VDD.n4674 VDD.n4673 0.0812292
R22018 VDD.n3889 VDD.n3888 0.0812292
R22019 VDD.n3086 VDD.n3085 0.0812292
R22020 VDD.n2270 VDD.n2269 0.0812292
R22021 VDD.n1499 VDD.n1498 0.0812292
R22022 VDD.n438 VDD.n437 0.0761154
R22023 VDD.n4615 VDD.n3895 0.0760208
R22024 VDD.n3828 VDD.n3092 0.0760208
R22025 VDD.n3030 VDD.n2276 0.0760208
R22026 VDD.n2142 VDD.n1505 0.0760208
R22027 VDD.n1374 VDD.n697 0.0760208
R22028 VDD.n4668 VDD.n4662 0.0708125
R22029 VDD.n3883 VDD.n3877 0.0708125
R22030 VDD.n3081 VDD.n3075 0.0708125
R22031 VDD.n2265 VDD.n2259 0.0708125
R22032 VDD.n1494 VDD.n1488 0.0708125
R22033 VDD.n4663 VDD.n3896 0.0680676
R22034 VDD.n4665 VDD.n4663 0.0680676
R22035 VDD.n3878 VDD.n3093 0.0680676
R22036 VDD.n3880 VDD.n3878 0.0680676
R22037 VDD.n3076 VDD.n2277 0.0680676
R22038 VDD.n3078 VDD.n3076 0.0680676
R22039 VDD.n2260 VDD.n1506 0.0680676
R22040 VDD.n2262 VDD.n2260 0.0680676
R22041 VDD.n1489 VDD.n698 0.0680676
R22042 VDD.n1491 VDD.n1489 0.0680676
R22043 VDD.n290 VDD.n197 0.0678077
R22044 VDD.n85 VDD.n82 0.0672614
R22045 VDD.n8 VDD.n5 0.0672614
R22046 VDD.n3117 VDD.n3116 0.065895
R22047 VDD.n344 VDD.n343 0.0656042
R22048 VDD.n435 VDD.n344 0.0656042
R22049 VDD.n4664 VDD.n3894 0.0574697
R22050 VDD.n3879 VDD.n3091 0.0574697
R22051 VDD.n3077 VDD.n2275 0.0574697
R22052 VDD.n2261 VDD.n1504 0.0574697
R22053 VDD.n1490 VDD.n696 0.0574697
R22054 VDD.n442 VDD.n339 0.0557885
R22055 VDD.n438 VDD.n339 0.0557885
R22056 VDD.n429 VDD.n343 0.0551875
R22057 VDD.n2760 VDD.n2450 0.0512937
R22058 VDD.n2769 VDD.n2448 0.0512937
R22059 VDD.n4669 VDD.n4668 0.0499792
R22060 VDD.n3884 VDD.n3883 0.0499792
R22061 VDD.n3082 VDD.n3081 0.0499792
R22062 VDD.n2266 VDD.n2265 0.0499792
R22063 VDD.n1495 VDD.n1494 0.0499792
R22064 VDD.n3897 VDD.n3895 0.0447708
R22065 VDD.n3094 VDD.n3092 0.0447708
R22066 VDD.n2278 VDD.n2276 0.0447708
R22067 VDD.n1507 VDD.n1505 0.0447708
R22068 VDD.n699 VDD.n697 0.0447708
R22069 VDD.n182 VDD.n88 0.0435147
R22070 VDD.n146 VDD.n89 0.0435147
R22071 VDD.n4675 VDD.n3896 0.0410405
R22072 VDD.n4666 VDD.n4665 0.0410405
R22073 VDD.n3890 VDD.n3093 0.0410405
R22074 VDD.n3881 VDD.n3880 0.0410405
R22075 VDD.n3087 VDD.n2277 0.0410405
R22076 VDD.n3079 VDD.n3078 0.0410405
R22077 VDD.n2271 VDD.n1506 0.0410405
R22078 VDD.n2263 VDD.n2262 0.0410405
R22079 VDD.n1500 VDD.n698 0.0410405
R22080 VDD.n1492 VDD.n1491 0.0410405
R22081 VDD.n156 VDD.n130 0.0405735
R22082 VDD.n4674 VDD.n3897 0.0395625
R22083 VDD.n3889 VDD.n3094 0.0395625
R22084 VDD.n3086 VDD.n2278 0.0395625
R22085 VDD.n2270 VDD.n1507 0.0395625
R22086 VDD.n1499 VDD.n699 0.0395625
R22087 VDD.n4669 VDD.n3902 0.0343542
R22088 VDD.n3884 VDD.n3099 0.0343542
R22089 VDD.n3082 VDD.n2283 0.0343542
R22090 VDD.n2266 VDD.n1511 0.0343542
R22091 VDD.n1495 VDD.n704 0.0343542
R22092 VDD.n43 VDD.n27 0.0330521
R22093 VDD.n408 VDD.n407 0.03175
R22094 VDD.n79 VDD.n78 0.03175
R22095 VDD.n4679 VDD 0.0297281
R22096 VDD.n1502 VDD.n696 0.0292489
R22097 VDD.n1490 VDD.n4 0.0292489
R22098 VDD.n2273 VDD.n1504 0.0292489
R22099 VDD.n2261 VDD.n3 0.0292489
R22100 VDD.n3089 VDD.n2275 0.0292489
R22101 VDD.n3077 VDD.n2 0.0292489
R22102 VDD.n3892 VDD.n3091 0.0292489
R22103 VDD.n3879 VDD.n1 0.0292489
R22104 VDD.n4677 VDD.n3894 0.0292489
R22105 VDD.n4664 VDD.n0 0.0292489
R22106 VDD.n443 VDD.n442 0.0287452
R22107 VDD VDD.n4679 0.027848
R22108 VDD.n443 VDD.n338 0.0275433
R22109 VDD VDD.n4678 0.0256491
R22110 VDD.n692 VDD.n606 0.0239375
R22111 VDD.n604 VDD.n525 0.0239375
R22112 VDD.n524 VDD.n445 0.0239375
R22113 VDD.n4679 VDD 0.00945938
R22114 VDD.n4679 VDD 0.00888304
R22115 VDD.n212 VDD.n187 0.00530769
R22116 VDD.n4673 VDD.n3898 0.00310417
R22117 VDD.n3888 VDD.n3095 0.00310417
R22118 VDD.n3085 VDD.n2279 0.00310417
R22119 VDD.n2269 VDD.n1508 0.00310417
R22120 VDD.n1498 VDD.n700 0.00310417
R22121 a_2324_44458.n43 a_2324_44458.n41 333.392
R22122 a_2324_44458.n43 a_2324_44458.n42 301.392
R22123 a_2324_44458.n45 a_2324_44458.n44 301.392
R22124 a_2324_44458.n47 a_2324_44458.n46 301.392
R22125 a_2324_44458.n38 a_2324_44458.n37 301.392
R22126 a_2324_44458.n40 a_2324_44458.n39 301.392
R22127 a_2324_44458.n49 a_2324_44458.n48 301.392
R22128 a_2324_44458.n36 a_2324_44458.n35 297.808
R22129 a_2324_44458.n2 a_2324_44458.n0 248.638
R22130 a_2324_44458.n2 a_2324_44458.n1 203.463
R22131 a_2324_44458.n4 a_2324_44458.n3 203.463
R22132 a_2324_44458.n8 a_2324_44458.n7 203.463
R22133 a_2324_44458.n32 a_2324_44458.n31 203.463
R22134 a_2324_44458.n18 a_2324_44458.n17 203.149
R22135 a_2324_44458.n6 a_2324_44458.n5 202.456
R22136 a_2324_44458.n34 a_2324_44458.n33 200.212
R22137 a_2324_44458.n27 a_2324_44458.n22 197.921
R22138 a_2324_44458.n18 a_2324_44458.n13 190.501
R22139 a_2324_44458.n29 a_2324_44458.n9 188.201
R22140 a_2324_44458.n10 a_2324_44458.t59 184.768
R22141 a_2324_44458.n11 a_2324_44458.t41 184.768
R22142 a_2324_44458.n12 a_2324_44458.t45 184.768
R22143 a_2324_44458.n13 a_2324_44458.t61 184.768
R22144 a_2324_44458.n14 a_2324_44458.t35 184.768
R22145 a_2324_44458.n15 a_2324_44458.t63 184.768
R22146 a_2324_44458.n16 a_2324_44458.t40 184.768
R22147 a_2324_44458.n17 a_2324_44458.t50 184.768
R22148 a_2324_44458.n22 a_2324_44458.t55 184.768
R22149 a_2324_44458.n21 a_2324_44458.t57 184.768
R22150 a_2324_44458.n20 a_2324_44458.t62 184.768
R22151 a_2324_44458.n19 a_2324_44458.t43 184.768
R22152 a_2324_44458.n23 a_2324_44458.t49 184.768
R22153 a_2324_44458.n24 a_2324_44458.t39 184.768
R22154 a_2324_44458.n25 a_2324_44458.t48 184.768
R22155 a_2324_44458.n26 a_2324_44458.t34 184.768
R22156 a_2324_44458.n27 a_2324_44458.n26 181.365
R22157 a_2324_44458.n10 a_2324_44458.t53 146.208
R22158 a_2324_44458.n11 a_2324_44458.t58 146.208
R22159 a_2324_44458.n12 a_2324_44458.t36 146.208
R22160 a_2324_44458.n13 a_2324_44458.t60 146.208
R22161 a_2324_44458.n14 a_2324_44458.t47 146.208
R22162 a_2324_44458.n15 a_2324_44458.t56 146.208
R22163 a_2324_44458.n16 a_2324_44458.t51 146.208
R22164 a_2324_44458.n17 a_2324_44458.t54 146.208
R22165 a_2324_44458.n22 a_2324_44458.t44 146.208
R22166 a_2324_44458.n21 a_2324_44458.t33 146.208
R22167 a_2324_44458.n20 a_2324_44458.t32 146.208
R22168 a_2324_44458.n19 a_2324_44458.t37 146.208
R22169 a_2324_44458.n23 a_2324_44458.t52 146.208
R22170 a_2324_44458.n24 a_2324_44458.t42 146.208
R22171 a_2324_44458.n25 a_2324_44458.t38 146.208
R22172 a_2324_44458.n26 a_2324_44458.t46 146.208
R22173 a_2324_44458.n4 a_2324_44458.n2 45.177
R22174 a_2324_44458.n30 a_2324_44458.n8 45.177
R22175 a_2324_44458.n32 a_2324_44458.n30 45.177
R22176 a_2324_44458.n6 a_2324_44458.n4 44.0476
R22177 a_2324_44458.n8 a_2324_44458.n6 44.0476
R22178 a_2324_44458.n11 a_2324_44458.n10 40.6397
R22179 a_2324_44458.n12 a_2324_44458.n11 40.6397
R22180 a_2324_44458.n13 a_2324_44458.n12 40.6397
R22181 a_2324_44458.n15 a_2324_44458.n14 40.6397
R22182 a_2324_44458.n16 a_2324_44458.n15 40.6397
R22183 a_2324_44458.n17 a_2324_44458.n16 40.6397
R22184 a_2324_44458.n22 a_2324_44458.n21 40.6397
R22185 a_2324_44458.n21 a_2324_44458.n20 40.6397
R22186 a_2324_44458.n20 a_2324_44458.n19 40.6397
R22187 a_2324_44458.n24 a_2324_44458.n23 40.6397
R22188 a_2324_44458.n25 a_2324_44458.n24 40.6397
R22189 a_2324_44458.n26 a_2324_44458.n25 40.6397
R22190 a_2324_44458.n0 a_2324_44458.t24 40.0005
R22191 a_2324_44458.n0 a_2324_44458.t22 40.0005
R22192 a_2324_44458.n1 a_2324_44458.t26 40.0005
R22193 a_2324_44458.n1 a_2324_44458.t30 40.0005
R22194 a_2324_44458.n3 a_2324_44458.t29 40.0005
R22195 a_2324_44458.n3 a_2324_44458.t25 40.0005
R22196 a_2324_44458.n5 a_2324_44458.t21 40.0005
R22197 a_2324_44458.n5 a_2324_44458.t28 40.0005
R22198 a_2324_44458.n7 a_2324_44458.t23 40.0005
R22199 a_2324_44458.n7 a_2324_44458.t16 40.0005
R22200 a_2324_44458.n9 a_2324_44458.t18 40.0005
R22201 a_2324_44458.n9 a_2324_44458.t31 40.0005
R22202 a_2324_44458.n31 a_2324_44458.t17 40.0005
R22203 a_2324_44458.n31 a_2324_44458.t19 40.0005
R22204 a_2324_44458.n33 a_2324_44458.t27 40.0005
R22205 a_2324_44458.n33 a_2324_44458.t20 40.0005
R22206 a_2324_44458.n45 a_2324_44458.n43 32.0005
R22207 a_2324_44458.n47 a_2324_44458.n45 32.0005
R22208 a_2324_44458.n40 a_2324_44458.n38 32.0005
R22209 a_2324_44458.n48 a_2324_44458.n40 32.0005
R22210 a_2324_44458.n48 a_2324_44458.n47 31.2005
R22211 a_2324_44458.n28 a_2324_44458.n18 29.3721
R22212 a_2324_44458.n41 a_2324_44458.t4 27.5805
R22213 a_2324_44458.n41 a_2324_44458.t13 27.5805
R22214 a_2324_44458.n42 a_2324_44458.t14 27.5805
R22215 a_2324_44458.n42 a_2324_44458.t12 27.5805
R22216 a_2324_44458.n44 a_2324_44458.t7 27.5805
R22217 a_2324_44458.n44 a_2324_44458.t6 27.5805
R22218 a_2324_44458.n46 a_2324_44458.t8 27.5805
R22219 a_2324_44458.n46 a_2324_44458.t11 27.5805
R22220 a_2324_44458.n37 a_2324_44458.t2 27.5805
R22221 a_2324_44458.n37 a_2324_44458.t9 27.5805
R22222 a_2324_44458.n35 a_2324_44458.t10 27.5805
R22223 a_2324_44458.n35 a_2324_44458.t3 27.5805
R22224 a_2324_44458.n39 a_2324_44458.t5 27.5805
R22225 a_2324_44458.n39 a_2324_44458.t0 27.5805
R22226 a_2324_44458.n49 a_2324_44458.t1 27.5805
R22227 a_2324_44458.t15 a_2324_44458.n49 27.5805
R22228 a_2324_44458.n28 a_2324_44458.n27 26.0403
R22229 a_2324_44458.n30 a_2324_44458.n29 15.262
R22230 a_2324_44458.n34 a_2324_44458.n32 13.177
R22231 a_2324_44458.n38 a_2324_44458.n36 10.2022
R22232 a_2324_44458.n29 a_2324_44458.n28 9.3005
R22233 a_2324_44458.n36 a_2324_44458.n34 8.68033
R22234 CAL_N.n6 CAL_N.n5 600.609
R22235 CAL_N.n6 CAL_N.t1 260.137
R22236 CAL_N CAL_N.t4 138.526
R22237 CAL_N.n5 CAL_N.t2 77.3934
R22238 CAL_N.n5 CAL_N.t0 77.3934
R22239 CAL_N.n1 CAL_N.t5 36.3712
R22240 CAL_N.n2 CAL_N.t5 36.3712
R22241 CAL_N.n3 CAL_N.t6 36.2721
R22242 CAL_N.t6 CAL_N.n0 36.2721
R22243 CAL_N.n2 CAL_N.t3 31.2287
R22244 CAL_N.t3 CAL_N.n1 31.2287
R22245 CAL_N CAL_N.n7 27.5511
R22246 CAL_N.n7 CAL_N.n6 10.1411
R22247 CAL_N.n4 CAL_N.n0 8.938
R22248 CAL_N.n4 CAL_N.n3 4.5005
R22249 CAL_N.n1 CAL_N.n0 0.0713333
R22250 CAL_N.n3 CAL_N.n2 0.0713333
R22251 CAL_N.n7 CAL_N.n4 0.0213333
R22252 a_3080_42308.n1 a_3080_42308.t6 580.173
R22253 a_3080_42308.n1 a_3080_42308.t7 579.144
R22254 a_3080_42308.n5 a_3080_42308.n4 380.32
R22255 a_3080_42308.n0 a_3080_42308.t5 260.322
R22256 a_3080_42308.n4 a_3080_42308.n3 185
R22257 a_3080_42308.n2 a_3080_42308.n0 177.798
R22258 a_3080_42308.n0 a_3080_42308.t4 175.169
R22259 a_3080_42308.n2 a_3080_42308.n1 103.156
R22260 a_3080_42308.t1 a_3080_42308.n5 26.5955
R22261 a_3080_42308.n5 a_3080_42308.t0 26.5955
R22262 a_3080_42308.n3 a_3080_42308.t3 24.9236
R22263 a_3080_42308.n3 a_3080_42308.t2 24.9236
R22264 a_3080_42308.n4 a_3080_42308.n2 21.4656
R22265 a_12861_44030.n27 a_12861_44030.n26 585
R22266 a_12861_44030.n12 a_12861_44030.t32 323.342
R22267 a_12861_44030.n13 a_12861_44030.t31 323.342
R22268 a_12861_44030.n1 a_12861_44030.t34 256.07
R22269 a_12861_44030.n30 a_12861_44030.n28 243.627
R22270 a_12861_44030.n17 a_12861_44030.t33 241.536
R22271 a_12861_44030.n0 a_12861_44030.t26 231.835
R22272 a_12861_44030.n19 a_12861_44030.t11 222.018
R22273 a_12861_44030.n5 a_12861_44030.t29 212.081
R22274 a_12861_44030.n9 a_12861_44030.t21 212.081
R22275 a_12861_44030.n8 a_12861_44030.t13 212.081
R22276 a_12861_44030.n7 a_12861_44030.t25 212.081
R22277 a_12861_44030.n21 a_12861_44030.t14 212.081
R22278 a_12861_44030.n22 a_12861_44030.t35 212.081
R22279 a_12861_44030.n30 a_12861_44030.n29 200.262
R22280 a_12861_44030.n12 a_12861_44030.t28 194.809
R22281 a_12861_44030.n13 a_12861_44030.t19 194.809
R22282 a_12861_44030.n32 a_12861_44030.n31 194.441
R22283 a_12861_44030.n18 a_12861_44030.n17 194.054
R22284 a_12861_44030.n23 a_12861_44030.n22 194.022
R22285 a_12861_44030.n15 a_12861_44030.n14 180.338
R22286 a_12861_44030.n2 a_12861_44030.n0 178.286
R22287 a_12861_44030.n4 a_12861_44030.n3 177.452
R22288 a_12861_44030.n2 a_12861_44030.n1 173.536
R22289 a_12861_44030.n17 a_12861_44030.t16 169.237
R22290 a_12861_44030.n16 a_12861_44030.n12 167.474
R22291 a_12861_44030.n15 a_12861_44030.n13 166.852
R22292 a_12861_44030.n11 a_12861_44030.n6 164.161
R22293 a_12861_44030.n0 a_12861_44030.t24 157.07
R22294 a_12861_44030.n1 a_12861_44030.t10 150.03
R22295 a_12861_44030.n3 a_12861_44030.t22 147.298
R22296 a_12861_44030.n14 a_12861_44030.t17 142.994
R22297 a_12861_44030.n19 a_12861_44030.t8 140.064
R22298 a_12861_44030.n5 a_12861_44030.t9 139.78
R22299 a_12861_44030.n9 a_12861_44030.t12 139.78
R22300 a_12861_44030.n8 a_12861_44030.t15 139.78
R22301 a_12861_44030.n7 a_12861_44030.t20 139.78
R22302 a_12861_44030.n21 a_12861_44030.t27 139.78
R22303 a_12861_44030.n22 a_12861_44030.t18 139.78
R22304 a_12861_44030.n3 a_12861_44030.t30 131.231
R22305 a_12861_44030.n14 a_12861_44030.t23 126.927
R22306 a_12861_44030.n20 a_12861_44030.n19 103.41
R22307 a_12861_44030.n10 a_12861_44030.n8 83.6
R22308 a_12861_44030.n31 a_12861_44030.n27 62.148
R22309 a_12861_44030.n8 a_12861_44030.n7 61.346
R22310 a_12861_44030.n22 a_12861_44030.n21 61.346
R22311 a_12861_44030.n11 a_12861_44030.n10 53.9823
R22312 a_12861_44030.n31 a_12861_44030.n30 50.5705
R22313 a_12861_44030.n9 a_12861_44030.n6 47.4702
R22314 a_12861_44030.n28 a_12861_44030.t6 40.0005
R22315 a_12861_44030.n28 a_12861_44030.t5 40.0005
R22316 a_12861_44030.n29 a_12861_44030.t4 40.0005
R22317 a_12861_44030.n29 a_12861_44030.t7 40.0005
R22318 a_12861_44030.n10 a_12861_44030.n9 36.3622
R22319 a_12861_44030.n26 a_12861_44030.t0 27.5805
R22320 a_12861_44030.n26 a_12861_44030.t1 27.5805
R22321 a_12861_44030.n32 a_12861_44030.t2 27.5805
R22322 a_12861_44030.t3 a_12861_44030.n32 27.5805
R22323 a_12861_44030.n20 a_12861_44030.n18 19.4085
R22324 a_12861_44030.n27 a_12861_44030.n25 19.1246
R22325 a_12861_44030.n6 a_12861_44030.n5 13.8763
R22326 a_12861_44030.n16 a_12861_44030.n15 12.8523
R22327 a_12861_44030.n25 a_12861_44030.n4 12.573
R22328 a_12861_44030.n18 a_12861_44030.n16 11.2024
R22329 a_12861_44030.n24 a_12861_44030.n11 9.3005
R22330 a_12861_44030.n23 a_12861_44030.n20 6.45533
R22331 a_12861_44030.n25 a_12861_44030.n24 5.8051
R22332 a_12861_44030.n24 a_12861_44030.n23 4.82775
R22333 a_12861_44030.n4 a_12861_44030.n2 4.4333
R22334 a_526_44458.n14 a_526_44458.t34 722.096
R22335 a_526_44458.n10 a_526_44458.t28 722.096
R22336 a_526_44458.n11 a_526_44458.t15 722.096
R22337 a_526_44458.n35 a_526_44458.n34 585
R22338 a_526_44458.n2 a_526_44458.n0 243.627
R22339 a_526_44458.n8 a_526_44458.t20 241.536
R22340 a_526_44458.n13 a_526_44458.t22 241.536
R22341 a_526_44458.n18 a_526_44458.t13 239.505
R22342 a_526_44458.n32 a_526_44458.t32 230.923
R22343 a_526_44458.n17 a_526_44458.t17 230.923
R22344 a_526_44458.n5 a_526_44458.t11 212.081
R22345 a_526_44458.n6 a_526_44458.t16 212.081
R22346 a_526_44458.n21 a_526_44458.t18 212.081
R22347 a_526_44458.n23 a_526_44458.t21 212.081
R22348 a_526_44458.n25 a_526_44458.t10 212.081
R22349 a_526_44458.n26 a_526_44458.t8 212.081
R22350 a_526_44458.n12 a_526_44458.n11 210.018
R22351 a_526_44458.n2 a_526_44458.n1 200.262
R22352 a_526_44458.n9 a_526_44458.n8 194.542
R22353 a_526_44458.n4 a_526_44458.n3 194.441
R22354 a_526_44458.n19 a_526_44458.n17 190.97
R22355 a_526_44458.n33 a_526_44458.n32 187.987
R22356 a_526_44458.n9 a_526_44458.n7 184.34
R22357 a_526_44458.n15 a_526_44458.n14 181.435
R22358 a_526_44458.n22 a_526_44458.n20 173.505
R22359 a_526_44458.n19 a_526_44458.n18 172.496
R22360 a_526_44458.n8 a_526_44458.t23 169.237
R22361 a_526_44458.n13 a_526_44458.t29 169.237
R22362 a_526_44458.n12 a_526_44458.n10 168.203
R22363 a_526_44458.n18 a_526_44458.t30 167.204
R22364 a_526_44458.n32 a_526_44458.t24 163.881
R22365 a_526_44458.n17 a_526_44458.t9 163.881
R22366 a_526_44458.n14 a_526_44458.t12 162.963
R22367 a_526_44458.n10 a_526_44458.t26 162.963
R22368 a_526_44458.n11 a_526_44458.t14 162.963
R22369 a_526_44458.n15 a_526_44458.n13 162.56
R22370 a_526_44458.n24 a_526_44458.n20 152
R22371 a_526_44458.n5 a_526_44458.t19 139.78
R22372 a_526_44458.n6 a_526_44458.t33 139.78
R22373 a_526_44458.n21 a_526_44458.t31 139.78
R22374 a_526_44458.n23 a_526_44458.t27 139.78
R22375 a_526_44458.n25 a_526_44458.t25 139.78
R22376 a_526_44458.n26 a_526_44458.t35 139.78
R22377 a_526_44458.n28 a_526_44458.n27 80.1844
R22378 a_526_44458.n34 a_526_44458.n4 62.148
R22379 a_526_44458.n4 a_526_44458.n2 50.5705
R22380 a_526_44458.n27 a_526_44458.n25 42.8185
R22381 a_526_44458.n0 a_526_44458.t6 40.0005
R22382 a_526_44458.n0 a_526_44458.t4 40.0005
R22383 a_526_44458.n1 a_526_44458.t7 40.0005
R22384 a_526_44458.n1 a_526_44458.t5 40.0005
R22385 a_526_44458.n7 a_526_44458.n5 30.6732
R22386 a_526_44458.n7 a_526_44458.n6 30.6732
R22387 a_526_44458.n22 a_526_44458.n21 30.6732
R22388 a_526_44458.n23 a_526_44458.n22 30.6732
R22389 a_526_44458.n24 a_526_44458.n23 30.6732
R22390 a_526_44458.n25 a_526_44458.n24 30.6732
R22391 a_526_44458.n3 a_526_44458.t0 27.5805
R22392 a_526_44458.n3 a_526_44458.t2 27.5805
R22393 a_526_44458.t3 a_526_44458.n35 27.5805
R22394 a_526_44458.n35 a_526_44458.t1 27.5805
R22395 a_526_44458.n28 a_526_44458.n20 20.9925
R22396 a_526_44458.n34 a_526_44458.n33 19.0174
R22397 a_526_44458.n29 a_526_44458.n28 17.8209
R22398 a_526_44458.n27 a_526_44458.n26 16.0782
R22399 a_526_44458.n31 a_526_44458.n30 9.48519
R22400 a_526_44458.n16 a_526_44458.n12 7.74861
R22401 a_526_44458.n16 a_526_44458.n15 6.51939
R22402 a_526_44458.n29 a_526_44458.n19 5.28725
R22403 a_526_44458.n33 a_526_44458.n31 4.82742
R22404 a_526_44458.n30 a_526_44458.n16 4.77889
R22405 a_526_44458.n31 a_526_44458.n9 4.5005
R22406 a_526_44458.n30 a_526_44458.n29 0.932667
R22407 a_n755_45592.t14 a_n755_45592.t20 378.255
R22408 a_n755_45592.n7 a_n755_45592.t14 335.993
R22409 a_n755_45592.n14 a_n755_45592.t21 334.723
R22410 a_n755_45592.n19 a_n755_45592.t13 256.726
R22411 a_n755_45592.n23 a_n755_45592.n0 248.088
R22412 a_n755_45592.n17 a_n755_45592.t23 241.536
R22413 a_n755_45592.n6 a_n755_45592.t8 236.18
R22414 a_n755_45592.n15 a_n755_45592.n14 232.254
R22415 a_n755_45592.n12 a_n755_45592.t10 231.835
R22416 a_n755_45592.n5 a_n755_45592.t11 229.369
R22417 a_n755_45592.n24 a_n755_45592.n23 208.507
R22418 a_n755_45592.n14 a_n755_45592.t9 206.19
R22419 a_n755_45592.n13 a_n755_45592.t26 201.369
R22420 a_n755_45592.n18 a_n755_45592.n17 178.436
R22421 a_n755_45592.n11 a_n755_45592.n4 176.713
R22422 a_n755_45592.n17 a_n755_45592.t16 169.237
R22423 a_n755_45592.n20 a_n755_45592.n19 166.964
R22424 a_n755_45592.n8 a_n755_45592.n5 164.893
R22425 a_n755_45592.n6 a_n755_45592.t18 163.881
R22426 a_n755_45592.n16 a_n755_45592.n12 163.84
R22427 a_n755_45592.n7 a_n755_45592.n6 163.168
R22428 a_n755_45592.n10 a_n755_45592.n9 162.837
R22429 a_n755_45592.n15 a_n755_45592.n13 162.315
R22430 a_n755_45592.n19 a_n755_45592.t24 161.275
R22431 a_n755_45592.n5 a_n755_45592.t25 157.07
R22432 a_n755_45592.n12 a_n755_45592.t27 157.07
R22433 a_n755_45592.n4 a_n755_45592.t17 142.994
R22434 a_n755_45592.n3 a_n755_45592.n1 137.575
R22435 a_n755_45592.n9 a_n755_45592.t15 137.177
R22436 a_n755_45592.n13 a_n755_45592.t12 132.282
R22437 a_n755_45592.n4 a_n755_45592.t19 126.927
R22438 a_n755_45592.n9 a_n755_45592.t22 121.109
R22439 a_n755_45592.n3 a_n755_45592.n2 99.1749
R22440 a_n755_45592.n22 a_n755_45592.n3 36.0958
R22441 a_n755_45592.n0 a_n755_45592.t2 26.5955
R22442 a_n755_45592.n0 a_n755_45592.t0 26.5955
R22443 a_n755_45592.n24 a_n755_45592.t1 26.5955
R22444 a_n755_45592.t3 a_n755_45592.n24 26.5955
R22445 a_n755_45592.n1 a_n755_45592.t7 24.9236
R22446 a_n755_45592.n1 a_n755_45592.t5 24.9236
R22447 a_n755_45592.n2 a_n755_45592.t4 24.9236
R22448 a_n755_45592.n2 a_n755_45592.t6 24.9236
R22449 a_n755_45592.n23 a_n755_45592.n22 17.2539
R22450 a_n755_45592.n21 a_n755_45592.n20 15.5609
R22451 a_n755_45592.n18 a_n755_45592.n16 15.1777
R22452 a_n755_45592.n22 a_n755_45592.n21 14.916
R22453 a_n755_45592.n8 a_n755_45592.n7 11.142
R22454 a_n755_45592.n10 a_n755_45592.n8 7.01389
R22455 a_n755_45592.n21 a_n755_45592.n11 5.02935
R22456 a_n755_45592.n11 a_n755_45592.n10 4.79462
R22457 a_n755_45592.n16 a_n755_45592.n15 3.46479
R22458 a_n755_45592.n20 a_n755_45592.n18 2.94963
R22459 a_5937_45572.n17 a_5937_45572.n16 365.022
R22460 a_5937_45572.n0 a_5937_45572.t14 256.07
R22461 a_5937_45572.n11 a_5937_45572.t11 241.536
R22462 a_5937_45572.n10 a_5937_45572.t17 241.536
R22463 a_5937_45572.n2 a_5937_45572.t6 240.484
R22464 a_5937_45572.n6 a_5937_45572.t10 236.18
R22465 a_5937_45572.n7 a_5937_45572.n6 235.887
R22466 a_5937_45572.n1 a_5937_45572.t13 234.483
R22467 a_5937_45572.n8 a_5937_45572.t4 230.155
R22468 a_5937_45572.n3 a_5937_45572.t8 229.369
R22469 a_5937_45572.n4 a_5937_45572.n2 205.026
R22470 a_5937_45572.n12 a_5937_45572.n11 198.696
R22471 a_5937_45572.n16 a_5937_45572.n15 185
R22472 a_5937_45572.n14 a_5937_45572.n0 182.036
R22473 a_5937_45572.n4 a_5937_45572.n3 175.464
R22474 a_5937_45572.n5 a_5937_45572.n1 171.472
R22475 a_5937_45572.n12 a_5937_45572.n10 170.111
R22476 a_5937_45572.n11 a_5937_45572.t18 169.237
R22477 a_5937_45572.n10 a_5937_45572.t5 169.237
R22478 a_5937_45572.n2 a_5937_45572.t19 168.185
R22479 a_5937_45572.n6 a_5937_45572.t12 163.881
R22480 a_5937_45572.n9 a_5937_45572.n8 163.605
R22481 a_5937_45572.n1 a_5937_45572.t7 162.184
R22482 a_5937_45572.n8 a_5937_45572.t15 157.856
R22483 a_5937_45572.n3 a_5937_45572.t16 157.07
R22484 a_5937_45572.n0 a_5937_45572.t9 150.03
R22485 a_5937_45572.n16 a_5937_45572.n14 28.4253
R22486 a_5937_45572.n17 a_5937_45572.t0 26.5955
R22487 a_5937_45572.t1 a_5937_45572.n17 26.5955
R22488 a_5937_45572.n15 a_5937_45572.t2 24.9236
R22489 a_5937_45572.n15 a_5937_45572.t3 24.9236
R22490 a_5937_45572.n13 a_5937_45572.n12 9.12704
R22491 a_5937_45572.n5 a_5937_45572.n4 8.01149
R22492 a_5937_45572.n9 a_5937_45572.n7 7.94796
R22493 a_5937_45572.n14 a_5937_45572.n13 7.30957
R22494 a_5937_45572.n7 a_5937_45572.n5 6.84819
R22495 a_5937_45572.n13 a_5937_45572.n9 4.97578
R22496 a_n1613_43370.n44 a_n1613_43370.n43 585
R22497 a_n1613_43370.n38 a_n1613_43370.t12 408.63
R22498 a_n1613_43370.n34 a_n1613_43370.t36 408.63
R22499 a_n1613_43370.n30 a_n1613_43370.t46 408.63
R22500 a_n1613_43370.n26 a_n1613_43370.t14 408.63
R22501 a_n1613_43370.n22 a_n1613_43370.t9 408.63
R22502 a_n1613_43370.n18 a_n1613_43370.t38 408.63
R22503 a_n1613_43370.n14 a_n1613_43370.t13 408.63
R22504 a_n1613_43370.n11 a_n1613_43370.t8 408.63
R22505 a_n1613_43370.n1 a_n1613_43370.t40 408.63
R22506 a_n1613_43370.n3 a_n1613_43370.t27 408.63
R22507 a_n1613_43370.n35 a_n1613_43370.t28 347.577
R22508 a_n1613_43370.n31 a_n1613_43370.t37 347.577
R22509 a_n1613_43370.n27 a_n1613_43370.t42 347.577
R22510 a_n1613_43370.n23 a_n1613_43370.t41 347.577
R22511 a_n1613_43370.n19 a_n1613_43370.t45 347.577
R22512 a_n1613_43370.n15 a_n1613_43370.t30 347.577
R22513 a_n1613_43370.n12 a_n1613_43370.t23 347.577
R22514 a_n1613_43370.n8 a_n1613_43370.t32 347.577
R22515 a_n1613_43370.n0 a_n1613_43370.t25 347.577
R22516 a_n1613_43370.n4 a_n1613_43370.t43 347.577
R22517 a_n1613_43370.n47 a_n1613_43370.n45 243.627
R22518 a_n1613_43370.n47 a_n1613_43370.n46 200.262
R22519 a_n1613_43370.n49 a_n1613_43370.n48 194.441
R22520 a_n1613_43370.n35 a_n1613_43370.t16 193.337
R22521 a_n1613_43370.n31 a_n1613_43370.t33 193.337
R22522 a_n1613_43370.n27 a_n1613_43370.t20 193.337
R22523 a_n1613_43370.n23 a_n1613_43370.t18 193.337
R22524 a_n1613_43370.n19 a_n1613_43370.t21 193.337
R22525 a_n1613_43370.n15 a_n1613_43370.t10 193.337
R22526 a_n1613_43370.n12 a_n1613_43370.t47 193.337
R22527 a_n1613_43370.n8 a_n1613_43370.t15 193.337
R22528 a_n1613_43370.n0 a_n1613_43370.t26 193.337
R22529 a_n1613_43370.n4 a_n1613_43370.t19 193.337
R22530 a_n1613_43370.n32 a_n1613_43370.n30 167.808
R22531 a_n1613_43370.n20 a_n1613_43370.n18 167.666
R22532 a_n1613_43370.n13 a_n1613_43370.n11 167.666
R22533 a_n1613_43370.n16 a_n1613_43370.n14 167.663
R22534 a_n1613_43370.n5 a_n1613_43370.n3 167.663
R22535 a_n1613_43370.n36 a_n1613_43370.n34 167.607
R22536 a_n1613_43370.n28 a_n1613_43370.n26 167.605
R22537 a_n1613_43370.n24 a_n1613_43370.n22 167.601
R22538 a_n1613_43370.n2 a_n1613_43370.n1 165.072
R22539 a_n1613_43370.n2 a_n1613_43370.n0 163.007
R22540 a_n1613_43370.n24 a_n1613_43370.n23 160.476
R22541 a_n1613_43370.n28 a_n1613_43370.n27 160.476
R22542 a_n1613_43370.n36 a_n1613_43370.n35 160.472
R22543 a_n1613_43370.n32 a_n1613_43370.n31 160.448
R22544 a_n1613_43370.n20 a_n1613_43370.n19 160.415
R22545 a_n1613_43370.n13 a_n1613_43370.n12 160.415
R22546 a_n1613_43370.n16 a_n1613_43370.n15 160.415
R22547 a_n1613_43370.n9 a_n1613_43370.n8 160.415
R22548 a_n1613_43370.n5 a_n1613_43370.n4 160.415
R22549 a_n1613_43370.n39 a_n1613_43370.n38 158.144
R22550 a_n1613_43370.n38 a_n1613_43370.t17 132.282
R22551 a_n1613_43370.n34 a_n1613_43370.t39 132.282
R22552 a_n1613_43370.n30 a_n1613_43370.t35 132.282
R22553 a_n1613_43370.n26 a_n1613_43370.t34 132.282
R22554 a_n1613_43370.n22 a_n1613_43370.t31 132.282
R22555 a_n1613_43370.n18 a_n1613_43370.t11 132.282
R22556 a_n1613_43370.n14 a_n1613_43370.t22 132.282
R22557 a_n1613_43370.n11 a_n1613_43370.t24 132.282
R22558 a_n1613_43370.n1 a_n1613_43370.t29 132.282
R22559 a_n1613_43370.n3 a_n1613_43370.t44 132.282
R22560 a_n1613_43370.n48 a_n1613_43370.n44 62.148
R22561 a_n1613_43370.n48 a_n1613_43370.n47 50.5705
R22562 a_n1613_43370.n45 a_n1613_43370.t4 40.0005
R22563 a_n1613_43370.n45 a_n1613_43370.t6 40.0005
R22564 a_n1613_43370.n46 a_n1613_43370.t7 40.0005
R22565 a_n1613_43370.n46 a_n1613_43370.t5 40.0005
R22566 a_n1613_43370.n7 a_n1613_43370.n6 37.2419
R22567 a_n1613_43370.n40 a_n1613_43370.n39 27.7325
R22568 a_n1613_43370.n43 a_n1613_43370.t1 27.5805
R22569 a_n1613_43370.n43 a_n1613_43370.t0 27.5805
R22570 a_n1613_43370.t3 a_n1613_43370.n49 27.5805
R22571 a_n1613_43370.n49 a_n1613_43370.t2 27.5805
R22572 a_n1613_43370.n33 a_n1613_43370.n29 20.2065
R22573 a_n1613_43370.n42 a_n1613_43370.n41 18.1475
R22574 a_n1613_43370.n44 a_n1613_43370.n42 17.4996
R22575 a_n1613_43370.n6 a_n1613_43370.n2 15.7922
R22576 a_n1613_43370.n17 a_n1613_43370.n16 15.1253
R22577 a_n1613_43370.n29 a_n1613_43370.n25 13.6063
R22578 a_n1613_43370.n37 a_n1613_43370.n33 11.2337
R22579 a_n1613_43370.n33 a_n1613_43370.n32 10.8046
R22580 a_n1613_43370.n39 a_n1613_43370.n10 9.3005
R22581 a_n1613_43370.n17 a_n1613_43370.n13 7.1494
R22582 a_n1613_43370.n40 a_n1613_43370.n37 6.47943
R22583 a_n1613_43370.n25 a_n1613_43370.n24 5.7653
R22584 a_n1613_43370.n42 a_n1613_43370.n7 5.27935
R22585 a_n1613_43370.n21 a_n1613_43370.n20 4.54912
R22586 a_n1613_43370.n10 a_n1613_43370.n9 2.54314
R22587 a_n1613_43370.n21 a_n1613_43370.n17 2.29171
R22588 a_n1613_43370.n25 a_n1613_43370.n21 1.69006
R22589 a_n1613_43370.n29 a_n1613_43370.n28 1.33124
R22590 a_n1613_43370.n9 a_n1613_43370.n7 0.62234
R22591 a_n1613_43370.n41 a_n1613_43370.n10 0.175249
R22592 a_n1613_43370.n37 a_n1613_43370.n36 0.141324
R22593 a_n1613_43370.n6 a_n1613_43370.n5 0.0498813
R22594 a_n1613_43370.n41 a_n1613_43370.n40 0.0101154
R22595 a_16327_47482.n44 a_16327_47482.n0 647.148
R22596 a_16327_47482.n38 a_16327_47482.t19 408.63
R22597 a_16327_47482.n33 a_16327_47482.t16 408.63
R22598 a_16327_47482.n23 a_16327_47482.t33 408.63
R22599 a_16327_47482.n18 a_16327_47482.t43 408.63
R22600 a_16327_47482.n11 a_16327_47482.t12 408.63
R22601 a_16327_47482.n14 a_16327_47482.t42 408.63
R22602 a_16327_47482.n28 a_16327_47482.t13 408.63
R22603 a_16327_47482.n8 a_16327_47482.t24 408.63
R22604 a_16327_47482.n4 a_16327_47482.t44 408.63
R22605 a_16327_47482.n39 a_16327_47482.t39 347.577
R22606 a_16327_47482.n34 a_16327_47482.t22 347.577
R22607 a_16327_47482.n24 a_16327_47482.t30 347.577
R22608 a_16327_47482.n19 a_16327_47482.t11 347.577
R22609 a_16327_47482.n12 a_16327_47482.t35 347.577
R22610 a_16327_47482.n15 a_16327_47482.t25 347.577
R22611 a_16327_47482.n29 a_16327_47482.t45 347.577
R22612 a_16327_47482.n7 a_16327_47482.t29 347.577
R22613 a_16327_47482.n5 a_16327_47482.t21 347.577
R22614 a_16327_47482.n10 a_16327_47482.t26 256.07
R22615 a_16327_47482.n3 a_16327_47482.n1 243.627
R22616 a_16327_47482.n3 a_16327_47482.n2 200.262
R22617 a_16327_47482.n45 a_16327_47482.n44 194.441
R22618 a_16327_47482.n39 a_16327_47482.t41 193.337
R22619 a_16327_47482.n34 a_16327_47482.t32 193.337
R22620 a_16327_47482.n24 a_16327_47482.t10 193.337
R22621 a_16327_47482.n19 a_16327_47482.t20 193.337
R22622 a_16327_47482.n12 a_16327_47482.t9 193.337
R22623 a_16327_47482.n15 a_16327_47482.t34 193.337
R22624 a_16327_47482.n29 a_16327_47482.t15 193.337
R22625 a_16327_47482.n7 a_16327_47482.t40 193.337
R22626 a_16327_47482.n5 a_16327_47482.t36 193.337
R22627 a_16327_47482.n22 a_16327_47482.n10 191.189
R22628 a_16327_47482.n16 a_16327_47482.n14 167.666
R22629 a_16327_47482.n6 a_16327_47482.n4 167.666
R22630 a_16327_47482.n20 a_16327_47482.n18 167.663
R22631 a_16327_47482.n40 a_16327_47482.n38 167.601
R22632 a_16327_47482.n35 a_16327_47482.n33 167.601
R22633 a_16327_47482.n9 a_16327_47482.n8 165.935
R22634 a_16327_47482.n25 a_16327_47482.n23 165.934
R22635 a_16327_47482.n13 a_16327_47482.n11 165.049
R22636 a_16327_47482.n13 a_16327_47482.n12 163.196
R22637 a_16327_47482.n30 a_16327_47482.n29 162.957
R22638 a_16327_47482.n9 a_16327_47482.n7 162.014
R22639 a_16327_47482.n25 a_16327_47482.n24 162.012
R22640 a_16327_47482.n40 a_16327_47482.n39 160.476
R22641 a_16327_47482.n35 a_16327_47482.n34 160.476
R22642 a_16327_47482.n16 a_16327_47482.n15 160.415
R22643 a_16327_47482.n6 a_16327_47482.n5 160.415
R22644 a_16327_47482.n20 a_16327_47482.n19 160.415
R22645 a_16327_47482.n31 a_16327_47482.n28 158.144
R22646 a_16327_47482.n10 a_16327_47482.t27 150.03
R22647 a_16327_47482.n38 a_16327_47482.t23 132.282
R22648 a_16327_47482.n33 a_16327_47482.t14 132.282
R22649 a_16327_47482.n23 a_16327_47482.t28 132.282
R22650 a_16327_47482.n18 a_16327_47482.t8 132.282
R22651 a_16327_47482.n11 a_16327_47482.t37 132.282
R22652 a_16327_47482.n14 a_16327_47482.t18 132.282
R22653 a_16327_47482.n28 a_16327_47482.t17 132.282
R22654 a_16327_47482.n8 a_16327_47482.t31 132.282
R22655 a_16327_47482.n4 a_16327_47482.t38 132.282
R22656 a_16327_47482.n1 a_16327_47482.t5 40.0005
R22657 a_16327_47482.n1 a_16327_47482.t6 40.0005
R22658 a_16327_47482.n2 a_16327_47482.t4 40.0005
R22659 a_16327_47482.n2 a_16327_47482.t7 40.0005
R22660 a_16327_47482.n43 a_16327_47482.n3 36.5217
R22661 a_16327_47482.n32 a_16327_47482.n31 27.7325
R22662 a_16327_47482.n0 a_16327_47482.t1 27.5805
R22663 a_16327_47482.n0 a_16327_47482.t0 27.5805
R22664 a_16327_47482.n45 a_16327_47482.t2 27.5805
R22665 a_16327_47482.t3 a_16327_47482.n45 27.5805
R22666 a_16327_47482.n21 a_16327_47482.n20 19.121
R22667 a_16327_47482.n17 a_16327_47482.n13 18.7214
R22668 a_16327_47482.n42 a_16327_47482.n41 17.2762
R22669 a_16327_47482.n44 a_16327_47482.n43 14.0492
R22670 a_16327_47482.n43 a_16327_47482.n42 12.5356
R22671 a_16327_47482.n22 a_16327_47482.n21 11.381
R22672 a_16327_47482.n31 a_16327_47482.n30 9.3005
R22673 a_16327_47482.n27 a_16327_47482.n26 9.22577
R22674 a_16327_47482.n41 a_16327_47482.n40 8.42977
R22675 a_16327_47482.n37 a_16327_47482.n9 7.53948
R22676 a_16327_47482.n26 a_16327_47482.n22 5.94006
R22677 a_16327_47482.n41 a_16327_47482.n37 5.49573
R22678 a_16327_47482.n37 a_16327_47482.n36 4.57639
R22679 a_16327_47482.n26 a_16327_47482.n25 4.5005
R22680 a_16327_47482.n36 a_16327_47482.n32 4.37513
R22681 a_16327_47482.n36 a_16327_47482.n35 0.854589
R22682 a_16327_47482.n42 a_16327_47482.n6 0.248745
R22683 a_16327_47482.n21 a_16327_47482.n17 0.200007
R22684 a_16327_47482.n30 a_16327_47482.n27 0.175249
R22685 a_16327_47482.n17 a_16327_47482.n16 0.0492375
R22686 a_16327_47482.n32 a_16327_47482.n27 0.0101154
R22687 a_n443_46116.n19 a_n443_46116.t12 414.432
R22688 a_n443_46116.n4 a_n443_46116.t20 414.432
R22689 a_n443_46116.n19 a_n443_46116.t16 300.349
R22690 a_n443_46116.n4 a_n443_46116.t23 300.349
R22691 a_n443_46116.n10 a_n443_46116.n8 261.344
R22692 a_n443_46116.n22 a_n443_46116.n0 248.088
R22693 a_n443_46116.n6 a_n443_46116.n5 246.228
R22694 a_n443_46116.n7 a_n443_46116.t14 241.536
R22695 a_n443_46116.n14 a_n443_46116.t11 241.536
R22696 a_n443_46116.n8 a_n443_46116.t21 236.18
R22697 a_n443_46116.n5 a_n443_46116.t24 236.18
R22698 a_n443_46116.n9 a_n443_46116.t18 234.392
R22699 a_n443_46116.n11 a_n443_46116.t9 230.155
R22700 a_n443_46116.n17 a_n443_46116.t25 229.369
R22701 a_n443_46116.n23 a_n443_46116.n22 208.507
R22702 a_n443_46116.n13 a_n443_46116.n7 208.482
R22703 a_n443_46116.n15 a_n443_46116.n14 175.294
R22704 a_n443_46116.n7 a_n443_46116.t17 169.237
R22705 a_n443_46116.n14 a_n443_46116.t8 169.237
R22706 a_n443_46116.n18 a_n443_46116.n17 167.459
R22707 a_n443_46116.n12 a_n443_46116.n11 163.899
R22708 a_n443_46116.n8 a_n443_46116.t10 163.881
R22709 a_n443_46116.n5 a_n443_46116.t15 163.881
R22710 a_n443_46116.n11 a_n443_46116.t19 157.856
R22711 a_n443_46116.n17 a_n443_46116.t22 157.07
R22712 a_n443_46116.n10 a_n443_46116.n9 153.165
R22713 a_n443_46116.n9 a_n443_46116.t13 150.442
R22714 a_n443_46116.n3 a_n443_46116.n1 137.575
R22715 a_n443_46116.n3 a_n443_46116.n2 99.1749
R22716 a_n443_46116.n20 a_n443_46116.n19 81.3745
R22717 a_n443_46116.n6 a_n443_46116.n4 64.1409
R22718 a_n443_46116.n21 a_n443_46116.n3 36.0958
R22719 a_n443_46116.n16 a_n443_46116.n6 27.6502
R22720 a_n443_46116.n0 a_n443_46116.t2 26.5955
R22721 a_n443_46116.n0 a_n443_46116.t1 26.5955
R22722 a_n443_46116.n23 a_n443_46116.t0 26.5955
R22723 a_n443_46116.t3 a_n443_46116.n23 26.5955
R22724 a_n443_46116.n1 a_n443_46116.t6 24.9236
R22725 a_n443_46116.n1 a_n443_46116.t4 24.9236
R22726 a_n443_46116.n2 a_n443_46116.t7 24.9236
R22727 a_n443_46116.n2 a_n443_46116.t5 24.9236
R22728 a_n443_46116.n21 a_n443_46116.n20 23.9628
R22729 a_n443_46116.n22 a_n443_46116.n21 17.2539
R22730 a_n443_46116.n16 a_n443_46116.n15 11.3542
R22731 a_n443_46116.n18 a_n443_46116.n16 10.2546
R22732 a_n443_46116.n12 a_n443_46116.n10 10.0053
R22733 a_n443_46116.n20 a_n443_46116.n18 9.36176
R22734 a_n443_46116.n13 a_n443_46116.n12 4.5005
R22735 a_n443_46116.n15 a_n443_46116.n13 3.21135
R22736 a_2437_43646.n1 a_2437_43646.t3 276.464
R22737 a_2437_43646.n2 a_2437_43646.n1 240.409
R22738 a_2437_43646.t0 a_2437_43646.n2 199.456
R22739 a_2437_43646.n1 a_2437_43646.t4 196.131
R22740 a_2437_43646.n2 a_2437_43646.n0 190.911
R22741 a_2437_43646.n0 a_2437_43646.t1 26.5955
R22742 a_2437_43646.n0 a_2437_43646.t2 26.5955
R22743 VDAC_Ni VDAC_Ni.t9 388.632
R22744 VDAC_Ni.n0 VDAC_Ni.t10 231.123
R22745 VDAC_Ni.n3 VDAC_Ni.n1 104.255
R22746 VDAC_Ni.n3 VDAC_Ni.n2 103.96
R22747 VDAC_Ni.n0 VDAC_Ni.t4 50.8513
R22748 VDAC_Ni.n8 VDAC_Ni.n7 37.3168
R22749 VDAC_Ni.n6 VDAC_Ni.n5 37.3168
R22750 VDAC_Ni.n1 VDAC_Ni.t1 16.253
R22751 VDAC_Ni.n1 VDAC_Ni.t2 16.253
R22752 VDAC_Ni.n2 VDAC_Ni.t0 16.253
R22753 VDAC_Ni.n2 VDAC_Ni.t3 16.253
R22754 VDAC_Ni.n7 VDAC_Ni.t7 9.9005
R22755 VDAC_Ni.n7 VDAC_Ni.t8 9.9005
R22756 VDAC_Ni.n5 VDAC_Ni.t5 9.9005
R22757 VDAC_Ni.n5 VDAC_Ni.t6 9.9005
R22758 VDAC_Ni.n9 VDAC_Ni.n8 1.89332
R22759 VDAC_Ni.n4 VDAC_Ni.n0 1.5005
R22760 VDAC_Ni.n4 VDAC_Ni.n3 1.5005
R22761 VDAC_Ni.n6 VDAC_Ni.n4 0.328625
R22762 VDAC_Ni.n8 VDAC_Ni.n6 0.313
R22763 VDAC_Ni.n9 VDAC_Ni 0.016125
R22764 VDAC_Ni VDAC_Ni.n9 0.0112759
R22765 a_n2810_45028.n3 a_n2810_45028.n2 380.32
R22766 a_n2810_45028.n2 a_n2810_45028.n0 263.298
R22767 a_n2810_45028.n0 a_n2810_45028.t5 228.649
R22768 a_n2810_45028.n2 a_n2810_45028.n1 185
R22769 a_n2810_45028.n0 a_n2810_45028.t4 156.35
R22770 a_n2810_45028.t1 a_n2810_45028.n3 26.5955
R22771 a_n2810_45028.n3 a_n2810_45028.t0 26.5955
R22772 a_n2810_45028.n1 a_n2810_45028.t2 24.9236
R22773 a_n2810_45028.n1 a_n2810_45028.t3 24.9236
R22774 a_3626_43646.n5 a_3626_43646.n4 677.66
R22775 a_3626_43646.n4 a_3626_43646.n0 291.856
R22776 a_3626_43646.n2 a_3626_43646.t6 276.464
R22777 a_3626_43646.n3 a_3626_43646.n2 206.565
R22778 a_3626_43646.n2 a_3626_43646.t7 196.131
R22779 a_3626_43646.n3 a_3626_43646.n1 190.487
R22780 a_3626_43646.n4 a_3626_43646.n3 54.5624
R22781 a_3626_43646.n0 a_3626_43646.t2 27.5805
R22782 a_3626_43646.n0 a_3626_43646.t5 27.5805
R22783 a_3626_43646.t1 a_3626_43646.n5 27.5805
R22784 a_3626_43646.n5 a_3626_43646.t0 27.5805
R22785 a_3626_43646.n1 a_3626_43646.t3 25.8467
R22786 a_3626_43646.n1 a_3626_43646.t4 25.8467
R22787 a_14021_43940.n1 a_14021_43940.t1 362.774
R22788 a_14021_43940.t0 a_14021_43940.n1 317.154
R22789 a_14021_43940.n0 a_14021_43940.t3 276.464
R22790 a_14021_43940.n1 a_14021_43940.n0 211.726
R22791 a_14021_43940.n0 a_14021_43940.t2 196.131
R22792 a_21076_30879.n0 a_21076_30879.t5 756.547
R22793 a_21076_30879.n2 a_21076_30879.t7 756.226
R22794 a_21076_30879.n0 a_21076_30879.t4 756.226
R22795 a_21076_30879.n1 a_21076_30879.t6 756.226
R22796 a_21076_30879.n5 a_21076_30879.n4 380.32
R22797 a_21076_30879.n4 a_21076_30879.n3 185
R22798 a_21076_30879.n4 a_21076_30879.n2 110.174
R22799 a_21076_30879.t1 a_21076_30879.n5 26.5955
R22800 a_21076_30879.n5 a_21076_30879.t0 26.5955
R22801 a_21076_30879.n3 a_21076_30879.t3 24.9236
R22802 a_21076_30879.n3 a_21076_30879.t2 24.9236
R22803 a_21076_30879.n1 a_21076_30879.n0 0.3205
R22804 a_21076_30879.n2 a_21076_30879.n1 0.304667
R22805 C8_N_btm C8_N_btm.n8 64.6984
R22806 C8_N_btm.n8 C8_N_btm.n7 43.4801
R22807 C8_N_btm.n2 C8_N_btm.n1 33.0333
R22808 C8_N_btm.n2 C8_N_btm.n0 32.3614
R22809 C8_N_btm.n4 C8_N_btm.n2 21.6828
R22810 C8_N_btm.n4 C8_N_btm.n3 20.8888
R22811 C8_N_btm.n6 C8_N_btm.n5 20.8766
R22812 C8_N_btm.n6 C8_N_btm.n4 11.2088
R22813 C8_N_btm.n7 C8_N_btm.t9 9.9005
R22814 C8_N_btm.n7 C8_N_btm.t8 9.9005
R22815 C8_N_btm.n8 C8_N_btm.n6 8.45883
R22816 C8_N_btm C8_N_btm.n250 5.75597
R22817 C8_N_btm.n0 C8_N_btm.t3 3.57113
R22818 C8_N_btm.n0 C8_N_btm.t2 3.57113
R22819 C8_N_btm.n1 C8_N_btm.t1 3.57113
R22820 C8_N_btm.n1 C8_N_btm.t0 3.57113
R22821 C8_N_btm.n3 C8_N_btm.t6 2.4755
R22822 C8_N_btm.n3 C8_N_btm.t7 2.4755
R22823 C8_N_btm.n5 C8_N_btm.t5 2.4755
R22824 C8_N_btm.n5 C8_N_btm.t4 2.4755
R22825 C8_N_btm.n207 C8_N_btm.n205 0.276161
R22826 C8_N_btm.n227 C8_N_btm.n226 0.276161
R22827 C8_N_btm.n122 C8_N_btm.n90 0.276161
R22828 C8_N_btm.n120 C8_N_btm.n117 0.276161
R22829 C8_N_btm.n94 C8_N_btm.n92 0.276161
R22830 C8_N_btm.n225 C8_N_btm.n195 0.228786
R22831 C8_N_btm.n196 C8_N_btm.n195 0.228786
R22832 C8_N_btm.n197 C8_N_btm.n196 0.228786
R22833 C8_N_btm.n198 C8_N_btm.n197 0.228786
R22834 C8_N_btm.n199 C8_N_btm.n198 0.228786
R22835 C8_N_btm.n200 C8_N_btm.n199 0.228786
R22836 C8_N_btm.n201 C8_N_btm.n200 0.228786
R22837 C8_N_btm.n202 C8_N_btm.n201 0.228786
R22838 C8_N_btm.n203 C8_N_btm.n202 0.228786
R22839 C8_N_btm.n204 C8_N_btm.n203 0.228786
R22840 C8_N_btm.n205 C8_N_btm.n204 0.228786
R22841 C8_N_btm.n226 C8_N_btm.n225 0.228786
R22842 C8_N_btm.n229 C8_N_btm.n228 0.228786
R22843 C8_N_btm.n194 C8_N_btm.n30 0.228786
R22844 C8_N_btm.n193 C8_N_btm.n192 0.228786
R22845 C8_N_btm.n191 C8_N_btm.n33 0.228786
R22846 C8_N_btm.n178 C8_N_btm.n34 0.228786
R22847 C8_N_btm.n90 C8_N_btm.n89 0.228786
R22848 C8_N_btm.n89 C8_N_btm.n88 0.228786
R22849 C8_N_btm.n88 C8_N_btm.n87 0.228786
R22850 C8_N_btm.n87 C8_N_btm.n79 0.228786
R22851 C8_N_btm.n79 C8_N_btm.n78 0.228786
R22852 C8_N_btm.n78 C8_N_btm.n76 0.228786
R22853 C8_N_btm.n76 C8_N_btm.n75 0.228786
R22854 C8_N_btm.n75 C8_N_btm.n74 0.228786
R22855 C8_N_btm.n74 C8_N_btm.n73 0.228786
R22856 C8_N_btm.n100 C8_N_btm.n99 0.228786
R22857 C8_N_btm.n98 C8_N_btm.n95 0.228786
R22858 C8_N_btm.n97 C8_N_btm.n96 0.228786
R22859 C8_N_btm.n59 C8_N_btm.n58 0.228786
R22860 C8_N_btm.n146 C8_N_btm.n145 0.228786
R22861 C8_N_btm.n147 C8_N_btm.n57 0.228786
R22862 C8_N_btm.n152 C8_N_btm.n151 0.228786
R22863 C8_N_btm.n150 C8_N_btm.n55 0.228786
R22864 C8_N_btm.n149 C8_N_btm.n148 0.228786
R22865 C8_N_btm.n50 C8_N_btm.n49 0.228786
R22866 C8_N_btm.n161 C8_N_btm.n160 0.228786
R22867 C8_N_btm.n162 C8_N_btm.n48 0.228786
R22868 C8_N_btm.n165 C8_N_btm.n46 0.228786
R22869 C8_N_btm.n164 C8_N_btm.n163 0.228786
R22870 C8_N_btm.n41 C8_N_btm.n40 0.228786
R22871 C8_N_btm.n176 C8_N_btm.n175 0.228786
R22872 C8_N_btm.n177 C8_N_btm.n39 0.228786
R22873 C8_N_btm.n183 C8_N_btm.n182 0.228786
R22874 C8_N_btm.n181 C8_N_btm.n37 0.228786
R22875 C8_N_btm.n206 C8_N_btm.n11 0.228786
R22876 C8_N_btm.n209 C8_N_btm.n208 0.228786
R22877 C8_N_btm.n12 C8_N_btm.n11 0.228786
R22878 C8_N_btm.n14 C8_N_btm.n12 0.228786
R22879 C8_N_btm.n210 C8_N_btm.n209 0.228786
R22880 C8_N_btm.n211 C8_N_btm.n210 0.228786
R22881 C8_N_btm.n15 C8_N_btm.n14 0.228786
R22882 C8_N_btm.n213 C8_N_btm.n15 0.228786
R22883 C8_N_btm.n212 C8_N_btm.n211 0.228786
R22884 C8_N_btm.n215 C8_N_btm.n212 0.228786
R22885 C8_N_btm.n214 C8_N_btm.n213 0.228786
R22886 C8_N_btm.n214 C8_N_btm.n19 0.228786
R22887 C8_N_btm.n216 C8_N_btm.n215 0.228786
R22888 C8_N_btm.n217 C8_N_btm.n216 0.228786
R22889 C8_N_btm.n20 C8_N_btm.n19 0.228786
R22890 C8_N_btm.n22 C8_N_btm.n20 0.228786
R22891 C8_N_btm.n218 C8_N_btm.n217 0.228786
R22892 C8_N_btm.n219 C8_N_btm.n218 0.228786
R22893 C8_N_btm.n23 C8_N_btm.n22 0.228786
R22894 C8_N_btm.n221 C8_N_btm.n23 0.228786
R22895 C8_N_btm.n220 C8_N_btm.n219 0.228786
R22896 C8_N_btm.n223 C8_N_btm.n220 0.228786
R22897 C8_N_btm.n222 C8_N_btm.n221 0.228786
R22898 C8_N_btm.n26 C8_N_btm.n24 0.228786
R22899 C8_N_btm.n190 C8_N_btm.n28 0.228786
R22900 C8_N_btm.n233 C8_N_btm.n27 0.228786
R22901 C8_N_btm.n234 C8_N_btm.n233 0.228786
R22902 C8_N_btm.n232 C8_N_btm.n26 0.228786
R22903 C8_N_btm.n232 C8_N_btm.n231 0.228786
R22904 C8_N_btm.n230 C8_N_btm.n29 0.228786
R22905 C8_N_btm.n222 C8_N_btm.n29 0.228786
R22906 C8_N_btm.n224 C8_N_btm.n223 0.228786
R22907 C8_N_btm.n224 C8_N_btm.n31 0.228786
R22908 C8_N_btm.n32 C8_N_btm.n31 0.228786
R22909 C8_N_btm.n230 C8_N_btm.n229 0.228786
R22910 C8_N_btm.n231 C8_N_btm.n30 0.228786
R22911 C8_N_btm.n192 C8_N_btm.n27 0.228786
R22912 C8_N_btm.n191 C8_N_btm.n190 0.228786
R22913 C8_N_btm.n189 C8_N_btm.n34 0.228786
R22914 C8_N_btm.n180 C8_N_btm.n179 0.228786
R22915 C8_N_btm.n186 C8_N_btm.n185 0.228786
R22916 C8_N_btm.n184 C8_N_btm.n36 0.228786
R22917 C8_N_btm.n43 C8_N_btm.n38 0.228786
R22918 C8_N_btm.n174 C8_N_btm.n173 0.228786
R22919 C8_N_btm.n172 C8_N_btm.n42 0.228786
R22920 C8_N_btm.n171 C8_N_btm.n44 0.228786
R22921 C8_N_btm.n170 C8_N_btm.n169 0.228786
R22922 C8_N_btm.n168 C8_N_btm.n45 0.228786
R22923 C8_N_btm.n52 C8_N_btm.n47 0.228786
R22924 C8_N_btm.n159 C8_N_btm.n158 0.228786
R22925 C8_N_btm.n157 C8_N_btm.n51 0.228786
R22926 C8_N_btm.n156 C8_N_btm.n53 0.228786
R22927 C8_N_btm.n155 C8_N_btm.n154 0.228786
R22928 C8_N_btm.n153 C8_N_btm.n54 0.228786
R22929 C8_N_btm.n61 C8_N_btm.n56 0.228786
R22930 C8_N_btm.n141 C8_N_btm.n60 0.228786
R22931 C8_N_btm.n144 C8_N_btm.n143 0.228786
R22932 C8_N_btm.n73 C8_N_btm.n62 0.228786
R22933 C8_N_btm.n140 C8_N_btm.n62 0.228786
R22934 C8_N_btm.n140 C8_N_btm.n63 0.228786
R22935 C8_N_btm.n139 C8_N_btm.n65 0.228786
R22936 C8_N_btm.n93 C8_N_btm.n64 0.228786
R22937 C8_N_btm.n137 C8_N_btm.n64 0.228786
R22938 C8_N_btm.n139 C8_N_btm.n138 0.228786
R22939 C8_N_btm.n138 C8_N_btm.n66 0.228786
R22940 C8_N_btm.n137 C8_N_btm.n136 0.228786
R22941 C8_N_btm.n136 C8_N_btm.n135 0.228786
R22942 C8_N_btm.n70 C8_N_btm.n66 0.228786
R22943 C8_N_btm.n133 C8_N_btm.n70 0.228786
R22944 C8_N_btm.n135 C8_N_btm.n134 0.228786
R22945 C8_N_btm.n134 C8_N_btm.n72 0.228786
R22946 C8_N_btm.n133 C8_N_btm.n132 0.228786
R22947 C8_N_btm.n132 C8_N_btm.n131 0.228786
R22948 C8_N_btm.n77 C8_N_btm.n72 0.228786
R22949 C8_N_btm.n129 C8_N_btm.n77 0.228786
R22950 C8_N_btm.n131 C8_N_btm.n130 0.228786
R22951 C8_N_btm.n130 C8_N_btm.n80 0.228786
R22952 C8_N_btm.n129 C8_N_btm.n128 0.228786
R22953 C8_N_btm.n128 C8_N_btm.n127 0.228786
R22954 C8_N_btm.n84 C8_N_btm.n80 0.228786
R22955 C8_N_btm.n125 C8_N_btm.n84 0.228786
R22956 C8_N_btm.n127 C8_N_btm.n126 0.228786
R22957 C8_N_btm.n126 C8_N_btm.n86 0.228786
R22958 C8_N_btm.n125 C8_N_btm.n124 0.228786
R22959 C8_N_btm.n124 C8_N_btm.n123 0.228786
R22960 C8_N_btm.n91 C8_N_btm.n86 0.228786
R22961 C8_N_btm.n121 C8_N_btm.n91 0.228786
R22962 C8_N_btm.n119 C8_N_btm.n118 0.228786
R22963 C8_N_btm.n117 C8_N_btm.n116 0.228786
R22964 C8_N_btm.n118 C8_N_btm.n85 0.228786
R22965 C8_N_btm.n85 C8_N_btm.n83 0.228786
R22966 C8_N_btm.n116 C8_N_btm.n115 0.228786
R22967 C8_N_btm.n115 C8_N_btm.n114 0.228786
R22968 C8_N_btm.n83 C8_N_btm.n82 0.228786
R22969 C8_N_btm.n82 C8_N_btm.n81 0.228786
R22970 C8_N_btm.n114 C8_N_btm.n113 0.228786
R22971 C8_N_btm.n113 C8_N_btm.n112 0.228786
R22972 C8_N_btm.n111 C8_N_btm.n81 0.228786
R22973 C8_N_btm.n111 C8_N_btm.n110 0.228786
R22974 C8_N_btm.n112 C8_N_btm.n109 0.228786
R22975 C8_N_btm.n109 C8_N_btm.n108 0.228786
R22976 C8_N_btm.n110 C8_N_btm.n71 0.228786
R22977 C8_N_btm.n71 C8_N_btm.n69 0.228786
R22978 C8_N_btm.n108 C8_N_btm.n107 0.228786
R22979 C8_N_btm.n107 C8_N_btm.n106 0.228786
R22980 C8_N_btm.n69 C8_N_btm.n68 0.228786
R22981 C8_N_btm.n68 C8_N_btm.n67 0.228786
R22982 C8_N_btm.n106 C8_N_btm.n105 0.228786
R22983 C8_N_btm.n105 C8_N_btm.n104 0.228786
R22984 C8_N_btm.n103 C8_N_btm.n67 0.228786
R22985 C8_N_btm.n103 C8_N_btm.n102 0.228786
R22986 C8_N_btm.n104 C8_N_btm.n92 0.228786
R22987 C8_N_btm.n102 C8_N_btm.n101 0.228786
R22988 C8_N_btm.n100 C8_N_btm.n93 0.228786
R22989 C8_N_btm.n95 C8_N_btm.n65 0.228786
R22990 C8_N_btm.n96 C8_N_btm.n63 0.228786
R22991 C8_N_btm.n60 C8_N_btm.n59 0.228786
R22992 C8_N_btm.n145 C8_N_btm.n144 0.228786
R22993 C8_N_btm.n57 C8_N_btm.n56 0.228786
R22994 C8_N_btm.n153 C8_N_btm.n152 0.228786
R22995 C8_N_btm.n154 C8_N_btm.n55 0.228786
R22996 C8_N_btm.n148 C8_N_btm.n53 0.228786
R22997 C8_N_btm.n51 C8_N_btm.n50 0.228786
R22998 C8_N_btm.n160 C8_N_btm.n159 0.228786
R22999 C8_N_btm.n48 C8_N_btm.n47 0.228786
R23000 C8_N_btm.n168 C8_N_btm.n167 0.228786
R23001 C8_N_btm.n167 C8_N_btm.n166 0.228786
R23002 C8_N_btm.n169 C8_N_btm.n46 0.228786
R23003 C8_N_btm.n163 C8_N_btm.n44 0.228786
R23004 C8_N_btm.n42 C8_N_btm.n41 0.228786
R23005 C8_N_btm.n175 C8_N_btm.n174 0.228786
R23006 C8_N_btm.n39 C8_N_btm.n38 0.228786
R23007 C8_N_btm.n184 C8_N_btm.n183 0.228786
R23008 C8_N_btm.n185 C8_N_btm.n37 0.228786
R23009 C8_N_btm.n179 C8_N_btm.n35 0.228786
R23010 C8_N_btm.n187 C8_N_btm.n35 0.228786
R23011 C8_N_btm.n189 C8_N_btm.n188 0.228786
R23012 C8_N_btm.n235 C8_N_btm.n234 0.228786
R23013 C8_N_btm.n236 C8_N_btm.n235 0.228786
R23014 C8_N_btm.n237 C8_N_btm.n24 0.228786
R23015 C8_N_btm.n238 C8_N_btm.n237 0.228786
R23016 C8_N_btm.n236 C8_N_btm.n21 0.228786
R23017 C8_N_btm.n21 C8_N_btm.n18 0.228786
R23018 C8_N_btm.n239 C8_N_btm.n238 0.228786
R23019 C8_N_btm.n240 C8_N_btm.n239 0.228786
R23020 C8_N_btm.n241 C8_N_btm.n18 0.228786
R23021 C8_N_btm.n242 C8_N_btm.n241 0.228786
R23022 C8_N_btm.n240 C8_N_btm.n17 0.228786
R23023 C8_N_btm.n17 C8_N_btm.n16 0.228786
R23024 C8_N_btm.n243 C8_N_btm.n242 0.228786
R23025 C8_N_btm.n244 C8_N_btm.n243 0.228786
R23026 C8_N_btm.n245 C8_N_btm.n16 0.228786
R23027 C8_N_btm.n246 C8_N_btm.n245 0.228786
R23028 C8_N_btm.n244 C8_N_btm.n13 0.228786
R23029 C8_N_btm.n13 C8_N_btm.n10 0.228786
R23030 C8_N_btm.n247 C8_N_btm.n246 0.228786
R23031 C8_N_btm.n248 C8_N_btm.n247 0.228786
R23032 C8_N_btm.n249 C8_N_btm.n10 0.228786
R23033 C8_N_btm.n250 C8_N_btm.n249 0.228786
R23034 C8_N_btm.n248 C8_N_btm.n9 0.228786
R23035 C8_N_btm.n207 C8_N_btm.n206 0.208893
R23036 C8_N_btm.n228 C8_N_btm.n227 0.208893
R23037 C8_N_btm.n122 C8_N_btm.n121 0.208893
R23038 C8_N_btm.n99 C8_N_btm.n94 0.208893
R23039 C8_N_btm.n142 C8_N_btm.n62 0.208893
R23040 C8_N_btm.n121 C8_N_btm.n120 0.208893
R23041 C8_N_btm.n234 C8_N_btm.n25 0.208893
R23042 C8_N_btm.n223 C8_N_btm.n195 0.09425
R23043 C8_N_btm.n219 C8_N_btm.n197 0.09425
R23044 C8_N_btm.n217 C8_N_btm.n199 0.09425
R23045 C8_N_btm.n215 C8_N_btm.n201 0.09425
R23046 C8_N_btm.n211 C8_N_btm.n203 0.09425
R23047 C8_N_btm.n209 C8_N_btm.n205 0.09425
R23048 C8_N_btm.n206 C8_N_btm.n9 0.09425
R23049 C8_N_btm.n208 C8_N_btm.n11 0.09425
R23050 C8_N_btm.n247 C8_N_btm.n12 0.09425
R23051 C8_N_btm.n209 C8_N_btm.n12 0.09425
R23052 C8_N_btm.n210 C8_N_btm.n14 0.09425
R23053 C8_N_btm.n210 C8_N_btm.n204 0.09425
R23054 C8_N_btm.n245 C8_N_btm.n15 0.09425
R23055 C8_N_btm.n211 C8_N_btm.n15 0.09425
R23056 C8_N_btm.n213 C8_N_btm.n212 0.09425
R23057 C8_N_btm.n212 C8_N_btm.n202 0.09425
R23058 C8_N_btm.n214 C8_N_btm.n17 0.09425
R23059 C8_N_btm.n215 C8_N_btm.n214 0.09425
R23060 C8_N_btm.n216 C8_N_btm.n19 0.09425
R23061 C8_N_btm.n216 C8_N_btm.n200 0.09425
R23062 C8_N_btm.n239 C8_N_btm.n20 0.09425
R23063 C8_N_btm.n217 C8_N_btm.n20 0.09425
R23064 C8_N_btm.n218 C8_N_btm.n22 0.09425
R23065 C8_N_btm.n218 C8_N_btm.n198 0.09425
R23066 C8_N_btm.n237 C8_N_btm.n23 0.09425
R23067 C8_N_btm.n219 C8_N_btm.n23 0.09425
R23068 C8_N_btm.n221 C8_N_btm.n220 0.09425
R23069 C8_N_btm.n220 C8_N_btm.n196 0.09425
R23070 C8_N_btm.n222 C8_N_btm.n26 0.09425
R23071 C8_N_btm.n223 C8_N_btm.n222 0.09425
R23072 C8_N_btm.n190 C8_N_btm.n27 0.09425
R23073 C8_N_btm.n231 C8_N_btm.n27 0.09425
R23074 C8_N_btm.n233 C8_N_btm.n232 0.09425
R23075 C8_N_btm.n232 C8_N_btm.n29 0.09425
R23076 C8_N_btm.n231 C8_N_btm.n230 0.09425
R23077 C8_N_btm.n230 C8_N_btm.n31 0.09425
R23078 C8_N_btm.n224 C8_N_btm.n29 0.09425
R23079 C8_N_btm.n225 C8_N_btm.n224 0.09425
R23080 C8_N_btm.n226 C8_N_btm.n31 0.09425
R23081 C8_N_btm.n229 C8_N_btm.n32 0.09425
R23082 C8_N_btm.n228 C8_N_btm.n194 0.09425
R23083 C8_N_btm.n192 C8_N_btm.n30 0.09425
R23084 C8_N_btm.n229 C8_N_btm.n30 0.09425
R23085 C8_N_btm.n193 C8_N_btm.n33 0.09425
R23086 C8_N_btm.n194 C8_N_btm.n193 0.09425
R23087 C8_N_btm.n191 C8_N_btm.n34 0.09425
R23088 C8_N_btm.n192 C8_N_btm.n191 0.09425
R23089 C8_N_btm.n178 C8_N_btm.n33 0.09425
R23090 C8_N_btm.n180 C8_N_btm.n178 0.09425
R23091 C8_N_btm.n123 C8_N_btm.n91 0.09425
R23092 C8_N_btm.n124 C8_N_btm.n90 0.09425
R23093 C8_N_btm.n88 C8_N_btm.n84 0.09425
R23094 C8_N_btm.n130 C8_N_btm.n79 0.09425
R23095 C8_N_btm.n132 C8_N_btm.n76 0.09425
R23096 C8_N_btm.n74 C8_N_btm.n70 0.09425
R23097 C8_N_btm.n185 C8_N_btm.n35 0.09425
R23098 C8_N_btm.n188 C8_N_btm.n187 0.09425
R23099 C8_N_btm.n186 C8_N_btm.n36 0.09425
R23100 C8_N_btm.n187 C8_N_btm.n186 0.09425
R23101 C8_N_btm.n184 C8_N_btm.n38 0.09425
R23102 C8_N_btm.n185 C8_N_btm.n184 0.09425
R23103 C8_N_btm.n173 C8_N_btm.n43 0.09425
R23104 C8_N_btm.n43 C8_N_btm.n36 0.09425
R23105 C8_N_btm.n174 C8_N_btm.n42 0.09425
R23106 C8_N_btm.n174 C8_N_btm.n38 0.09425
R23107 C8_N_btm.n172 C8_N_btm.n171 0.09425
R23108 C8_N_btm.n173 C8_N_btm.n172 0.09425
R23109 C8_N_btm.n169 C8_N_btm.n44 0.09425
R23110 C8_N_btm.n44 C8_N_btm.n42 0.09425
R23111 C8_N_btm.n170 C8_N_btm.n45 0.09425
R23112 C8_N_btm.n171 C8_N_btm.n170 0.09425
R23113 C8_N_btm.n168 C8_N_btm.n47 0.09425
R23114 C8_N_btm.n169 C8_N_btm.n168 0.09425
R23115 C8_N_btm.n158 C8_N_btm.n52 0.09425
R23116 C8_N_btm.n52 C8_N_btm.n45 0.09425
R23117 C8_N_btm.n159 C8_N_btm.n51 0.09425
R23118 C8_N_btm.n159 C8_N_btm.n47 0.09425
R23119 C8_N_btm.n157 C8_N_btm.n156 0.09425
R23120 C8_N_btm.n158 C8_N_btm.n157 0.09425
R23121 C8_N_btm.n154 C8_N_btm.n53 0.09425
R23122 C8_N_btm.n53 C8_N_btm.n51 0.09425
R23123 C8_N_btm.n155 C8_N_btm.n54 0.09425
R23124 C8_N_btm.n156 C8_N_btm.n155 0.09425
R23125 C8_N_btm.n153 C8_N_btm.n56 0.09425
R23126 C8_N_btm.n154 C8_N_btm.n153 0.09425
R23127 C8_N_btm.n143 C8_N_btm.n61 0.09425
R23128 C8_N_btm.n61 C8_N_btm.n54 0.09425
R23129 C8_N_btm.n63 C8_N_btm.n60 0.09425
R23130 C8_N_btm.n144 C8_N_btm.n60 0.09425
R23131 C8_N_btm.n144 C8_N_btm.n56 0.09425
R23132 C8_N_btm.n141 C8_N_btm.n140 0.09425
R23133 C8_N_btm.n138 C8_N_btm.n62 0.09425
R23134 C8_N_btm.n65 C8_N_btm.n63 0.09425
R23135 C8_N_btm.n102 C8_N_btm.n93 0.09425
R23136 C8_N_btm.n93 C8_N_btm.n65 0.09425
R23137 C8_N_btm.n139 C8_N_btm.n64 0.09425
R23138 C8_N_btm.n140 C8_N_btm.n139 0.09425
R23139 C8_N_btm.n137 C8_N_btm.n67 0.09425
R23140 C8_N_btm.n138 C8_N_btm.n137 0.09425
R23141 C8_N_btm.n136 C8_N_btm.n66 0.09425
R23142 C8_N_btm.n73 C8_N_btm.n66 0.09425
R23143 C8_N_btm.n135 C8_N_btm.n69 0.09425
R23144 C8_N_btm.n135 C8_N_btm.n70 0.09425
R23145 C8_N_btm.n134 C8_N_btm.n133 0.09425
R23146 C8_N_btm.n133 C8_N_btm.n75 0.09425
R23147 C8_N_btm.n110 C8_N_btm.n72 0.09425
R23148 C8_N_btm.n132 C8_N_btm.n72 0.09425
R23149 C8_N_btm.n131 C8_N_btm.n77 0.09425
R23150 C8_N_btm.n131 C8_N_btm.n78 0.09425
R23151 C8_N_btm.n129 C8_N_btm.n81 0.09425
R23152 C8_N_btm.n130 C8_N_btm.n129 0.09425
R23153 C8_N_btm.n128 C8_N_btm.n80 0.09425
R23154 C8_N_btm.n87 C8_N_btm.n80 0.09425
R23155 C8_N_btm.n127 C8_N_btm.n83 0.09425
R23156 C8_N_btm.n127 C8_N_btm.n84 0.09425
R23157 C8_N_btm.n126 C8_N_btm.n125 0.09425
R23158 C8_N_btm.n125 C8_N_btm.n89 0.09425
R23159 C8_N_btm.n118 C8_N_btm.n86 0.09425
R23160 C8_N_btm.n124 C8_N_btm.n86 0.09425
R23161 C8_N_btm.n119 C8_N_btm.n91 0.09425
R23162 C8_N_btm.n118 C8_N_btm.n117 0.09425
R23163 C8_N_btm.n116 C8_N_btm.n85 0.09425
R23164 C8_N_btm.n126 C8_N_btm.n85 0.09425
R23165 C8_N_btm.n115 C8_N_btm.n83 0.09425
R23166 C8_N_btm.n114 C8_N_btm.n82 0.09425
R23167 C8_N_btm.n128 C8_N_btm.n82 0.09425
R23168 C8_N_btm.n113 C8_N_btm.n81 0.09425
R23169 C8_N_btm.n112 C8_N_btm.n111 0.09425
R23170 C8_N_btm.n111 C8_N_btm.n77 0.09425
R23171 C8_N_btm.n110 C8_N_btm.n109 0.09425
R23172 C8_N_btm.n108 C8_N_btm.n71 0.09425
R23173 C8_N_btm.n134 C8_N_btm.n71 0.09425
R23174 C8_N_btm.n107 C8_N_btm.n69 0.09425
R23175 C8_N_btm.n106 C8_N_btm.n68 0.09425
R23176 C8_N_btm.n136 C8_N_btm.n68 0.09425
R23177 C8_N_btm.n105 C8_N_btm.n67 0.09425
R23178 C8_N_btm.n104 C8_N_btm.n103 0.09425
R23179 C8_N_btm.n103 C8_N_btm.n64 0.09425
R23180 C8_N_btm.n102 C8_N_btm.n92 0.09425
R23181 C8_N_btm.n101 C8_N_btm.n100 0.09425
R23182 C8_N_btm.n100 C8_N_btm.n95 0.09425
R23183 C8_N_btm.n99 C8_N_btm.n98 0.09425
R23184 C8_N_btm.n98 C8_N_btm.n97 0.09425
R23185 C8_N_btm.n96 C8_N_btm.n95 0.09425
R23186 C8_N_btm.n96 C8_N_btm.n59 0.09425
R23187 C8_N_btm.n97 C8_N_btm.n58 0.09425
R23188 C8_N_btm.n146 C8_N_btm.n58 0.09425
R23189 C8_N_btm.n145 C8_N_btm.n59 0.09425
R23190 C8_N_btm.n145 C8_N_btm.n57 0.09425
R23191 C8_N_btm.n147 C8_N_btm.n146 0.09425
R23192 C8_N_btm.n151 C8_N_btm.n147 0.09425
R23193 C8_N_btm.n152 C8_N_btm.n57 0.09425
R23194 C8_N_btm.n152 C8_N_btm.n55 0.09425
R23195 C8_N_btm.n151 C8_N_btm.n150 0.09425
R23196 C8_N_btm.n150 C8_N_btm.n149 0.09425
R23197 C8_N_btm.n148 C8_N_btm.n55 0.09425
R23198 C8_N_btm.n148 C8_N_btm.n50 0.09425
R23199 C8_N_btm.n149 C8_N_btm.n49 0.09425
R23200 C8_N_btm.n161 C8_N_btm.n49 0.09425
R23201 C8_N_btm.n160 C8_N_btm.n50 0.09425
R23202 C8_N_btm.n160 C8_N_btm.n48 0.09425
R23203 C8_N_btm.n162 C8_N_btm.n161 0.09425
R23204 C8_N_btm.n166 C8_N_btm.n162 0.09425
R23205 C8_N_btm.n167 C8_N_btm.n48 0.09425
R23206 C8_N_btm.n167 C8_N_btm.n46 0.09425
R23207 C8_N_btm.n165 C8_N_btm.n164 0.09425
R23208 C8_N_btm.n163 C8_N_btm.n46 0.09425
R23209 C8_N_btm.n163 C8_N_btm.n41 0.09425
R23210 C8_N_btm.n164 C8_N_btm.n40 0.09425
R23211 C8_N_btm.n176 C8_N_btm.n40 0.09425
R23212 C8_N_btm.n175 C8_N_btm.n41 0.09425
R23213 C8_N_btm.n175 C8_N_btm.n39 0.09425
R23214 C8_N_btm.n177 C8_N_btm.n176 0.09425
R23215 C8_N_btm.n182 C8_N_btm.n177 0.09425
R23216 C8_N_btm.n183 C8_N_btm.n39 0.09425
R23217 C8_N_btm.n183 C8_N_btm.n37 0.09425
R23218 C8_N_btm.n182 C8_N_btm.n181 0.09425
R23219 C8_N_btm.n181 C8_N_btm.n180 0.09425
R23220 C8_N_btm.n179 C8_N_btm.n37 0.09425
R23221 C8_N_btm.n179 C8_N_btm.n34 0.09425
R23222 C8_N_btm.n189 C8_N_btm.n35 0.09425
R23223 C8_N_btm.n190 C8_N_btm.n189 0.09425
R23224 C8_N_btm.n233 C8_N_btm.n28 0.09425
R23225 C8_N_btm.n234 C8_N_btm.n26 0.09425
R23226 C8_N_btm.n235 C8_N_btm.n24 0.09425
R23227 C8_N_btm.n221 C8_N_btm.n24 0.09425
R23228 C8_N_btm.n237 C8_N_btm.n236 0.09425
R23229 C8_N_btm.n238 C8_N_btm.n21 0.09425
R23230 C8_N_btm.n238 C8_N_btm.n22 0.09425
R23231 C8_N_btm.n239 C8_N_btm.n18 0.09425
R23232 C8_N_btm.n241 C8_N_btm.n240 0.09425
R23233 C8_N_btm.n240 C8_N_btm.n19 0.09425
R23234 C8_N_btm.n242 C8_N_btm.n17 0.09425
R23235 C8_N_btm.n243 C8_N_btm.n16 0.09425
R23236 C8_N_btm.n213 C8_N_btm.n16 0.09425
R23237 C8_N_btm.n245 C8_N_btm.n244 0.09425
R23238 C8_N_btm.n246 C8_N_btm.n13 0.09425
R23239 C8_N_btm.n246 C8_N_btm.n14 0.09425
R23240 C8_N_btm.n247 C8_N_btm.n10 0.09425
R23241 C8_N_btm.n249 C8_N_btm.n248 0.09425
R23242 C8_N_btm.n248 C8_N_btm.n11 0.09425
R23243 C8_N_btm.n250 C8_N_btm.n9 0.09425
R23244 C8_N_btm.n166 C8_N_btm.n165 0.0816039
R23245 C8_N_btm.n143 C8_N_btm.n142 0.047875
R23246 C8_N_btm.n188 C8_N_btm.n25 0.047875
R23247 C8_N_btm.n208 C8_N_btm.n207 0.0342289
R23248 C8_N_btm.n227 C8_N_btm.n32 0.0342289
R23249 C8_N_btm.n123 C8_N_btm.n122 0.0342289
R23250 C8_N_btm.n142 C8_N_btm.n141 0.0342289
R23251 C8_N_btm.n120 C8_N_btm.n119 0.0342289
R23252 C8_N_btm.n101 C8_N_btm.n94 0.0342289
R23253 C8_N_btm.n28 C8_N_btm.n25 0.0342289
R23254 VREF.n0 VREF.t64 67.0515
R23255 VREF.n36 VREF.t53 67.0515
R23256 VREF.n4 VREF.t50 66.3952
R23257 VREF.n3 VREF.t51 66.3952
R23258 VREF.n2 VREF.t33 66.3952
R23259 VREF.n1 VREF.t71 66.3952
R23260 VREF.n0 VREF.t70 66.3952
R23261 VREF.n40 VREF.t52 66.3952
R23262 VREF.n39 VREF.t63 66.3952
R23263 VREF.n38 VREF.t62 66.3952
R23264 VREF.n37 VREF.t73 66.3952
R23265 VREF.n36 VREF.t72 66.3952
R23266 VREF VREF.n71 38.4352
R23267 VREF VREF.n35 38.2723
R23268 VREF.n35 VREF.t14 34.2201
R23269 VREF.n71 VREF.t34 34.2201
R23270 VREF.n34 VREF.n33 30.6495
R23271 VREF.n32 VREF.n31 30.6495
R23272 VREF.n30 VREF.n29 30.6495
R23273 VREF.n28 VREF.n27 30.6495
R23274 VREF.n26 VREF.n25 30.6495
R23275 VREF.n24 VREF.n23 30.6495
R23276 VREF.n22 VREF.n21 30.6495
R23277 VREF.n20 VREF.n19 30.6495
R23278 VREF.n18 VREF.n17 30.6495
R23279 VREF.n16 VREF.n15 30.6495
R23280 VREF.n14 VREF.n13 30.6495
R23281 VREF.n12 VREF.n11 30.6495
R23282 VREF.n10 VREF.n9 30.6495
R23283 VREF.n8 VREF.n7 30.6495
R23284 VREF.n6 VREF.n5 30.6495
R23285 VREF.n70 VREF.n69 30.6495
R23286 VREF.n68 VREF.n67 30.6495
R23287 VREF.n66 VREF.n65 30.6495
R23288 VREF.n64 VREF.n63 30.6495
R23289 VREF.n62 VREF.n61 30.6495
R23290 VREF.n60 VREF.n59 30.6495
R23291 VREF.n58 VREF.n57 30.6495
R23292 VREF.n56 VREF.n55 30.6495
R23293 VREF.n54 VREF.n53 30.6495
R23294 VREF.n52 VREF.n51 30.6495
R23295 VREF.n50 VREF.n49 30.6495
R23296 VREF.n48 VREF.n47 30.6495
R23297 VREF.n46 VREF.n45 30.6495
R23298 VREF.n44 VREF.n43 30.6495
R23299 VREF.n42 VREF.n41 30.6495
R23300 VREF.n33 VREF.t13 3.57113
R23301 VREF.n33 VREF.t26 3.57113
R23302 VREF.n31 VREF.t21 3.57113
R23303 VREF.n31 VREF.t17 3.57113
R23304 VREF.n29 VREF.t20 3.57113
R23305 VREF.n29 VREF.t27 3.57113
R23306 VREF.n27 VREF.t23 3.57113
R23307 VREF.n27 VREF.t15 3.57113
R23308 VREF.n25 VREF.t25 3.57113
R23309 VREF.n25 VREF.t19 3.57113
R23310 VREF.n23 VREF.t12 3.57113
R23311 VREF.n23 VREF.t22 3.57113
R23312 VREF.n21 VREF.t24 3.57113
R23313 VREF.n21 VREF.t16 3.57113
R23314 VREF.n19 VREF.t18 3.57113
R23315 VREF.n19 VREF.t6 3.57113
R23316 VREF.n17 VREF.t5 3.57113
R23317 VREF.n17 VREF.t10 3.57113
R23318 VREF.n15 VREF.t9 3.57113
R23319 VREF.n15 VREF.t7 3.57113
R23320 VREF.n13 VREF.t11 3.57113
R23321 VREF.n13 VREF.t4 3.57113
R23322 VREF.n11 VREF.t8 3.57113
R23323 VREF.n11 VREF.t3 3.57113
R23324 VREF.n9 VREF.t2 3.57113
R23325 VREF.n9 VREF.t1 3.57113
R23326 VREF.n7 VREF.t0 3.57113
R23327 VREF.n7 VREF.t29 3.57113
R23328 VREF.n5 VREF.t28 3.57113
R23329 VREF.n5 VREF.t32 3.57113
R23330 VREF.n69 VREF.t46 3.57113
R23331 VREF.n69 VREF.t44 3.57113
R23332 VREF.n67 VREF.t36 3.57113
R23333 VREF.n67 VREF.t42 3.57113
R23334 VREF.n65 VREF.t47 3.57113
R23335 VREF.n65 VREF.t43 3.57113
R23336 VREF.n63 VREF.t45 3.57113
R23337 VREF.n63 VREF.t41 3.57113
R23338 VREF.n61 VREF.t37 3.57113
R23339 VREF.n61 VREF.t49 3.57113
R23340 VREF.n59 VREF.t35 3.57113
R23341 VREF.n59 VREF.t48 3.57113
R23342 VREF.n57 VREF.t39 3.57113
R23343 VREF.n57 VREF.t40 3.57113
R23344 VREF.n55 VREF.t56 3.57113
R23345 VREF.n55 VREF.t38 3.57113
R23346 VREF.n53 VREF.t58 3.57113
R23347 VREF.n53 VREF.t59 3.57113
R23348 VREF.n51 VREF.t61 3.57113
R23349 VREF.n51 VREF.t57 3.57113
R23350 VREF.n49 VREF.t60 3.57113
R23351 VREF.n49 VREF.t55 3.57113
R23352 VREF.n47 VREF.t69 3.57113
R23353 VREF.n47 VREF.t54 3.57113
R23354 VREF.n45 VREF.t68 3.57113
R23355 VREF.n45 VREF.t67 3.57113
R23356 VREF.n43 VREF.t30 3.57113
R23357 VREF.n43 VREF.t66 3.57113
R23358 VREF.n41 VREF.t65 3.57113
R23359 VREF.n41 VREF.t31 3.57113
R23360 VREF.n8 VREF.n6 0.71925
R23361 VREF.n10 VREF.n8 0.71925
R23362 VREF.n14 VREF.n12 0.71925
R23363 VREF.n16 VREF.n14 0.71925
R23364 VREF.n20 VREF.n18 0.71925
R23365 VREF.n24 VREF.n22 0.71925
R23366 VREF.n26 VREF.n24 0.71925
R23367 VREF.n30 VREF.n28 0.71925
R23368 VREF.n34 VREF.n32 0.71925
R23369 VREF.n35 VREF.n34 0.71925
R23370 VREF.n44 VREF.n42 0.71925
R23371 VREF.n46 VREF.n44 0.71925
R23372 VREF.n50 VREF.n48 0.71925
R23373 VREF.n52 VREF.n50 0.71925
R23374 VREF.n56 VREF.n54 0.71925
R23375 VREF.n60 VREF.n58 0.71925
R23376 VREF.n62 VREF.n60 0.71925
R23377 VREF.n66 VREF.n64 0.71925
R23378 VREF.n70 VREF.n68 0.71925
R23379 VREF.n71 VREF.n70 0.71925
R23380 VREF.n2 VREF.n1 0.688
R23381 VREF.n12 VREF.n10 0.688
R23382 VREF.n18 VREF.n16 0.688
R23383 VREF.n22 VREF.n20 0.688
R23384 VREF.n28 VREF.n26 0.688
R23385 VREF.n32 VREF.n30 0.688
R23386 VREF.n38 VREF.n37 0.688
R23387 VREF.n48 VREF.n46 0.688
R23388 VREF.n54 VREF.n52 0.688
R23389 VREF.n58 VREF.n56 0.688
R23390 VREF.n64 VREF.n62 0.688
R23391 VREF.n68 VREF.n66 0.688
R23392 VREF.n1 VREF.n0 0.65675
R23393 VREF.n3 VREF.n2 0.65675
R23394 VREF.n4 VREF.n3 0.65675
R23395 VREF.n6 VREF.n4 0.65675
R23396 VREF.n37 VREF.n36 0.65675
R23397 VREF.n39 VREF.n38 0.65675
R23398 VREF.n40 VREF.n39 0.65675
R23399 VREF.n42 VREF.n40 0.65675
R23400 a_n3565_37414.n4 a_n3565_37414.t8 556.423
R23401 a_n3565_37414.n8 a_n3565_37414.n7 340.637
R23402 a_n3565_37414.n3 a_n3565_37414.t9 241.536
R23403 a_n3565_37414.n7 a_n3565_37414.n6 195.577
R23404 a_n3565_37414.n3 a_n3565_37414.t10 169.237
R23405 a_n3565_37414.n4 a_n3565_37414.n3 168.505
R23406 a_n3565_37414.n2 a_n3565_37414.n0 137.189
R23407 a_n3565_37414.n2 a_n3565_37414.n1 98.788
R23408 a_n3565_37414.n7 a_n3565_37414.n5 39.0246
R23409 a_n3565_37414.n6 a_n3565_37414.t1 26.5955
R23410 a_n3565_37414.n6 a_n3565_37414.t0 26.5955
R23411 a_n3565_37414.t3 a_n3565_37414.n8 26.5955
R23412 a_n3565_37414.n8 a_n3565_37414.t2 26.5955
R23413 a_n3565_37414.n5 a_n3565_37414.n2 25.9824
R23414 a_n3565_37414.n0 a_n3565_37414.t7 24.9236
R23415 a_n3565_37414.n0 a_n3565_37414.t5 24.9236
R23416 a_n3565_37414.n1 a_n3565_37414.t4 24.9236
R23417 a_n3565_37414.n1 a_n3565_37414.t6 24.9236
R23418 a_n3565_37414.n5 a_n3565_37414.n4 9.38613
R23419 a_1307_43914.n33 a_1307_43914.n32 647.148
R23420 a_1307_43914.n24 a_1307_43914.n22 459.668
R23421 a_1307_43914.n23 a_1307_43914.t28 329.902
R23422 a_1307_43914.n22 a_1307_43914.t27 272.062
R23423 a_1307_43914.n30 a_1307_43914.n0 243.627
R23424 a_1307_43914.n17 a_1307_43914.t9 241.536
R23425 a_1307_43914.n2 a_1307_43914.t29 236.552
R23426 a_1307_43914.n1 a_1307_43914.t33 236.552
R23427 a_1307_43914.n18 a_1307_43914.t15 236.552
R23428 a_1307_43914.n16 a_1307_43914.t34 231.835
R23429 a_1307_43914.n14 a_1307_43914.t32 231.835
R23430 a_1307_43914.n15 a_1307_43914.t23 231.017
R23431 a_1307_43914.n4 a_1307_43914.t26 212.081
R23432 a_1307_43914.n6 a_1307_43914.t24 212.081
R23433 a_1307_43914.n8 a_1307_43914.t14 212.081
R23434 a_1307_43914.n7 a_1307_43914.t20 212.081
R23435 a_1307_43914.n22 a_1307_43914.t25 206.19
R23436 a_1307_43914.n11 a_1307_43914.n3 203.839
R23437 a_1307_43914.n3 a_1307_43914.t18 196.549
R23438 a_1307_43914.n19 a_1307_43914.n17 196.37
R23439 a_1307_43914.n32 a_1307_43914.n31 194.441
R23440 a_1307_43914.n29 a_1307_43914.n28 185
R23441 a_1307_43914.n13 a_1307_43914.n1 176.852
R23442 a_1307_43914.n19 a_1307_43914.n18 170.905
R23443 a_1307_43914.n17 a_1307_43914.t17 169.237
R23444 a_1307_43914.n12 a_1307_43914.n2 167.966
R23445 a_1307_43914.n2 a_1307_43914.t12 164.251
R23446 a_1307_43914.n1 a_1307_43914.t22 164.251
R23447 a_1307_43914.n18 a_1307_43914.t35 164.251
R23448 a_1307_43914.n20 a_1307_43914.n16 163.84
R23449 a_1307_43914.n26 a_1307_43914.n14 163.84
R23450 a_1307_43914.n21 a_1307_43914.n15 163.435
R23451 a_1307_43914.n10 a_1307_43914.n5 162.752
R23452 a_1307_43914.n10 a_1307_43914.n9 162.752
R23453 a_1307_43914.n15 a_1307_43914.t30 158.716
R23454 a_1307_43914.n16 a_1307_43914.t11 157.07
R23455 a_1307_43914.n14 a_1307_43914.t16 157.07
R23456 a_1307_43914.n24 a_1307_43914.n23 152
R23457 a_1307_43914.n3 a_1307_43914.t13 148.35
R23458 a_1307_43914.n23 a_1307_43914.t31 148.35
R23459 a_1307_43914.n4 a_1307_43914.t10 139.78
R23460 a_1307_43914.n6 a_1307_43914.t19 139.78
R23461 a_1307_43914.n8 a_1307_43914.t21 139.78
R23462 a_1307_43914.n7 a_1307_43914.t8 139.78
R23463 a_1307_43914.n8 a_1307_43914.n7 61.346
R23464 a_1307_43914.n32 a_1307_43914.n30 50.5705
R23465 a_1307_43914.n0 a_1307_43914.t7 40.0005
R23466 a_1307_43914.n0 a_1307_43914.t4 40.0005
R23467 a_1307_43914.n28 a_1307_43914.t6 40.0005
R23468 a_1307_43914.n28 a_1307_43914.t5 40.0005
R23469 a_1307_43914.n5 a_1307_43914.n4 30.6732
R23470 a_1307_43914.n6 a_1307_43914.n5 30.6732
R23471 a_1307_43914.n9 a_1307_43914.n6 30.6732
R23472 a_1307_43914.n9 a_1307_43914.n8 30.6732
R23473 a_1307_43914.n31 a_1307_43914.t2 27.5805
R23474 a_1307_43914.n31 a_1307_43914.t1 27.5805
R23475 a_1307_43914.t3 a_1307_43914.n33 27.5805
R23476 a_1307_43914.n33 a_1307_43914.t0 27.5805
R23477 a_1307_43914.n25 a_1307_43914.n24 27.4285
R23478 a_1307_43914.n29 a_1307_43914.n27 20.2936
R23479 a_1307_43914.n11 a_1307_43914.n10 17.6235
R23480 a_1307_43914.n30 a_1307_43914.n29 15.262
R23481 a_1307_43914.n20 a_1307_43914.n19 10.4738
R23482 a_1307_43914.n13 a_1307_43914.n12 4.5005
R23483 a_1307_43914.n21 a_1307_43914.n20 3.28621
R23484 a_1307_43914.n27 a_1307_43914.n26 2.80957
R23485 a_1307_43914.n25 a_1307_43914.n21 2.57742
R23486 a_1307_43914.n27 a_1307_43914.n13 2.11314
R23487 a_1307_43914.n12 a_1307_43914.n11 1.68457
R23488 a_1307_43914.n26 a_1307_43914.n25 0.934566
R23489 a_n913_45002.n5 a_n913_45002.n4 256.104
R23490 a_n913_45002.n2 a_n913_45002.n0 241.847
R23491 a_n913_45002.n26 a_n913_45002.t27 230.363
R23492 a_n913_45002.n9 a_n913_45002.t28 230.363
R23493 a_n913_45002.n10 a_n913_45002.t31 230.363
R23494 a_n913_45002.n11 a_n913_45002.t13 230.363
R23495 a_n913_45002.n21 a_n913_45002.t21 230.363
R23496 a_n913_45002.n19 a_n913_45002.t22 230.363
R23497 a_n913_45002.n17 a_n913_45002.t14 230.363
R23498 a_n913_45002.n15 a_n913_45002.t23 230.363
R23499 a_n913_45002.n12 a_n913_45002.t30 230.363
R23500 a_n913_45002.n13 a_n913_45002.t17 230.363
R23501 a_n913_45002.n28 a_n913_45002.t15 230.363
R23502 a_n913_45002.n8 a_n913_45002.n7 205.28
R23503 a_n913_45002.n5 a_n913_45002.n3 202.094
R23504 a_n913_45002.n29 a_n913_45002.n28 196.138
R23505 a_n913_45002.n31 a_n913_45002.n30 190.911
R23506 a_n913_45002.n2 a_n913_45002.n1 185
R23507 a_n913_45002.n18 a_n913_45002.n17 175.252
R23508 a_n913_45002.n20 a_n913_45002.n19 174.038
R23509 a_n913_45002.n14 a_n913_45002.n13 168.998
R23510 a_n913_45002.n27 a_n913_45002.n26 163.84
R23511 a_n913_45002.n25 a_n913_45002.n9 163.536
R23512 a_n913_45002.n24 a_n913_45002.n10 163.536
R23513 a_n913_45002.n23 a_n913_45002.n11 163.536
R23514 a_n913_45002.n22 a_n913_45002.n21 163.349
R23515 a_n913_45002.n16 a_n913_45002.n15 163.349
R23516 a_n913_45002.n14 a_n913_45002.n12 163.349
R23517 a_n913_45002.n26 a_n913_45002.t25 158.064
R23518 a_n913_45002.n9 a_n913_45002.t19 158.064
R23519 a_n913_45002.n10 a_n913_45002.t18 158.064
R23520 a_n913_45002.n11 a_n913_45002.t32 158.064
R23521 a_n913_45002.n21 a_n913_45002.t24 158.064
R23522 a_n913_45002.n19 a_n913_45002.t33 158.064
R23523 a_n913_45002.n17 a_n913_45002.t20 158.064
R23524 a_n913_45002.n15 a_n913_45002.t26 158.064
R23525 a_n913_45002.n12 a_n913_45002.t29 158.064
R23526 a_n913_45002.n13 a_n913_45002.t16 158.064
R23527 a_n913_45002.n28 a_n913_45002.t12 158.064
R23528 a_n913_45002.n16 a_n913_45002.n14 53.212
R23529 a_n913_45002.n30 a_n913_45002.n8 52.7703
R23530 a_n913_45002.n8 a_n913_45002.n6 36.8946
R23531 a_n913_45002.n6 a_n913_45002.n2 28.2251
R23532 a_n913_45002.n3 a_n913_45002.t7 26.5955
R23533 a_n913_45002.n3 a_n913_45002.t4 26.5955
R23534 a_n913_45002.n4 a_n913_45002.t6 26.5955
R23535 a_n913_45002.n4 a_n913_45002.t5 26.5955
R23536 a_n913_45002.n7 a_n913_45002.t0 26.5955
R23537 a_n913_45002.n7 a_n913_45002.t2 26.5955
R23538 a_n913_45002.t3 a_n913_45002.n31 26.5955
R23539 a_n913_45002.n31 a_n913_45002.t1 26.5955
R23540 a_n913_45002.n1 a_n913_45002.t9 24.9236
R23541 a_n913_45002.n1 a_n913_45002.t11 24.9236
R23542 a_n913_45002.n0 a_n913_45002.t8 24.9236
R23543 a_n913_45002.n0 a_n913_45002.t10 24.9236
R23544 a_n913_45002.n22 a_n913_45002.n20 20.3535
R23545 a_n913_45002.n30 a_n913_45002.n29 18.9814
R23546 a_n913_45002.n6 a_n913_45002.n5 13.9299
R23547 a_n913_45002.n29 a_n913_45002.n27 12.892
R23548 a_n913_45002.n18 a_n913_45002.n16 11.1461
R23549 a_n913_45002.n27 a_n913_45002.n25 10.5184
R23550 a_n913_45002.n20 a_n913_45002.n18 7.6722
R23551 a_n913_45002.n23 a_n913_45002.n22 7.64057
R23552 a_n913_45002.n25 a_n913_45002.n24 7.1255
R23553 a_n913_45002.n24 a_n913_45002.n23 2.05407
R23554 a_n2661_43370.n0 a_n2661_43370.t4 276.464
R23555 a_n2661_43370.n1 a_n2661_43370.n0 208.779
R23556 a_n2661_43370.n2 a_n2661_43370.n1 196.846
R23557 a_n2661_43370.n0 a_n2661_43370.t3 196.131
R23558 a_n2661_43370.n1 a_n2661_43370.t2 193.519
R23559 a_n2661_43370.n2 a_n2661_43370.t1 26.5955
R23560 a_n2661_43370.t0 a_n2661_43370.n2 26.5955
R23561 a_584_46384.n4 a_584_46384.t17 414.432
R23562 a_584_46384.n5 a_584_46384.t15 414.432
R23563 a_584_46384.n4 a_584_46384.t10 300.349
R23564 a_584_46384.n5 a_584_46384.t21 300.349
R23565 a_584_46384.n11 a_584_46384.n9 259.221
R23566 a_584_46384.n19 a_584_46384.n0 248.087
R23567 a_584_46384.n14 a_584_46384.t9 241.536
R23568 a_584_46384.n6 a_584_46384.t20 241.536
R23569 a_584_46384.n10 a_584_46384.t13 236.18
R23570 a_584_46384.n9 a_584_46384.t16 234.392
R23571 a_584_46384.n12 a_584_46384.n8 212.248
R23572 a_584_46384.n7 a_584_46384.t22 212.081
R23573 a_584_46384.n8 a_584_46384.t19 212.081
R23574 a_584_46384.n20 a_584_46384.n19 208.506
R23575 a_584_46384.n13 a_584_46384.n6 174.275
R23576 a_584_46384.n15 a_584_46384.n14 170.581
R23577 a_584_46384.n14 a_584_46384.t18 169.237
R23578 a_584_46384.n6 a_584_46384.t12 169.237
R23579 a_584_46384.n10 a_584_46384.t8 163.881
R23580 a_584_46384.n11 a_584_46384.n10 152
R23581 a_584_46384.n9 a_584_46384.t11 150.442
R23582 a_584_46384.n7 a_584_46384.t23 139.78
R23583 a_584_46384.n8 a_584_46384.t14 139.78
R23584 a_584_46384.n3 a_584_46384.n1 137.576
R23585 a_584_46384.n3 a_584_46384.n2 99.1759
R23586 a_584_46384.n8 a_584_46384.n7 61.346
R23587 a_584_46384.n19 a_584_46384.n18 38.4831
R23588 a_584_46384.n0 a_584_46384.t2 26.5955
R23589 a_584_46384.n0 a_584_46384.t0 26.5955
R23590 a_584_46384.t3 a_584_46384.n20 26.5955
R23591 a_584_46384.n20 a_584_46384.t1 26.5955
R23592 a_584_46384.n1 a_584_46384.t7 24.9236
R23593 a_584_46384.n1 a_584_46384.t4 24.9236
R23594 a_584_46384.n2 a_584_46384.t6 24.9236
R23595 a_584_46384.n2 a_584_46384.t5 24.9236
R23596 a_584_46384.n16 a_584_46384.n15 23.4466
R23597 a_584_46384.n17 a_584_46384.n4 20.0626
R23598 a_584_46384.n12 a_584_46384.n11 18.6598
R23599 a_584_46384.n18 a_584_46384.n3 14.8665
R23600 a_584_46384.n18 a_584_46384.n17 14.3332
R23601 a_584_46384.n17 a_584_46384.n16 11.767
R23602 a_584_46384.n16 a_584_46384.n5 10.499
R23603 a_584_46384.n13 a_584_46384.n12 9.28846
R23604 a_584_46384.n15 a_584_46384.n13 6.02676
R23605 a_2107_46812.n0 a_2107_46812.t3 236.18
R23606 a_2107_46812.t0 a_2107_46812.n1 235.673
R23607 a_2107_46812.n1 a_2107_46812.n0 208.721
R23608 a_2107_46812.n1 a_2107_46812.t1 185.165
R23609 a_2107_46812.n0 a_2107_46812.t2 163.881
R23610 a_n1059_45260.n9 a_n1059_45260.t21 657.383
R23611 a_n1059_45260.t21 a_n1059_45260.t12 378.255
R23612 a_n1059_45260.n4 a_n1059_45260.t16 327.99
R23613 a_n1059_45260.n6 a_n1059_45260.t22 256.728
R23614 a_n1059_45260.n20 a_n1059_45260.n19 248.085
R23615 a_n1059_45260.n7 a_n1059_45260.t9 241.536
R23616 a_n1059_45260.n3 a_n1059_45260.t8 241.536
R23617 a_n1059_45260.n8 a_n1059_45260.t20 231.835
R23618 a_n1059_45260.n19 a_n1059_45260.n18 208.507
R23619 a_n1059_45260.n13 a_n1059_45260.n12 201.16
R23620 a_n1059_45260.n4 a_n1059_45260.t17 199.457
R23621 a_n1059_45260.n9 a_n1059_45260.n8 190.814
R23622 a_n1059_45260.n14 a_n1059_45260.n7 180.369
R23623 a_n1059_45260.n5 a_n1059_45260.n4 178.679
R23624 a_n1059_45260.n12 a_n1059_45260.t19 173.34
R23625 a_n1059_45260.n11 a_n1059_45260.n10 169.498
R23626 a_n1059_45260.n7 a_n1059_45260.t15 169.237
R23627 a_n1059_45260.n3 a_n1059_45260.t13 169.237
R23628 a_n1059_45260.n5 a_n1059_45260.n3 163.912
R23629 a_n1059_45260.n12 a_n1059_45260.t14 162.81
R23630 a_n1059_45260.n15 a_n1059_45260.n6 162.653
R23631 a_n1059_45260.n6 a_n1059_45260.t23 161.275
R23632 a_n1059_45260.n8 a_n1059_45260.t11 157.07
R23633 a_n1059_45260.n2 a_n1059_45260.n0 137.576
R23634 a_n1059_45260.n10 a_n1059_45260.t18 137.177
R23635 a_n1059_45260.n10 a_n1059_45260.t10 121.109
R23636 a_n1059_45260.n2 a_n1059_45260.n1 99.1759
R23637 a_n1059_45260.n19 a_n1059_45260.n17 38.4831
R23638 a_n1059_45260.n18 a_n1059_45260.t1 26.5955
R23639 a_n1059_45260.n18 a_n1059_45260.t2 26.5955
R23640 a_n1059_45260.n20 a_n1059_45260.t0 26.5955
R23641 a_n1059_45260.t3 a_n1059_45260.n20 26.5955
R23642 a_n1059_45260.n0 a_n1059_45260.t6 24.9236
R23643 a_n1059_45260.n0 a_n1059_45260.t5 24.9236
R23644 a_n1059_45260.n1 a_n1059_45260.t4 24.9236
R23645 a_n1059_45260.n1 a_n1059_45260.t7 24.9236
R23646 a_n1059_45260.n14 a_n1059_45260.n13 19.0335
R23647 a_n1059_45260.n17 a_n1059_45260.n16 16.6056
R23648 a_n1059_45260.n17 a_n1059_45260.n2 14.8665
R23649 a_n1059_45260.n13 a_n1059_45260.n11 9.8918
R23650 a_n1059_45260.n16 a_n1059_45260.n15 8.72028
R23651 a_n1059_45260.n16 a_n1059_45260.n5 8.26149
R23652 a_n1059_45260.n11 a_n1059_45260.n9 4.57639
R23653 a_n1059_45260.n15 a_n1059_45260.n14 3.58979
R23654 a_n1794_35082.n23 a_n1794_35082.n22 296.139
R23655 a_n1794_35082.n22 a_n1794_35082.n0 269.182
R23656 a_n1794_35082.n13 a_n1794_35082.t8 212.081
R23657 a_n1794_35082.n15 a_n1794_35082.t16 212.081
R23658 a_n1794_35082.n17 a_n1794_35082.t5 212.081
R23659 a_n1794_35082.n11 a_n1794_35082.t6 212.081
R23660 a_n1794_35082.n1 a_n1794_35082.t10 212.081
R23661 a_n1794_35082.n7 a_n1794_35082.t17 212.081
R23662 a_n1794_35082.n5 a_n1794_35082.t13 212.081
R23663 a_n1794_35082.n3 a_n1794_35082.t18 212.081
R23664 a_n1794_35082.n20 a_n1794_35082.n11 194.47
R23665 a_n1794_35082.n10 a_n1794_35082.n1 194.47
R23666 a_n1794_35082.n14 a_n1794_35082.n12 173.505
R23667 a_n1794_35082.n4 a_n1794_35082.n2 173.505
R23668 a_n1794_35082.n19 a_n1794_35082.n18 152
R23669 a_n1794_35082.n16 a_n1794_35082.n12 152
R23670 a_n1794_35082.n6 a_n1794_35082.n2 152
R23671 a_n1794_35082.n9 a_n1794_35082.n8 152
R23672 a_n1794_35082.n13 a_n1794_35082.t12 139.78
R23673 a_n1794_35082.n15 a_n1794_35082.t4 139.78
R23674 a_n1794_35082.n17 a_n1794_35082.t19 139.78
R23675 a_n1794_35082.n11 a_n1794_35082.t9 139.78
R23676 a_n1794_35082.n1 a_n1794_35082.t11 139.78
R23677 a_n1794_35082.n7 a_n1794_35082.t7 139.78
R23678 a_n1794_35082.n5 a_n1794_35082.t14 139.78
R23679 a_n1794_35082.n3 a_n1794_35082.t15 139.78
R23680 a_n1794_35082.n21 a_n1794_35082.n10 106.132
R23681 a_n1794_35082.n22 a_n1794_35082.n21 71.8985
R23682 a_n1794_35082.n14 a_n1794_35082.n13 30.6732
R23683 a_n1794_35082.n15 a_n1794_35082.n14 30.6732
R23684 a_n1794_35082.n16 a_n1794_35082.n15 30.6732
R23685 a_n1794_35082.n17 a_n1794_35082.n16 30.6732
R23686 a_n1794_35082.n18 a_n1794_35082.n17 30.6732
R23687 a_n1794_35082.n18 a_n1794_35082.n11 30.6732
R23688 a_n1794_35082.n8 a_n1794_35082.n1 30.6732
R23689 a_n1794_35082.n8 a_n1794_35082.n7 30.6732
R23690 a_n1794_35082.n7 a_n1794_35082.n6 30.6732
R23691 a_n1794_35082.n6 a_n1794_35082.n5 30.6732
R23692 a_n1794_35082.n5 a_n1794_35082.n4 30.6732
R23693 a_n1794_35082.n4 a_n1794_35082.n3 30.6732
R23694 a_n1794_35082.n21 a_n1794_35082.n20 29.3278
R23695 a_n1794_35082.t1 a_n1794_35082.n23 26.5955
R23696 a_n1794_35082.n23 a_n1794_35082.t0 26.5955
R23697 a_n1794_35082.n0 a_n1794_35082.t2 24.9236
R23698 a_n1794_35082.n0 a_n1794_35082.t3 24.9236
R23699 a_n1794_35082.n19 a_n1794_35082.n12 21.5045
R23700 a_n1794_35082.n9 a_n1794_35082.n2 21.5045
R23701 a_n1794_35082.n20 a_n1794_35082.n19 8.07753
R23702 a_n1794_35082.n10 a_n1794_35082.n9 8.07752
R23703 a_n1696_34930.n3 a_n1696_34930.t14 749.612
R23704 a_n1696_34930.n9 a_n1696_34930.t15 748.122
R23705 a_n1696_34930.n7 a_n1696_34930.t11 748.122
R23706 a_n1696_34930.n3 a_n1696_34930.t8 684.441
R23707 a_n1696_34930.n5 a_n1696_34930.t9 684.441
R23708 a_n1696_34930.n4 a_n1696_34930.t10 684.441
R23709 a_n1696_34930.n9 a_n1696_34930.t13 678.014
R23710 a_n1696_34930.n7 a_n1696_34930.t12 678.014
R23711 a_n1696_34930.n14 a_n1696_34930.n13 244.069
R23712 a_n1696_34930.n2 a_n1696_34930.n0 236.589
R23713 a_n1696_34930.n13 a_n1696_34930.n12 204.893
R23714 a_n1696_34930.n2 a_n1696_34930.n1 200.321
R23715 a_n1696_34930.n8 a_n1696_34930.n7 163.538
R23716 a_n1696_34930.n10 a_n1696_34930.n9 163.538
R23717 a_n1696_34930.n6 a_n1696_34930.n5 161.512
R23718 a_n1696_34930.n6 a_n1696_34930.n3 161.488
R23719 a_n1696_34930.n4 a_n1696_34930.n3 65.1723
R23720 a_n1696_34930.n5 a_n1696_34930.n4 65.1723
R23721 a_n1696_34930.n11 a_n1696_34930.n2 26.8022
R23722 a_n1696_34930.n12 a_n1696_34930.t0 26.5955
R23723 a_n1696_34930.n12 a_n1696_34930.t2 26.5955
R23724 a_n1696_34930.t3 a_n1696_34930.n14 26.5955
R23725 a_n1696_34930.n14 a_n1696_34930.t1 26.5955
R23726 a_n1696_34930.n13 a_n1696_34930.n11 25.4552
R23727 a_n1696_34930.n0 a_n1696_34930.t4 24.9236
R23728 a_n1696_34930.n0 a_n1696_34930.t6 24.9236
R23729 a_n1696_34930.n1 a_n1696_34930.t5 24.9236
R23730 a_n1696_34930.n1 a_n1696_34930.t7 24.9236
R23731 a_n1696_34930.n8 a_n1696_34930.n6 8.34135
R23732 a_n1696_34930.n11 a_n1696_34930.n10 6.02253
R23733 a_n1696_34930.n10 a_n1696_34930.n8 2.47042
R23734 a_n1925_42282.n0 a_n1925_42282.t4 276.464
R23735 a_n1925_42282.n1 a_n1925_42282.n0 249.421
R23736 a_n1925_42282.n1 a_n1925_42282.t1 199.456
R23737 a_n1925_42282.n0 a_n1925_42282.t3 196.131
R23738 a_n1925_42282.n2 a_n1925_42282.n1 190.911
R23739 a_n1925_42282.n2 a_n1925_42282.t2 26.5955
R23740 a_n1925_42282.t0 a_n1925_42282.n2 26.5955
R23741 a_12549_44172.t9 a_12549_44172.t4 403.274
R23742 a_12549_44172.n10 a_12549_44172.n6 337.009
R23743 a_12549_44172.n3 a_12549_44172.t31 328.659
R23744 a_12549_44172.n16 a_12549_44172.t9 325.175
R23745 a_12549_44172.n2 a_12549_44172.t29 295.432
R23746 a_12549_44172.n12 a_12549_44172.t19 295.432
R23747 a_12549_44172.n23 a_12549_44172.t21 293.969
R23748 a_12549_44172.n28 a_12549_44172.n27 287.752
R23749 a_12549_44172.n27 a_12549_44172.n0 277.568
R23750 a_12549_44172.n17 a_12549_44172.t8 261.887
R23751 a_12549_44172.n1 a_12549_44172.t14 241.536
R23752 a_12549_44172.n2 a_12549_44172.t25 237.591
R23753 a_12549_44172.n12 a_12549_44172.t22 237.591
R23754 a_12549_44172.n22 a_12549_44172.t28 230.363
R23755 a_12549_44172.n19 a_12549_44172.t5 212.081
R23756 a_12549_44172.n20 a_12549_44172.t18 212.081
R23757 a_12549_44172.n7 a_12549_44172.t11 212.081
R23758 a_12549_44172.n8 a_12549_44172.t20 212.081
R23759 a_12549_44172.n4 a_12549_44172.t24 212.081
R23760 a_12549_44172.n5 a_12549_44172.t15 212.081
R23761 a_12549_44172.n10 a_12549_44172.n9 211.035
R23762 a_12549_44172.n14 a_12549_44172.n2 200.619
R23763 a_12549_44172.n11 a_12549_44172.n3 195.167
R23764 a_12549_44172.n24 a_12549_44172.n22 176.358
R23765 a_12549_44172.n18 a_12549_44172.n17 172.165
R23766 a_12549_44172.n13 a_12549_44172.n12 169.751
R23767 a_12549_44172.n1 a_12549_44172.t26 169.237
R23768 a_12549_44172.n15 a_12549_44172.n1 166.696
R23769 a_12549_44172.n24 a_12549_44172.n23 163.879
R23770 a_12549_44172.n22 a_12549_44172.t13 158.064
R23771 a_12549_44172.n17 a_12549_44172.t27 155.847
R23772 a_12549_44172.n19 a_12549_44172.t30 139.78
R23773 a_12549_44172.n20 a_12549_44172.t10 139.78
R23774 a_12549_44172.n7 a_12549_44172.t7 139.78
R23775 a_12549_44172.n8 a_12549_44172.t16 139.78
R23776 a_12549_44172.n4 a_12549_44172.t17 139.78
R23777 a_12549_44172.n5 a_12549_44172.t23 139.78
R23778 a_12549_44172.n23 a_12549_44172.t6 138.338
R23779 a_12549_44172.n3 a_12549_44172.t12 126.219
R23780 a_12549_44172.n25 a_12549_44172.n21 101.695
R23781 a_12549_44172.n21 a_12549_44172.n19 52.4879
R23782 a_12549_44172.n9 a_12549_44172.n8 38.7066
R23783 a_12549_44172.n6 a_12549_44172.n5 37.246
R23784 a_12549_44172.n27 a_12549_44172.n26 31.9964
R23785 a_12549_44172.n9 a_12549_44172.n7 27.752
R23786 a_12549_44172.t1 a_12549_44172.n28 26.5955
R23787 a_12549_44172.n28 a_12549_44172.t0 26.5955
R23788 a_12549_44172.n0 a_12549_44172.t3 24.9236
R23789 a_12549_44172.n0 a_12549_44172.t2 24.9236
R23790 a_12549_44172.n11 a_12549_44172.n10 24.223
R23791 a_12549_44172.n6 a_12549_44172.n4 24.1005
R23792 a_12549_44172.n21 a_12549_44172.n20 9.34851
R23793 a_12549_44172.n25 a_12549_44172.n24 8.26939
R23794 a_12549_44172.n14 a_12549_44172.n13 8.07481
R23795 a_12549_44172.n15 a_12549_44172.n14 6.21255
R23796 a_12549_44172.n16 a_12549_44172.n15 6.0002
R23797 a_12549_44172.n13 a_12549_44172.n11 5.16448
R23798 a_12549_44172.n26 a_12549_44172.n25 4.32448
R23799 a_12549_44172.n18 a_12549_44172.n16 2.95053
R23800 a_12549_44172.n26 a_12549_44172.n18 0.500267
R23801 a_743_42282.n2 a_743_42282.n1 336.675
R23802 a_743_42282.n4 a_743_42282.t9 276.464
R23803 a_743_42282.n8 a_743_42282.n7 273.32
R23804 a_743_42282.n5 a_743_42282.n4 206.931
R23805 a_743_42282.n4 a_743_42282.t8 196.131
R23806 a_743_42282.n7 a_743_42282.n0 190.726
R23807 a_743_42282.n5 a_743_42282.n3 189.431
R23808 a_743_42282.n3 a_743_42282.n2 185
R23809 a_743_42282.n7 a_743_42282.n6 47.6805
R23810 a_743_42282.n1 a_743_42282.t6 27.5805
R23811 a_743_42282.n1 a_743_42282.t4 27.5805
R23812 a_743_42282.n3 a_743_42282.t5 25.8467
R23813 a_743_42282.n3 a_743_42282.t7 25.8467
R23814 a_743_42282.n0 a_743_42282.t3 25.8467
R23815 a_743_42282.n0 a_743_42282.t2 25.8467
R23816 a_743_42282.t1 a_743_42282.n8 25.8467
R23817 a_743_42282.n8 a_743_42282.t0 25.8467
R23818 a_743_42282.n6 a_743_42282.n5 11.7104
R23819 a_743_42282.n6 a_743_42282.n2 0.229071
R23820 a_n4064_39616.n6 a_n4064_39616.t9 1415.15
R23821 a_n4064_39616.n5 a_n4064_39616.t11 1330.32
R23822 a_n4064_39616.n4 a_n4064_39616.t8 1320.68
R23823 a_n4064_39616.n6 a_n4064_39616.t13 1320.68
R23824 a_n4064_39616.n11 a_n4064_39616.n10 360.399
R23825 a_n4064_39616.n3 a_n4064_39616.t12 241.536
R23826 a_n4064_39616.n2 a_n4064_39616.n1 232.862
R23827 a_n4064_39616.n12 a_n4064_39616.n11 203.161
R23828 a_n4064_39616.n8 a_n4064_39616.n3 172.543
R23829 a_n4064_39616.n3 a_n4064_39616.t10 169.237
R23830 a_n4064_39616.n7 a_n4064_39616.n4 161.764
R23831 a_n4064_39616.n7 a_n4064_39616.n6 161.3
R23832 a_n4064_39616.n2 a_n4064_39616.n0 95.6721
R23833 a_n4064_39616.n6 a_n4064_39616.n5 84.8325
R23834 a_n4064_39616.n5 a_n4064_39616.n4 84.8325
R23835 a_n4064_39616.n8 a_n4064_39616.n7 79.6846
R23836 a_n4064_39616.n9 a_n4064_39616.n2 61.9632
R23837 a_n4064_39616.n10 a_n4064_39616.t2 27.5805
R23838 a_n4064_39616.n10 a_n4064_39616.t1 27.5805
R23839 a_n4064_39616.n12 a_n4064_39616.t0 27.5805
R23840 a_n4064_39616.t3 a_n4064_39616.n12 27.5805
R23841 a_n4064_39616.n1 a_n4064_39616.t7 25.8467
R23842 a_n4064_39616.n1 a_n4064_39616.t6 25.8467
R23843 a_n4064_39616.n0 a_n4064_39616.t4 25.8467
R23844 a_n4064_39616.n0 a_n4064_39616.t5 25.8467
R23845 a_n4064_39616.n11 a_n4064_39616.n9 21.2775
R23846 a_n4064_39616.n9 a_n4064_39616.n8 9.3005
R23847 a_n2293_43922.n1 a_n2293_43922.n0 282.245
R23848 a_n2293_43922.n0 a_n2293_43922.t3 276.464
R23849 a_n2293_43922.n2 a_n2293_43922.n1 259.06
R23850 a_n2293_43922.n0 a_n2293_43922.t4 196.131
R23851 a_n2293_43922.n1 a_n2293_43922.t2 131.308
R23852 a_n2293_43922.t0 a_n2293_43922.n2 26.5955
R23853 a_n2293_43922.n2 a_n2293_43922.t1 26.5955
R23854 a_3232_43370.n3 a_3232_43370.t7 265.101
R23855 a_3232_43370.n4 a_3232_43370.t20 263.493
R23856 a_3232_43370.n1 a_3232_43370.t23 263.493
R23857 a_3232_43370.n14 a_3232_43370.t15 254.256
R23858 a_3232_43370.n21 a_3232_43370.n20 243.679
R23859 a_3232_43370.n12 a_3232_43370.t19 240.484
R23860 a_3232_43370.n8 a_3232_43370.t11 239.505
R23861 a_3232_43370.n10 a_3232_43370.t10 230.155
R23862 a_3232_43370.n6 a_3232_43370.t6 230.155
R23863 a_3232_43370.n13 a_3232_43370.n12 227.15
R23864 a_3232_43370.n9 a_3232_43370.t8 212.081
R23865 a_3232_43370.n18 a_3232_43370.n0 209.448
R23866 a_3232_43370.n11 a_3232_43370.n9 207.758
R23867 a_3232_43370.n20 a_3232_43370.n19 205.28
R23868 a_3232_43370.n7 a_3232_43370.n3 186.225
R23869 a_3232_43370.n14 a_3232_43370.t14 181.956
R23870 a_3232_43370.n16 a_3232_43370.n8 177.665
R23871 a_3232_43370.n7 a_3232_43370.n6 174.191
R23872 a_3232_43370.n11 a_3232_43370.n10 168.851
R23873 a_3232_43370.n12 a_3232_43370.t12 168.185
R23874 a_3232_43370.n8 a_3232_43370.t13 167.204
R23875 a_3232_43370.n9 a_3232_43370.t9 165.341
R23876 a_3232_43370.n15 a_3232_43370.n14 164.958
R23877 a_3232_43370.n2 a_3232_43370.t21 160.667
R23878 a_3232_43370.n10 a_3232_43370.t17 157.856
R23879 a_3232_43370.n5 a_3232_43370.t16 133.353
R23880 a_3232_43370.n4 a_3232_43370.t18 128.534
R23881 a_3232_43370.n1 a_3232_43370.t22 128.534
R23882 a_3232_43370.n5 a_3232_43370.n4 83.4688
R23883 a_3232_43370.n2 a_3232_43370.n1 83.4688
R23884 a_3232_43370.n20 a_3232_43370.n18 52.1955
R23885 a_3232_43370.n16 a_3232_43370.n15 39.1045
R23886 a_3232_43370.n3 a_3232_43370.n2 32.1338
R23887 a_3232_43370.n19 a_3232_43370.t2 26.5955
R23888 a_3232_43370.n19 a_3232_43370.t3 26.5955
R23889 a_3232_43370.n21 a_3232_43370.t0 26.5955
R23890 a_3232_43370.t1 a_3232_43370.n21 26.5955
R23891 a_3232_43370.n0 a_3232_43370.t4 24.9236
R23892 a_3232_43370.n0 a_3232_43370.t5 24.9236
R23893 a_3232_43370.n17 a_3232_43370.n16 21.7546
R23894 a_3232_43370.n18 a_3232_43370.n17 14.8829
R23895 a_3232_43370.n15 a_3232_43370.n13 10.1087
R23896 a_3232_43370.n17 a_3232_43370.n7 9.00599
R23897 a_3232_43370.n6 a_3232_43370.n5 8.76414
R23898 a_3232_43370.n13 a_3232_43370.n11 5.43457
R23899 a_1666_39043.n2 a_1666_39043.t5 440.13
R23900 a_1666_39043.n0 a_1666_39043.t2 239.113
R23901 a_1666_39043.n1 a_1666_39043.t6 230.576
R23902 a_1666_39043.n2 a_1666_39043.t4 192.331
R23903 a_1666_39043.n3 a_1666_39043.n1 170.291
R23904 a_1666_39043.n1 a_1666_39043.t3 158.275
R23905 a_1666_39043.t0 a_1666_39043.n4 85.6451
R23906 a_1666_39043.n0 a_1666_39043.t1 61.169
R23907 a_1666_39043.n4 a_1666_39043.n3 5.84425
R23908 a_1666_39043.n3 a_1666_39043.n2 4.5005
R23909 a_1666_39043.n4 a_1666_39043.n0 1.59495
R23910 a_n3420_39072.n3 a_n3420_39072.t10 444.502
R23911 a_n3420_39072.n8 a_n3420_39072.n7 360.399
R23912 a_n3420_39072.n3 a_n3420_39072.t9 356.68
R23913 a_n3420_39072.n5 a_n3420_39072.n3 257.639
R23914 a_n3420_39072.n4 a_n3420_39072.t8 241.536
R23915 a_n3420_39072.n2 a_n3420_39072.n1 232.862
R23916 a_n3420_39072.n9 a_n3420_39072.n8 203.161
R23917 a_n3420_39072.n4 a_n3420_39072.t11 169.237
R23918 a_n3420_39072.n5 a_n3420_39072.n4 167.149
R23919 a_n3420_39072.n2 a_n3420_39072.n0 95.6721
R23920 a_n3420_39072.n6 a_n3420_39072.n2 60.5918
R23921 a_n3420_39072.n7 a_n3420_39072.t2 27.5805
R23922 a_n3420_39072.n7 a_n3420_39072.t1 27.5805
R23923 a_n3420_39072.t3 a_n3420_39072.n9 27.5805
R23924 a_n3420_39072.n9 a_n3420_39072.t0 27.5805
R23925 a_n3420_39072.n1 a_n3420_39072.t6 25.8467
R23926 a_n3420_39072.n1 a_n3420_39072.t4 25.8467
R23927 a_n3420_39072.n0 a_n3420_39072.t5 25.8467
R23928 a_n3420_39072.n0 a_n3420_39072.t7 25.8467
R23929 a_n3420_39072.n8 a_n3420_39072.n6 22.6489
R23930 a_n3420_39072.n6 a_n3420_39072.n5 9.3012
R23931 a_19237_31679.n1 a_19237_31679.t4 602.944
R23932 a_19237_31679.n2 a_19237_31679.n1 287.752
R23933 a_19237_31679.n1 a_19237_31679.n0 277.568
R23934 a_19237_31679.t1 a_19237_31679.n2 26.5955
R23935 a_19237_31679.n2 a_19237_31679.t0 26.5955
R23936 a_19237_31679.n0 a_19237_31679.t3 24.9236
R23937 a_19237_31679.n0 a_19237_31679.t2 24.9236
R23938 a_n2312_39304.n3 a_n2312_39304.n2 287.752
R23939 a_n2312_39304.n2 a_n2312_39304.n0 277.568
R23940 a_n2312_39304.n2 a_n2312_39304.n1 271.13
R23941 a_n2312_39304.n1 a_n2312_39304.t4 228.649
R23942 a_n2312_39304.n1 a_n2312_39304.t5 156.35
R23943 a_n2312_39304.t1 a_n2312_39304.n3 26.5955
R23944 a_n2312_39304.n3 a_n2312_39304.t0 26.5955
R23945 a_n2312_39304.n0 a_n2312_39304.t3 24.9236
R23946 a_n2312_39304.n0 a_n2312_39304.t2 24.9236
R23947 a_10193_42453.n3 a_10193_42453.t5 722.096
R23948 a_10193_42453.n13 a_10193_42453.t8 722.096
R23949 a_10193_42453.n11 a_10193_42453.t12 722.096
R23950 a_10193_42453.n9 a_10193_42453.t4 722.096
R23951 a_10193_42453.n21 a_10193_42453.n20 380.32
R23952 a_10193_42453.n4 a_10193_42453.t18 241.536
R23953 a_10193_42453.n15 a_10193_42453.t7 241.536
R23954 a_10193_42453.n7 a_10193_42453.t14 241.536
R23955 a_10193_42453.n6 a_10193_42453.t23 241.536
R23956 a_10193_42453.n1 a_10193_42453.t20 241.536
R23957 a_10193_42453.n0 a_10193_42453.t13 230.155
R23958 a_10193_42453.n5 a_10193_42453.n4 199.482
R23959 a_10193_42453.n8 a_10193_42453.n6 187.677
R23960 a_10193_42453.n20 a_10193_42453.n19 185
R23961 a_10193_42453.n12 a_10193_42453.n11 180.619
R23962 a_10193_42453.n16 a_10193_42453.n15 180.496
R23963 a_10193_42453.n14 a_10193_42453.n13 179.311
R23964 a_10193_42453.n5 a_10193_42453.n3 175.577
R23965 a_10193_42453.n10 a_10193_42453.n9 172.516
R23966 a_10193_42453.n2 a_10193_42453.n1 171.775
R23967 a_10193_42453.n4 a_10193_42453.t9 169.237
R23968 a_10193_42453.n15 a_10193_42453.t21 169.237
R23969 a_10193_42453.n7 a_10193_42453.t17 169.237
R23970 a_10193_42453.n6 a_10193_42453.t6 169.237
R23971 a_10193_42453.n1 a_10193_42453.t11 169.237
R23972 a_10193_42453.n8 a_10193_42453.n7 168.183
R23973 a_10193_42453.n3 a_10193_42453.t10 162.963
R23974 a_10193_42453.n13 a_10193_42453.t22 162.963
R23975 a_10193_42453.n11 a_10193_42453.t19 162.963
R23976 a_10193_42453.n9 a_10193_42453.t15 162.963
R23977 a_10193_42453.n2 a_10193_42453.n0 162.868
R23978 a_10193_42453.n0 a_10193_42453.t16 157.856
R23979 a_10193_42453.t1 a_10193_42453.n21 26.5955
R23980 a_10193_42453.n21 a_10193_42453.t0 26.5955
R23981 a_10193_42453.n16 a_10193_42453.n14 25.6653
R23982 a_10193_42453.n19 a_10193_42453.t3 24.9236
R23983 a_10193_42453.n19 a_10193_42453.t2 24.9236
R23984 a_10193_42453.n20 a_10193_42453.n18 16.6197
R23985 a_10193_42453.n10 a_10193_42453.n8 15.5506
R23986 a_10193_42453.n14 a_10193_42453.n12 15.0939
R23987 a_10193_42453.n18 a_10193_42453.n17 8.68953
R23988 a_10193_42453.n17 a_10193_42453.n5 6.07519
R23989 a_10193_42453.n18 a_10193_42453.n2 6.02162
R23990 a_10193_42453.n17 a_10193_42453.n16 1.21805
R23991 a_10193_42453.n12 a_10193_42453.n10 0.475775
R23992 a_6151_47436.n6 a_6151_47436.t12 408.63
R23993 a_6151_47436.n2 a_6151_47436.t9 408.63
R23994 a_6151_47436.t0 a_6151_47436.n11 375.046
R23995 a_6151_47436.n7 a_6151_47436.t2 347.577
R23996 a_6151_47436.n3 a_6151_47436.t7 347.577
R23997 a_6151_47436.n11 a_6151_47436.t1 299.062
R23998 a_6151_47436.n0 a_6151_47436.t3 276.464
R23999 a_6151_47436.n1 a_6151_47436.t8 238.59
R24000 a_6151_47436.n1 a_6151_47436.t6 203.244
R24001 a_6151_47436.n0 a_6151_47436.t4 196.131
R24002 a_6151_47436.n7 a_6151_47436.t13 193.337
R24003 a_6151_47436.n3 a_6151_47436.t10 193.337
R24004 a_6151_47436.n5 a_6151_47436.n1 179.07
R24005 a_6151_47436.n8 a_6151_47436.n6 167.607
R24006 a_6151_47436.n4 a_6151_47436.n2 165.179
R24007 a_6151_47436.n10 a_6151_47436.n0 165.179
R24008 a_6151_47436.n4 a_6151_47436.n3 162.834
R24009 a_6151_47436.n8 a_6151_47436.n7 160.472
R24010 a_6151_47436.n6 a_6151_47436.t11 132.282
R24011 a_6151_47436.n2 a_6151_47436.t5 132.282
R24012 a_6151_47436.n10 a_6151_47436.n9 36.5102
R24013 a_6151_47436.n5 a_6151_47436.n4 14.9401
R24014 a_6151_47436.n9 a_6151_47436.n5 10.0194
R24015 a_6151_47436.n11 a_6151_47436.n10 9.3005
R24016 a_6151_47436.n9 a_6151_47436.n8 0.141324
R24017 a_4190_30871.n19 a_4190_30871.t21 1421.83
R24018 a_4190_30871.n9 a_4190_30871.t16 1421.83
R24019 a_4190_30871.n12 a_4190_30871.t8 1327.11
R24020 a_4190_30871.n16 a_4190_30871.t19 1327.11
R24021 a_4190_30871.n18 a_4190_30871.t20 1327.11
R24022 a_4190_30871.n8 a_4190_30871.t4 1327.11
R24023 a_4190_30871.n6 a_4190_30871.t15 1327.11
R24024 a_4190_30871.n2 a_4190_30871.t5 1327.11
R24025 a_4190_30871.n19 a_4190_30871.t10 1320.68
R24026 a_4190_30871.n17 a_4190_30871.t12 1320.68
R24027 a_4190_30871.n15 a_4190_30871.t13 1320.68
R24028 a_4190_30871.n13 a_4190_30871.t6 1320.68
R24029 a_4190_30871.n3 a_4190_30871.t14 1320.68
R24030 a_4190_30871.n5 a_4190_30871.t11 1320.68
R24031 a_4190_30871.n7 a_4190_30871.t7 1320.68
R24032 a_4190_30871.n9 a_4190_30871.t18 1320.68
R24033 a_4190_30871.n25 a_4190_30871.n24 287.752
R24034 a_4190_30871.n24 a_4190_30871.n0 277.568
R24035 a_4190_30871.n22 a_4190_30871.t17 260.322
R24036 a_4190_30871.n23 a_4190_30871.n22 189.659
R24037 a_4190_30871.n22 a_4190_30871.t9 175.169
R24038 a_4190_30871.n14 a_4190_30871.n13 161.701
R24039 a_4190_30871.n4 a_4190_30871.n3 161.701
R24040 a_4190_30871.n20 a_4190_30871.n19 161.3
R24041 a_4190_30871.n15 a_4190_30871.n14 161.3
R24042 a_4190_30871.n17 a_4190_30871.n11 161.3
R24043 a_4190_30871.n10 a_4190_30871.n9 161.3
R24044 a_4190_30871.n7 a_4190_30871.n1 161.3
R24045 a_4190_30871.n5 a_4190_30871.n4 161.3
R24046 a_4190_30871.n13 a_4190_30871.n12 94.7191
R24047 a_4190_30871.n15 a_4190_30871.n12 94.7191
R24048 a_4190_30871.n16 a_4190_30871.n15 94.7191
R24049 a_4190_30871.n17 a_4190_30871.n16 94.7191
R24050 a_4190_30871.n18 a_4190_30871.n17 94.7191
R24051 a_4190_30871.n19 a_4190_30871.n18 94.7191
R24052 a_4190_30871.n9 a_4190_30871.n8 94.7191
R24053 a_4190_30871.n8 a_4190_30871.n7 94.7191
R24054 a_4190_30871.n7 a_4190_30871.n6 94.7191
R24055 a_4190_30871.n6 a_4190_30871.n5 94.7191
R24056 a_4190_30871.n5 a_4190_30871.n2 94.7191
R24057 a_4190_30871.n3 a_4190_30871.n2 94.7191
R24058 a_4190_30871.n23 a_4190_30871.n21 77.1582
R24059 a_4190_30871.n21 a_4190_30871.n20 38.8203
R24060 a_4190_30871.n21 a_4190_30871.n10 35.3495
R24061 a_4190_30871.n24 a_4190_30871.n23 33.2329
R24062 a_4190_30871.t1 a_4190_30871.n25 26.5955
R24063 a_4190_30871.n25 a_4190_30871.t0 26.5955
R24064 a_4190_30871.n0 a_4190_30871.t3 24.9236
R24065 a_4190_30871.n0 a_4190_30871.t2 24.9236
R24066 a_4190_30871.n14 a_4190_30871.n11 0.4005
R24067 a_4190_30871.n20 a_4190_30871.n11 0.4005
R24068 a_4190_30871.n10 a_4190_30871.n1 0.4005
R24069 a_4190_30871.n4 a_4190_30871.n1 0.4005
R24070 C10_N_btm C10_N_btm.n32 90.5213
R24071 C10_N_btm.n2 C10_N_btm.n0 33.0802
R24072 C10_N_btm.n14 C10_N_btm.n13 32.3614
R24073 C10_N_btm.n12 C10_N_btm.n11 32.3614
R24074 C10_N_btm.n10 C10_N_btm.n9 32.3614
R24075 C10_N_btm.n8 C10_N_btm.n7 32.3614
R24076 C10_N_btm.n6 C10_N_btm.n5 32.3614
R24077 C10_N_btm.n4 C10_N_btm.n3 32.3614
R24078 C10_N_btm.n2 C10_N_btm.n1 32.3614
R24079 C10_N_btm.n22 C10_N_btm.n14 29.1203
R24080 C10_N_btm.n24 C10_N_btm.n23 20.3263
R24081 C10_N_btm.n28 C10_N_btm.n26 15.4755
R24082 C10_N_btm.n17 C10_N_btm.n15 15.394
R24083 C10_N_btm.n30 C10_N_btm.n29 14.9755
R24084 C10_N_btm.n31 C10_N_btm.n25 14.9755
R24085 C10_N_btm.n28 C10_N_btm.n27 14.9755
R24086 C10_N_btm.n21 C10_N_btm.n20 14.894
R24087 C10_N_btm.n19 C10_N_btm.n18 14.894
R24088 C10_N_btm.n17 C10_N_btm.n16 14.894
R24089 C10_N_btm.n24 C10_N_btm.n22 6.29217
R24090 C10_N_btm.n22 C10_N_btm.n21 5.43279
R24091 C10_N_btm C10_N_btm.n1044 5.34972
R24092 C10_N_btm.n32 C10_N_btm.n31 5.33904
R24093 C10_N_btm.n32 C10_N_btm.n24 4.7505
R24094 C10_N_btm.n13 C10_N_btm.t10 3.57113
R24095 C10_N_btm.n13 C10_N_btm.t9 3.57113
R24096 C10_N_btm.n11 C10_N_btm.t22 3.57113
R24097 C10_N_btm.n11 C10_N_btm.t17 3.57113
R24098 C10_N_btm.n9 C10_N_btm.t13 3.57113
R24099 C10_N_btm.n9 C10_N_btm.t16 3.57113
R24100 C10_N_btm.n7 C10_N_btm.t23 3.57113
R24101 C10_N_btm.n7 C10_N_btm.t19 3.57113
R24102 C10_N_btm.n5 C10_N_btm.t11 3.57113
R24103 C10_N_btm.n5 C10_N_btm.t21 3.57113
R24104 C10_N_btm.n3 C10_N_btm.t15 3.57113
R24105 C10_N_btm.n3 C10_N_btm.t8 3.57113
R24106 C10_N_btm.n1 C10_N_btm.t18 3.57113
R24107 C10_N_btm.n1 C10_N_btm.t20 3.57113
R24108 C10_N_btm.n0 C10_N_btm.t12 3.57113
R24109 C10_N_btm.n0 C10_N_btm.t14 3.57113
R24110 C10_N_btm.n26 C10_N_btm.t1 2.4755
R24111 C10_N_btm.n26 C10_N_btm.t7 2.4755
R24112 C10_N_btm.n29 C10_N_btm.t2 2.4755
R24113 C10_N_btm.n29 C10_N_btm.t5 2.4755
R24114 C10_N_btm.n25 C10_N_btm.t6 2.4755
R24115 C10_N_btm.n25 C10_N_btm.t3 2.4755
R24116 C10_N_btm.n23 C10_N_btm.t32 2.4755
R24117 C10_N_btm.n23 C10_N_btm.t33 2.4755
R24118 C10_N_btm.n20 C10_N_btm.t31 2.4755
R24119 C10_N_btm.n20 C10_N_btm.t28 2.4755
R24120 C10_N_btm.n18 C10_N_btm.t25 2.4755
R24121 C10_N_btm.n18 C10_N_btm.t26 2.4755
R24122 C10_N_btm.n16 C10_N_btm.t29 2.4755
R24123 C10_N_btm.n16 C10_N_btm.t24 2.4755
R24124 C10_N_btm.n15 C10_N_btm.t27 2.4755
R24125 C10_N_btm.n15 C10_N_btm.t30 2.4755
R24126 C10_N_btm.n27 C10_N_btm.t0 2.4755
R24127 C10_N_btm.n27 C10_N_btm.t4 2.4755
R24128 C10_N_btm.n4 C10_N_btm.n2 0.71925
R24129 C10_N_btm.n8 C10_N_btm.n6 0.71925
R24130 C10_N_btm.n12 C10_N_btm.n10 0.71925
R24131 C10_N_btm.n6 C10_N_btm.n4 0.688
R24132 C10_N_btm.n10 C10_N_btm.n8 0.688
R24133 C10_N_btm.n14 C10_N_btm.n12 0.672375
R24134 C10_N_btm.n19 C10_N_btm.n17 0.5005
R24135 C10_N_btm.n30 C10_N_btm.n28 0.5005
R24136 C10_N_btm.n31 C10_N_btm.n30 0.484875
R24137 C10_N_btm.n21 C10_N_btm.n19 0.453625
R24138 C10_N_btm.n182 C10_N_btm.n181 0.276161
R24139 C10_N_btm.n217 C10_N_btm.n216 0.276161
R24140 C10_N_btm.n645 C10_N_btm.n644 0.276161
R24141 C10_N_btm.n429 C10_N_btm.n424 0.276161
R24142 C10_N_btm.n598 C10_N_btm.n597 0.276161
R24143 C10_N_btm.n185 C10_N_btm.n183 0.228786
R24144 C10_N_btm.n183 C10_N_btm.n182 0.228786
R24145 C10_N_btm.n186 C10_N_btm.n185 0.228786
R24146 C10_N_btm.n187 C10_N_btm.n186 0.228786
R24147 C10_N_btm.n190 C10_N_btm.n188 0.228786
R24148 C10_N_btm.n188 C10_N_btm.n187 0.228786
R24149 C10_N_btm.n191 C10_N_btm.n190 0.228786
R24150 C10_N_btm.n192 C10_N_btm.n191 0.228786
R24151 C10_N_btm.n195 C10_N_btm.n193 0.228786
R24152 C10_N_btm.n193 C10_N_btm.n192 0.228786
R24153 C10_N_btm.n196 C10_N_btm.n195 0.228786
R24154 C10_N_btm.n197 C10_N_btm.n196 0.228786
R24155 C10_N_btm.n200 C10_N_btm.n198 0.228786
R24156 C10_N_btm.n198 C10_N_btm.n197 0.228786
R24157 C10_N_btm.n201 C10_N_btm.n200 0.228786
R24158 C10_N_btm.n202 C10_N_btm.n201 0.228786
R24159 C10_N_btm.n205 C10_N_btm.n203 0.228786
R24160 C10_N_btm.n203 C10_N_btm.n202 0.228786
R24161 C10_N_btm.n206 C10_N_btm.n205 0.228786
R24162 C10_N_btm.n207 C10_N_btm.n206 0.228786
R24163 C10_N_btm.n210 C10_N_btm.n208 0.228786
R24164 C10_N_btm.n208 C10_N_btm.n207 0.228786
R24165 C10_N_btm.n211 C10_N_btm.n210 0.228786
R24166 C10_N_btm.n212 C10_N_btm.n211 0.228786
R24167 C10_N_btm.n215 C10_N_btm.n213 0.228786
R24168 C10_N_btm.n213 C10_N_btm.n212 0.228786
R24169 C10_N_btm.n216 C10_N_btm.n215 0.228786
R24170 C10_N_btm.n924 C10_N_btm.n923 0.228786
R24171 C10_N_btm.n922 C10_N_btm.n178 0.228786
R24172 C10_N_btm.n921 C10_N_btm.n218 0.228786
R24173 C10_N_btm.n920 C10_N_btm.n919 0.228786
R24174 C10_N_btm.n918 C10_N_btm.n219 0.228786
R24175 C10_N_btm.n236 C10_N_btm.n221 0.228786
R24176 C10_N_btm.n903 C10_N_btm.n902 0.228786
R24177 C10_N_btm.n901 C10_N_btm.n235 0.228786
R24178 C10_N_btm.n900 C10_N_btm.n237 0.228786
R24179 C10_N_btm.n899 C10_N_btm.n898 0.228786
R24180 C10_N_btm.n897 C10_N_btm.n238 0.228786
R24181 C10_N_btm.n255 C10_N_btm.n240 0.228786
R24182 C10_N_btm.n879 C10_N_btm.n878 0.228786
R24183 C10_N_btm.n877 C10_N_btm.n254 0.228786
R24184 C10_N_btm.n644 C10_N_btm.n409 0.228786
R24185 C10_N_btm.n408 C10_N_btm.n407 0.228786
R24186 C10_N_btm.n409 C10_N_btm.n408 0.228786
R24187 C10_N_btm.n407 C10_N_btm.n406 0.228786
R24188 C10_N_btm.n406 C10_N_btm.n400 0.228786
R24189 C10_N_btm.n399 C10_N_btm.n398 0.228786
R24190 C10_N_btm.n400 C10_N_btm.n399 0.228786
R24191 C10_N_btm.n398 C10_N_btm.n397 0.228786
R24192 C10_N_btm.n397 C10_N_btm.n391 0.228786
R24193 C10_N_btm.n390 C10_N_btm.n389 0.228786
R24194 C10_N_btm.n391 C10_N_btm.n390 0.228786
R24195 C10_N_btm.n389 C10_N_btm.n388 0.228786
R24196 C10_N_btm.n388 C10_N_btm.n382 0.228786
R24197 C10_N_btm.n671 C10_N_btm.n379 0.228786
R24198 C10_N_btm.n382 C10_N_btm.n379 0.228786
R24199 C10_N_btm.n672 C10_N_btm.n671 0.228786
R24200 C10_N_btm.n673 C10_N_btm.n672 0.228786
R24201 C10_N_btm.n675 C10_N_btm.n375 0.228786
R24202 C10_N_btm.n675 C10_N_btm.n674 0.228786
R24203 C10_N_btm.n674 C10_N_btm.n673 0.228786
R24204 C10_N_btm.n375 C10_N_btm.n374 0.228786
R24205 C10_N_btm.n596 C10_N_btm.n595 0.228786
R24206 C10_N_btm.n594 C10_N_btm.n465 0.228786
R24207 C10_N_btm.n516 C10_N_btm.n466 0.228786
R24208 C10_N_btm.n517 C10_N_btm.n515 0.228786
R24209 C10_N_btm.n519 C10_N_btm.n518 0.228786
R24210 C10_N_btm.n351 C10_N_btm.n350 0.228786
R24211 C10_N_btm.n689 C10_N_btm.n688 0.228786
R24212 C10_N_btm.n690 C10_N_btm.n349 0.228786
R24213 C10_N_btm.n713 C10_N_btm.n712 0.228786
R24214 C10_N_btm.n711 C10_N_btm.n347 0.228786
R24215 C10_N_btm.n710 C10_N_btm.n709 0.228786
R24216 C10_N_btm.n708 C10_N_btm.n691 0.228786
R24217 C10_N_btm.n695 C10_N_btm.n692 0.228786
R24218 C10_N_btm.n698 C10_N_btm.n697 0.228786
R24219 C10_N_btm.n696 C10_N_btm.n694 0.228786
R24220 C10_N_btm.n317 C10_N_btm.n316 0.228786
R24221 C10_N_btm.n734 C10_N_btm.n733 0.228786
R24222 C10_N_btm.n735 C10_N_btm.n315 0.228786
R24223 C10_N_btm.n816 C10_N_btm.n815 0.228786
R24224 C10_N_btm.n814 C10_N_btm.n313 0.228786
R24225 C10_N_btm.n813 C10_N_btm.n812 0.228786
R24226 C10_N_btm.n811 C10_N_btm.n736 0.228786
R24227 C10_N_btm.n744 C10_N_btm.n737 0.228786
R24228 C10_N_btm.n745 C10_N_btm.n743 0.228786
R24229 C10_N_btm.n802 C10_N_btm.n746 0.228786
R24230 C10_N_btm.n801 C10_N_btm.n800 0.228786
R24231 C10_N_btm.n799 C10_N_btm.n747 0.228786
R24232 C10_N_btm.n798 C10_N_btm.n748 0.228786
R24233 C10_N_btm.n797 C10_N_btm.n796 0.228786
R24234 C10_N_btm.n795 C10_N_btm.n749 0.228786
R24235 C10_N_btm.n768 C10_N_btm.n751 0.228786
R24236 C10_N_btm.n769 C10_N_btm.n767 0.228786
R24237 C10_N_btm.n786 C10_N_btm.n770 0.228786
R24238 C10_N_btm.n785 C10_N_btm.n784 0.228786
R24239 C10_N_btm.n783 C10_N_btm.n771 0.228786
R24240 C10_N_btm.n782 C10_N_btm.n772 0.228786
R24241 C10_N_btm.n781 C10_N_btm.n780 0.228786
R24242 C10_N_btm.n284 C10_N_btm.n283 0.228786
R24243 C10_N_btm.n848 C10_N_btm.n847 0.228786
R24244 C10_N_btm.n849 C10_N_btm.n282 0.228786
R24245 C10_N_btm.n856 C10_N_btm.n850 0.228786
R24246 C10_N_btm.n855 C10_N_btm.n854 0.228786
R24247 C10_N_btm.n853 C10_N_btm.n852 0.228786
R24248 C10_N_btm.n258 C10_N_btm.n257 0.228786
R24249 C10_N_btm.n875 C10_N_btm.n874 0.228786
R24250 C10_N_btm.n128 C10_N_btm.n35 0.228786
R24251 C10_N_btm.n129 C10_N_btm.n127 0.228786
R24252 C10_N_btm.n973 C10_N_btm.n972 0.228786
R24253 C10_N_btm.n971 C10_N_btm.n124 0.228786
R24254 C10_N_btm.n970 C10_N_btm.n130 0.228786
R24255 C10_N_btm.n969 C10_N_btm.n968 0.228786
R24256 C10_N_btm.n967 C10_N_btm.n131 0.228786
R24257 C10_N_btm.n135 C10_N_btm.n134 0.228786
R24258 C10_N_btm.n134 C10_N_btm.n133 0.228786
R24259 C10_N_btm.n967 C10_N_btm.n966 0.228786
R24260 C10_N_btm.n966 C10_N_btm.n965 0.228786
R24261 C10_N_btm.n964 C10_N_btm.n132 0.228786
R24262 C10_N_btm.n968 C10_N_btm.n132 0.228786
R24263 C10_N_btm.n130 C10_N_btm.n123 0.228786
R24264 C10_N_btm.n123 C10_N_btm.n122 0.228786
R24265 C10_N_btm.n976 C10_N_btm.n975 0.228786
R24266 C10_N_btm.n975 C10_N_btm.n124 0.228786
R24267 C10_N_btm.n974 C10_N_btm.n973 0.228786
R24268 C10_N_btm.n974 C10_N_btm.n120 0.228786
R24269 C10_N_btm.n126 C10_N_btm.n125 0.228786
R24270 C10_N_btm.n127 C10_N_btm.n126 0.228786
R24271 C10_N_btm.n36 C10_N_btm.n35 0.228786
R24272 C10_N_btm.n38 C10_N_btm.n36 0.228786
R24273 C10_N_btm.n117 C10_N_btm.n39 0.228786
R24274 C10_N_btm.n39 C10_N_btm.n38 0.228786
R24275 C10_N_btm.n125 C10_N_btm.n119 0.228786
R24276 C10_N_btm.n119 C10_N_btm.n118 0.228786
R24277 C10_N_btm.n979 C10_N_btm.n978 0.228786
R24278 C10_N_btm.n978 C10_N_btm.n120 0.228786
R24279 C10_N_btm.n977 C10_N_btm.n976 0.228786
R24280 C10_N_btm.n977 C10_N_btm.n113 0.228786
R24281 C10_N_btm.n137 C10_N_btm.n121 0.228786
R24282 C10_N_btm.n122 C10_N_btm.n121 0.228786
R24283 C10_N_btm.n964 C10_N_btm.n963 0.228786
R24284 C10_N_btm.n963 C10_N_btm.n962 0.228786
R24285 C10_N_btm.n961 C10_N_btm.n136 0.228786
R24286 C10_N_btm.n965 C10_N_btm.n136 0.228786
R24287 C10_N_btm.n184 C10_N_btm.n135 0.228786
R24288 C10_N_btm.n184 C10_N_btm.n139 0.228786
R24289 C10_N_btm.n141 C10_N_btm.n140 0.228786
R24290 C10_N_btm.n140 C10_N_btm.n139 0.228786
R24291 C10_N_btm.n961 C10_N_btm.n960 0.228786
R24292 C10_N_btm.n960 C10_N_btm.n959 0.228786
R24293 C10_N_btm.n958 C10_N_btm.n138 0.228786
R24294 C10_N_btm.n962 C10_N_btm.n138 0.228786
R24295 C10_N_btm.n137 C10_N_btm.n112 0.228786
R24296 C10_N_btm.n112 C10_N_btm.n111 0.228786
R24297 C10_N_btm.n982 C10_N_btm.n981 0.228786
R24298 C10_N_btm.n981 C10_N_btm.n113 0.228786
R24299 C10_N_btm.n980 C10_N_btm.n979 0.228786
R24300 C10_N_btm.n980 C10_N_btm.n109 0.228786
R24301 C10_N_btm.n115 C10_N_btm.n114 0.228786
R24302 C10_N_btm.n118 C10_N_btm.n115 0.228786
R24303 C10_N_btm.n117 C10_N_btm.n116 0.228786
R24304 C10_N_btm.n116 C10_N_btm.n43 0.228786
R24305 C10_N_btm.n46 C10_N_btm.n44 0.228786
R24306 C10_N_btm.n44 C10_N_btm.n43 0.228786
R24307 C10_N_btm.n114 C10_N_btm.n108 0.228786
R24308 C10_N_btm.n108 C10_N_btm.n107 0.228786
R24309 C10_N_btm.n985 C10_N_btm.n984 0.228786
R24310 C10_N_btm.n984 C10_N_btm.n109 0.228786
R24311 C10_N_btm.n983 C10_N_btm.n982 0.228786
R24312 C10_N_btm.n983 C10_N_btm.n102 0.228786
R24313 C10_N_btm.n143 C10_N_btm.n110 0.228786
R24314 C10_N_btm.n111 C10_N_btm.n110 0.228786
R24315 C10_N_btm.n958 C10_N_btm.n957 0.228786
R24316 C10_N_btm.n957 C10_N_btm.n956 0.228786
R24317 C10_N_btm.n955 C10_N_btm.n142 0.228786
R24318 C10_N_btm.n959 C10_N_btm.n142 0.228786
R24319 C10_N_btm.n189 C10_N_btm.n141 0.228786
R24320 C10_N_btm.n189 C10_N_btm.n145 0.228786
R24321 C10_N_btm.n147 C10_N_btm.n146 0.228786
R24322 C10_N_btm.n146 C10_N_btm.n145 0.228786
R24323 C10_N_btm.n955 C10_N_btm.n954 0.228786
R24324 C10_N_btm.n954 C10_N_btm.n953 0.228786
R24325 C10_N_btm.n952 C10_N_btm.n144 0.228786
R24326 C10_N_btm.n956 C10_N_btm.n144 0.228786
R24327 C10_N_btm.n143 C10_N_btm.n101 0.228786
R24328 C10_N_btm.n101 C10_N_btm.n100 0.228786
R24329 C10_N_btm.n988 C10_N_btm.n987 0.228786
R24330 C10_N_btm.n987 C10_N_btm.n102 0.228786
R24331 C10_N_btm.n986 C10_N_btm.n985 0.228786
R24332 C10_N_btm.n986 C10_N_btm.n98 0.228786
R24333 C10_N_btm.n106 C10_N_btm.n105 0.228786
R24334 C10_N_btm.n107 C10_N_btm.n106 0.228786
R24335 C10_N_btm.n47 C10_N_btm.n46 0.228786
R24336 C10_N_btm.n104 C10_N_btm.n47 0.228786
R24337 C10_N_btm.n103 C10_N_btm.n51 0.228786
R24338 C10_N_btm.n104 C10_N_btm.n103 0.228786
R24339 C10_N_btm.n105 C10_N_btm.n97 0.228786
R24340 C10_N_btm.n97 C10_N_btm.n96 0.228786
R24341 C10_N_btm.n991 C10_N_btm.n990 0.228786
R24342 C10_N_btm.n990 C10_N_btm.n98 0.228786
R24343 C10_N_btm.n989 C10_N_btm.n988 0.228786
R24344 C10_N_btm.n989 C10_N_btm.n93 0.228786
R24345 C10_N_btm.n149 C10_N_btm.n99 0.228786
R24346 C10_N_btm.n100 C10_N_btm.n99 0.228786
R24347 C10_N_btm.n952 C10_N_btm.n951 0.228786
R24348 C10_N_btm.n951 C10_N_btm.n950 0.228786
R24349 C10_N_btm.n949 C10_N_btm.n148 0.228786
R24350 C10_N_btm.n953 C10_N_btm.n148 0.228786
R24351 C10_N_btm.n194 C10_N_btm.n147 0.228786
R24352 C10_N_btm.n194 C10_N_btm.n151 0.228786
R24353 C10_N_btm.n153 C10_N_btm.n152 0.228786
R24354 C10_N_btm.n152 C10_N_btm.n151 0.228786
R24355 C10_N_btm.n949 C10_N_btm.n948 0.228786
R24356 C10_N_btm.n948 C10_N_btm.n947 0.228786
R24357 C10_N_btm.n946 C10_N_btm.n150 0.228786
R24358 C10_N_btm.n950 C10_N_btm.n150 0.228786
R24359 C10_N_btm.n149 C10_N_btm.n92 0.228786
R24360 C10_N_btm.n92 C10_N_btm.n91 0.228786
R24361 C10_N_btm.n994 C10_N_btm.n993 0.228786
R24362 C10_N_btm.n993 C10_N_btm.n93 0.228786
R24363 C10_N_btm.n992 C10_N_btm.n991 0.228786
R24364 C10_N_btm.n992 C10_N_btm.n89 0.228786
R24365 C10_N_btm.n95 C10_N_btm.n94 0.228786
R24366 C10_N_btm.n96 C10_N_btm.n95 0.228786
R24367 C10_N_btm.n52 C10_N_btm.n51 0.228786
R24368 C10_N_btm.n54 C10_N_btm.n52 0.228786
R24369 C10_N_btm.n86 C10_N_btm.n55 0.228786
R24370 C10_N_btm.n55 C10_N_btm.n54 0.228786
R24371 C10_N_btm.n94 C10_N_btm.n88 0.228786
R24372 C10_N_btm.n88 C10_N_btm.n87 0.228786
R24373 C10_N_btm.n997 C10_N_btm.n996 0.228786
R24374 C10_N_btm.n996 C10_N_btm.n89 0.228786
R24375 C10_N_btm.n995 C10_N_btm.n994 0.228786
R24376 C10_N_btm.n995 C10_N_btm.n82 0.228786
R24377 C10_N_btm.n155 C10_N_btm.n90 0.228786
R24378 C10_N_btm.n91 C10_N_btm.n90 0.228786
R24379 C10_N_btm.n946 C10_N_btm.n945 0.228786
R24380 C10_N_btm.n945 C10_N_btm.n944 0.228786
R24381 C10_N_btm.n943 C10_N_btm.n154 0.228786
R24382 C10_N_btm.n947 C10_N_btm.n154 0.228786
R24383 C10_N_btm.n199 C10_N_btm.n153 0.228786
R24384 C10_N_btm.n199 C10_N_btm.n157 0.228786
R24385 C10_N_btm.n159 C10_N_btm.n158 0.228786
R24386 C10_N_btm.n158 C10_N_btm.n157 0.228786
R24387 C10_N_btm.n943 C10_N_btm.n942 0.228786
R24388 C10_N_btm.n942 C10_N_btm.n941 0.228786
R24389 C10_N_btm.n940 C10_N_btm.n156 0.228786
R24390 C10_N_btm.n944 C10_N_btm.n156 0.228786
R24391 C10_N_btm.n155 C10_N_btm.n81 0.228786
R24392 C10_N_btm.n81 C10_N_btm.n80 0.228786
R24393 C10_N_btm.n1000 C10_N_btm.n999 0.228786
R24394 C10_N_btm.n999 C10_N_btm.n82 0.228786
R24395 C10_N_btm.n998 C10_N_btm.n997 0.228786
R24396 C10_N_btm.n998 C10_N_btm.n78 0.228786
R24397 C10_N_btm.n84 C10_N_btm.n83 0.228786
R24398 C10_N_btm.n87 C10_N_btm.n84 0.228786
R24399 C10_N_btm.n86 C10_N_btm.n85 0.228786
R24400 C10_N_btm.n85 C10_N_btm.n59 0.228786
R24401 C10_N_btm.n62 C10_N_btm.n60 0.228786
R24402 C10_N_btm.n60 C10_N_btm.n59 0.228786
R24403 C10_N_btm.n83 C10_N_btm.n76 0.228786
R24404 C10_N_btm.n1004 C10_N_btm.n76 0.228786
R24405 C10_N_btm.n1003 C10_N_btm.n1002 0.228786
R24406 C10_N_btm.n1002 C10_N_btm.n78 0.228786
R24407 C10_N_btm.n1001 C10_N_btm.n1000 0.228786
R24408 C10_N_btm.n1001 C10_N_btm.n77 0.228786
R24409 C10_N_btm.n161 C10_N_btm.n79 0.228786
R24410 C10_N_btm.n80 C10_N_btm.n79 0.228786
R24411 C10_N_btm.n940 C10_N_btm.n939 0.228786
R24412 C10_N_btm.n939 C10_N_btm.n938 0.228786
R24413 C10_N_btm.n937 C10_N_btm.n160 0.228786
R24414 C10_N_btm.n941 C10_N_btm.n160 0.228786
R24415 C10_N_btm.n204 C10_N_btm.n159 0.228786
R24416 C10_N_btm.n204 C10_N_btm.n163 0.228786
R24417 C10_N_btm.n165 C10_N_btm.n164 0.228786
R24418 C10_N_btm.n164 C10_N_btm.n163 0.228786
R24419 C10_N_btm.n937 C10_N_btm.n936 0.228786
R24420 C10_N_btm.n936 C10_N_btm.n935 0.228786
R24421 C10_N_btm.n934 C10_N_btm.n162 0.228786
R24422 C10_N_btm.n938 C10_N_btm.n162 0.228786
R24423 C10_N_btm.n226 C10_N_btm.n161 0.228786
R24424 C10_N_btm.n226 C10_N_btm.n167 0.228786
R24425 C10_N_btm.n228 C10_N_btm.n227 0.228786
R24426 C10_N_btm.n227 C10_N_btm.n77 0.228786
R24427 C10_N_btm.n1003 C10_N_btm.n75 0.228786
R24428 C10_N_btm.n75 C10_N_btm.n74 0.228786
R24429 C10_N_btm.n1006 C10_N_btm.n1005 0.228786
R24430 C10_N_btm.n1005 C10_N_btm.n1004 0.228786
R24431 C10_N_btm.n63 C10_N_btm.n62 0.228786
R24432 C10_N_btm.n72 C10_N_btm.n63 0.228786
R24433 C10_N_btm.n1012 C10_N_btm.n1011 0.228786
R24434 C10_N_btm.n66 C10_N_btm.n64 0.228786
R24435 C10_N_btm.n1010 C10_N_btm.n66 0.228786
R24436 C10_N_btm.n1009 C10_N_btm.n1008 0.228786
R24437 C10_N_btm.n1008 C10_N_btm.n72 0.228786
R24438 C10_N_btm.n1007 C10_N_btm.n1006 0.228786
R24439 C10_N_btm.n1007 C10_N_btm.n70 0.228786
R24440 C10_N_btm.n911 C10_N_btm.n73 0.228786
R24441 C10_N_btm.n74 C10_N_btm.n73 0.228786
R24442 C10_N_btm.n229 C10_N_btm.n228 0.228786
R24443 C10_N_btm.n230 C10_N_btm.n229 0.228786
R24444 C10_N_btm.n169 C10_N_btm.n168 0.228786
R24445 C10_N_btm.n168 C10_N_btm.n167 0.228786
R24446 C10_N_btm.n934 C10_N_btm.n933 0.228786
R24447 C10_N_btm.n933 C10_N_btm.n932 0.228786
R24448 C10_N_btm.n931 C10_N_btm.n166 0.228786
R24449 C10_N_btm.n935 C10_N_btm.n166 0.228786
R24450 C10_N_btm.n209 C10_N_btm.n165 0.228786
R24451 C10_N_btm.n209 C10_N_btm.n171 0.228786
R24452 C10_N_btm.n173 C10_N_btm.n172 0.228786
R24453 C10_N_btm.n172 C10_N_btm.n171 0.228786
R24454 C10_N_btm.n931 C10_N_btm.n930 0.228786
R24455 C10_N_btm.n930 C10_N_btm.n929 0.228786
R24456 C10_N_btm.n928 C10_N_btm.n170 0.228786
R24457 C10_N_btm.n932 C10_N_btm.n170 0.228786
R24458 C10_N_btm.n225 C10_N_btm.n169 0.228786
R24459 C10_N_btm.n225 C10_N_btm.n175 0.228786
R24460 C10_N_btm.n914 C10_N_btm.n913 0.228786
R24461 C10_N_btm.n913 C10_N_btm.n230 0.228786
R24462 C10_N_btm.n912 C10_N_btm.n911 0.228786
R24463 C10_N_btm.n912 C10_N_btm.n224 0.228786
R24464 C10_N_btm.n910 C10_N_btm.n909 0.228786
R24465 C10_N_btm.n910 C10_N_btm.n70 0.228786
R24466 C10_N_btm.n1009 C10_N_btm.n71 0.228786
R24467 C10_N_btm.n908 C10_N_btm.n71 0.228786
R24468 C10_N_btm.n907 C10_N_btm.n69 0.228786
R24469 C10_N_btm.n1010 C10_N_btm.n69 0.228786
R24470 C10_N_btm.n892 C10_N_btm.n68 0.228786
R24471 C10_N_btm.n1011 C10_N_btm.n67 0.228786
R24472 C10_N_btm.n232 C10_N_btm.n67 0.228786
R24473 C10_N_btm.n893 C10_N_btm.n892 0.228786
R24474 C10_N_btm.n891 C10_N_btm.n243 0.228786
R24475 C10_N_btm.n881 C10_N_btm.n880 0.228786
R24476 C10_N_btm.n248 C10_N_btm.n242 0.228786
R24477 C10_N_btm.n242 C10_N_btm.n241 0.228786
R24478 C10_N_btm.n896 C10_N_btm.n895 0.228786
R24479 C10_N_btm.n895 C10_N_btm.n243 0.228786
R24480 C10_N_btm.n894 C10_N_btm.n893 0.228786
R24481 C10_N_btm.n894 C10_N_btm.n239 0.228786
R24482 C10_N_btm.n234 C10_N_btm.n233 0.228786
R24483 C10_N_btm.n233 C10_N_btm.n232 0.228786
R24484 C10_N_btm.n907 C10_N_btm.n906 0.228786
R24485 C10_N_btm.n906 C10_N_btm.n905 0.228786
R24486 C10_N_btm.n904 C10_N_btm.n231 0.228786
R24487 C10_N_btm.n908 C10_N_btm.n231 0.228786
R24488 C10_N_btm.n909 C10_N_btm.n223 0.228786
R24489 C10_N_btm.n223 C10_N_btm.n222 0.228786
R24490 C10_N_btm.n917 C10_N_btm.n916 0.228786
R24491 C10_N_btm.n916 C10_N_btm.n224 0.228786
R24492 C10_N_btm.n915 C10_N_btm.n914 0.228786
R24493 C10_N_btm.n915 C10_N_btm.n220 0.228786
R24494 C10_N_btm.n177 C10_N_btm.n176 0.228786
R24495 C10_N_btm.n176 C10_N_btm.n175 0.228786
R24496 C10_N_btm.n928 C10_N_btm.n927 0.228786
R24497 C10_N_btm.n927 C10_N_btm.n926 0.228786
R24498 C10_N_btm.n925 C10_N_btm.n174 0.228786
R24499 C10_N_btm.n929 C10_N_btm.n174 0.228786
R24500 C10_N_btm.n214 C10_N_btm.n173 0.228786
R24501 C10_N_btm.n214 C10_N_btm.n179 0.228786
R24502 C10_N_btm.n180 C10_N_btm.n179 0.228786
R24503 C10_N_btm.n925 C10_N_btm.n924 0.228786
R24504 C10_N_btm.n926 C10_N_btm.n178 0.228786
R24505 C10_N_btm.n218 C10_N_btm.n177 0.228786
R24506 C10_N_btm.n919 C10_N_btm.n220 0.228786
R24507 C10_N_btm.n918 C10_N_btm.n917 0.228786
R24508 C10_N_btm.n222 C10_N_btm.n221 0.228786
R24509 C10_N_btm.n904 C10_N_btm.n903 0.228786
R24510 C10_N_btm.n905 C10_N_btm.n235 0.228786
R24511 C10_N_btm.n237 C10_N_btm.n234 0.228786
R24512 C10_N_btm.n898 C10_N_btm.n239 0.228786
R24513 C10_N_btm.n897 C10_N_btm.n896 0.228786
R24514 C10_N_btm.n241 C10_N_btm.n240 0.228786
R24515 C10_N_btm.n880 C10_N_btm.n879 0.228786
R24516 C10_N_btm.n254 C10_N_btm.n253 0.228786
R24517 C10_N_btm.n876 C10_N_btm.n256 0.228786
R24518 C10_N_btm.n638 C10_N_btm.n637 0.228786
R24519 C10_N_btm.n639 C10_N_btm.n638 0.228786
R24520 C10_N_btm.n640 C10_N_btm.n415 0.228786
R24521 C10_N_btm.n418 C10_N_btm.n415 0.228786
R24522 C10_N_btm.n555 C10_N_btm.n414 0.228786
R24523 C10_N_btm.n641 C10_N_btm.n414 0.228786
R24524 C10_N_btm.n642 C10_N_btm.n413 0.228786
R24525 C10_N_btm.n413 C10_N_btm.n412 0.228786
R24526 C10_N_btm.n648 C10_N_btm.n647 0.228786
R24527 C10_N_btm.n647 C10_N_btm.n643 0.228786
R24528 C10_N_btm.n646 C10_N_btm.n410 0.228786
R24529 C10_N_btm.n651 C10_N_btm.n650 0.228786
R24530 C10_N_btm.n650 C10_N_btm.n410 0.228786
R24531 C10_N_btm.n649 C10_N_btm.n648 0.228786
R24532 C10_N_btm.n649 C10_N_btm.n405 0.228786
R24533 C10_N_btm.n553 C10_N_btm.n411 0.228786
R24534 C10_N_btm.n412 C10_N_btm.n411 0.228786
R24535 C10_N_btm.n556 C10_N_btm.n555 0.228786
R24536 C10_N_btm.n556 C10_N_btm.n554 0.228786
R24537 C10_N_btm.n558 C10_N_btm.n557 0.228786
R24538 C10_N_btm.n557 C10_N_btm.n418 0.228786
R24539 C10_N_btm.n637 C10_N_btm.n419 0.228786
R24540 C10_N_btm.n491 C10_N_btm.n419 0.228786
R24541 C10_N_btm.n560 C10_N_btm.n490 0.228786
R24542 C10_N_btm.n560 C10_N_btm.n491 0.228786
R24543 C10_N_btm.n559 C10_N_btm.n558 0.228786
R24544 C10_N_btm.n559 C10_N_btm.n552 0.228786
R24545 C10_N_btm.n551 C10_N_btm.n492 0.228786
R24546 C10_N_btm.n554 C10_N_btm.n492 0.228786
R24547 C10_N_btm.n553 C10_N_btm.n404 0.228786
R24548 C10_N_btm.n404 C10_N_btm.n403 0.228786
R24549 C10_N_btm.n654 C10_N_btm.n653 0.228786
R24550 C10_N_btm.n653 C10_N_btm.n405 0.228786
R24551 C10_N_btm.n652 C10_N_btm.n651 0.228786
R24552 C10_N_btm.n652 C10_N_btm.n401 0.228786
R24553 C10_N_btm.n657 C10_N_btm.n656 0.228786
R24554 C10_N_btm.n656 C10_N_btm.n401 0.228786
R24555 C10_N_btm.n655 C10_N_btm.n654 0.228786
R24556 C10_N_btm.n655 C10_N_btm.n396 0.228786
R24557 C10_N_btm.n494 C10_N_btm.n402 0.228786
R24558 C10_N_btm.n403 C10_N_btm.n402 0.228786
R24559 C10_N_btm.n551 C10_N_btm.n550 0.228786
R24560 C10_N_btm.n550 C10_N_btm.n549 0.228786
R24561 C10_N_btm.n548 C10_N_btm.n493 0.228786
R24562 C10_N_btm.n552 C10_N_btm.n493 0.228786
R24563 C10_N_btm.n490 C10_N_btm.n489 0.228786
R24564 C10_N_btm.n489 C10_N_btm.n488 0.228786
R24565 C10_N_btm.n487 C10_N_btm.n486 0.228786
R24566 C10_N_btm.n488 C10_N_btm.n487 0.228786
R24567 C10_N_btm.n548 C10_N_btm.n547 0.228786
R24568 C10_N_btm.n547 C10_N_btm.n546 0.228786
R24569 C10_N_btm.n545 C10_N_btm.n495 0.228786
R24570 C10_N_btm.n549 C10_N_btm.n495 0.228786
R24571 C10_N_btm.n494 C10_N_btm.n395 0.228786
R24572 C10_N_btm.n395 C10_N_btm.n394 0.228786
R24573 C10_N_btm.n660 C10_N_btm.n659 0.228786
R24574 C10_N_btm.n659 C10_N_btm.n396 0.228786
R24575 C10_N_btm.n658 C10_N_btm.n657 0.228786
R24576 C10_N_btm.n658 C10_N_btm.n392 0.228786
R24577 C10_N_btm.n663 C10_N_btm.n662 0.228786
R24578 C10_N_btm.n662 C10_N_btm.n392 0.228786
R24579 C10_N_btm.n661 C10_N_btm.n660 0.228786
R24580 C10_N_btm.n661 C10_N_btm.n387 0.228786
R24581 C10_N_btm.n497 C10_N_btm.n393 0.228786
R24582 C10_N_btm.n394 C10_N_btm.n393 0.228786
R24583 C10_N_btm.n545 C10_N_btm.n544 0.228786
R24584 C10_N_btm.n544 C10_N_btm.n543 0.228786
R24585 C10_N_btm.n542 C10_N_btm.n496 0.228786
R24586 C10_N_btm.n546 C10_N_btm.n496 0.228786
R24587 C10_N_btm.n486 C10_N_btm.n485 0.228786
R24588 C10_N_btm.n485 C10_N_btm.n484 0.228786
R24589 C10_N_btm.n483 C10_N_btm.n482 0.228786
R24590 C10_N_btm.n484 C10_N_btm.n483 0.228786
R24591 C10_N_btm.n542 C10_N_btm.n541 0.228786
R24592 C10_N_btm.n541 C10_N_btm.n540 0.228786
R24593 C10_N_btm.n539 C10_N_btm.n498 0.228786
R24594 C10_N_btm.n543 C10_N_btm.n498 0.228786
R24595 C10_N_btm.n497 C10_N_btm.n386 0.228786
R24596 C10_N_btm.n386 C10_N_btm.n385 0.228786
R24597 C10_N_btm.n666 C10_N_btm.n665 0.228786
R24598 C10_N_btm.n665 C10_N_btm.n387 0.228786
R24599 C10_N_btm.n664 C10_N_btm.n663 0.228786
R24600 C10_N_btm.n664 C10_N_btm.n383 0.228786
R24601 C10_N_btm.n669 C10_N_btm.n668 0.228786
R24602 C10_N_btm.n668 C10_N_btm.n383 0.228786
R24603 C10_N_btm.n667 C10_N_btm.n666 0.228786
R24604 C10_N_btm.n667 C10_N_btm.n381 0.228786
R24605 C10_N_btm.n500 C10_N_btm.n384 0.228786
R24606 C10_N_btm.n385 C10_N_btm.n384 0.228786
R24607 C10_N_btm.n539 C10_N_btm.n538 0.228786
R24608 C10_N_btm.n538 C10_N_btm.n537 0.228786
R24609 C10_N_btm.n536 C10_N_btm.n499 0.228786
R24610 C10_N_btm.n540 C10_N_btm.n499 0.228786
R24611 C10_N_btm.n482 C10_N_btm.n481 0.228786
R24612 C10_N_btm.n481 C10_N_btm.n480 0.228786
R24613 C10_N_btm.n479 C10_N_btm.n478 0.228786
R24614 C10_N_btm.n480 C10_N_btm.n479 0.228786
R24615 C10_N_btm.n536 C10_N_btm.n535 0.228786
R24616 C10_N_btm.n535 C10_N_btm.n534 0.228786
R24617 C10_N_btm.n533 C10_N_btm.n501 0.228786
R24618 C10_N_btm.n537 C10_N_btm.n501 0.228786
R24619 C10_N_btm.n503 C10_N_btm.n500 0.228786
R24620 C10_N_btm.n504 C10_N_btm.n503 0.228786
R24621 C10_N_btm.n506 C10_N_btm.n380 0.228786
R24622 C10_N_btm.n381 C10_N_btm.n380 0.228786
R24623 C10_N_btm.n670 C10_N_btm.n669 0.228786
R24624 C10_N_btm.n670 C10_N_btm.n378 0.228786
R24625 C10_N_btm.n676 C10_N_btm.n376 0.228786
R24626 C10_N_btm.n377 C10_N_btm.n376 0.228786
R24627 C10_N_btm.n378 C10_N_btm.n377 0.228786
R24628 C10_N_btm.n507 C10_N_btm.n506 0.228786
R24629 C10_N_btm.n508 C10_N_btm.n507 0.228786
R24630 C10_N_btm.n509 C10_N_btm.n505 0.228786
R24631 C10_N_btm.n505 C10_N_btm.n504 0.228786
R24632 C10_N_btm.n533 C10_N_btm.n532 0.228786
R24633 C10_N_btm.n532 C10_N_btm.n531 0.228786
R24634 C10_N_btm.n530 C10_N_btm.n502 0.228786
R24635 C10_N_btm.n534 C10_N_btm.n502 0.228786
R24636 C10_N_btm.n478 C10_N_btm.n477 0.228786
R24637 C10_N_btm.n477 C10_N_btm.n476 0.228786
R24638 C10_N_btm.n476 C10_N_btm.n475 0.228786
R24639 C10_N_btm.n475 C10_N_btm.n474 0.228786
R24640 C10_N_btm.n529 C10_N_btm.n528 0.228786
R24641 C10_N_btm.n530 C10_N_btm.n529 0.228786
R24642 C10_N_btm.n531 C10_N_btm.n511 0.228786
R24643 C10_N_btm.n512 C10_N_btm.n511 0.228786
R24644 C10_N_btm.n510 C10_N_btm.n365 0.228786
R24645 C10_N_btm.n510 C10_N_btm.n509 0.228786
R24646 C10_N_btm.n508 C10_N_btm.n366 0.228786
R24647 C10_N_btm.n679 C10_N_btm.n678 0.228786
R24648 C10_N_btm.n678 C10_N_btm.n366 0.228786
R24649 C10_N_btm.n677 C10_N_btm.n676 0.228786
R24650 C10_N_btm.n677 C10_N_btm.n364 0.228786
R24651 C10_N_btm.n884 C10_N_btm.n883 0.228786
R24652 C10_N_btm.n888 C10_N_btm.n245 0.228786
R24653 C10_N_btm.n887 C10_N_btm.n886 0.228786
R24654 C10_N_btm.n886 C10_N_btm.n885 0.228786
R24655 C10_N_btm.n252 C10_N_btm.n251 0.228786
R24656 C10_N_btm.n251 C10_N_btm.n250 0.228786
R24657 C10_N_btm.n268 C10_N_btm.n250 0.228786
R24658 C10_N_btm.n884 C10_N_btm.n247 0.228786
R24659 C10_N_btm.n247 C10_N_btm.n246 0.228786
R24660 C10_N_btm.n269 C10_N_btm.n268 0.228786
R24661 C10_N_btm.n267 C10_N_btm.n265 0.228786
R24662 C10_N_btm.n270 C10_N_btm.n267 0.228786
R24663 C10_N_btm.n868 C10_N_btm.n867 0.228786
R24664 C10_N_btm.n866 C10_N_btm.n266 0.228786
R24665 C10_N_btm.n865 C10_N_btm.n271 0.228786
R24666 C10_N_btm.n864 C10_N_btm.n863 0.228786
R24667 C10_N_btm.n306 C10_N_btm.n305 0.228786
R24668 C10_N_btm.n327 C10_N_btm.n326 0.228786
R24669 C10_N_btm.n333 C10_N_btm.n332 0.228786
R24670 C10_N_btm.n334 C10_N_btm.n325 0.228786
R24671 C10_N_btm.n727 C10_N_btm.n335 0.228786
R24672 C10_N_btm.n726 C10_N_btm.n725 0.228786
R24673 C10_N_btm.n724 C10_N_btm.n336 0.228786
R24674 C10_N_btm.n723 C10_N_btm.n337 0.228786
R24675 C10_N_btm.n722 C10_N_btm.n721 0.228786
R24676 C10_N_btm.n720 C10_N_btm.n338 0.228786
R24677 C10_N_btm.n367 C10_N_btm.n340 0.228786
R24678 C10_N_btm.n373 C10_N_btm.n372 0.228786
R24679 C10_N_btm.n374 C10_N_btm.n373 0.228786
R24680 C10_N_btm.n364 C10_N_btm.n362 0.228786
R24681 C10_N_btm.n362 C10_N_btm.n361 0.228786
R24682 C10_N_btm.n682 C10_N_btm.n360 0.228786
R24683 C10_N_btm.n681 C10_N_btm.n680 0.228786
R24684 C10_N_btm.n680 C10_N_btm.n679 0.228786
R24685 C10_N_btm.n363 C10_N_btm.n360 0.228786
R24686 C10_N_btm.n365 C10_N_btm.n363 0.228786
R24687 C10_N_btm.n513 C10_N_btm.n512 0.228786
R24688 C10_N_btm.n514 C10_N_btm.n513 0.228786
R24689 C10_N_btm.n527 C10_N_btm.n526 0.228786
R24690 C10_N_btm.n528 C10_N_btm.n527 0.228786
R24691 C10_N_btm.n474 C10_N_btm.n473 0.228786
R24692 C10_N_btm.n473 C10_N_btm.n472 0.228786
R24693 C10_N_btm.n472 C10_N_btm.n471 0.228786
R24694 C10_N_btm.n471 C10_N_btm.n470 0.228786
R24695 C10_N_btm.n525 C10_N_btm.n524 0.228786
R24696 C10_N_btm.n526 C10_N_btm.n525 0.228786
R24697 C10_N_btm.n514 C10_N_btm.n359 0.228786
R24698 C10_N_btm.n357 C10_N_btm.n356 0.228786
R24699 C10_N_btm.n359 C10_N_btm.n357 0.228786
R24700 C10_N_btm.n683 C10_N_btm.n682 0.228786
R24701 C10_N_btm.n684 C10_N_btm.n683 0.228786
R24702 C10_N_btm.n358 C10_N_btm.n354 0.228786
R24703 C10_N_btm.n681 C10_N_btm.n358 0.228786
R24704 C10_N_btm.n368 C10_N_btm.n361 0.228786
R24705 C10_N_btm.n369 C10_N_btm.n368 0.228786
R24706 C10_N_btm.n371 C10_N_btm.n370 0.228786
R24707 C10_N_btm.n372 C10_N_btm.n371 0.228786
R24708 C10_N_btm.n341 C10_N_btm.n340 0.228786
R24709 C10_N_btm.n342 C10_N_btm.n341 0.228786
R24710 C10_N_btm.n719 C10_N_btm.n718 0.228786
R24711 C10_N_btm.n720 C10_N_btm.n719 0.228786
R24712 C10_N_btm.n721 C10_N_btm.n339 0.228786
R24713 C10_N_btm.n343 C10_N_btm.n339 0.228786
R24714 C10_N_btm.n704 C10_N_btm.n703 0.228786
R24715 C10_N_btm.n703 C10_N_btm.n337 0.228786
R24716 C10_N_btm.n702 C10_N_btm.n336 0.228786
R24717 C10_N_btm.n702 C10_N_btm.n701 0.228786
R24718 C10_N_btm.n323 C10_N_btm.n322 0.228786
R24719 C10_N_btm.n726 C10_N_btm.n323 0.228786
R24720 C10_N_btm.n728 C10_N_btm.n727 0.228786
R24721 C10_N_btm.n729 C10_N_btm.n728 0.228786
R24722 C10_N_btm.n324 C10_N_btm.n320 0.228786
R24723 C10_N_btm.n325 C10_N_btm.n324 0.228786
R24724 C10_N_btm.n332 C10_N_btm.n331 0.228786
R24725 C10_N_btm.n331 C10_N_btm.n330 0.228786
R24726 C10_N_btm.n329 C10_N_btm.n328 0.228786
R24727 C10_N_btm.n328 C10_N_btm.n327 0.228786
R24728 C10_N_btm.n307 C10_N_btm.n306 0.228786
R24729 C10_N_btm.n308 C10_N_btm.n307 0.228786
R24730 C10_N_btm.n822 C10_N_btm.n821 0.228786
R24731 C10_N_btm.n823 C10_N_btm.n822 0.228786
R24732 C10_N_btm.n825 C10_N_btm.n304 0.228786
R24733 C10_N_btm.n309 C10_N_btm.n304 0.228786
R24734 C10_N_btm.n807 C10_N_btm.n303 0.228786
R24735 C10_N_btm.n826 C10_N_btm.n303 0.228786
R24736 C10_N_btm.n827 C10_N_btm.n302 0.228786
R24737 C10_N_btm.n806 C10_N_btm.n302 0.228786
R24738 C10_N_btm.n805 C10_N_btm.n301 0.228786
R24739 C10_N_btm.n828 C10_N_btm.n301 0.228786
R24740 C10_N_btm.n829 C10_N_btm.n300 0.228786
R24741 C10_N_btm.n740 C10_N_btm.n300 0.228786
R24742 C10_N_btm.n755 C10_N_btm.n299 0.228786
R24743 C10_N_btm.n830 C10_N_btm.n299 0.228786
R24744 C10_N_btm.n831 C10_N_btm.n298 0.228786
R24745 C10_N_btm.n760 C10_N_btm.n298 0.228786
R24746 C10_N_btm.n761 C10_N_btm.n297 0.228786
R24747 C10_N_btm.n832 C10_N_btm.n297 0.228786
R24748 C10_N_btm.n833 C10_N_btm.n296 0.228786
R24749 C10_N_btm.n792 C10_N_btm.n296 0.228786
R24750 C10_N_btm.n791 C10_N_btm.n295 0.228786
R24751 C10_N_btm.n834 C10_N_btm.n295 0.228786
R24752 C10_N_btm.n835 C10_N_btm.n294 0.228786
R24753 C10_N_btm.n790 C10_N_btm.n294 0.228786
R24754 C10_N_btm.n789 C10_N_btm.n293 0.228786
R24755 C10_N_btm.n836 C10_N_btm.n293 0.228786
R24756 C10_N_btm.n837 C10_N_btm.n292 0.228786
R24757 C10_N_btm.n763 C10_N_btm.n292 0.228786
R24758 C10_N_btm.n775 C10_N_btm.n291 0.228786
R24759 C10_N_btm.n838 C10_N_btm.n291 0.228786
R24760 C10_N_btm.n839 C10_N_btm.n290 0.228786
R24761 C10_N_btm.n774 C10_N_btm.n290 0.228786
R24762 C10_N_btm.n288 C10_N_btm.n287 0.228786
R24763 C10_N_btm.n840 C10_N_btm.n288 0.228786
R24764 C10_N_btm.n842 C10_N_btm.n841 0.228786
R24765 C10_N_btm.n843 C10_N_btm.n842 0.228786
R24766 C10_N_btm.n275 C10_N_btm.n274 0.228786
R24767 C10_N_btm.n289 C10_N_btm.n274 0.228786
R24768 C10_N_btm.n862 C10_N_btm.n861 0.228786
R24769 C10_N_btm.n861 C10_N_btm.n860 0.228786
R24770 C10_N_btm.n859 C10_N_btm.n273 0.228786
R24771 C10_N_btm.n863 C10_N_btm.n273 0.228786
R24772 C10_N_btm.n277 C10_N_btm.n271 0.228786
R24773 C10_N_btm.n278 C10_N_btm.n277 0.228786
R24774 C10_N_btm.n264 C10_N_btm.n263 0.228786
R24775 C10_N_btm.n266 C10_N_btm.n264 0.228786
R24776 C10_N_btm.n869 C10_N_btm.n868 0.228786
R24777 C10_N_btm.n870 C10_N_btm.n869 0.228786
R24778 C10_N_btm.n265 C10_N_btm.n261 0.228786
R24779 C10_N_btm.n873 C10_N_btm.n872 0.228786
R24780 C10_N_btm.n872 C10_N_btm.n261 0.228786
R24781 C10_N_btm.n871 C10_N_btm.n870 0.228786
R24782 C10_N_btm.n871 C10_N_btm.n259 0.228786
R24783 C10_N_btm.n851 C10_N_btm.n262 0.228786
R24784 C10_N_btm.n263 C10_N_btm.n262 0.228786
R24785 C10_N_btm.n279 C10_N_btm.n278 0.228786
R24786 C10_N_btm.n281 C10_N_btm.n279 0.228786
R24787 C10_N_btm.n858 C10_N_btm.n857 0.228786
R24788 C10_N_btm.n859 C10_N_btm.n858 0.228786
R24789 C10_N_btm.n860 C10_N_btm.n276 0.228786
R24790 C10_N_btm.n280 C10_N_btm.n276 0.228786
R24791 C10_N_btm.n846 C10_N_btm.n845 0.228786
R24792 C10_N_btm.n845 C10_N_btm.n275 0.228786
R24793 C10_N_btm.n844 C10_N_btm.n843 0.228786
R24794 C10_N_btm.n844 C10_N_btm.n285 0.228786
R24795 C10_N_btm.n779 C10_N_btm.n286 0.228786
R24796 C10_N_btm.n287 C10_N_btm.n286 0.228786
R24797 C10_N_btm.n774 C10_N_btm.n773 0.228786
R24798 C10_N_btm.n778 C10_N_btm.n773 0.228786
R24799 C10_N_btm.n777 C10_N_btm.n776 0.228786
R24800 C10_N_btm.n776 C10_N_btm.n775 0.228786
R24801 C10_N_btm.n764 C10_N_btm.n763 0.228786
R24802 C10_N_btm.n766 C10_N_btm.n764 0.228786
R24803 C10_N_btm.n788 C10_N_btm.n787 0.228786
R24804 C10_N_btm.n789 C10_N_btm.n788 0.228786
R24805 C10_N_btm.n790 C10_N_btm.n762 0.228786
R24806 C10_N_btm.n765 C10_N_btm.n762 0.228786
R24807 C10_N_btm.n754 C10_N_btm.n752 0.228786
R24808 C10_N_btm.n791 C10_N_btm.n754 0.228786
R24809 C10_N_btm.n793 C10_N_btm.n792 0.228786
R24810 C10_N_btm.n794 C10_N_btm.n793 0.228786
R24811 C10_N_btm.n753 C10_N_btm.n750 0.228786
R24812 C10_N_btm.n761 C10_N_btm.n753 0.228786
R24813 C10_N_btm.n760 C10_N_btm.n759 0.228786
R24814 C10_N_btm.n759 C10_N_btm.n758 0.228786
R24815 C10_N_btm.n757 C10_N_btm.n756 0.228786
R24816 C10_N_btm.n756 C10_N_btm.n755 0.228786
R24817 C10_N_btm.n741 C10_N_btm.n740 0.228786
R24818 C10_N_btm.n742 C10_N_btm.n741 0.228786
R24819 C10_N_btm.n804 C10_N_btm.n803 0.228786
R24820 C10_N_btm.n805 C10_N_btm.n804 0.228786
R24821 C10_N_btm.n806 C10_N_btm.n739 0.228786
R24822 C10_N_btm.n739 C10_N_btm.n738 0.228786
R24823 C10_N_btm.n809 C10_N_btm.n808 0.228786
R24824 C10_N_btm.n808 C10_N_btm.n807 0.228786
R24825 C10_N_btm.n310 C10_N_btm.n309 0.228786
R24826 C10_N_btm.n810 C10_N_btm.n310 0.228786
R24827 C10_N_btm.n820 C10_N_btm.n311 0.228786
R24828 C10_N_btm.n821 C10_N_btm.n820 0.228786
R24829 C10_N_btm.n819 C10_N_btm.n308 0.228786
R24830 C10_N_btm.n819 C10_N_btm.n818 0.228786
R24831 C10_N_btm.n817 C10_N_btm.n312 0.228786
R24832 C10_N_btm.n329 C10_N_btm.n312 0.228786
R24833 C10_N_btm.n330 C10_N_btm.n319 0.228786
R24834 C10_N_btm.n319 C10_N_btm.n314 0.228786
R24835 C10_N_btm.n732 C10_N_btm.n731 0.228786
R24836 C10_N_btm.n731 C10_N_btm.n320 0.228786
R24837 C10_N_btm.n730 C10_N_btm.n729 0.228786
R24838 C10_N_btm.n730 C10_N_btm.n318 0.228786
R24839 C10_N_btm.n693 C10_N_btm.n321 0.228786
R24840 C10_N_btm.n322 C10_N_btm.n321 0.228786
R24841 C10_N_btm.n701 C10_N_btm.n700 0.228786
R24842 C10_N_btm.n700 C10_N_btm.n699 0.228786
R24843 C10_N_btm.n706 C10_N_btm.n705 0.228786
R24844 C10_N_btm.n705 C10_N_btm.n704 0.228786
R24845 C10_N_btm.n344 C10_N_btm.n343 0.228786
R24846 C10_N_btm.n707 C10_N_btm.n344 0.228786
R24847 C10_N_btm.n717 C10_N_btm.n345 0.228786
R24848 C10_N_btm.n718 C10_N_btm.n717 0.228786
R24849 C10_N_btm.n716 C10_N_btm.n342 0.228786
R24850 C10_N_btm.n716 C10_N_btm.n715 0.228786
R24851 C10_N_btm.n714 C10_N_btm.n346 0.228786
R24852 C10_N_btm.n370 C10_N_btm.n346 0.228786
R24853 C10_N_btm.n369 C10_N_btm.n353 0.228786
R24854 C10_N_btm.n353 C10_N_btm.n348 0.228786
R24855 C10_N_btm.n687 C10_N_btm.n686 0.228786
R24856 C10_N_btm.n686 C10_N_btm.n354 0.228786
R24857 C10_N_btm.n685 C10_N_btm.n684 0.228786
R24858 C10_N_btm.n685 C10_N_btm.n352 0.228786
R24859 C10_N_btm.n522 C10_N_btm.n521 0.228786
R24860 C10_N_btm.n520 C10_N_btm.n355 0.228786
R24861 C10_N_btm.n356 C10_N_btm.n355 0.228786
R24862 C10_N_btm.n523 C10_N_btm.n522 0.228786
R24863 C10_N_btm.n524 C10_N_btm.n523 0.228786
R24864 C10_N_btm.n470 C10_N_btm.n469 0.228786
R24865 C10_N_btm.n469 C10_N_btm.n468 0.228786
R24866 C10_N_btm.n468 C10_N_btm.n467 0.228786
R24867 C10_N_btm.n593 C10_N_btm.n592 0.228786
R24868 C10_N_btm.n463 C10_N_btm.n462 0.228786
R24869 C10_N_btm.n462 C10_N_btm.n460 0.228786
R24870 C10_N_btm.n592 C10_N_btm.n591 0.228786
R24871 C10_N_btm.n591 C10_N_btm.n590 0.228786
R24872 C10_N_btm.n460 C10_N_btm.n459 0.228786
R24873 C10_N_btm.n588 C10_N_btm.n459 0.228786
R24874 C10_N_btm.n590 C10_N_btm.n589 0.228786
R24875 C10_N_btm.n589 C10_N_btm.n586 0.228786
R24876 C10_N_btm.n588 C10_N_btm.n587 0.228786
R24877 C10_N_btm.n587 C10_N_btm.n455 0.228786
R24878 C10_N_btm.n586 C10_N_btm.n585 0.228786
R24879 C10_N_btm.n585 C10_N_btm.n584 0.228786
R24880 C10_N_btm.n455 C10_N_btm.n454 0.228786
R24881 C10_N_btm.n454 C10_N_btm.n452 0.228786
R24882 C10_N_btm.n584 C10_N_btm.n583 0.228786
R24883 C10_N_btm.n583 C10_N_btm.n582 0.228786
R24884 C10_N_btm.n452 C10_N_btm.n451 0.228786
R24885 C10_N_btm.n580 C10_N_btm.n451 0.228786
R24886 C10_N_btm.n582 C10_N_btm.n581 0.228786
R24887 C10_N_btm.n581 C10_N_btm.n578 0.228786
R24888 C10_N_btm.n580 C10_N_btm.n579 0.228786
R24889 C10_N_btm.n579 C10_N_btm.n447 0.228786
R24890 C10_N_btm.n578 C10_N_btm.n577 0.228786
R24891 C10_N_btm.n577 C10_N_btm.n576 0.228786
R24892 C10_N_btm.n447 C10_N_btm.n446 0.228786
R24893 C10_N_btm.n446 C10_N_btm.n444 0.228786
R24894 C10_N_btm.n576 C10_N_btm.n575 0.228786
R24895 C10_N_btm.n575 C10_N_btm.n574 0.228786
R24896 C10_N_btm.n444 C10_N_btm.n443 0.228786
R24897 C10_N_btm.n572 C10_N_btm.n443 0.228786
R24898 C10_N_btm.n574 C10_N_btm.n573 0.228786
R24899 C10_N_btm.n573 C10_N_btm.n570 0.228786
R24900 C10_N_btm.n572 C10_N_btm.n571 0.228786
R24901 C10_N_btm.n571 C10_N_btm.n439 0.228786
R24902 C10_N_btm.n570 C10_N_btm.n569 0.228786
R24903 C10_N_btm.n569 C10_N_btm.n568 0.228786
R24904 C10_N_btm.n439 C10_N_btm.n438 0.228786
R24905 C10_N_btm.n438 C10_N_btm.n436 0.228786
R24906 C10_N_btm.n568 C10_N_btm.n567 0.228786
R24907 C10_N_btm.n567 C10_N_btm.n566 0.228786
R24908 C10_N_btm.n436 C10_N_btm.n435 0.228786
R24909 C10_N_btm.n564 C10_N_btm.n435 0.228786
R24910 C10_N_btm.n566 C10_N_btm.n565 0.228786
R24911 C10_N_btm.n565 C10_N_btm.n562 0.228786
R24912 C10_N_btm.n564 C10_N_btm.n563 0.228786
R24913 C10_N_btm.n563 C10_N_btm.n423 0.228786
R24914 C10_N_btm.n562 C10_N_btm.n561 0.228786
R24915 C10_N_btm.n561 C10_N_btm.n421 0.228786
R24916 C10_N_btm.n633 C10_N_btm.n423 0.228786
R24917 C10_N_btm.n634 C10_N_btm.n633 0.228786
R24918 C10_N_btm.n635 C10_N_btm.n421 0.228786
R24919 C10_N_btm.n636 C10_N_btm.n635 0.228786
R24920 C10_N_btm.n634 C10_N_btm.n420 0.228786
R24921 C10_N_btm.n426 C10_N_btm.n420 0.228786
R24922 C10_N_btm.n636 C10_N_btm.n417 0.228786
R24923 C10_N_btm.n417 C10_N_btm.n416 0.228786
R24924 C10_N_btm.n426 C10_N_btm.n425 0.228786
R24925 C10_N_btm.n428 C10_N_btm.n427 0.228786
R24926 C10_N_btm.n428 C10_N_btm.n422 0.228786
R24927 C10_N_btm.n430 C10_N_btm.n429 0.228786
R24928 C10_N_btm.n431 C10_N_btm.n430 0.228786
R24929 C10_N_btm.n632 C10_N_btm.n422 0.228786
R24930 C10_N_btm.n632 C10_N_btm.n631 0.228786
R24931 C10_N_btm.n630 C10_N_btm.n431 0.228786
R24932 C10_N_btm.n630 C10_N_btm.n629 0.228786
R24933 C10_N_btm.n631 C10_N_btm.n432 0.228786
R24934 C10_N_btm.n433 C10_N_btm.n432 0.228786
R24935 C10_N_btm.n629 C10_N_btm.n628 0.228786
R24936 C10_N_btm.n628 C10_N_btm.n627 0.228786
R24937 C10_N_btm.n626 C10_N_btm.n433 0.228786
R24938 C10_N_btm.n626 C10_N_btm.n625 0.228786
R24939 C10_N_btm.n627 C10_N_btm.n434 0.228786
R24940 C10_N_btm.n437 C10_N_btm.n434 0.228786
R24941 C10_N_btm.n625 C10_N_btm.n624 0.228786
R24942 C10_N_btm.n624 C10_N_btm.n623 0.228786
R24943 C10_N_btm.n622 C10_N_btm.n437 0.228786
R24944 C10_N_btm.n622 C10_N_btm.n621 0.228786
R24945 C10_N_btm.n623 C10_N_btm.n440 0.228786
R24946 C10_N_btm.n441 C10_N_btm.n440 0.228786
R24947 C10_N_btm.n621 C10_N_btm.n620 0.228786
R24948 C10_N_btm.n620 C10_N_btm.n619 0.228786
R24949 C10_N_btm.n618 C10_N_btm.n441 0.228786
R24950 C10_N_btm.n618 C10_N_btm.n617 0.228786
R24951 C10_N_btm.n619 C10_N_btm.n442 0.228786
R24952 C10_N_btm.n445 C10_N_btm.n442 0.228786
R24953 C10_N_btm.n617 C10_N_btm.n616 0.228786
R24954 C10_N_btm.n616 C10_N_btm.n615 0.228786
R24955 C10_N_btm.n614 C10_N_btm.n445 0.228786
R24956 C10_N_btm.n614 C10_N_btm.n613 0.228786
R24957 C10_N_btm.n615 C10_N_btm.n448 0.228786
R24958 C10_N_btm.n449 C10_N_btm.n448 0.228786
R24959 C10_N_btm.n613 C10_N_btm.n612 0.228786
R24960 C10_N_btm.n612 C10_N_btm.n611 0.228786
R24961 C10_N_btm.n610 C10_N_btm.n449 0.228786
R24962 C10_N_btm.n610 C10_N_btm.n609 0.228786
R24963 C10_N_btm.n611 C10_N_btm.n450 0.228786
R24964 C10_N_btm.n453 C10_N_btm.n450 0.228786
R24965 C10_N_btm.n609 C10_N_btm.n608 0.228786
R24966 C10_N_btm.n608 C10_N_btm.n607 0.228786
R24967 C10_N_btm.n606 C10_N_btm.n453 0.228786
R24968 C10_N_btm.n606 C10_N_btm.n605 0.228786
R24969 C10_N_btm.n607 C10_N_btm.n456 0.228786
R24970 C10_N_btm.n457 C10_N_btm.n456 0.228786
R24971 C10_N_btm.n605 C10_N_btm.n604 0.228786
R24972 C10_N_btm.n604 C10_N_btm.n603 0.228786
R24973 C10_N_btm.n602 C10_N_btm.n457 0.228786
R24974 C10_N_btm.n602 C10_N_btm.n601 0.228786
R24975 C10_N_btm.n603 C10_N_btm.n458 0.228786
R24976 C10_N_btm.n461 C10_N_btm.n458 0.228786
R24977 C10_N_btm.n601 C10_N_btm.n600 0.228786
R24978 C10_N_btm.n600 C10_N_btm.n599 0.228786
R24979 C10_N_btm.n598 C10_N_btm.n461 0.228786
R24980 C10_N_btm.n599 C10_N_btm.n464 0.228786
R24981 C10_N_btm.n595 C10_N_btm.n463 0.228786
R24982 C10_N_btm.n594 C10_N_btm.n593 0.228786
R24983 C10_N_btm.n467 C10_N_btm.n466 0.228786
R24984 C10_N_btm.n521 C10_N_btm.n515 0.228786
R24985 C10_N_btm.n520 C10_N_btm.n519 0.228786
R24986 C10_N_btm.n352 C10_N_btm.n351 0.228786
R24987 C10_N_btm.n688 C10_N_btm.n687 0.228786
R24988 C10_N_btm.n349 C10_N_btm.n348 0.228786
R24989 C10_N_btm.n714 C10_N_btm.n713 0.228786
R24990 C10_N_btm.n715 C10_N_btm.n347 0.228786
R24991 C10_N_btm.n709 C10_N_btm.n345 0.228786
R24992 C10_N_btm.n708 C10_N_btm.n707 0.228786
R24993 C10_N_btm.n706 C10_N_btm.n692 0.228786
R24994 C10_N_btm.n699 C10_N_btm.n698 0.228786
R24995 C10_N_btm.n694 C10_N_btm.n693 0.228786
R24996 C10_N_btm.n318 C10_N_btm.n317 0.228786
R24997 C10_N_btm.n733 C10_N_btm.n732 0.228786
R24998 C10_N_btm.n315 C10_N_btm.n314 0.228786
R24999 C10_N_btm.n817 C10_N_btm.n816 0.228786
R25000 C10_N_btm.n818 C10_N_btm.n313 0.228786
R25001 C10_N_btm.n812 C10_N_btm.n311 0.228786
R25002 C10_N_btm.n811 C10_N_btm.n810 0.228786
R25003 C10_N_btm.n809 C10_N_btm.n737 0.228786
R25004 C10_N_btm.n743 C10_N_btm.n738 0.228786
R25005 C10_N_btm.n803 C10_N_btm.n802 0.228786
R25006 C10_N_btm.n801 C10_N_btm.n742 0.228786
R25007 C10_N_btm.n757 C10_N_btm.n747 0.228786
R25008 C10_N_btm.n758 C10_N_btm.n748 0.228786
R25009 C10_N_btm.n796 C10_N_btm.n750 0.228786
R25010 C10_N_btm.n795 C10_N_btm.n794 0.228786
R25011 C10_N_btm.n752 C10_N_btm.n751 0.228786
R25012 C10_N_btm.n767 C10_N_btm.n765 0.228786
R25013 C10_N_btm.n787 C10_N_btm.n786 0.228786
R25014 C10_N_btm.n785 C10_N_btm.n766 0.228786
R25015 C10_N_btm.n777 C10_N_btm.n771 0.228786
R25016 C10_N_btm.n778 C10_N_btm.n772 0.228786
R25017 C10_N_btm.n780 C10_N_btm.n779 0.228786
R25018 C10_N_btm.n285 C10_N_btm.n284 0.228786
R25019 C10_N_btm.n847 C10_N_btm.n846 0.228786
R25020 C10_N_btm.n282 C10_N_btm.n280 0.228786
R25021 C10_N_btm.n857 C10_N_btm.n856 0.228786
R25022 C10_N_btm.n855 C10_N_btm.n281 0.228786
R25023 C10_N_btm.n852 C10_N_btm.n851 0.228786
R25024 C10_N_btm.n259 C10_N_btm.n258 0.228786
R25025 C10_N_btm.n874 C10_N_btm.n873 0.228786
R25026 C10_N_btm.n260 C10_N_btm.n256 0.228786
R25027 C10_N_btm.n260 C10_N_btm.n252 0.228786
R25028 C10_N_btm.n882 C10_N_btm.n253 0.228786
R25029 C10_N_btm.n883 C10_N_btm.n882 0.228786
R25030 C10_N_btm.n881 C10_N_btm.n249 0.228786
R25031 C10_N_btm.n885 C10_N_btm.n249 0.228786
R25032 C10_N_btm.n248 C10_N_btm.n244 0.228786
R25033 C10_N_btm.n245 C10_N_btm.n244 0.228786
R25034 C10_N_btm.n891 C10_N_btm.n890 0.228786
R25035 C10_N_btm.n890 C10_N_btm.n889 0.228786
R25036 C10_N_btm.n68 C10_N_btm.n65 0.228786
R25037 C10_N_btm.n1013 C10_N_btm.n1012 0.228786
R25038 C10_N_btm.n1014 C10_N_btm.n1013 0.228786
R25039 C10_N_btm.n1015 C10_N_btm.n64 0.228786
R25040 C10_N_btm.n1016 C10_N_btm.n1015 0.228786
R25041 C10_N_btm.n1014 C10_N_btm.n61 0.228786
R25042 C10_N_btm.n61 C10_N_btm.n58 0.228786
R25043 C10_N_btm.n1017 C10_N_btm.n1016 0.228786
R25044 C10_N_btm.n1018 C10_N_btm.n1017 0.228786
R25045 C10_N_btm.n1019 C10_N_btm.n58 0.228786
R25046 C10_N_btm.n1020 C10_N_btm.n1019 0.228786
R25047 C10_N_btm.n1018 C10_N_btm.n57 0.228786
R25048 C10_N_btm.n57 C10_N_btm.n56 0.228786
R25049 C10_N_btm.n1021 C10_N_btm.n1020 0.228786
R25050 C10_N_btm.n1022 C10_N_btm.n1021 0.228786
R25051 C10_N_btm.n1023 C10_N_btm.n56 0.228786
R25052 C10_N_btm.n1024 C10_N_btm.n1023 0.228786
R25053 C10_N_btm.n1022 C10_N_btm.n53 0.228786
R25054 C10_N_btm.n53 C10_N_btm.n50 0.228786
R25055 C10_N_btm.n1025 C10_N_btm.n1024 0.228786
R25056 C10_N_btm.n1026 C10_N_btm.n1025 0.228786
R25057 C10_N_btm.n1027 C10_N_btm.n50 0.228786
R25058 C10_N_btm.n1028 C10_N_btm.n1027 0.228786
R25059 C10_N_btm.n1026 C10_N_btm.n49 0.228786
R25060 C10_N_btm.n49 C10_N_btm.n48 0.228786
R25061 C10_N_btm.n1029 C10_N_btm.n1028 0.228786
R25062 C10_N_btm.n1030 C10_N_btm.n1029 0.228786
R25063 C10_N_btm.n1031 C10_N_btm.n48 0.228786
R25064 C10_N_btm.n1032 C10_N_btm.n1031 0.228786
R25065 C10_N_btm.n1030 C10_N_btm.n45 0.228786
R25066 C10_N_btm.n45 C10_N_btm.n42 0.228786
R25067 C10_N_btm.n1033 C10_N_btm.n1032 0.228786
R25068 C10_N_btm.n1034 C10_N_btm.n1033 0.228786
R25069 C10_N_btm.n1035 C10_N_btm.n42 0.228786
R25070 C10_N_btm.n1036 C10_N_btm.n1035 0.228786
R25071 C10_N_btm.n1034 C10_N_btm.n41 0.228786
R25072 C10_N_btm.n41 C10_N_btm.n40 0.228786
R25073 C10_N_btm.n1037 C10_N_btm.n1036 0.228786
R25074 C10_N_btm.n1038 C10_N_btm.n1037 0.228786
R25075 C10_N_btm.n1039 C10_N_btm.n40 0.228786
R25076 C10_N_btm.n1040 C10_N_btm.n1039 0.228786
R25077 C10_N_btm.n1038 C10_N_btm.n37 0.228786
R25078 C10_N_btm.n37 C10_N_btm.n34 0.228786
R25079 C10_N_btm.n1041 C10_N_btm.n1040 0.228786
R25080 C10_N_btm.n1042 C10_N_btm.n1041 0.228786
R25081 C10_N_btm.n1043 C10_N_btm.n34 0.228786
R25082 C10_N_btm.n1044 C10_N_btm.n1043 0.228786
R25083 C10_N_btm.n1042 C10_N_btm.n33 0.228786
R25084 C10_N_btm.n181 C10_N_btm.n131 0.208893
R25085 C10_N_btm.n923 C10_N_btm.n217 0.208893
R25086 C10_N_btm.n645 C10_N_btm.n643 0.208893
R25087 C10_N_btm.n597 C10_N_btm.n596 0.208893
R25088 C10_N_btm.n864 C10_N_btm.n272 0.208893
R25089 C10_N_btm.n824 C10_N_btm.n305 0.208893
R25090 C10_N_btm.n425 C10_N_btm.n424 0.208893
R25091 C10_N_btm.n1008 C10_N_btm.n66 0.09425
R25092 C10_N_btm.n1004 C10_N_btm.n62 0.09425
R25093 C10_N_btm.n1017 C10_N_btm.n60 0.09425
R25094 C10_N_btm.n87 C10_N_btm.n86 0.09425
R25095 C10_N_btm.n1023 C10_N_btm.n55 0.09425
R25096 C10_N_btm.n96 C10_N_btm.n51 0.09425
R25097 C10_N_btm.n103 C10_N_btm.n49 0.09425
R25098 C10_N_btm.n107 C10_N_btm.n46 0.09425
R25099 C10_N_btm.n1033 C10_N_btm.n44 0.09425
R25100 C10_N_btm.n118 C10_N_btm.n117 0.09425
R25101 C10_N_btm.n1039 C10_N_btm.n39 0.09425
R25102 C10_N_btm.n127 C10_N_btm.n35 0.09425
R25103 C10_N_btm.n128 C10_N_btm.n33 0.09425
R25104 C10_N_btm.n129 C10_N_btm.n128 0.09425
R25105 C10_N_btm.n972 C10_N_btm.n129 0.09425
R25106 C10_N_btm.n973 C10_N_btm.n127 0.09425
R25107 C10_N_btm.n973 C10_N_btm.n124 0.09425
R25108 C10_N_btm.n972 C10_N_btm.n971 0.09425
R25109 C10_N_btm.n971 C10_N_btm.n970 0.09425
R25110 C10_N_btm.n130 C10_N_btm.n124 0.09425
R25111 C10_N_btm.n968 C10_N_btm.n130 0.09425
R25112 C10_N_btm.n970 C10_N_btm.n969 0.09425
R25113 C10_N_btm.n969 C10_N_btm.n131 0.09425
R25114 C10_N_btm.n968 C10_N_btm.n967 0.09425
R25115 C10_N_btm.n967 C10_N_btm.n133 0.09425
R25116 C10_N_btm.n182 C10_N_btm.n134 0.09425
R25117 C10_N_btm.n965 C10_N_btm.n135 0.09425
R25118 C10_N_btm.n183 C10_N_btm.n135 0.09425
R25119 C10_N_btm.n966 C10_N_btm.n132 0.09425
R25120 C10_N_btm.n966 C10_N_btm.n134 0.09425
R25121 C10_N_btm.n964 C10_N_btm.n122 0.09425
R25122 C10_N_btm.n965 C10_N_btm.n964 0.09425
R25123 C10_N_btm.n975 C10_N_btm.n123 0.09425
R25124 C10_N_btm.n132 C10_N_btm.n123 0.09425
R25125 C10_N_btm.n976 C10_N_btm.n120 0.09425
R25126 C10_N_btm.n976 C10_N_btm.n122 0.09425
R25127 C10_N_btm.n974 C10_N_btm.n126 0.09425
R25128 C10_N_btm.n975 C10_N_btm.n974 0.09425
R25129 C10_N_btm.n125 C10_N_btm.n38 0.09425
R25130 C10_N_btm.n125 C10_N_btm.n120 0.09425
R25131 C10_N_btm.n1041 C10_N_btm.n36 0.09425
R25132 C10_N_btm.n126 C10_N_btm.n36 0.09425
R25133 C10_N_btm.n119 C10_N_btm.n39 0.09425
R25134 C10_N_btm.n978 C10_N_btm.n119 0.09425
R25135 C10_N_btm.n979 C10_N_btm.n118 0.09425
R25136 C10_N_btm.n979 C10_N_btm.n113 0.09425
R25137 C10_N_btm.n978 C10_N_btm.n977 0.09425
R25138 C10_N_btm.n977 C10_N_btm.n121 0.09425
R25139 C10_N_btm.n137 C10_N_btm.n113 0.09425
R25140 C10_N_btm.n962 C10_N_btm.n137 0.09425
R25141 C10_N_btm.n963 C10_N_btm.n121 0.09425
R25142 C10_N_btm.n963 C10_N_btm.n136 0.09425
R25143 C10_N_btm.n962 C10_N_btm.n961 0.09425
R25144 C10_N_btm.n961 C10_N_btm.n139 0.09425
R25145 C10_N_btm.n184 C10_N_btm.n136 0.09425
R25146 C10_N_btm.n185 C10_N_btm.n184 0.09425
R25147 C10_N_btm.n186 C10_N_btm.n139 0.09425
R25148 C10_N_btm.n187 C10_N_btm.n140 0.09425
R25149 C10_N_btm.n959 C10_N_btm.n141 0.09425
R25150 C10_N_btm.n188 C10_N_btm.n141 0.09425
R25151 C10_N_btm.n960 C10_N_btm.n138 0.09425
R25152 C10_N_btm.n960 C10_N_btm.n140 0.09425
R25153 C10_N_btm.n958 C10_N_btm.n111 0.09425
R25154 C10_N_btm.n959 C10_N_btm.n958 0.09425
R25155 C10_N_btm.n981 C10_N_btm.n112 0.09425
R25156 C10_N_btm.n138 C10_N_btm.n112 0.09425
R25157 C10_N_btm.n982 C10_N_btm.n109 0.09425
R25158 C10_N_btm.n982 C10_N_btm.n111 0.09425
R25159 C10_N_btm.n980 C10_N_btm.n115 0.09425
R25160 C10_N_btm.n981 C10_N_btm.n980 0.09425
R25161 C10_N_btm.n114 C10_N_btm.n43 0.09425
R25162 C10_N_btm.n114 C10_N_btm.n109 0.09425
R25163 C10_N_btm.n116 C10_N_btm.n41 0.09425
R25164 C10_N_btm.n116 C10_N_btm.n115 0.09425
R25165 C10_N_btm.n108 C10_N_btm.n44 0.09425
R25166 C10_N_btm.n984 C10_N_btm.n108 0.09425
R25167 C10_N_btm.n985 C10_N_btm.n107 0.09425
R25168 C10_N_btm.n985 C10_N_btm.n102 0.09425
R25169 C10_N_btm.n984 C10_N_btm.n983 0.09425
R25170 C10_N_btm.n983 C10_N_btm.n110 0.09425
R25171 C10_N_btm.n143 C10_N_btm.n102 0.09425
R25172 C10_N_btm.n956 C10_N_btm.n143 0.09425
R25173 C10_N_btm.n957 C10_N_btm.n110 0.09425
R25174 C10_N_btm.n957 C10_N_btm.n142 0.09425
R25175 C10_N_btm.n956 C10_N_btm.n955 0.09425
R25176 C10_N_btm.n955 C10_N_btm.n145 0.09425
R25177 C10_N_btm.n189 C10_N_btm.n142 0.09425
R25178 C10_N_btm.n190 C10_N_btm.n189 0.09425
R25179 C10_N_btm.n191 C10_N_btm.n145 0.09425
R25180 C10_N_btm.n192 C10_N_btm.n146 0.09425
R25181 C10_N_btm.n953 C10_N_btm.n147 0.09425
R25182 C10_N_btm.n193 C10_N_btm.n147 0.09425
R25183 C10_N_btm.n954 C10_N_btm.n144 0.09425
R25184 C10_N_btm.n954 C10_N_btm.n146 0.09425
R25185 C10_N_btm.n952 C10_N_btm.n100 0.09425
R25186 C10_N_btm.n953 C10_N_btm.n952 0.09425
R25187 C10_N_btm.n987 C10_N_btm.n101 0.09425
R25188 C10_N_btm.n144 C10_N_btm.n101 0.09425
R25189 C10_N_btm.n988 C10_N_btm.n98 0.09425
R25190 C10_N_btm.n988 C10_N_btm.n100 0.09425
R25191 C10_N_btm.n986 C10_N_btm.n106 0.09425
R25192 C10_N_btm.n987 C10_N_btm.n986 0.09425
R25193 C10_N_btm.n105 C10_N_btm.n104 0.09425
R25194 C10_N_btm.n105 C10_N_btm.n98 0.09425
R25195 C10_N_btm.n1031 C10_N_btm.n47 0.09425
R25196 C10_N_btm.n106 C10_N_btm.n47 0.09425
R25197 C10_N_btm.n103 C10_N_btm.n97 0.09425
R25198 C10_N_btm.n990 C10_N_btm.n97 0.09425
R25199 C10_N_btm.n991 C10_N_btm.n96 0.09425
R25200 C10_N_btm.n991 C10_N_btm.n93 0.09425
R25201 C10_N_btm.n990 C10_N_btm.n989 0.09425
R25202 C10_N_btm.n989 C10_N_btm.n99 0.09425
R25203 C10_N_btm.n149 C10_N_btm.n93 0.09425
R25204 C10_N_btm.n950 C10_N_btm.n149 0.09425
R25205 C10_N_btm.n951 C10_N_btm.n99 0.09425
R25206 C10_N_btm.n951 C10_N_btm.n148 0.09425
R25207 C10_N_btm.n950 C10_N_btm.n949 0.09425
R25208 C10_N_btm.n949 C10_N_btm.n151 0.09425
R25209 C10_N_btm.n194 C10_N_btm.n148 0.09425
R25210 C10_N_btm.n195 C10_N_btm.n194 0.09425
R25211 C10_N_btm.n196 C10_N_btm.n151 0.09425
R25212 C10_N_btm.n197 C10_N_btm.n152 0.09425
R25213 C10_N_btm.n947 C10_N_btm.n153 0.09425
R25214 C10_N_btm.n198 C10_N_btm.n153 0.09425
R25215 C10_N_btm.n948 C10_N_btm.n150 0.09425
R25216 C10_N_btm.n948 C10_N_btm.n152 0.09425
R25217 C10_N_btm.n946 C10_N_btm.n91 0.09425
R25218 C10_N_btm.n947 C10_N_btm.n946 0.09425
R25219 C10_N_btm.n993 C10_N_btm.n92 0.09425
R25220 C10_N_btm.n150 C10_N_btm.n92 0.09425
R25221 C10_N_btm.n994 C10_N_btm.n89 0.09425
R25222 C10_N_btm.n994 C10_N_btm.n91 0.09425
R25223 C10_N_btm.n992 C10_N_btm.n95 0.09425
R25224 C10_N_btm.n993 C10_N_btm.n992 0.09425
R25225 C10_N_btm.n94 C10_N_btm.n54 0.09425
R25226 C10_N_btm.n94 C10_N_btm.n89 0.09425
R25227 C10_N_btm.n1025 C10_N_btm.n52 0.09425
R25228 C10_N_btm.n95 C10_N_btm.n52 0.09425
R25229 C10_N_btm.n88 C10_N_btm.n55 0.09425
R25230 C10_N_btm.n996 C10_N_btm.n88 0.09425
R25231 C10_N_btm.n997 C10_N_btm.n87 0.09425
R25232 C10_N_btm.n997 C10_N_btm.n82 0.09425
R25233 C10_N_btm.n996 C10_N_btm.n995 0.09425
R25234 C10_N_btm.n995 C10_N_btm.n90 0.09425
R25235 C10_N_btm.n155 C10_N_btm.n82 0.09425
R25236 C10_N_btm.n944 C10_N_btm.n155 0.09425
R25237 C10_N_btm.n945 C10_N_btm.n90 0.09425
R25238 C10_N_btm.n945 C10_N_btm.n154 0.09425
R25239 C10_N_btm.n944 C10_N_btm.n943 0.09425
R25240 C10_N_btm.n943 C10_N_btm.n157 0.09425
R25241 C10_N_btm.n199 C10_N_btm.n154 0.09425
R25242 C10_N_btm.n200 C10_N_btm.n199 0.09425
R25243 C10_N_btm.n201 C10_N_btm.n157 0.09425
R25244 C10_N_btm.n202 C10_N_btm.n158 0.09425
R25245 C10_N_btm.n941 C10_N_btm.n159 0.09425
R25246 C10_N_btm.n203 C10_N_btm.n159 0.09425
R25247 C10_N_btm.n942 C10_N_btm.n156 0.09425
R25248 C10_N_btm.n942 C10_N_btm.n158 0.09425
R25249 C10_N_btm.n940 C10_N_btm.n80 0.09425
R25250 C10_N_btm.n941 C10_N_btm.n940 0.09425
R25251 C10_N_btm.n999 C10_N_btm.n81 0.09425
R25252 C10_N_btm.n156 C10_N_btm.n81 0.09425
R25253 C10_N_btm.n1000 C10_N_btm.n78 0.09425
R25254 C10_N_btm.n1000 C10_N_btm.n80 0.09425
R25255 C10_N_btm.n998 C10_N_btm.n84 0.09425
R25256 C10_N_btm.n999 C10_N_btm.n998 0.09425
R25257 C10_N_btm.n83 C10_N_btm.n59 0.09425
R25258 C10_N_btm.n83 C10_N_btm.n78 0.09425
R25259 C10_N_btm.n85 C10_N_btm.n57 0.09425
R25260 C10_N_btm.n85 C10_N_btm.n84 0.09425
R25261 C10_N_btm.n76 C10_N_btm.n60 0.09425
R25262 C10_N_btm.n1002 C10_N_btm.n76 0.09425
R25263 C10_N_btm.n1004 C10_N_btm.n1003 0.09425
R25264 C10_N_btm.n1003 C10_N_btm.n77 0.09425
R25265 C10_N_btm.n1002 C10_N_btm.n1001 0.09425
R25266 C10_N_btm.n1001 C10_N_btm.n79 0.09425
R25267 C10_N_btm.n161 C10_N_btm.n77 0.09425
R25268 C10_N_btm.n938 C10_N_btm.n161 0.09425
R25269 C10_N_btm.n939 C10_N_btm.n79 0.09425
R25270 C10_N_btm.n939 C10_N_btm.n160 0.09425
R25271 C10_N_btm.n938 C10_N_btm.n937 0.09425
R25272 C10_N_btm.n937 C10_N_btm.n163 0.09425
R25273 C10_N_btm.n204 C10_N_btm.n160 0.09425
R25274 C10_N_btm.n205 C10_N_btm.n204 0.09425
R25275 C10_N_btm.n206 C10_N_btm.n163 0.09425
R25276 C10_N_btm.n207 C10_N_btm.n164 0.09425
R25277 C10_N_btm.n935 C10_N_btm.n165 0.09425
R25278 C10_N_btm.n208 C10_N_btm.n165 0.09425
R25279 C10_N_btm.n936 C10_N_btm.n162 0.09425
R25280 C10_N_btm.n936 C10_N_btm.n164 0.09425
R25281 C10_N_btm.n934 C10_N_btm.n167 0.09425
R25282 C10_N_btm.n935 C10_N_btm.n934 0.09425
R25283 C10_N_btm.n227 C10_N_btm.n226 0.09425
R25284 C10_N_btm.n226 C10_N_btm.n162 0.09425
R25285 C10_N_btm.n228 C10_N_btm.n74 0.09425
R25286 C10_N_btm.n228 C10_N_btm.n167 0.09425
R25287 C10_N_btm.n1005 C10_N_btm.n75 0.09425
R25288 C10_N_btm.n227 C10_N_btm.n75 0.09425
R25289 C10_N_btm.n1006 C10_N_btm.n72 0.09425
R25290 C10_N_btm.n1006 C10_N_btm.n74 0.09425
R25291 C10_N_btm.n1015 C10_N_btm.n63 0.09425
R25292 C10_N_btm.n1005 C10_N_btm.n63 0.09425
R25293 C10_N_btm.n1011 C10_N_btm.n1010 0.09425
R25294 C10_N_btm.n1010 C10_N_btm.n1009 0.09425
R25295 C10_N_btm.n1009 C10_N_btm.n70 0.09425
R25296 C10_N_btm.n1008 C10_N_btm.n1007 0.09425
R25297 C10_N_btm.n1007 C10_N_btm.n73 0.09425
R25298 C10_N_btm.n911 C10_N_btm.n70 0.09425
R25299 C10_N_btm.n911 C10_N_btm.n230 0.09425
R25300 C10_N_btm.n229 C10_N_btm.n73 0.09425
R25301 C10_N_btm.n229 C10_N_btm.n168 0.09425
R25302 C10_N_btm.n230 C10_N_btm.n169 0.09425
R25303 C10_N_btm.n932 C10_N_btm.n169 0.09425
R25304 C10_N_btm.n933 C10_N_btm.n168 0.09425
R25305 C10_N_btm.n933 C10_N_btm.n166 0.09425
R25306 C10_N_btm.n932 C10_N_btm.n931 0.09425
R25307 C10_N_btm.n931 C10_N_btm.n171 0.09425
R25308 C10_N_btm.n209 C10_N_btm.n166 0.09425
R25309 C10_N_btm.n210 C10_N_btm.n209 0.09425
R25310 C10_N_btm.n211 C10_N_btm.n171 0.09425
R25311 C10_N_btm.n212 C10_N_btm.n172 0.09425
R25312 C10_N_btm.n929 C10_N_btm.n173 0.09425
R25313 C10_N_btm.n213 C10_N_btm.n173 0.09425
R25314 C10_N_btm.n930 C10_N_btm.n170 0.09425
R25315 C10_N_btm.n930 C10_N_btm.n172 0.09425
R25316 C10_N_btm.n928 C10_N_btm.n175 0.09425
R25317 C10_N_btm.n929 C10_N_btm.n928 0.09425
R25318 C10_N_btm.n913 C10_N_btm.n225 0.09425
R25319 C10_N_btm.n225 C10_N_btm.n170 0.09425
R25320 C10_N_btm.n914 C10_N_btm.n224 0.09425
R25321 C10_N_btm.n914 C10_N_btm.n175 0.09425
R25322 C10_N_btm.n912 C10_N_btm.n910 0.09425
R25323 C10_N_btm.n913 C10_N_btm.n912 0.09425
R25324 C10_N_btm.n909 C10_N_btm.n908 0.09425
R25325 C10_N_btm.n909 C10_N_btm.n224 0.09425
R25326 C10_N_btm.n71 C10_N_btm.n69 0.09425
R25327 C10_N_btm.n910 C10_N_btm.n71 0.09425
R25328 C10_N_btm.n907 C10_N_btm.n232 0.09425
R25329 C10_N_btm.n908 C10_N_btm.n907 0.09425
R25330 C10_N_btm.n892 C10_N_btm.n67 0.09425
R25331 C10_N_btm.n69 C10_N_btm.n67 0.09425
R25332 C10_N_btm.n893 C10_N_btm.n243 0.09425
R25333 C10_N_btm.n893 C10_N_btm.n232 0.09425
R25334 C10_N_btm.n895 C10_N_btm.n242 0.09425
R25335 C10_N_btm.n880 C10_N_btm.n241 0.09425
R25336 C10_N_btm.n896 C10_N_btm.n241 0.09425
R25337 C10_N_btm.n896 C10_N_btm.n239 0.09425
R25338 C10_N_btm.n895 C10_N_btm.n894 0.09425
R25339 C10_N_btm.n894 C10_N_btm.n233 0.09425
R25340 C10_N_btm.n239 C10_N_btm.n234 0.09425
R25341 C10_N_btm.n905 C10_N_btm.n234 0.09425
R25342 C10_N_btm.n906 C10_N_btm.n233 0.09425
R25343 C10_N_btm.n906 C10_N_btm.n231 0.09425
R25344 C10_N_btm.n905 C10_N_btm.n904 0.09425
R25345 C10_N_btm.n904 C10_N_btm.n222 0.09425
R25346 C10_N_btm.n231 C10_N_btm.n223 0.09425
R25347 C10_N_btm.n916 C10_N_btm.n223 0.09425
R25348 C10_N_btm.n917 C10_N_btm.n222 0.09425
R25349 C10_N_btm.n917 C10_N_btm.n220 0.09425
R25350 C10_N_btm.n916 C10_N_btm.n915 0.09425
R25351 C10_N_btm.n915 C10_N_btm.n176 0.09425
R25352 C10_N_btm.n220 C10_N_btm.n177 0.09425
R25353 C10_N_btm.n926 C10_N_btm.n177 0.09425
R25354 C10_N_btm.n927 C10_N_btm.n176 0.09425
R25355 C10_N_btm.n927 C10_N_btm.n174 0.09425
R25356 C10_N_btm.n926 C10_N_btm.n925 0.09425
R25357 C10_N_btm.n925 C10_N_btm.n179 0.09425
R25358 C10_N_btm.n214 C10_N_btm.n174 0.09425
R25359 C10_N_btm.n215 C10_N_btm.n214 0.09425
R25360 C10_N_btm.n216 C10_N_btm.n179 0.09425
R25361 C10_N_btm.n924 C10_N_btm.n178 0.09425
R25362 C10_N_btm.n924 C10_N_btm.n180 0.09425
R25363 C10_N_btm.n922 C10_N_btm.n921 0.09425
R25364 C10_N_btm.n923 C10_N_btm.n922 0.09425
R25365 C10_N_btm.n919 C10_N_btm.n218 0.09425
R25366 C10_N_btm.n218 C10_N_btm.n178 0.09425
R25367 C10_N_btm.n920 C10_N_btm.n219 0.09425
R25368 C10_N_btm.n921 C10_N_btm.n920 0.09425
R25369 C10_N_btm.n918 C10_N_btm.n221 0.09425
R25370 C10_N_btm.n919 C10_N_btm.n918 0.09425
R25371 C10_N_btm.n902 C10_N_btm.n236 0.09425
R25372 C10_N_btm.n236 C10_N_btm.n219 0.09425
R25373 C10_N_btm.n903 C10_N_btm.n235 0.09425
R25374 C10_N_btm.n903 C10_N_btm.n221 0.09425
R25375 C10_N_btm.n901 C10_N_btm.n900 0.09425
R25376 C10_N_btm.n902 C10_N_btm.n901 0.09425
R25377 C10_N_btm.n898 C10_N_btm.n237 0.09425
R25378 C10_N_btm.n237 C10_N_btm.n235 0.09425
R25379 C10_N_btm.n899 C10_N_btm.n238 0.09425
R25380 C10_N_btm.n900 C10_N_btm.n899 0.09425
R25381 C10_N_btm.n897 C10_N_btm.n240 0.09425
R25382 C10_N_btm.n898 C10_N_btm.n897 0.09425
R25383 C10_N_btm.n878 C10_N_btm.n255 0.09425
R25384 C10_N_btm.n255 C10_N_btm.n238 0.09425
R25385 C10_N_btm.n879 C10_N_btm.n254 0.09425
R25386 C10_N_btm.n879 C10_N_btm.n240 0.09425
R25387 C10_N_btm.n878 C10_N_btm.n877 0.09425
R25388 C10_N_btm.n877 C10_N_btm.n876 0.09425
R25389 C10_N_btm.n534 C10_N_btm.n478 0.09425
R25390 C10_N_btm.n577 C10_N_btm.n479 0.09425
R25391 C10_N_btm.n540 C10_N_btm.n482 0.09425
R25392 C10_N_btm.n573 C10_N_btm.n483 0.09425
R25393 C10_N_btm.n546 C10_N_btm.n486 0.09425
R25394 C10_N_btm.n567 C10_N_btm.n487 0.09425
R25395 C10_N_btm.n552 C10_N_btm.n490 0.09425
R25396 C10_N_btm.n561 C10_N_btm.n560 0.09425
R25397 C10_N_btm.n637 C10_N_btm.n418 0.09425
R25398 C10_N_btm.n638 C10_N_btm.n417 0.09425
R25399 C10_N_btm.n643 C10_N_btm.n642 0.09425
R25400 C10_N_btm.n642 C10_N_btm.n641 0.09425
R25401 C10_N_btm.n641 C10_N_btm.n640 0.09425
R25402 C10_N_btm.n425 C10_N_btm.n416 0.09425
R25403 C10_N_btm.n639 C10_N_btm.n416 0.09425
R25404 C10_N_btm.n640 C10_N_btm.n639 0.09425
R25405 C10_N_btm.n638 C10_N_btm.n415 0.09425
R25406 C10_N_btm.n415 C10_N_btm.n414 0.09425
R25407 C10_N_btm.n555 C10_N_btm.n418 0.09425
R25408 C10_N_btm.n555 C10_N_btm.n412 0.09425
R25409 C10_N_btm.n414 C10_N_btm.n413 0.09425
R25410 C10_N_btm.n647 C10_N_btm.n413 0.09425
R25411 C10_N_btm.n648 C10_N_btm.n412 0.09425
R25412 C10_N_btm.n648 C10_N_btm.n410 0.09425
R25413 C10_N_btm.n647 C10_N_btm.n646 0.09425
R25414 C10_N_btm.n644 C10_N_btm.n410 0.09425
R25415 C10_N_btm.n650 C10_N_btm.n409 0.09425
R25416 C10_N_btm.n651 C10_N_btm.n405 0.09425
R25417 C10_N_btm.n651 C10_N_btm.n408 0.09425
R25418 C10_N_btm.n649 C10_N_btm.n411 0.09425
R25419 C10_N_btm.n650 C10_N_btm.n649 0.09425
R25420 C10_N_btm.n554 C10_N_btm.n553 0.09425
R25421 C10_N_btm.n553 C10_N_btm.n405 0.09425
R25422 C10_N_btm.n557 C10_N_btm.n556 0.09425
R25423 C10_N_btm.n556 C10_N_btm.n411 0.09425
R25424 C10_N_btm.n558 C10_N_btm.n491 0.09425
R25425 C10_N_btm.n558 C10_N_btm.n554 0.09425
R25426 C10_N_btm.n635 C10_N_btm.n419 0.09425
R25427 C10_N_btm.n557 C10_N_btm.n419 0.09425
R25428 C10_N_btm.n560 C10_N_btm.n559 0.09425
R25429 C10_N_btm.n559 C10_N_btm.n492 0.09425
R25430 C10_N_btm.n552 C10_N_btm.n551 0.09425
R25431 C10_N_btm.n551 C10_N_btm.n403 0.09425
R25432 C10_N_btm.n492 C10_N_btm.n404 0.09425
R25433 C10_N_btm.n653 C10_N_btm.n404 0.09425
R25434 C10_N_btm.n654 C10_N_btm.n403 0.09425
R25435 C10_N_btm.n654 C10_N_btm.n401 0.09425
R25436 C10_N_btm.n653 C10_N_btm.n652 0.09425
R25437 C10_N_btm.n652 C10_N_btm.n407 0.09425
R25438 C10_N_btm.n406 C10_N_btm.n401 0.09425
R25439 C10_N_btm.n656 C10_N_btm.n400 0.09425
R25440 C10_N_btm.n657 C10_N_btm.n396 0.09425
R25441 C10_N_btm.n657 C10_N_btm.n399 0.09425
R25442 C10_N_btm.n655 C10_N_btm.n402 0.09425
R25443 C10_N_btm.n656 C10_N_btm.n655 0.09425
R25444 C10_N_btm.n549 C10_N_btm.n494 0.09425
R25445 C10_N_btm.n494 C10_N_btm.n396 0.09425
R25446 C10_N_btm.n550 C10_N_btm.n493 0.09425
R25447 C10_N_btm.n550 C10_N_btm.n402 0.09425
R25448 C10_N_btm.n548 C10_N_btm.n488 0.09425
R25449 C10_N_btm.n549 C10_N_btm.n548 0.09425
R25450 C10_N_btm.n565 C10_N_btm.n489 0.09425
R25451 C10_N_btm.n493 C10_N_btm.n489 0.09425
R25452 C10_N_btm.n547 C10_N_btm.n487 0.09425
R25453 C10_N_btm.n547 C10_N_btm.n495 0.09425
R25454 C10_N_btm.n546 C10_N_btm.n545 0.09425
R25455 C10_N_btm.n545 C10_N_btm.n394 0.09425
R25456 C10_N_btm.n495 C10_N_btm.n395 0.09425
R25457 C10_N_btm.n659 C10_N_btm.n395 0.09425
R25458 C10_N_btm.n660 C10_N_btm.n394 0.09425
R25459 C10_N_btm.n660 C10_N_btm.n392 0.09425
R25460 C10_N_btm.n659 C10_N_btm.n658 0.09425
R25461 C10_N_btm.n658 C10_N_btm.n398 0.09425
R25462 C10_N_btm.n397 C10_N_btm.n392 0.09425
R25463 C10_N_btm.n662 C10_N_btm.n391 0.09425
R25464 C10_N_btm.n663 C10_N_btm.n387 0.09425
R25465 C10_N_btm.n663 C10_N_btm.n390 0.09425
R25466 C10_N_btm.n661 C10_N_btm.n393 0.09425
R25467 C10_N_btm.n662 C10_N_btm.n661 0.09425
R25468 C10_N_btm.n543 C10_N_btm.n497 0.09425
R25469 C10_N_btm.n497 C10_N_btm.n387 0.09425
R25470 C10_N_btm.n544 C10_N_btm.n496 0.09425
R25471 C10_N_btm.n544 C10_N_btm.n393 0.09425
R25472 C10_N_btm.n542 C10_N_btm.n484 0.09425
R25473 C10_N_btm.n543 C10_N_btm.n542 0.09425
R25474 C10_N_btm.n569 C10_N_btm.n485 0.09425
R25475 C10_N_btm.n496 C10_N_btm.n485 0.09425
R25476 C10_N_btm.n541 C10_N_btm.n483 0.09425
R25477 C10_N_btm.n541 C10_N_btm.n498 0.09425
R25478 C10_N_btm.n540 C10_N_btm.n539 0.09425
R25479 C10_N_btm.n539 C10_N_btm.n385 0.09425
R25480 C10_N_btm.n498 C10_N_btm.n386 0.09425
R25481 C10_N_btm.n665 C10_N_btm.n386 0.09425
R25482 C10_N_btm.n666 C10_N_btm.n385 0.09425
R25483 C10_N_btm.n666 C10_N_btm.n383 0.09425
R25484 C10_N_btm.n665 C10_N_btm.n664 0.09425
R25485 C10_N_btm.n664 C10_N_btm.n389 0.09425
R25486 C10_N_btm.n388 C10_N_btm.n383 0.09425
R25487 C10_N_btm.n668 C10_N_btm.n382 0.09425
R25488 C10_N_btm.n669 C10_N_btm.n381 0.09425
R25489 C10_N_btm.n669 C10_N_btm.n379 0.09425
R25490 C10_N_btm.n667 C10_N_btm.n384 0.09425
R25491 C10_N_btm.n668 C10_N_btm.n667 0.09425
R25492 C10_N_btm.n537 C10_N_btm.n500 0.09425
R25493 C10_N_btm.n500 C10_N_btm.n381 0.09425
R25494 C10_N_btm.n538 C10_N_btm.n499 0.09425
R25495 C10_N_btm.n538 C10_N_btm.n384 0.09425
R25496 C10_N_btm.n536 C10_N_btm.n480 0.09425
R25497 C10_N_btm.n537 C10_N_btm.n536 0.09425
R25498 C10_N_btm.n575 C10_N_btm.n481 0.09425
R25499 C10_N_btm.n499 C10_N_btm.n481 0.09425
R25500 C10_N_btm.n535 C10_N_btm.n479 0.09425
R25501 C10_N_btm.n535 C10_N_btm.n501 0.09425
R25502 C10_N_btm.n534 C10_N_btm.n533 0.09425
R25503 C10_N_btm.n533 C10_N_btm.n504 0.09425
R25504 C10_N_btm.n503 C10_N_btm.n501 0.09425
R25505 C10_N_btm.n503 C10_N_btm.n380 0.09425
R25506 C10_N_btm.n506 C10_N_btm.n504 0.09425
R25507 C10_N_btm.n506 C10_N_btm.n378 0.09425
R25508 C10_N_btm.n670 C10_N_btm.n380 0.09425
R25509 C10_N_btm.n671 C10_N_btm.n670 0.09425
R25510 C10_N_btm.n672 C10_N_btm.n378 0.09425
R25511 C10_N_btm.n673 C10_N_btm.n377 0.09425
R25512 C10_N_btm.n676 C10_N_btm.n675 0.09425
R25513 C10_N_btm.n508 C10_N_btm.n376 0.09425
R25514 C10_N_btm.n674 C10_N_btm.n376 0.09425
R25515 C10_N_btm.n507 C10_N_btm.n505 0.09425
R25516 C10_N_btm.n507 C10_N_btm.n377 0.09425
R25517 C10_N_btm.n531 C10_N_btm.n509 0.09425
R25518 C10_N_btm.n509 C10_N_btm.n508 0.09425
R25519 C10_N_btm.n532 C10_N_btm.n502 0.09425
R25520 C10_N_btm.n532 C10_N_btm.n505 0.09425
R25521 C10_N_btm.n530 C10_N_btm.n476 0.09425
R25522 C10_N_btm.n531 C10_N_btm.n530 0.09425
R25523 C10_N_btm.n581 C10_N_btm.n477 0.09425
R25524 C10_N_btm.n502 C10_N_btm.n477 0.09425
R25525 C10_N_btm.n583 C10_N_btm.n475 0.09425
R25526 C10_N_btm.n529 C10_N_btm.n475 0.09425
R25527 C10_N_btm.n528 C10_N_btm.n474 0.09425
R25528 C10_N_btm.n528 C10_N_btm.n512 0.09425
R25529 C10_N_btm.n529 C10_N_btm.n511 0.09425
R25530 C10_N_btm.n511 C10_N_btm.n510 0.09425
R25531 C10_N_btm.n512 C10_N_btm.n365 0.09425
R25532 C10_N_btm.n678 C10_N_btm.n365 0.09425
R25533 C10_N_btm.n510 C10_N_btm.n366 0.09425
R25534 C10_N_btm.n676 C10_N_btm.n366 0.09425
R25535 C10_N_btm.n679 C10_N_btm.n363 0.09425
R25536 C10_N_btm.n679 C10_N_btm.n364 0.09425
R25537 C10_N_btm.n678 C10_N_btm.n677 0.09425
R25538 C10_N_btm.n677 C10_N_btm.n375 0.09425
R25539 C10_N_btm.n374 C10_N_btm.n364 0.09425
R25540 C10_N_btm.n883 C10_N_btm.n251 0.09425
R25541 C10_N_btm.n883 C10_N_btm.n249 0.09425
R25542 C10_N_btm.n885 C10_N_btm.n244 0.09425
R25543 C10_N_btm.n890 C10_N_btm.n245 0.09425
R25544 C10_N_btm.n889 C10_N_btm.n65 0.09425
R25545 C10_N_btm.n269 C10_N_btm.n246 0.09425
R25546 C10_N_btm.n887 C10_N_btm.n246 0.09425
R25547 C10_N_btm.n888 C10_N_btm.n887 0.09425
R25548 C10_N_btm.n889 C10_N_btm.n888 0.09425
R25549 C10_N_btm.n886 C10_N_btm.n247 0.09425
R25550 C10_N_btm.n886 C10_N_btm.n245 0.09425
R25551 C10_N_btm.n265 C10_N_btm.n250 0.09425
R25552 C10_N_btm.n872 C10_N_btm.n252 0.09425
R25553 C10_N_btm.n882 C10_N_btm.n252 0.09425
R25554 C10_N_btm.n884 C10_N_btm.n250 0.09425
R25555 C10_N_btm.n885 C10_N_btm.n884 0.09425
R25556 C10_N_btm.n268 C10_N_btm.n267 0.09425
R25557 C10_N_btm.n268 C10_N_btm.n247 0.09425
R25558 C10_N_btm.n867 C10_N_btm.n270 0.09425
R25559 C10_N_btm.n270 C10_N_btm.n269 0.09425
R25560 C10_N_btm.n868 C10_N_btm.n266 0.09425
R25561 C10_N_btm.n868 C10_N_btm.n267 0.09425
R25562 C10_N_btm.n866 C10_N_btm.n865 0.09425
R25563 C10_N_btm.n867 C10_N_btm.n866 0.09425
R25564 C10_N_btm.n863 C10_N_btm.n271 0.09425
R25565 C10_N_btm.n271 C10_N_btm.n266 0.09425
R25566 C10_N_btm.n865 C10_N_btm.n864 0.09425
R25567 C10_N_btm.n863 C10_N_btm.n862 0.09425
R25568 C10_N_btm.n841 C10_N_btm.n289 0.09425
R25569 C10_N_btm.n841 C10_N_btm.n840 0.09425
R25570 C10_N_btm.n840 C10_N_btm.n839 0.09425
R25571 C10_N_btm.n839 C10_N_btm.n838 0.09425
R25572 C10_N_btm.n838 C10_N_btm.n837 0.09425
R25573 C10_N_btm.n837 C10_N_btm.n836 0.09425
R25574 C10_N_btm.n836 C10_N_btm.n835 0.09425
R25575 C10_N_btm.n835 C10_N_btm.n834 0.09425
R25576 C10_N_btm.n834 C10_N_btm.n833 0.09425
R25577 C10_N_btm.n833 C10_N_btm.n832 0.09425
R25578 C10_N_btm.n832 C10_N_btm.n831 0.09425
R25579 C10_N_btm.n831 C10_N_btm.n830 0.09425
R25580 C10_N_btm.n830 C10_N_btm.n829 0.09425
R25581 C10_N_btm.n829 C10_N_btm.n828 0.09425
R25582 C10_N_btm.n828 C10_N_btm.n827 0.09425
R25583 C10_N_btm.n827 C10_N_btm.n826 0.09425
R25584 C10_N_btm.n826 C10_N_btm.n825 0.09425
R25585 C10_N_btm.n823 C10_N_btm.n306 0.09425
R25586 C10_N_btm.n326 C10_N_btm.n305 0.09425
R25587 C10_N_btm.n332 C10_N_btm.n327 0.09425
R25588 C10_N_btm.n327 C10_N_btm.n306 0.09425
R25589 C10_N_btm.n334 C10_N_btm.n333 0.09425
R25590 C10_N_btm.n333 C10_N_btm.n326 0.09425
R25591 C10_N_btm.n727 C10_N_btm.n325 0.09425
R25592 C10_N_btm.n332 C10_N_btm.n325 0.09425
R25593 C10_N_btm.n725 C10_N_btm.n335 0.09425
R25594 C10_N_btm.n335 C10_N_btm.n334 0.09425
R25595 C10_N_btm.n726 C10_N_btm.n336 0.09425
R25596 C10_N_btm.n727 C10_N_btm.n726 0.09425
R25597 C10_N_btm.n724 C10_N_btm.n723 0.09425
R25598 C10_N_btm.n725 C10_N_btm.n724 0.09425
R25599 C10_N_btm.n721 C10_N_btm.n337 0.09425
R25600 C10_N_btm.n337 C10_N_btm.n336 0.09425
R25601 C10_N_btm.n722 C10_N_btm.n338 0.09425
R25602 C10_N_btm.n723 C10_N_btm.n722 0.09425
R25603 C10_N_btm.n720 C10_N_btm.n340 0.09425
R25604 C10_N_btm.n721 C10_N_btm.n720 0.09425
R25605 C10_N_btm.n373 C10_N_btm.n367 0.09425
R25606 C10_N_btm.n367 C10_N_btm.n338 0.09425
R25607 C10_N_btm.n372 C10_N_btm.n361 0.09425
R25608 C10_N_btm.n372 C10_N_btm.n340 0.09425
R25609 C10_N_btm.n680 C10_N_btm.n362 0.09425
R25610 C10_N_btm.n373 C10_N_btm.n362 0.09425
R25611 C10_N_btm.n682 C10_N_btm.n681 0.09425
R25612 C10_N_btm.n681 C10_N_btm.n361 0.09425
R25613 C10_N_btm.n514 C10_N_btm.n360 0.09425
R25614 C10_N_btm.n680 C10_N_btm.n360 0.09425
R25615 C10_N_btm.n527 C10_N_btm.n513 0.09425
R25616 C10_N_btm.n513 C10_N_btm.n363 0.09425
R25617 C10_N_btm.n526 C10_N_btm.n472 0.09425
R25618 C10_N_btm.n526 C10_N_btm.n514 0.09425
R25619 C10_N_btm.n585 C10_N_btm.n473 0.09425
R25620 C10_N_btm.n527 C10_N_btm.n473 0.09425
R25621 C10_N_btm.n589 C10_N_btm.n471 0.09425
R25622 C10_N_btm.n525 C10_N_btm.n471 0.09425
R25623 C10_N_btm.n524 C10_N_btm.n470 0.09425
R25624 C10_N_btm.n524 C10_N_btm.n357 0.09425
R25625 C10_N_btm.n525 C10_N_btm.n359 0.09425
R25626 C10_N_btm.n682 C10_N_btm.n359 0.09425
R25627 C10_N_btm.n523 C10_N_btm.n356 0.09425
R25628 C10_N_btm.n684 C10_N_btm.n356 0.09425
R25629 C10_N_btm.n683 C10_N_btm.n357 0.09425
R25630 C10_N_btm.n683 C10_N_btm.n358 0.09425
R25631 C10_N_btm.n684 C10_N_btm.n354 0.09425
R25632 C10_N_btm.n369 C10_N_btm.n354 0.09425
R25633 C10_N_btm.n368 C10_N_btm.n358 0.09425
R25634 C10_N_btm.n371 C10_N_btm.n368 0.09425
R25635 C10_N_btm.n370 C10_N_btm.n369 0.09425
R25636 C10_N_btm.n370 C10_N_btm.n342 0.09425
R25637 C10_N_btm.n371 C10_N_btm.n341 0.09425
R25638 C10_N_btm.n719 C10_N_btm.n341 0.09425
R25639 C10_N_btm.n718 C10_N_btm.n342 0.09425
R25640 C10_N_btm.n718 C10_N_btm.n343 0.09425
R25641 C10_N_btm.n719 C10_N_btm.n339 0.09425
R25642 C10_N_btm.n703 C10_N_btm.n339 0.09425
R25643 C10_N_btm.n704 C10_N_btm.n343 0.09425
R25644 C10_N_btm.n704 C10_N_btm.n701 0.09425
R25645 C10_N_btm.n703 C10_N_btm.n702 0.09425
R25646 C10_N_btm.n702 C10_N_btm.n323 0.09425
R25647 C10_N_btm.n701 C10_N_btm.n322 0.09425
R25648 C10_N_btm.n729 C10_N_btm.n322 0.09425
R25649 C10_N_btm.n728 C10_N_btm.n323 0.09425
R25650 C10_N_btm.n728 C10_N_btm.n324 0.09425
R25651 C10_N_btm.n729 C10_N_btm.n320 0.09425
R25652 C10_N_btm.n330 C10_N_btm.n320 0.09425
R25653 C10_N_btm.n331 C10_N_btm.n324 0.09425
R25654 C10_N_btm.n331 C10_N_btm.n328 0.09425
R25655 C10_N_btm.n330 C10_N_btm.n329 0.09425
R25656 C10_N_btm.n329 C10_N_btm.n308 0.09425
R25657 C10_N_btm.n328 C10_N_btm.n307 0.09425
R25658 C10_N_btm.n822 C10_N_btm.n307 0.09425
R25659 C10_N_btm.n821 C10_N_btm.n308 0.09425
R25660 C10_N_btm.n821 C10_N_btm.n309 0.09425
R25661 C10_N_btm.n822 C10_N_btm.n304 0.09425
R25662 C10_N_btm.n304 C10_N_btm.n303 0.09425
R25663 C10_N_btm.n807 C10_N_btm.n309 0.09425
R25664 C10_N_btm.n807 C10_N_btm.n806 0.09425
R25665 C10_N_btm.n303 C10_N_btm.n302 0.09425
R25666 C10_N_btm.n302 C10_N_btm.n301 0.09425
R25667 C10_N_btm.n806 C10_N_btm.n805 0.09425
R25668 C10_N_btm.n805 C10_N_btm.n740 0.09425
R25669 C10_N_btm.n301 C10_N_btm.n300 0.09425
R25670 C10_N_btm.n300 C10_N_btm.n299 0.09425
R25671 C10_N_btm.n755 C10_N_btm.n740 0.09425
R25672 C10_N_btm.n760 C10_N_btm.n755 0.09425
R25673 C10_N_btm.n299 C10_N_btm.n298 0.09425
R25674 C10_N_btm.n298 C10_N_btm.n297 0.09425
R25675 C10_N_btm.n761 C10_N_btm.n760 0.09425
R25676 C10_N_btm.n792 C10_N_btm.n761 0.09425
R25677 C10_N_btm.n297 C10_N_btm.n296 0.09425
R25678 C10_N_btm.n296 C10_N_btm.n295 0.09425
R25679 C10_N_btm.n792 C10_N_btm.n791 0.09425
R25680 C10_N_btm.n791 C10_N_btm.n790 0.09425
R25681 C10_N_btm.n295 C10_N_btm.n294 0.09425
R25682 C10_N_btm.n294 C10_N_btm.n293 0.09425
R25683 C10_N_btm.n790 C10_N_btm.n789 0.09425
R25684 C10_N_btm.n789 C10_N_btm.n763 0.09425
R25685 C10_N_btm.n293 C10_N_btm.n292 0.09425
R25686 C10_N_btm.n292 C10_N_btm.n291 0.09425
R25687 C10_N_btm.n775 C10_N_btm.n763 0.09425
R25688 C10_N_btm.n775 C10_N_btm.n774 0.09425
R25689 C10_N_btm.n291 C10_N_btm.n290 0.09425
R25690 C10_N_btm.n290 C10_N_btm.n288 0.09425
R25691 C10_N_btm.n774 C10_N_btm.n287 0.09425
R25692 C10_N_btm.n843 C10_N_btm.n287 0.09425
R25693 C10_N_btm.n842 C10_N_btm.n288 0.09425
R25694 C10_N_btm.n842 C10_N_btm.n274 0.09425
R25695 C10_N_btm.n843 C10_N_btm.n275 0.09425
R25696 C10_N_btm.n860 C10_N_btm.n275 0.09425
R25697 C10_N_btm.n861 C10_N_btm.n274 0.09425
R25698 C10_N_btm.n861 C10_N_btm.n273 0.09425
R25699 C10_N_btm.n860 C10_N_btm.n859 0.09425
R25700 C10_N_btm.n859 C10_N_btm.n278 0.09425
R25701 C10_N_btm.n277 C10_N_btm.n273 0.09425
R25702 C10_N_btm.n277 C10_N_btm.n264 0.09425
R25703 C10_N_btm.n278 C10_N_btm.n263 0.09425
R25704 C10_N_btm.n870 C10_N_btm.n263 0.09425
R25705 C10_N_btm.n869 C10_N_btm.n264 0.09425
R25706 C10_N_btm.n869 C10_N_btm.n265 0.09425
R25707 C10_N_btm.n870 C10_N_btm.n261 0.09425
R25708 C10_N_btm.n261 C10_N_btm.n251 0.09425
R25709 C10_N_btm.n873 C10_N_btm.n259 0.09425
R25710 C10_N_btm.n873 C10_N_btm.n260 0.09425
R25711 C10_N_btm.n871 C10_N_btm.n262 0.09425
R25712 C10_N_btm.n872 C10_N_btm.n871 0.09425
R25713 C10_N_btm.n851 C10_N_btm.n281 0.09425
R25714 C10_N_btm.n851 C10_N_btm.n259 0.09425
R25715 C10_N_btm.n858 C10_N_btm.n279 0.09425
R25716 C10_N_btm.n279 C10_N_btm.n262 0.09425
R25717 C10_N_btm.n857 C10_N_btm.n280 0.09425
R25718 C10_N_btm.n857 C10_N_btm.n281 0.09425
R25719 C10_N_btm.n845 C10_N_btm.n276 0.09425
R25720 C10_N_btm.n858 C10_N_btm.n276 0.09425
R25721 C10_N_btm.n846 C10_N_btm.n285 0.09425
R25722 C10_N_btm.n846 C10_N_btm.n280 0.09425
R25723 C10_N_btm.n844 C10_N_btm.n286 0.09425
R25724 C10_N_btm.n845 C10_N_btm.n844 0.09425
R25725 C10_N_btm.n779 C10_N_btm.n778 0.09425
R25726 C10_N_btm.n779 C10_N_btm.n285 0.09425
R25727 C10_N_btm.n776 C10_N_btm.n773 0.09425
R25728 C10_N_btm.n773 C10_N_btm.n286 0.09425
R25729 C10_N_btm.n777 C10_N_btm.n766 0.09425
R25730 C10_N_btm.n778 C10_N_btm.n777 0.09425
R25731 C10_N_btm.n788 C10_N_btm.n764 0.09425
R25732 C10_N_btm.n776 C10_N_btm.n764 0.09425
R25733 C10_N_btm.n787 C10_N_btm.n765 0.09425
R25734 C10_N_btm.n787 C10_N_btm.n766 0.09425
R25735 C10_N_btm.n762 C10_N_btm.n754 0.09425
R25736 C10_N_btm.n788 C10_N_btm.n762 0.09425
R25737 C10_N_btm.n794 C10_N_btm.n752 0.09425
R25738 C10_N_btm.n765 C10_N_btm.n752 0.09425
R25739 C10_N_btm.n793 C10_N_btm.n753 0.09425
R25740 C10_N_btm.n793 C10_N_btm.n754 0.09425
R25741 C10_N_btm.n758 C10_N_btm.n750 0.09425
R25742 C10_N_btm.n794 C10_N_btm.n750 0.09425
R25743 C10_N_btm.n759 C10_N_btm.n756 0.09425
R25744 C10_N_btm.n759 C10_N_btm.n753 0.09425
R25745 C10_N_btm.n757 C10_N_btm.n742 0.09425
R25746 C10_N_btm.n758 C10_N_btm.n757 0.09425
R25747 C10_N_btm.n804 C10_N_btm.n741 0.09425
R25748 C10_N_btm.n756 C10_N_btm.n741 0.09425
R25749 C10_N_btm.n803 C10_N_btm.n738 0.09425
R25750 C10_N_btm.n803 C10_N_btm.n742 0.09425
R25751 C10_N_btm.n808 C10_N_btm.n739 0.09425
R25752 C10_N_btm.n804 C10_N_btm.n739 0.09425
R25753 C10_N_btm.n810 C10_N_btm.n809 0.09425
R25754 C10_N_btm.n809 C10_N_btm.n738 0.09425
R25755 C10_N_btm.n820 C10_N_btm.n310 0.09425
R25756 C10_N_btm.n808 C10_N_btm.n310 0.09425
R25757 C10_N_btm.n818 C10_N_btm.n311 0.09425
R25758 C10_N_btm.n810 C10_N_btm.n311 0.09425
R25759 C10_N_btm.n819 C10_N_btm.n312 0.09425
R25760 C10_N_btm.n820 C10_N_btm.n819 0.09425
R25761 C10_N_btm.n817 C10_N_btm.n314 0.09425
R25762 C10_N_btm.n818 C10_N_btm.n817 0.09425
R25763 C10_N_btm.n731 C10_N_btm.n319 0.09425
R25764 C10_N_btm.n319 C10_N_btm.n312 0.09425
R25765 C10_N_btm.n732 C10_N_btm.n318 0.09425
R25766 C10_N_btm.n732 C10_N_btm.n314 0.09425
R25767 C10_N_btm.n730 C10_N_btm.n321 0.09425
R25768 C10_N_btm.n731 C10_N_btm.n730 0.09425
R25769 C10_N_btm.n699 C10_N_btm.n693 0.09425
R25770 C10_N_btm.n693 C10_N_btm.n318 0.09425
R25771 C10_N_btm.n705 C10_N_btm.n700 0.09425
R25772 C10_N_btm.n700 C10_N_btm.n321 0.09425
R25773 C10_N_btm.n707 C10_N_btm.n706 0.09425
R25774 C10_N_btm.n706 C10_N_btm.n699 0.09425
R25775 C10_N_btm.n717 C10_N_btm.n344 0.09425
R25776 C10_N_btm.n705 C10_N_btm.n344 0.09425
R25777 C10_N_btm.n715 C10_N_btm.n345 0.09425
R25778 C10_N_btm.n707 C10_N_btm.n345 0.09425
R25779 C10_N_btm.n716 C10_N_btm.n346 0.09425
R25780 C10_N_btm.n717 C10_N_btm.n716 0.09425
R25781 C10_N_btm.n714 C10_N_btm.n348 0.09425
R25782 C10_N_btm.n715 C10_N_btm.n714 0.09425
R25783 C10_N_btm.n686 C10_N_btm.n353 0.09425
R25784 C10_N_btm.n353 C10_N_btm.n346 0.09425
R25785 C10_N_btm.n687 C10_N_btm.n352 0.09425
R25786 C10_N_btm.n687 C10_N_btm.n348 0.09425
R25787 C10_N_btm.n685 C10_N_btm.n355 0.09425
R25788 C10_N_btm.n686 C10_N_btm.n685 0.09425
R25789 C10_N_btm.n521 C10_N_btm.n467 0.09425
R25790 C10_N_btm.n521 C10_N_btm.n520 0.09425
R25791 C10_N_btm.n520 C10_N_btm.n352 0.09425
R25792 C10_N_btm.n522 C10_N_btm.n468 0.09425
R25793 C10_N_btm.n522 C10_N_btm.n355 0.09425
R25794 C10_N_btm.n591 C10_N_btm.n469 0.09425
R25795 C10_N_btm.n523 C10_N_btm.n469 0.09425
R25796 C10_N_btm.n593 C10_N_btm.n467 0.09425
R25797 C10_N_btm.n599 C10_N_btm.n463 0.09425
R25798 C10_N_btm.n593 C10_N_btm.n463 0.09425
R25799 C10_N_btm.n592 C10_N_btm.n462 0.09425
R25800 C10_N_btm.n592 C10_N_btm.n468 0.09425
R25801 C10_N_btm.n601 C10_N_btm.n460 0.09425
R25802 C10_N_btm.n591 C10_N_btm.n460 0.09425
R25803 C10_N_btm.n590 C10_N_btm.n459 0.09425
R25804 C10_N_btm.n590 C10_N_btm.n470 0.09425
R25805 C10_N_btm.n588 C10_N_btm.n457 0.09425
R25806 C10_N_btm.n589 C10_N_btm.n588 0.09425
R25807 C10_N_btm.n587 C10_N_btm.n586 0.09425
R25808 C10_N_btm.n586 C10_N_btm.n472 0.09425
R25809 C10_N_btm.n607 C10_N_btm.n455 0.09425
R25810 C10_N_btm.n585 C10_N_btm.n455 0.09425
R25811 C10_N_btm.n584 C10_N_btm.n454 0.09425
R25812 C10_N_btm.n584 C10_N_btm.n474 0.09425
R25813 C10_N_btm.n609 C10_N_btm.n452 0.09425
R25814 C10_N_btm.n583 C10_N_btm.n452 0.09425
R25815 C10_N_btm.n582 C10_N_btm.n451 0.09425
R25816 C10_N_btm.n582 C10_N_btm.n476 0.09425
R25817 C10_N_btm.n580 C10_N_btm.n449 0.09425
R25818 C10_N_btm.n581 C10_N_btm.n580 0.09425
R25819 C10_N_btm.n579 C10_N_btm.n578 0.09425
R25820 C10_N_btm.n578 C10_N_btm.n478 0.09425
R25821 C10_N_btm.n615 C10_N_btm.n447 0.09425
R25822 C10_N_btm.n577 C10_N_btm.n447 0.09425
R25823 C10_N_btm.n576 C10_N_btm.n446 0.09425
R25824 C10_N_btm.n576 C10_N_btm.n480 0.09425
R25825 C10_N_btm.n617 C10_N_btm.n444 0.09425
R25826 C10_N_btm.n575 C10_N_btm.n444 0.09425
R25827 C10_N_btm.n574 C10_N_btm.n443 0.09425
R25828 C10_N_btm.n574 C10_N_btm.n482 0.09425
R25829 C10_N_btm.n572 C10_N_btm.n441 0.09425
R25830 C10_N_btm.n573 C10_N_btm.n572 0.09425
R25831 C10_N_btm.n571 C10_N_btm.n570 0.09425
R25832 C10_N_btm.n570 C10_N_btm.n484 0.09425
R25833 C10_N_btm.n623 C10_N_btm.n439 0.09425
R25834 C10_N_btm.n569 C10_N_btm.n439 0.09425
R25835 C10_N_btm.n568 C10_N_btm.n438 0.09425
R25836 C10_N_btm.n568 C10_N_btm.n486 0.09425
R25837 C10_N_btm.n625 C10_N_btm.n436 0.09425
R25838 C10_N_btm.n567 C10_N_btm.n436 0.09425
R25839 C10_N_btm.n566 C10_N_btm.n435 0.09425
R25840 C10_N_btm.n566 C10_N_btm.n488 0.09425
R25841 C10_N_btm.n564 C10_N_btm.n433 0.09425
R25842 C10_N_btm.n565 C10_N_btm.n564 0.09425
R25843 C10_N_btm.n563 C10_N_btm.n562 0.09425
R25844 C10_N_btm.n562 C10_N_btm.n490 0.09425
R25845 C10_N_btm.n631 C10_N_btm.n423 0.09425
R25846 C10_N_btm.n561 C10_N_btm.n423 0.09425
R25847 C10_N_btm.n633 C10_N_btm.n421 0.09425
R25848 C10_N_btm.n491 C10_N_btm.n421 0.09425
R25849 C10_N_btm.n634 C10_N_btm.n422 0.09425
R25850 C10_N_btm.n635 C10_N_btm.n634 0.09425
R25851 C10_N_btm.n636 C10_N_btm.n420 0.09425
R25852 C10_N_btm.n637 C10_N_btm.n636 0.09425
R25853 C10_N_btm.n427 C10_N_btm.n426 0.09425
R25854 C10_N_btm.n426 C10_N_btm.n417 0.09425
R25855 C10_N_btm.n429 C10_N_btm.n428 0.09425
R25856 C10_N_btm.n428 C10_N_btm.n420 0.09425
R25857 C10_N_btm.n430 C10_N_btm.n422 0.09425
R25858 C10_N_btm.n632 C10_N_btm.n431 0.09425
R25859 C10_N_btm.n633 C10_N_btm.n632 0.09425
R25860 C10_N_btm.n631 C10_N_btm.n630 0.09425
R25861 C10_N_btm.n629 C10_N_btm.n432 0.09425
R25862 C10_N_btm.n563 C10_N_btm.n432 0.09425
R25863 C10_N_btm.n628 C10_N_btm.n433 0.09425
R25864 C10_N_btm.n627 C10_N_btm.n626 0.09425
R25865 C10_N_btm.n626 C10_N_btm.n435 0.09425
R25866 C10_N_btm.n625 C10_N_btm.n434 0.09425
R25867 C10_N_btm.n624 C10_N_btm.n437 0.09425
R25868 C10_N_btm.n624 C10_N_btm.n438 0.09425
R25869 C10_N_btm.n623 C10_N_btm.n622 0.09425
R25870 C10_N_btm.n621 C10_N_btm.n440 0.09425
R25871 C10_N_btm.n571 C10_N_btm.n440 0.09425
R25872 C10_N_btm.n620 C10_N_btm.n441 0.09425
R25873 C10_N_btm.n619 C10_N_btm.n618 0.09425
R25874 C10_N_btm.n618 C10_N_btm.n443 0.09425
R25875 C10_N_btm.n617 C10_N_btm.n442 0.09425
R25876 C10_N_btm.n616 C10_N_btm.n445 0.09425
R25877 C10_N_btm.n616 C10_N_btm.n446 0.09425
R25878 C10_N_btm.n615 C10_N_btm.n614 0.09425
R25879 C10_N_btm.n613 C10_N_btm.n448 0.09425
R25880 C10_N_btm.n579 C10_N_btm.n448 0.09425
R25881 C10_N_btm.n612 C10_N_btm.n449 0.09425
R25882 C10_N_btm.n611 C10_N_btm.n610 0.09425
R25883 C10_N_btm.n610 C10_N_btm.n451 0.09425
R25884 C10_N_btm.n609 C10_N_btm.n450 0.09425
R25885 C10_N_btm.n608 C10_N_btm.n453 0.09425
R25886 C10_N_btm.n608 C10_N_btm.n454 0.09425
R25887 C10_N_btm.n607 C10_N_btm.n606 0.09425
R25888 C10_N_btm.n605 C10_N_btm.n456 0.09425
R25889 C10_N_btm.n587 C10_N_btm.n456 0.09425
R25890 C10_N_btm.n604 C10_N_btm.n457 0.09425
R25891 C10_N_btm.n603 C10_N_btm.n602 0.09425
R25892 C10_N_btm.n602 C10_N_btm.n459 0.09425
R25893 C10_N_btm.n601 C10_N_btm.n458 0.09425
R25894 C10_N_btm.n600 C10_N_btm.n461 0.09425
R25895 C10_N_btm.n600 C10_N_btm.n462 0.09425
R25896 C10_N_btm.n599 C10_N_btm.n598 0.09425
R25897 C10_N_btm.n595 C10_N_btm.n464 0.09425
R25898 C10_N_btm.n596 C10_N_btm.n465 0.09425
R25899 C10_N_btm.n595 C10_N_btm.n594 0.09425
R25900 C10_N_btm.n594 C10_N_btm.n466 0.09425
R25901 C10_N_btm.n516 C10_N_btm.n465 0.09425
R25902 C10_N_btm.n517 C10_N_btm.n516 0.09425
R25903 C10_N_btm.n515 C10_N_btm.n466 0.09425
R25904 C10_N_btm.n519 C10_N_btm.n515 0.09425
R25905 C10_N_btm.n518 C10_N_btm.n517 0.09425
R25906 C10_N_btm.n518 C10_N_btm.n350 0.09425
R25907 C10_N_btm.n519 C10_N_btm.n351 0.09425
R25908 C10_N_btm.n688 C10_N_btm.n351 0.09425
R25909 C10_N_btm.n689 C10_N_btm.n350 0.09425
R25910 C10_N_btm.n690 C10_N_btm.n689 0.09425
R25911 C10_N_btm.n688 C10_N_btm.n349 0.09425
R25912 C10_N_btm.n713 C10_N_btm.n349 0.09425
R25913 C10_N_btm.n712 C10_N_btm.n690 0.09425
R25914 C10_N_btm.n712 C10_N_btm.n711 0.09425
R25915 C10_N_btm.n713 C10_N_btm.n347 0.09425
R25916 C10_N_btm.n709 C10_N_btm.n347 0.09425
R25917 C10_N_btm.n711 C10_N_btm.n710 0.09425
R25918 C10_N_btm.n710 C10_N_btm.n691 0.09425
R25919 C10_N_btm.n709 C10_N_btm.n708 0.09425
R25920 C10_N_btm.n708 C10_N_btm.n692 0.09425
R25921 C10_N_btm.n695 C10_N_btm.n691 0.09425
R25922 C10_N_btm.n697 C10_N_btm.n695 0.09425
R25923 C10_N_btm.n698 C10_N_btm.n692 0.09425
R25924 C10_N_btm.n698 C10_N_btm.n694 0.09425
R25925 C10_N_btm.n697 C10_N_btm.n696 0.09425
R25926 C10_N_btm.n696 C10_N_btm.n316 0.09425
R25927 C10_N_btm.n694 C10_N_btm.n317 0.09425
R25928 C10_N_btm.n733 C10_N_btm.n317 0.09425
R25929 C10_N_btm.n734 C10_N_btm.n316 0.09425
R25930 C10_N_btm.n735 C10_N_btm.n734 0.09425
R25931 C10_N_btm.n733 C10_N_btm.n315 0.09425
R25932 C10_N_btm.n816 C10_N_btm.n315 0.09425
R25933 C10_N_btm.n815 C10_N_btm.n735 0.09425
R25934 C10_N_btm.n815 C10_N_btm.n814 0.09425
R25935 C10_N_btm.n816 C10_N_btm.n313 0.09425
R25936 C10_N_btm.n812 C10_N_btm.n313 0.09425
R25937 C10_N_btm.n814 C10_N_btm.n813 0.09425
R25938 C10_N_btm.n813 C10_N_btm.n736 0.09425
R25939 C10_N_btm.n812 C10_N_btm.n811 0.09425
R25940 C10_N_btm.n811 C10_N_btm.n737 0.09425
R25941 C10_N_btm.n744 C10_N_btm.n736 0.09425
R25942 C10_N_btm.n745 C10_N_btm.n744 0.09425
R25943 C10_N_btm.n743 C10_N_btm.n737 0.09425
R25944 C10_N_btm.n802 C10_N_btm.n743 0.09425
R25945 C10_N_btm.n746 C10_N_btm.n745 0.09425
R25946 C10_N_btm.n800 C10_N_btm.n746 0.09425
R25947 C10_N_btm.n802 C10_N_btm.n801 0.09425
R25948 C10_N_btm.n801 C10_N_btm.n747 0.09425
R25949 C10_N_btm.n800 C10_N_btm.n799 0.09425
R25950 C10_N_btm.n799 C10_N_btm.n798 0.09425
R25951 C10_N_btm.n748 C10_N_btm.n747 0.09425
R25952 C10_N_btm.n796 C10_N_btm.n748 0.09425
R25953 C10_N_btm.n798 C10_N_btm.n797 0.09425
R25954 C10_N_btm.n797 C10_N_btm.n749 0.09425
R25955 C10_N_btm.n796 C10_N_btm.n795 0.09425
R25956 C10_N_btm.n795 C10_N_btm.n751 0.09425
R25957 C10_N_btm.n768 C10_N_btm.n749 0.09425
R25958 C10_N_btm.n769 C10_N_btm.n768 0.09425
R25959 C10_N_btm.n767 C10_N_btm.n751 0.09425
R25960 C10_N_btm.n786 C10_N_btm.n767 0.09425
R25961 C10_N_btm.n770 C10_N_btm.n769 0.09425
R25962 C10_N_btm.n784 C10_N_btm.n770 0.09425
R25963 C10_N_btm.n786 C10_N_btm.n785 0.09425
R25964 C10_N_btm.n785 C10_N_btm.n771 0.09425
R25965 C10_N_btm.n784 C10_N_btm.n783 0.09425
R25966 C10_N_btm.n783 C10_N_btm.n782 0.09425
R25967 C10_N_btm.n772 C10_N_btm.n771 0.09425
R25968 C10_N_btm.n780 C10_N_btm.n772 0.09425
R25969 C10_N_btm.n782 C10_N_btm.n781 0.09425
R25970 C10_N_btm.n781 C10_N_btm.n283 0.09425
R25971 C10_N_btm.n780 C10_N_btm.n284 0.09425
R25972 C10_N_btm.n847 C10_N_btm.n284 0.09425
R25973 C10_N_btm.n848 C10_N_btm.n283 0.09425
R25974 C10_N_btm.n849 C10_N_btm.n848 0.09425
R25975 C10_N_btm.n847 C10_N_btm.n282 0.09425
R25976 C10_N_btm.n856 C10_N_btm.n282 0.09425
R25977 C10_N_btm.n850 C10_N_btm.n849 0.09425
R25978 C10_N_btm.n854 C10_N_btm.n850 0.09425
R25979 C10_N_btm.n856 C10_N_btm.n855 0.09425
R25980 C10_N_btm.n855 C10_N_btm.n852 0.09425
R25981 C10_N_btm.n854 C10_N_btm.n853 0.09425
R25982 C10_N_btm.n853 C10_N_btm.n257 0.09425
R25983 C10_N_btm.n852 C10_N_btm.n258 0.09425
R25984 C10_N_btm.n874 C10_N_btm.n258 0.09425
R25985 C10_N_btm.n875 C10_N_btm.n257 0.09425
R25986 C10_N_btm.n876 C10_N_btm.n875 0.09425
R25987 C10_N_btm.n874 C10_N_btm.n256 0.09425
R25988 C10_N_btm.n256 C10_N_btm.n254 0.09425
R25989 C10_N_btm.n260 C10_N_btm.n253 0.09425
R25990 C10_N_btm.n880 C10_N_btm.n253 0.09425
R25991 C10_N_btm.n882 C10_N_btm.n881 0.09425
R25992 C10_N_btm.n881 C10_N_btm.n242 0.09425
R25993 C10_N_btm.n249 C10_N_btm.n248 0.09425
R25994 C10_N_btm.n248 C10_N_btm.n243 0.09425
R25995 C10_N_btm.n891 C10_N_btm.n244 0.09425
R25996 C10_N_btm.n892 C10_N_btm.n891 0.09425
R25997 C10_N_btm.n890 C10_N_btm.n68 0.09425
R25998 C10_N_btm.n1011 C10_N_btm.n68 0.09425
R25999 C10_N_btm.n1012 C10_N_btm.n65 0.09425
R26000 C10_N_btm.n1012 C10_N_btm.n66 0.09425
R26001 C10_N_btm.n1013 C10_N_btm.n64 0.09425
R26002 C10_N_btm.n72 C10_N_btm.n64 0.09425
R26003 C10_N_btm.n1015 C10_N_btm.n1014 0.09425
R26004 C10_N_btm.n1016 C10_N_btm.n61 0.09425
R26005 C10_N_btm.n1016 C10_N_btm.n62 0.09425
R26006 C10_N_btm.n1017 C10_N_btm.n58 0.09425
R26007 C10_N_btm.n1019 C10_N_btm.n1018 0.09425
R26008 C10_N_btm.n1018 C10_N_btm.n59 0.09425
R26009 C10_N_btm.n1020 C10_N_btm.n57 0.09425
R26010 C10_N_btm.n1021 C10_N_btm.n56 0.09425
R26011 C10_N_btm.n86 C10_N_btm.n56 0.09425
R26012 C10_N_btm.n1023 C10_N_btm.n1022 0.09425
R26013 C10_N_btm.n1024 C10_N_btm.n53 0.09425
R26014 C10_N_btm.n1024 C10_N_btm.n54 0.09425
R26015 C10_N_btm.n1025 C10_N_btm.n50 0.09425
R26016 C10_N_btm.n1027 C10_N_btm.n1026 0.09425
R26017 C10_N_btm.n1026 C10_N_btm.n51 0.09425
R26018 C10_N_btm.n1028 C10_N_btm.n49 0.09425
R26019 C10_N_btm.n1029 C10_N_btm.n48 0.09425
R26020 C10_N_btm.n104 C10_N_btm.n48 0.09425
R26021 C10_N_btm.n1031 C10_N_btm.n1030 0.09425
R26022 C10_N_btm.n1032 C10_N_btm.n45 0.09425
R26023 C10_N_btm.n1032 C10_N_btm.n46 0.09425
R26024 C10_N_btm.n1033 C10_N_btm.n42 0.09425
R26025 C10_N_btm.n1035 C10_N_btm.n1034 0.09425
R26026 C10_N_btm.n1034 C10_N_btm.n43 0.09425
R26027 C10_N_btm.n1036 C10_N_btm.n41 0.09425
R26028 C10_N_btm.n1037 C10_N_btm.n40 0.09425
R26029 C10_N_btm.n117 C10_N_btm.n40 0.09425
R26030 C10_N_btm.n1039 C10_N_btm.n1038 0.09425
R26031 C10_N_btm.n1040 C10_N_btm.n37 0.09425
R26032 C10_N_btm.n1040 C10_N_btm.n38 0.09425
R26033 C10_N_btm.n1041 C10_N_btm.n34 0.09425
R26034 C10_N_btm.n1043 C10_N_btm.n1042 0.09425
R26035 C10_N_btm.n1042 C10_N_btm.n35 0.09425
R26036 C10_N_btm.n1044 C10_N_btm.n33 0.09425
R26037 C10_N_btm.n289 C10_N_btm.n272 0.047875
R26038 C10_N_btm.n825 C10_N_btm.n824 0.047875
R26039 C10_N_btm.n181 C10_N_btm.n133 0.0342289
R26040 C10_N_btm.n217 C10_N_btm.n180 0.0342289
R26041 C10_N_btm.n646 C10_N_btm.n645 0.0342289
R26042 C10_N_btm.n862 C10_N_btm.n272 0.0342289
R26043 C10_N_btm.n824 C10_N_btm.n823 0.0342289
R26044 C10_N_btm.n427 C10_N_btm.n424 0.0342289
R26045 C10_N_btm.n597 C10_N_btm.n464 0.0342289
R26046 VCM VCM.n59 62.1408
R26047 VCM VCM.n29 61.9779
R26048 VCM.n0 VCM.t22 47.8989
R26049 VCM.n31 VCM.t23 47.8989
R26050 VCM.n0 VCM.t61 47.4614
R26051 VCM.n1 VCM.t19 47.4614
R26052 VCM.n2 VCM.t0 47.4614
R26053 VCM.n3 VCM.t20 47.4614
R26054 VCM.n4 VCM.t43 47.4614
R26055 VCM.n7 VCM.t27 47.4614
R26056 VCM.n38 VCM.t26 47.4614
R26057 VCM.n35 VCM.t42 47.4614
R26058 VCM.n34 VCM.t21 47.4614
R26059 VCM.n33 VCM.t1 47.4614
R26060 VCM.n32 VCM.t18 47.4614
R26061 VCM.n31 VCM.t60 47.4614
R26062 VCM.n6 VCM.n5 37.5614
R26063 VCM.n37 VCM.n36 37.5614
R26064 VCM.n29 VCM.t54 17.4125
R26065 VCM.n59 VCM.t53 17.4125
R26066 VCM.n10 VCM.n8 15.4323
R26067 VCM.n40 VCM.n30 15.4323
R26068 VCM.n28 VCM.n27 14.9375
R26069 VCM.n26 VCM.n25 14.9375
R26070 VCM.n24 VCM.n23 14.9375
R26071 VCM.n22 VCM.n21 14.9375
R26072 VCM.n20 VCM.n19 14.9375
R26073 VCM.n18 VCM.n17 14.9375
R26074 VCM.n16 VCM.n15 14.9375
R26075 VCM.n14 VCM.n13 14.9375
R26076 VCM.n12 VCM.n11 14.9375
R26077 VCM.n10 VCM.n9 14.9375
R26078 VCM.n58 VCM.n57 14.9375
R26079 VCM.n56 VCM.n55 14.9375
R26080 VCM.n54 VCM.n53 14.9375
R26081 VCM.n52 VCM.n51 14.9375
R26082 VCM.n50 VCM.n49 14.9375
R26083 VCM.n48 VCM.n47 14.9375
R26084 VCM.n46 VCM.n45 14.9375
R26085 VCM.n44 VCM.n43 14.9375
R26086 VCM.n42 VCM.n41 14.9375
R26087 VCM.n40 VCM.n39 14.9375
R26088 VCM.n5 VCM.t25 9.9005
R26089 VCM.n5 VCM.t62 9.9005
R26090 VCM.n36 VCM.t63 9.9005
R26091 VCM.n36 VCM.t24 9.9005
R26092 VCM.n10 VCM.n7 8.35002
R26093 VCM.n40 VCM.n38 8.35002
R26094 VCM.n27 VCM.t50 2.4755
R26095 VCM.n27 VCM.t51 2.4755
R26096 VCM.n25 VCM.t59 2.4755
R26097 VCM.n25 VCM.t45 2.4755
R26098 VCM.n23 VCM.t46 2.4755
R26099 VCM.n23 VCM.t52 2.4755
R26100 VCM.n21 VCM.t47 2.4755
R26101 VCM.n21 VCM.t8 2.4755
R26102 VCM.n19 VCM.t5 2.4755
R26103 VCM.n19 VCM.t4 2.4755
R26104 VCM.n17 VCM.t7 2.4755
R26105 VCM.n17 VCM.t2 2.4755
R26106 VCM.n15 VCM.t6 2.4755
R26107 VCM.n15 VCM.t3 2.4755
R26108 VCM.n13 VCM.t9 2.4755
R26109 VCM.n13 VCM.t38 2.4755
R26110 VCM.n11 VCM.t32 2.4755
R26111 VCM.n11 VCM.t39 2.4755
R26112 VCM.n9 VCM.t33 2.4755
R26113 VCM.n9 VCM.t29 2.4755
R26114 VCM.n8 VCM.t28 2.4755
R26115 VCM.n8 VCM.t41 2.4755
R26116 VCM.n57 VCM.t49 2.4755
R26117 VCM.n57 VCM.t48 2.4755
R26118 VCM.n55 VCM.t44 2.4755
R26119 VCM.n55 VCM.t56 2.4755
R26120 VCM.n53 VCM.t55 2.4755
R26121 VCM.n53 VCM.t57 2.4755
R26122 VCM.n51 VCM.t16 2.4755
R26123 VCM.n51 VCM.t58 2.4755
R26124 VCM.n49 VCM.t14 2.4755
R26125 VCM.n49 VCM.t17 2.4755
R26126 VCM.n47 VCM.t13 2.4755
R26127 VCM.n47 VCM.t11 2.4755
R26128 VCM.n45 VCM.t12 2.4755
R26129 VCM.n45 VCM.t10 2.4755
R26130 VCM.n43 VCM.t35 2.4755
R26131 VCM.n43 VCM.t15 2.4755
R26132 VCM.n41 VCM.t37 2.4755
R26133 VCM.n41 VCM.t34 2.4755
R26134 VCM.n39 VCM.t30 2.4755
R26135 VCM.n39 VCM.t36 2.4755
R26136 VCM.n30 VCM.t40 2.4755
R26137 VCM.n30 VCM.t31 2.4755
R26138 VCM.n16 VCM.n14 0.53175
R26139 VCM.n24 VCM.n22 0.53175
R26140 VCM.n46 VCM.n44 0.53175
R26141 VCM.n54 VCM.n52 0.53175
R26142 VCM.n14 VCM.n12 0.5005
R26143 VCM.n18 VCM.n16 0.5005
R26144 VCM.n20 VCM.n18 0.5005
R26145 VCM.n22 VCM.n20 0.5005
R26146 VCM.n26 VCM.n24 0.5005
R26147 VCM.n28 VCM.n26 0.5005
R26148 VCM.n29 VCM.n28 0.5005
R26149 VCM.n44 VCM.n42 0.5005
R26150 VCM.n48 VCM.n46 0.5005
R26151 VCM.n50 VCM.n48 0.5005
R26152 VCM.n52 VCM.n50 0.5005
R26153 VCM.n56 VCM.n54 0.5005
R26154 VCM.n58 VCM.n56 0.5005
R26155 VCM.n59 VCM.n58 0.5005
R26156 VCM.n12 VCM.n10 0.495292
R26157 VCM.n42 VCM.n40 0.495292
R26158 VCM.n6 VCM.n4 0.438
R26159 VCM.n4 VCM.n3 0.438
R26160 VCM.n3 VCM.n2 0.438
R26161 VCM.n2 VCM.n1 0.438
R26162 VCM.n1 VCM.n0 0.438
R26163 VCM.n32 VCM.n31 0.438
R26164 VCM.n33 VCM.n32 0.438
R26165 VCM.n34 VCM.n33 0.438
R26166 VCM.n35 VCM.n34 0.438
R26167 VCM.n37 VCM.n35 0.438
R26168 VCM.n7 VCM.n6 0.396333
R26169 VCM.n38 VCM.n37 0.396333
R26170 a_11967_42832.n46 a_11967_42832.n45 333.392
R26171 a_11967_42832.n35 a_11967_42832.n34 301.392
R26172 a_11967_42832.n37 a_11967_42832.n36 301.392
R26173 a_11967_42832.n39 a_11967_42832.n38 301.392
R26174 a_11967_42832.n41 a_11967_42832.n40 301.392
R26175 a_11967_42832.n43 a_11967_42832.n42 301.392
R26176 a_11967_42832.n45 a_11967_42832.n44 301.392
R26177 a_11967_42832.n33 a_11967_42832.n32 297.808
R26178 a_11967_42832.n19 a_11967_42832.t41 294.557
R26179 a_11967_42832.n17 a_11967_42832.t40 294.557
R26180 a_11967_42832.n27 a_11967_42832.t45 294.557
R26181 a_11967_42832.n22 a_11967_42832.t44 294.557
R26182 a_11967_42832.n23 a_11967_42832.t38 294.557
R26183 a_11967_42832.n24 a_11967_42832.t43 294.557
R26184 a_11967_42832.n21 a_11967_42832.t32 294.557
R26185 a_11967_42832.n2 a_11967_42832.n0 248.638
R26186 a_11967_42832.n15 a_11967_42832.t33 212.081
R26187 a_11967_42832.n16 a_11967_42832.t47 212.081
R26188 a_11967_42832.n19 a_11967_42832.t34 211.01
R26189 a_11967_42832.n17 a_11967_42832.t46 211.01
R26190 a_11967_42832.n27 a_11967_42832.t35 211.01
R26191 a_11967_42832.n22 a_11967_42832.t37 211.01
R26192 a_11967_42832.n23 a_11967_42832.t42 211.01
R26193 a_11967_42832.n24 a_11967_42832.t49 211.01
R26194 a_11967_42832.n21 a_11967_42832.t36 211.01
R26195 a_11967_42832.n2 a_11967_42832.n1 203.463
R26196 a_11967_42832.n4 a_11967_42832.n3 203.463
R26197 a_11967_42832.n8 a_11967_42832.n7 203.463
R26198 a_11967_42832.n10 a_11967_42832.n9 203.463
R26199 a_11967_42832.n12 a_11967_42832.n11 203.463
R26200 a_11967_42832.n6 a_11967_42832.n5 202.456
R26201 a_11967_42832.n14 a_11967_42832.n13 200.212
R26202 a_11967_42832.n18 a_11967_42832.n16 194.331
R26203 a_11967_42832.n28 a_11967_42832.n27 187.893
R26204 a_11967_42832.n20 a_11967_42832.n19 174.832
R26205 a_11967_42832.n26 a_11967_42832.n22 172.784
R26206 a_11967_42832.n25 a_11967_42832.n24 163.94
R26207 a_11967_42832.n29 a_11967_42832.n21 162.585
R26208 a_11967_42832.n18 a_11967_42832.n17 162.398
R26209 a_11967_42832.n25 a_11967_42832.n23 162.398
R26210 a_11967_42832.n15 a_11967_42832.t39 139.78
R26211 a_11967_42832.n16 a_11967_42832.t48 139.78
R26212 a_11967_42832.n16 a_11967_42832.n15 61.346
R26213 a_11967_42832.n4 a_11967_42832.n2 45.177
R26214 a_11967_42832.n10 a_11967_42832.n8 45.177
R26215 a_11967_42832.n12 a_11967_42832.n10 45.177
R26216 a_11967_42832.n6 a_11967_42832.n4 44.0476
R26217 a_11967_42832.n8 a_11967_42832.n6 44.0476
R26218 a_11967_42832.n0 a_11967_42832.t26 40.0005
R26219 a_11967_42832.n0 a_11967_42832.t19 40.0005
R26220 a_11967_42832.n1 a_11967_42832.t21 40.0005
R26221 a_11967_42832.n1 a_11967_42832.t28 40.0005
R26222 a_11967_42832.n3 a_11967_42832.t17 40.0005
R26223 a_11967_42832.n3 a_11967_42832.t23 40.0005
R26224 a_11967_42832.n5 a_11967_42832.t27 40.0005
R26225 a_11967_42832.n5 a_11967_42832.t22 40.0005
R26226 a_11967_42832.n7 a_11967_42832.t20 40.0005
R26227 a_11967_42832.n7 a_11967_42832.t29 40.0005
R26228 a_11967_42832.n9 a_11967_42832.t24 40.0005
R26229 a_11967_42832.n9 a_11967_42832.t25 40.0005
R26230 a_11967_42832.n11 a_11967_42832.t30 40.0005
R26231 a_11967_42832.n11 a_11967_42832.t18 40.0005
R26232 a_11967_42832.n13 a_11967_42832.t31 40.0005
R26233 a_11967_42832.n13 a_11967_42832.t16 40.0005
R26234 a_11967_42832.n37 a_11967_42832.n35 32.0005
R26235 a_11967_42832.n39 a_11967_42832.n37 32.0005
R26236 a_11967_42832.n43 a_11967_42832.n41 32.0005
R26237 a_11967_42832.n45 a_11967_42832.n43 32.0005
R26238 a_11967_42832.n41 a_11967_42832.n39 31.2005
R26239 a_11967_42832.n34 a_11967_42832.t7 27.5805
R26240 a_11967_42832.n34 a_11967_42832.t6 27.5805
R26241 a_11967_42832.n32 a_11967_42832.t5 27.5805
R26242 a_11967_42832.n32 a_11967_42832.t10 27.5805
R26243 a_11967_42832.n36 a_11967_42832.t2 27.5805
R26244 a_11967_42832.n36 a_11967_42832.t0 27.5805
R26245 a_11967_42832.n38 a_11967_42832.t3 27.5805
R26246 a_11967_42832.n38 a_11967_42832.t14 27.5805
R26247 a_11967_42832.n40 a_11967_42832.t11 27.5805
R26248 a_11967_42832.n40 a_11967_42832.t1 27.5805
R26249 a_11967_42832.n42 a_11967_42832.t4 27.5805
R26250 a_11967_42832.n42 a_11967_42832.t12 27.5805
R26251 a_11967_42832.n44 a_11967_42832.t8 27.5805
R26252 a_11967_42832.n44 a_11967_42832.t9 27.5805
R26253 a_11967_42832.n46 a_11967_42832.t13 27.5805
R26254 a_11967_42832.t15 a_11967_42832.n46 27.5805
R26255 a_11967_42832.n31 a_11967_42832.n30 19.2018
R26256 a_11967_42832.n26 a_11967_42832.n25 17.6265
R26257 a_11967_42832.n14 a_11967_42832.n12 13.177
R26258 a_11967_42832.n30 a_11967_42832.n29 11.1063
R26259 a_11967_42832.n20 a_11967_42832.n18 10.7668
R26260 a_11967_42832.n30 a_11967_42832.n20 10.5913
R26261 a_11967_42832.n35 a_11967_42832.n33 10.2022
R26262 a_11967_42832.n33 a_11967_42832.n31 8.35071
R26263 a_11967_42832.n28 a_11967_42832.n26 4.98814
R26264 a_11967_42832.n29 a_11967_42832.n28 3.22028
R26265 a_11967_42832.n31 a_11967_42832.n14 0.330114
R26266 a_n4209_39590.n4 a_n4209_39590.t8 756.547
R26267 a_n4209_39590.n10 a_n4209_39590.t11 756.231
R26268 a_n4209_39590.n9 a_n4209_39590.t15 756.226
R26269 a_n4209_39590.n8 a_n4209_39590.t13 756.226
R26270 a_n4209_39590.n7 a_n4209_39590.t12 756.226
R26271 a_n4209_39590.n6 a_n4209_39590.t17 756.226
R26272 a_n4209_39590.n5 a_n4209_39590.t9 756.226
R26273 a_n4209_39590.n4 a_n4209_39590.t16 756.226
R26274 a_n4209_39590.n15 a_n4209_39590.n14 340.637
R26275 a_n4209_39590.n3 a_n4209_39590.t14 241.536
R26276 a_n4209_39590.n14 a_n4209_39590.n13 195.577
R26277 a_n4209_39590.n11 a_n4209_39590.n3 173.952
R26278 a_n4209_39590.n3 a_n4209_39590.t10 169.237
R26279 a_n4209_39590.n2 a_n4209_39590.n0 137.189
R26280 a_n4209_39590.n2 a_n4209_39590.n1 98.788
R26281 a_n4209_39590.n11 a_n4209_39590.n10 69.0005
R26282 a_n4209_39590.n14 a_n4209_39590.n12 37.1695
R26283 a_n4209_39590.n12 a_n4209_39590.n2 27.8375
R26284 a_n4209_39590.n13 a_n4209_39590.t2 26.5955
R26285 a_n4209_39590.n13 a_n4209_39590.t0 26.5955
R26286 a_n4209_39590.n15 a_n4209_39590.t1 26.5955
R26287 a_n4209_39590.t3 a_n4209_39590.n15 26.5955
R26288 a_n4209_39590.n0 a_n4209_39590.t7 24.9236
R26289 a_n4209_39590.n0 a_n4209_39590.t6 24.9236
R26290 a_n4209_39590.n1 a_n4209_39590.t5 24.9236
R26291 a_n4209_39590.n1 a_n4209_39590.t4 24.9236
R26292 a_n4209_39590.n12 a_n4209_39590.n11 9.30997
R26293 a_n4209_39590.n5 a_n4209_39590.n4 0.3205
R26294 a_n4209_39590.n6 a_n4209_39590.n5 0.3205
R26295 a_n4209_39590.n7 a_n4209_39590.n6 0.3205
R26296 a_n4209_39590.n8 a_n4209_39590.n7 0.3205
R26297 a_n4209_39590.n9 a_n4209_39590.n8 0.3205
R26298 a_n4209_39590.n10 a_n4209_39590.n9 0.298833
R26299 a_11599_46634.n2 a_11599_46634.n0 333.392
R26300 a_11599_46634.n39 a_11599_46634.n38 301.392
R26301 a_11599_46634.n41 a_11599_46634.n40 301.392
R26302 a_11599_46634.n43 a_11599_46634.n42 301.392
R26303 a_11599_46634.n45 a_11599_46634.n44 301.392
R26304 a_11599_46634.n2 a_11599_46634.n1 301.392
R26305 a_11599_46634.n47 a_11599_46634.n46 301.392
R26306 a_11599_46634.n35 a_11599_46634.n34 296.8
R26307 a_11599_46634.n25 a_11599_46634.t40 294.557
R26308 a_11599_46634.n26 a_11599_46634.t45 294.557
R26309 a_11599_46634.n24 a_11599_46634.t37 294.557
R26310 a_11599_46634.n29 a_11599_46634.t42 294.557
R26311 a_11599_46634.n30 a_11599_46634.t48 294.557
R26312 a_11599_46634.n18 a_11599_46634.t34 294.557
R26313 a_11599_46634.n19 a_11599_46634.t47 294.557
R26314 a_11599_46634.n20 a_11599_46634.t36 294.557
R26315 a_11599_46634.n17 a_11599_46634.t35 294.557
R26316 a_11599_46634.n5 a_11599_46634.n3 248.638
R26317 a_11599_46634.n25 a_11599_46634.t46 211.01
R26318 a_11599_46634.n26 a_11599_46634.t44 211.01
R26319 a_11599_46634.n24 a_11599_46634.t39 211.01
R26320 a_11599_46634.n29 a_11599_46634.t38 211.01
R26321 a_11599_46634.n30 a_11599_46634.t33 211.01
R26322 a_11599_46634.n18 a_11599_46634.t49 211.01
R26323 a_11599_46634.n19 a_11599_46634.t43 211.01
R26324 a_11599_46634.n20 a_11599_46634.t41 211.01
R26325 a_11599_46634.n17 a_11599_46634.t32 211.01
R26326 a_11599_46634.n5 a_11599_46634.n4 203.463
R26327 a_11599_46634.n7 a_11599_46634.n6 203.463
R26328 a_11599_46634.n11 a_11599_46634.n10 203.463
R26329 a_11599_46634.n13 a_11599_46634.n12 203.463
R26330 a_11599_46634.n15 a_11599_46634.n14 203.463
R26331 a_11599_46634.n9 a_11599_46634.n8 202.456
R26332 a_11599_46634.n36 a_11599_46634.n16 199.278
R26333 a_11599_46634.n31 a_11599_46634.n29 184.709
R26334 a_11599_46634.n21 a_11599_46634.n20 183.34
R26335 a_11599_46634.n28 a_11599_46634.n24 175.602
R26336 a_11599_46634.n23 a_11599_46634.n17 175.019
R26337 a_11599_46634.n21 a_11599_46634.n19 174.832
R26338 a_11599_46634.n22 a_11599_46634.n18 169.802
R26339 a_11599_46634.n31 a_11599_46634.n30 168.891
R26340 a_11599_46634.n27 a_11599_46634.n26 162.691
R26341 a_11599_46634.n27 a_11599_46634.n25 162.398
R26342 a_11599_46634.n7 a_11599_46634.n5 45.177
R26343 a_11599_46634.n13 a_11599_46634.n11 45.177
R26344 a_11599_46634.n15 a_11599_46634.n13 45.177
R26345 a_11599_46634.n9 a_11599_46634.n7 44.0476
R26346 a_11599_46634.n11 a_11599_46634.n9 44.0476
R26347 a_11599_46634.n3 a_11599_46634.t20 40.0005
R26348 a_11599_46634.n3 a_11599_46634.t26 40.0005
R26349 a_11599_46634.n4 a_11599_46634.t30 40.0005
R26350 a_11599_46634.n4 a_11599_46634.t16 40.0005
R26351 a_11599_46634.n6 a_11599_46634.t31 40.0005
R26352 a_11599_46634.n6 a_11599_46634.t29 40.0005
R26353 a_11599_46634.n8 a_11599_46634.t21 40.0005
R26354 a_11599_46634.n8 a_11599_46634.t19 40.0005
R26355 a_11599_46634.n10 a_11599_46634.t27 40.0005
R26356 a_11599_46634.n10 a_11599_46634.t24 40.0005
R26357 a_11599_46634.n12 a_11599_46634.t17 40.0005
R26358 a_11599_46634.n12 a_11599_46634.t22 40.0005
R26359 a_11599_46634.n14 a_11599_46634.t28 40.0005
R26360 a_11599_46634.n14 a_11599_46634.t23 40.0005
R26361 a_11599_46634.n16 a_11599_46634.t18 40.0005
R26362 a_11599_46634.n16 a_11599_46634.t25 40.0005
R26363 a_11599_46634.n41 a_11599_46634.n39 32.0005
R26364 a_11599_46634.n43 a_11599_46634.n41 32.0005
R26365 a_11599_46634.n46 a_11599_46634.n2 32.0005
R26366 a_11599_46634.n46 a_11599_46634.n45 32.0005
R26367 a_11599_46634.n45 a_11599_46634.n43 31.2005
R26368 a_11599_46634.n38 a_11599_46634.t5 27.5805
R26369 a_11599_46634.n38 a_11599_46634.t1 27.5805
R26370 a_11599_46634.n34 a_11599_46634.t3 27.5805
R26371 a_11599_46634.n34 a_11599_46634.t10 27.5805
R26372 a_11599_46634.n40 a_11599_46634.t6 27.5805
R26373 a_11599_46634.n40 a_11599_46634.t13 27.5805
R26374 a_11599_46634.n42 a_11599_46634.t11 27.5805
R26375 a_11599_46634.n42 a_11599_46634.t0 27.5805
R26376 a_11599_46634.n44 a_11599_46634.t8 27.5805
R26377 a_11599_46634.n44 a_11599_46634.t14 27.5805
R26378 a_11599_46634.n0 a_11599_46634.t2 27.5805
R26379 a_11599_46634.n0 a_11599_46634.t9 27.5805
R26380 a_11599_46634.n1 a_11599_46634.t7 27.5805
R26381 a_11599_46634.n1 a_11599_46634.t12 27.5805
R26382 a_11599_46634.n47 a_11599_46634.t4 27.5805
R26383 a_11599_46634.t15 a_11599_46634.n47 27.5805
R26384 a_11599_46634.n28 a_11599_46634.n27 19.4456
R26385 a_11599_46634.n35 a_11599_46634.n33 16.4752
R26386 a_11599_46634.n37 a_11599_46634.n15 13.177
R26387 a_11599_46634.n23 a_11599_46634.n22 10.3631
R26388 a_11599_46634.n39 a_11599_46634.n37 10.2022
R26389 a_11599_46634.n32 a_11599_46634.n28 9.64336
R26390 a_11599_46634.n33 a_11599_46634.n32 7.73814
R26391 a_11599_46634.n37 a_11599_46634.n36 7.34263
R26392 a_11599_46634.n33 a_11599_46634.n23 6.57193
R26393 a_11599_46634.n22 a_11599_46634.n21 5.88649
R26394 a_11599_46634.n32 a_11599_46634.n31 4.5005
R26395 a_11599_46634.n36 a_11599_46634.n35 0.0969973
R26396 a_n971_45724.n17 a_n971_45724.n15 459.668
R26397 a_n971_45724.n13 a_n971_45724.n11 459.668
R26398 a_n971_45724.n3 a_n971_45724.n1 459.668
R26399 a_n971_45724.n27 a_n971_45724.n26 380.32
R26400 a_n971_45724.n0 a_n971_45724.t24 330.12
R26401 a_n971_45724.n16 a_n971_45724.t23 329.902
R26402 a_n971_45724.n12 a_n971_45724.t13 329.902
R26403 a_n971_45724.n2 a_n971_45724.t26 329.902
R26404 a_n971_45724.n15 a_n971_45724.t8 272.062
R26405 a_n971_45724.n11 a_n971_45724.t22 272.062
R26406 a_n971_45724.n1 a_n971_45724.t28 272.062
R26407 a_n971_45724.n21 a_n971_45724.t16 256.716
R26408 a_n971_45724.n23 a_n971_45724.t10 241.536
R26409 a_n971_45724.n5 a_n971_45724.t27 241.536
R26410 a_n971_45724.n19 a_n971_45724.t25 236.18
R26411 a_n971_45724.n4 a_n971_45724.n0 222.053
R26412 a_n971_45724.n15 a_n971_45724.t29 206.19
R26413 a_n971_45724.n11 a_n971_45724.t19 206.19
R26414 a_n971_45724.n1 a_n971_45724.t15 206.19
R26415 a_n971_45724.n0 a_n971_45724.t18 201.587
R26416 a_n971_45724.n24 a_n971_45724.n23 198.696
R26417 a_n971_45724.n26 a_n971_45724.n25 185
R26418 a_n971_45724.n22 a_n971_45724.n21 175.931
R26419 a_n971_45724.n23 a_n971_45724.t11 169.237
R26420 a_n971_45724.n5 a_n971_45724.t4 169.237
R26421 a_n971_45724.n7 a_n971_45724.n6 168.282
R26422 a_n971_45724.n7 a_n971_45724.n5 168.064
R26423 a_n971_45724.n9 a_n971_45724.n8 167.631
R26424 a_n971_45724.n19 a_n971_45724.t6 163.881
R26425 a_n971_45724.n20 a_n971_45724.n19 162.464
R26426 a_n971_45724.n21 a_n971_45724.t21 161.275
R26427 a_n971_45724.n17 a_n971_45724.n16 152
R26428 a_n971_45724.n13 a_n971_45724.n12 152
R26429 a_n971_45724.n3 a_n971_45724.n2 152
R26430 a_n971_45724.n16 a_n971_45724.t20 148.35
R26431 a_n971_45724.n12 a_n971_45724.t14 148.35
R26432 a_n971_45724.n2 a_n971_45724.t7 148.35
R26433 a_n971_45724.n6 a_n971_45724.t9 142.994
R26434 a_n971_45724.n8 a_n971_45724.t12 137.177
R26435 a_n971_45724.n6 a_n971_45724.t17 126.927
R26436 a_n971_45724.n8 a_n971_45724.t5 121.109
R26437 a_n971_45724.n22 a_n971_45724.n20 27.9336
R26438 a_n971_45724.n10 a_n971_45724.n4 27.2452
R26439 a_n971_45724.n27 a_n971_45724.t0 26.5955
R26440 a_n971_45724.t1 a_n971_45724.n27 26.5955
R26441 a_n971_45724.n25 a_n971_45724.t3 24.9236
R26442 a_n971_45724.n25 a_n971_45724.t2 24.9236
R26443 a_n971_45724.n20 a_n971_45724.n18 20.6734
R26444 a_n971_45724.n14 a_n971_45724.n13 18.5163
R26445 a_n971_45724.n18 a_n971_45724.n14 16.8413
R26446 a_n971_45724.n18 a_n971_45724.n17 14.0163
R26447 a_n971_45724.n4 a_n971_45724.n3 14.0163
R26448 a_n971_45724.n10 a_n971_45724.n9 13.7793
R26449 a_n971_45724.n14 a_n971_45724.n10 11.701
R26450 a_n971_45724.n26 a_n971_45724.n24 11.4352
R26451 a_n971_45724.n9 a_n971_45724.n7 7.19847
R26452 a_n971_45724.n24 a_n971_45724.n22 0.705335
R26453 CLK_DATA.n5 CLK_DATA.n4 647.148
R26454 CLK_DATA.n2 CLK_DATA.n0 243.627
R26455 CLK_DATA.n2 CLK_DATA.n1 200.262
R26456 CLK_DATA.n5 CLK_DATA.n3 194.441
R26457 CLK_DATA.n6 CLK_DATA.n5 42.8458
R26458 CLK_DATA.n0 CLK_DATA.t5 40.0005
R26459 CLK_DATA.n0 CLK_DATA.t7 40.0005
R26460 CLK_DATA.n1 CLK_DATA.t6 40.0005
R26461 CLK_DATA.n1 CLK_DATA.t4 40.0005
R26462 CLK_DATA.n3 CLK_DATA.t0 27.5805
R26463 CLK_DATA.n3 CLK_DATA.t2 27.5805
R26464 CLK_DATA.n4 CLK_DATA.t3 27.5805
R26465 CLK_DATA.n4 CLK_DATA.t1 27.5805
R26466 CLK_DATA CLK_DATA.n6 15.6872
R26467 CLK_DATA.n6 CLK_DATA.n2 7.72512
R26468 a_4958_30871.n7 a_4958_30871.t8 1421.83
R26469 a_4958_30871.n1 a_4958_30871.t12 1421.83
R26470 a_4958_30871.n6 a_4958_30871.t11 1327.11
R26471 a_4958_30871.n2 a_4958_30871.t13 1327.11
R26472 a_4958_30871.n7 a_4958_30871.t7 1320.68
R26473 a_4958_30871.n5 a_4958_30871.t10 1320.68
R26474 a_4958_30871.n3 a_4958_30871.t6 1320.68
R26475 a_4958_30871.n1 a_4958_30871.t4 1320.68
R26476 a_4958_30871.n13 a_4958_30871.n12 287.752
R26477 a_4958_30871.n12 a_4958_30871.n0 277.568
R26478 a_4958_30871.n10 a_4958_30871.t9 260.322
R26479 a_4958_30871.n11 a_4958_30871.n10 175.754
R26480 a_4958_30871.n10 a_4958_30871.t5 175.169
R26481 a_4958_30871.n8 a_4958_30871.n5 161.698
R26482 a_4958_30871.n4 a_4958_30871.n3 161.698
R26483 a_4958_30871.n8 a_4958_30871.n7 161.303
R26484 a_4958_30871.n4 a_4958_30871.n1 161.303
R26485 a_4958_30871.n6 a_4958_30871.n5 94.7191
R26486 a_4958_30871.n7 a_4958_30871.n6 94.7191
R26487 a_4958_30871.n2 a_4958_30871.n1 94.7191
R26488 a_4958_30871.n3 a_4958_30871.n2 94.7191
R26489 a_4958_30871.n11 a_4958_30871.n9 70.4551
R26490 a_4958_30871.n9 a_4958_30871.n8 34.9536
R26491 a_4958_30871.n9 a_4958_30871.n4 32.2328
R26492 a_4958_30871.n12 a_4958_30871.n11 31.4561
R26493 a_4958_30871.t1 a_4958_30871.n13 26.5955
R26494 a_4958_30871.n13 a_4958_30871.t0 26.5955
R26495 a_4958_30871.n0 a_4958_30871.t3 24.9236
R26496 a_4958_30871.n0 a_4958_30871.t2 24.9236
R26497 C9_P_btm C9_P_btm.n15 80.5005
R26498 C9_P_btm.n2 C9_P_btm.n0 33.0802
R26499 C9_P_btm.n6 C9_P_btm.n5 32.3614
R26500 C9_P_btm.n4 C9_P_btm.n3 32.3614
R26501 C9_P_btm.n2 C9_P_btm.n1 32.3614
R26502 C9_P_btm.n10 C9_P_btm.n6 24.0265
R26503 C9_P_btm.n11 C9_P_btm.t16 23.0826
R26504 C9_P_btm.n14 C9_P_btm.n12 15.4287
R26505 C9_P_btm.n9 C9_P_btm.n8 15.3784
R26506 C9_P_btm.n14 C9_P_btm.n13 14.9755
R26507 C9_P_btm.n9 C9_P_btm.n7 14.894
R26508 C9_P_btm.n15 C9_P_btm.n11 7.16717
R26509 C9_P_btm.n10 C9_P_btm.n9 5.71404
R26510 C9_P_btm.n15 C9_P_btm.n14 5.62029
R26511 C9_P_btm C9_P_btm.n513 5.56847
R26512 C9_P_btm.n11 C9_P_btm.n10 3.91717
R26513 C9_P_btm.n5 C9_P_btm.t10 3.57113
R26514 C9_P_btm.n5 C9_P_btm.t8 3.57113
R26515 C9_P_btm.n3 C9_P_btm.t13 3.57113
R26516 C9_P_btm.n3 C9_P_btm.t15 3.57113
R26517 C9_P_btm.n1 C9_P_btm.t14 3.57113
R26518 C9_P_btm.n1 C9_P_btm.t9 3.57113
R26519 C9_P_btm.n0 C9_P_btm.t12 3.57113
R26520 C9_P_btm.n0 C9_P_btm.t11 3.57113
R26521 C9_P_btm.n7 C9_P_btm.t2 2.4755
R26522 C9_P_btm.n7 C9_P_btm.t1 2.4755
R26523 C9_P_btm.n13 C9_P_btm.t7 2.4755
R26524 C9_P_btm.n13 C9_P_btm.t5 2.4755
R26525 C9_P_btm.n12 C9_P_btm.t6 2.4755
R26526 C9_P_btm.n12 C9_P_btm.t4 2.4755
R26527 C9_P_btm.n8 C9_P_btm.t3 2.4755
R26528 C9_P_btm.n8 C9_P_btm.t0 2.4755
R26529 C9_P_btm.n4 C9_P_btm.n2 0.688
R26530 C9_P_btm.n6 C9_P_btm.n4 0.672375
R26531 C9_P_btm.n289 C9_P_btm.n286 0.276161
R26532 C9_P_btm.n83 C9_P_btm.n82 0.276161
R26533 C9_P_btm.n105 C9_P_btm.n104 0.276161
R26534 C9_P_btm.n265 C9_P_btm.n264 0.276161
R26535 C9_P_btm.n332 C9_P_btm.n291 0.276161
R26536 C9_P_btm.n84 C9_P_btm.n77 0.228786
R26537 C9_P_btm.n81 C9_P_btm.n78 0.228786
R26538 C9_P_btm.n145 C9_P_btm.n144 0.228786
R26539 C9_P_btm.n169 C9_P_btm.n168 0.228786
R26540 C9_P_btm.n167 C9_P_btm.n166 0.228786
R26541 C9_P_btm.n177 C9_P_btm.n165 0.228786
R26542 C9_P_btm.n175 C9_P_btm.n174 0.228786
R26543 C9_P_btm.n174 C9_P_btm.n158 0.228786
R26544 C9_P_btm.n173 C9_P_btm.n172 0.228786
R26545 C9_P_btm.n171 C9_P_btm.n170 0.228786
R26546 C9_P_btm.n147 C9_P_btm.n146 0.228786
R26547 C9_P_btm.n473 C9_P_btm.n472 0.228786
R26548 C9_P_btm.n148 C9_P_btm.n143 0.228786
R26549 C9_P_btm.n458 C9_P_btm.n142 0.228786
R26550 C9_P_btm.n457 C9_P_btm.n141 0.228786
R26551 C9_P_btm.n456 C9_P_btm.n140 0.228786
R26552 C9_P_btm.n439 C9_P_btm.n139 0.228786
R26553 C9_P_btm.n49 C9_P_btm.n48 0.228786
R26554 C9_P_btm.n484 C9_P_btm.n483 0.228786
R26555 C9_P_btm.n50 C9_P_btm.n46 0.228786
R26556 C9_P_btm.n136 C9_P_btm.n135 0.228786
R26557 C9_P_btm.n134 C9_P_btm.n52 0.228786
R26558 C9_P_btm.n79 C9_P_btm.n53 0.228786
R26559 C9_P_btm.n132 C9_P_btm.n53 0.228786
R26560 C9_P_btm.n76 C9_P_btm.n54 0.228786
R26561 C9_P_btm.n55 C9_P_btm.n54 0.228786
R26562 C9_P_btm.n86 C9_P_btm.n85 0.228786
R26563 C9_P_btm.n87 C9_P_btm.n57 0.228786
R26564 C9_P_btm.n59 C9_P_btm.n58 0.228786
R26565 C9_P_btm.n61 C9_P_btm.n60 0.228786
R26566 C9_P_btm.n63 C9_P_btm.n62 0.228786
R26567 C9_P_btm.n65 C9_P_btm.n64 0.228786
R26568 C9_P_btm.n67 C9_P_btm.n66 0.228786
R26569 C9_P_btm.n69 C9_P_btm.n68 0.228786
R26570 C9_P_btm.n71 C9_P_btm.n70 0.228786
R26571 C9_P_btm.n73 C9_P_btm.n72 0.228786
R26572 C9_P_btm.n106 C9_P_btm.n18 0.228786
R26573 C9_P_btm.n108 C9_P_btm.n107 0.228786
R26574 C9_P_btm.n109 C9_P_btm.n108 0.228786
R26575 C9_P_btm.n19 C9_P_btm.n18 0.228786
R26576 C9_P_btm.n21 C9_P_btm.n19 0.228786
R26577 C9_P_btm.n110 C9_P_btm.n109 0.228786
R26578 C9_P_btm.n111 C9_P_btm.n110 0.228786
R26579 C9_P_btm.n22 C9_P_btm.n21 0.228786
R26580 C9_P_btm.n113 C9_P_btm.n22 0.228786
R26581 C9_P_btm.n112 C9_P_btm.n111 0.228786
R26582 C9_P_btm.n115 C9_P_btm.n112 0.228786
R26583 C9_P_btm.n114 C9_P_btm.n113 0.228786
R26584 C9_P_btm.n114 C9_P_btm.n26 0.228786
R26585 C9_P_btm.n116 C9_P_btm.n115 0.228786
R26586 C9_P_btm.n117 C9_P_btm.n116 0.228786
R26587 C9_P_btm.n27 C9_P_btm.n26 0.228786
R26588 C9_P_btm.n29 C9_P_btm.n27 0.228786
R26589 C9_P_btm.n118 C9_P_btm.n117 0.228786
R26590 C9_P_btm.n119 C9_P_btm.n118 0.228786
R26591 C9_P_btm.n30 C9_P_btm.n29 0.228786
R26592 C9_P_btm.n121 C9_P_btm.n30 0.228786
R26593 C9_P_btm.n120 C9_P_btm.n119 0.228786
R26594 C9_P_btm.n123 C9_P_btm.n120 0.228786
R26595 C9_P_btm.n122 C9_P_btm.n121 0.228786
R26596 C9_P_btm.n122 C9_P_btm.n34 0.228786
R26597 C9_P_btm.n124 C9_P_btm.n123 0.228786
R26598 C9_P_btm.n125 C9_P_btm.n124 0.228786
R26599 C9_P_btm.n35 C9_P_btm.n34 0.228786
R26600 C9_P_btm.n37 C9_P_btm.n35 0.228786
R26601 C9_P_btm.n126 C9_P_btm.n125 0.228786
R26602 C9_P_btm.n127 C9_P_btm.n126 0.228786
R26603 C9_P_btm.n38 C9_P_btm.n37 0.228786
R26604 C9_P_btm.n129 C9_P_btm.n38 0.228786
R26605 C9_P_btm.n128 C9_P_btm.n127 0.228786
R26606 C9_P_btm.n128 C9_P_btm.n56 0.228786
R26607 C9_P_btm.n130 C9_P_btm.n129 0.228786
R26608 C9_P_btm.n131 C9_P_btm.n130 0.228786
R26609 C9_P_btm.n43 C9_P_btm.n42 0.228786
R26610 C9_P_btm.n133 C9_P_btm.n43 0.228786
R26611 C9_P_btm.n488 C9_P_btm.n44 0.228786
R26612 C9_P_btm.n487 C9_P_btm.n486 0.228786
R26613 C9_P_btm.n485 C9_P_btm.n45 0.228786
R26614 C9_P_btm.n446 C9_P_btm.n47 0.228786
R26615 C9_P_btm.n441 C9_P_btm.n440 0.228786
R26616 C9_P_btm.n455 C9_P_btm.n454 0.228786
R26617 C9_P_btm.n438 C9_P_btm.n437 0.228786
R26618 C9_P_btm.n460 C9_P_btm.n459 0.228786
R26619 C9_P_btm.n461 C9_P_btm.n149 0.228786
R26620 C9_P_btm.n471 C9_P_btm.n150 0.228786
R26621 C9_P_btm.n470 C9_P_btm.n469 0.228786
R26622 C9_P_btm.n468 C9_P_btm.n151 0.228786
R26623 C9_P_btm.n157 C9_P_btm.n153 0.228786
R26624 C9_P_btm.n431 C9_P_btm.n430 0.228786
R26625 C9_P_btm.n429 C9_P_btm.n156 0.228786
R26626 C9_P_btm.n428 C9_P_btm.n427 0.228786
R26627 C9_P_btm.n429 C9_P_btm.n159 0.228786
R26628 C9_P_btm.n164 C9_P_btm.n159 0.228786
R26629 C9_P_btm.n427 C9_P_btm.n426 0.228786
R26630 C9_P_btm.n426 C9_P_btm.n425 0.228786
R26631 C9_P_btm.n424 C9_P_btm.n163 0.228786
R26632 C9_P_btm.n424 C9_P_btm.n423 0.228786
R26633 C9_P_btm.n422 C9_P_btm.n179 0.228786
R26634 C9_P_btm.n421 C9_P_btm.n180 0.228786
R26635 C9_P_btm.n420 C9_P_btm.n419 0.228786
R26636 C9_P_btm.n418 C9_P_btm.n181 0.228786
R26637 C9_P_btm.n202 C9_P_btm.n183 0.228786
R26638 C9_P_btm.n246 C9_P_btm.n245 0.228786
R26639 C9_P_btm.n212 C9_P_btm.n211 0.228786
R26640 C9_P_btm.n379 C9_P_btm.n378 0.228786
R26641 C9_P_btm.n380 C9_P_btm.n200 0.228786
R26642 C9_P_btm.n200 C9_P_btm.n199 0.228786
R26643 C9_P_btm.n383 C9_P_btm.n382 0.228786
R26644 C9_P_btm.n201 C9_P_btm.n197 0.228786
R26645 C9_P_btm.n208 C9_P_btm.n207 0.228786
R26646 C9_P_btm.n206 C9_P_btm.n205 0.228786
R26647 C9_P_btm.n185 C9_P_btm.n184 0.228786
R26648 C9_P_btm.n417 C9_P_btm.n416 0.228786
R26649 C9_P_btm.n186 C9_P_btm.n182 0.228786
R26650 C9_P_btm.n402 C9_P_btm.n401 0.228786
R26651 C9_P_btm.n400 C9_P_btm.n399 0.228786
R26652 C9_P_btm.n162 C9_P_btm.n160 0.228786
R26653 C9_P_btm.n398 C9_P_btm.n397 0.228786
R26654 C9_P_btm.n404 C9_P_btm.n403 0.228786
R26655 C9_P_btm.n392 C9_P_btm.n187 0.228786
R26656 C9_P_btm.n415 C9_P_btm.n188 0.228786
R26657 C9_P_btm.n414 C9_P_btm.n413 0.228786
R26658 C9_P_btm.n412 C9_P_btm.n189 0.228786
R26659 C9_P_btm.n196 C9_P_btm.n191 0.228786
R26660 C9_P_btm.n386 C9_P_btm.n385 0.228786
R26661 C9_P_btm.n384 C9_P_btm.n195 0.228786
R26662 C9_P_btm.n364 C9_P_btm.n198 0.228786
R26663 C9_P_btm.n363 C9_P_btm.n213 0.228786
R26664 C9_P_btm.n377 C9_P_btm.n213 0.228786
R26665 C9_P_btm.n376 C9_P_btm.n375 0.228786
R26666 C9_P_btm.n375 C9_P_btm.n215 0.228786
R26667 C9_P_btm.n372 C9_P_btm.n216 0.228786
R26668 C9_P_btm.n374 C9_P_btm.n373 0.228786
R26669 C9_P_btm.n374 C9_P_btm.n214 0.228786
R26670 C9_P_btm.n242 C9_P_btm.n216 0.228786
R26671 C9_P_btm.n244 C9_P_btm.n242 0.228786
R26672 C9_P_btm.n247 C9_P_btm.n244 0.228786
R26673 C9_P_btm.n239 C9_P_btm.n238 0.228786
R26674 C9_P_btm.n248 C9_P_btm.n243 0.228786
R26675 C9_P_btm.n251 C9_P_btm.n250 0.228786
R26676 C9_P_btm.n253 C9_P_btm.n241 0.228786
R26677 C9_P_btm.n252 C9_P_btm.n218 0.228786
R26678 C9_P_btm.n255 C9_P_btm.n254 0.228786
R26679 C9_P_btm.n231 C9_P_btm.n230 0.228786
R26680 C9_P_btm.n233 C9_P_btm.n231 0.228786
R26681 C9_P_btm.n257 C9_P_btm.n256 0.228786
R26682 C9_P_btm.n258 C9_P_btm.n257 0.228786
R26683 C9_P_btm.n234 C9_P_btm.n233 0.228786
R26684 C9_P_btm.n260 C9_P_btm.n234 0.228786
R26685 C9_P_btm.n259 C9_P_btm.n258 0.228786
R26686 C9_P_btm.n259 C9_P_btm.n240 0.228786
R26687 C9_P_btm.n261 C9_P_btm.n260 0.228786
R26688 C9_P_btm.n262 C9_P_btm.n261 0.228786
R26689 C9_P_btm.n263 C9_P_btm.n262 0.228786
R26690 C9_P_btm.n237 C9_P_btm.n236 0.228786
R26691 C9_P_btm.n266 C9_P_btm.n265 0.228786
R26692 C9_P_btm.n268 C9_P_btm.n235 0.228786
R26693 C9_P_btm.n267 C9_P_btm.n232 0.228786
R26694 C9_P_btm.n270 C9_P_btm.n269 0.228786
R26695 C9_P_btm.n272 C9_P_btm.n229 0.228786
R26696 C9_P_btm.n271 C9_P_btm.n228 0.228786
R26697 C9_P_btm.n274 C9_P_btm.n273 0.228786
R26698 C9_P_btm.n275 C9_P_btm.n274 0.228786
R26699 C9_P_btm.n314 C9_P_btm.n223 0.228786
R26700 C9_P_btm.n312 C9_P_btm.n225 0.228786
R26701 C9_P_btm.n353 C9_P_btm.n227 0.228786
R26702 C9_P_btm.n310 C9_P_btm.n227 0.228786
R26703 C9_P_btm.n312 C9_P_btm.n311 0.228786
R26704 C9_P_btm.n319 C9_P_btm.n313 0.228786
R26705 C9_P_btm.n321 C9_P_btm.n320 0.228786
R26706 C9_P_btm.n307 C9_P_btm.n301 0.228786
R26707 C9_P_btm.n309 C9_P_btm.n279 0.228786
R26708 C9_P_btm.n280 C9_P_btm.n279 0.228786
R26709 C9_P_btm.n282 C9_P_btm.n280 0.228786
R26710 C9_P_btm.n324 C9_P_btm.n323 0.228786
R26711 C9_P_btm.n322 C9_P_btm.n300 0.228786
R26712 C9_P_btm.n299 C9_P_btm.n296 0.228786
R26713 C9_P_btm.n328 C9_P_btm.n296 0.228786
R26714 C9_P_btm.n326 C9_P_btm.n325 0.228786
R26715 C9_P_btm.n298 C9_P_btm.n283 0.228786
R26716 C9_P_btm.n298 C9_P_btm.n297 0.228786
R26717 C9_P_btm.n297 C9_P_btm.n287 0.228786
R26718 C9_P_btm.n327 C9_P_btm.n293 0.228786
R26719 C9_P_btm.n330 C9_P_btm.n329 0.228786
R26720 C9_P_btm.n333 C9_P_btm.n290 0.228786
R26721 C9_P_btm.n292 C9_P_btm.n290 0.228786
R26722 C9_P_btm.n335 C9_P_btm.n288 0.228786
R26723 C9_P_btm.n335 C9_P_btm.n334 0.228786
R26724 C9_P_btm.n337 C9_P_btm.n336 0.228786
R26725 C9_P_btm.n339 C9_P_btm.n286 0.228786
R26726 C9_P_btm.n338 C9_P_btm.n337 0.228786
R26727 C9_P_btm.n338 C9_P_btm.n285 0.228786
R26728 C9_P_btm.n340 C9_P_btm.n339 0.228786
R26729 C9_P_btm.n341 C9_P_btm.n340 0.228786
R26730 C9_P_btm.n285 C9_P_btm.n284 0.228786
R26731 C9_P_btm.n343 C9_P_btm.n284 0.228786
R26732 C9_P_btm.n342 C9_P_btm.n341 0.228786
R26733 C9_P_btm.n342 C9_P_btm.n281 0.228786
R26734 C9_P_btm.n344 C9_P_btm.n343 0.228786
R26735 C9_P_btm.n345 C9_P_btm.n344 0.228786
R26736 C9_P_btm.n281 C9_P_btm.n278 0.228786
R26737 C9_P_btm.n347 C9_P_btm.n278 0.228786
R26738 C9_P_btm.n346 C9_P_btm.n345 0.228786
R26739 C9_P_btm.n346 C9_P_btm.n277 0.228786
R26740 C9_P_btm.n348 C9_P_btm.n347 0.228786
R26741 C9_P_btm.n349 C9_P_btm.n348 0.228786
R26742 C9_P_btm.n277 C9_P_btm.n276 0.228786
R26743 C9_P_btm.n351 C9_P_btm.n276 0.228786
R26744 C9_P_btm.n350 C9_P_btm.n349 0.228786
R26745 C9_P_btm.n350 C9_P_btm.n275 0.228786
R26746 C9_P_btm.n352 C9_P_btm.n351 0.228786
R26747 C9_P_btm.n352 C9_P_btm.n226 0.228786
R26748 C9_P_btm.n354 C9_P_btm.n353 0.228786
R26749 C9_P_btm.n354 C9_P_btm.n224 0.228786
R26750 C9_P_btm.n356 C9_P_btm.n355 0.228786
R26751 C9_P_btm.n356 C9_P_btm.n222 0.228786
R26752 C9_P_btm.n358 C9_P_btm.n357 0.228786
R26753 C9_P_btm.n358 C9_P_btm.n220 0.228786
R26754 C9_P_btm.n360 C9_P_btm.n219 0.228786
R26755 C9_P_btm.n371 C9_P_btm.n370 0.228786
R26756 C9_P_btm.n369 C9_P_btm.n217 0.228786
R26757 C9_P_btm.n368 C9_P_btm.n361 0.228786
R26758 C9_P_btm.n367 C9_P_btm.n366 0.228786
R26759 C9_P_btm.n365 C9_P_btm.n362 0.228786
R26760 C9_P_btm.n194 C9_P_btm.n193 0.228786
R26761 C9_P_btm.n388 C9_P_btm.n387 0.228786
R26762 C9_P_btm.n389 C9_P_btm.n192 0.228786
R26763 C9_P_btm.n411 C9_P_btm.n410 0.228786
R26764 C9_P_btm.n409 C9_P_btm.n190 0.228786
R26765 C9_P_btm.n408 C9_P_btm.n390 0.228786
R26766 C9_P_btm.n407 C9_P_btm.n406 0.228786
R26767 C9_P_btm.n395 C9_P_btm.n393 0.228786
R26768 C9_P_btm.n394 C9_P_btm.n161 0.228786
R26769 C9_P_btm.n434 C9_P_btm.n154 0.228786
R26770 C9_P_btm.n467 C9_P_btm.n466 0.228786
R26771 C9_P_btm.n465 C9_P_btm.n152 0.228786
R26772 C9_P_btm.n464 C9_P_btm.n463 0.228786
R26773 C9_P_btm.n462 C9_P_btm.n435 0.228786
R26774 C9_P_btm.n443 C9_P_btm.n436 0.228786
R26775 C9_P_btm.n444 C9_P_btm.n442 0.228786
R26776 C9_P_btm.n453 C9_P_btm.n445 0.228786
R26777 C9_P_btm.n452 C9_P_btm.n451 0.228786
R26778 C9_P_btm.n450 C9_P_btm.n447 0.228786
R26779 C9_P_btm.n449 C9_P_btm.n448 0.228786
R26780 C9_P_btm.n41 C9_P_btm.n40 0.228786
R26781 C9_P_btm.n490 C9_P_btm.n489 0.228786
R26782 C9_P_btm.n492 C9_P_btm.n39 0.228786
R26783 C9_P_btm.n491 C9_P_btm.n36 0.228786
R26784 C9_P_btm.n494 C9_P_btm.n493 0.228786
R26785 C9_P_btm.n496 C9_P_btm.n33 0.228786
R26786 C9_P_btm.n495 C9_P_btm.n32 0.228786
R26787 C9_P_btm.n498 C9_P_btm.n497 0.228786
R26788 C9_P_btm.n500 C9_P_btm.n31 0.228786
R26789 C9_P_btm.n499 C9_P_btm.n28 0.228786
R26790 C9_P_btm.n502 C9_P_btm.n501 0.228786
R26791 C9_P_btm.n504 C9_P_btm.n25 0.228786
R26792 C9_P_btm.n503 C9_P_btm.n24 0.228786
R26793 C9_P_btm.n506 C9_P_btm.n505 0.228786
R26794 C9_P_btm.n508 C9_P_btm.n23 0.228786
R26795 C9_P_btm.n507 C9_P_btm.n20 0.228786
R26796 C9_P_btm.n510 C9_P_btm.n509 0.228786
R26797 C9_P_btm.n512 C9_P_btm.n17 0.228786
R26798 C9_P_btm.n511 C9_P_btm.n16 0.228786
R26799 C9_P_btm.n75 C9_P_btm.n74 0.228786
R26800 C9_P_btm.n83 C9_P_btm.n75 0.228786
R26801 C9_P_btm.n85 C9_P_btm.n84 0.228786
R26802 C9_P_btm.n78 C9_P_btm.n76 0.228786
R26803 C9_P_btm.n80 C9_P_btm.n79 0.228786
R26804 C9_P_btm.n52 C9_P_btm.n51 0.228786
R26805 C9_P_btm.n137 C9_P_btm.n136 0.228786
R26806 C9_P_btm.n138 C9_P_btm.n50 0.228786
R26807 C9_P_btm.n483 C9_P_btm.n482 0.228786
R26808 C9_P_btm.n481 C9_P_btm.n49 0.228786
R26809 C9_P_btm.n480 C9_P_btm.n139 0.228786
R26810 C9_P_btm.n479 C9_P_btm.n140 0.228786
R26811 C9_P_btm.n478 C9_P_btm.n141 0.228786
R26812 C9_P_btm.n477 C9_P_btm.n142 0.228786
R26813 C9_P_btm.n476 C9_P_btm.n143 0.228786
R26814 C9_P_btm.n474 C9_P_btm.n473 0.228786
R26815 C9_P_btm.n146 C9_P_btm.n145 0.228786
R26816 C9_P_btm.n170 C9_P_btm.n169 0.228786
R26817 C9_P_btm.n173 C9_P_btm.n167 0.228786
R26818 C9_P_btm.n176 C9_P_btm.n175 0.228786
R26819 C9_P_btm.n425 C9_P_btm.n178 0.228786
R26820 C9_P_btm.n165 C9_P_btm.n164 0.228786
R26821 C9_P_btm.n430 C9_P_btm.n158 0.228786
R26822 C9_P_btm.n172 C9_P_btm.n157 0.228786
R26823 C9_P_btm.n171 C9_P_btm.n151 0.228786
R26824 C9_P_btm.n470 C9_P_btm.n147 0.228786
R26825 C9_P_btm.n472 C9_P_btm.n471 0.228786
R26826 C9_P_btm.n149 C9_P_btm.n148 0.228786
R26827 C9_P_btm.n459 C9_P_btm.n458 0.228786
R26828 C9_P_btm.n457 C9_P_btm.n438 0.228786
R26829 C9_P_btm.n456 C9_P_btm.n455 0.228786
R26830 C9_P_btm.n440 C9_P_btm.n439 0.228786
R26831 C9_P_btm.n48 C9_P_btm.n47 0.228786
R26832 C9_P_btm.n485 C9_P_btm.n484 0.228786
R26833 C9_P_btm.n486 C9_P_btm.n46 0.228786
R26834 C9_P_btm.n135 C9_P_btm.n44 0.228786
R26835 C9_P_btm.n134 C9_P_btm.n133 0.228786
R26836 C9_P_btm.n132 C9_P_btm.n131 0.228786
R26837 C9_P_btm.n56 C9_P_btm.n55 0.228786
R26838 C9_P_btm.n87 C9_P_btm.n86 0.228786
R26839 C9_P_btm.n88 C9_P_btm.n74 0.228786
R26840 C9_P_btm.n89 C9_P_btm.n88 0.228786
R26841 C9_P_btm.n58 C9_P_btm.n57 0.228786
R26842 C9_P_btm.n90 C9_P_btm.n89 0.228786
R26843 C9_P_btm.n91 C9_P_btm.n90 0.228786
R26844 C9_P_btm.n60 C9_P_btm.n59 0.228786
R26845 C9_P_btm.n92 C9_P_btm.n91 0.228786
R26846 C9_P_btm.n93 C9_P_btm.n92 0.228786
R26847 C9_P_btm.n62 C9_P_btm.n61 0.228786
R26848 C9_P_btm.n94 C9_P_btm.n93 0.228786
R26849 C9_P_btm.n95 C9_P_btm.n94 0.228786
R26850 C9_P_btm.n64 C9_P_btm.n63 0.228786
R26851 C9_P_btm.n96 C9_P_btm.n95 0.228786
R26852 C9_P_btm.n97 C9_P_btm.n96 0.228786
R26853 C9_P_btm.n66 C9_P_btm.n65 0.228786
R26854 C9_P_btm.n98 C9_P_btm.n97 0.228786
R26855 C9_P_btm.n99 C9_P_btm.n98 0.228786
R26856 C9_P_btm.n68 C9_P_btm.n67 0.228786
R26857 C9_P_btm.n100 C9_P_btm.n99 0.228786
R26858 C9_P_btm.n101 C9_P_btm.n100 0.228786
R26859 C9_P_btm.n70 C9_P_btm.n69 0.228786
R26860 C9_P_btm.n102 C9_P_btm.n101 0.228786
R26861 C9_P_btm.n103 C9_P_btm.n102 0.228786
R26862 C9_P_btm.n72 C9_P_btm.n71 0.228786
R26863 C9_P_btm.n104 C9_P_btm.n103 0.228786
R26864 C9_P_btm.n42 C9_P_btm.n39 0.228786
R26865 C9_P_btm.n489 C9_P_btm.n488 0.228786
R26866 C9_P_btm.n487 C9_P_btm.n41 0.228786
R26867 C9_P_btm.n448 C9_P_btm.n45 0.228786
R26868 C9_P_btm.n447 C9_P_btm.n446 0.228786
R26869 C9_P_btm.n452 C9_P_btm.n441 0.228786
R26870 C9_P_btm.n454 C9_P_btm.n453 0.228786
R26871 C9_P_btm.n442 C9_P_btm.n437 0.228786
R26872 C9_P_btm.n460 C9_P_btm.n436 0.228786
R26873 C9_P_btm.n462 C9_P_btm.n461 0.228786
R26874 C9_P_btm.n463 C9_P_btm.n150 0.228786
R26875 C9_P_btm.n469 C9_P_btm.n152 0.228786
R26876 C9_P_btm.n468 C9_P_btm.n467 0.228786
R26877 C9_P_btm.n154 C9_P_btm.n153 0.228786
R26878 C9_P_btm.n432 C9_P_btm.n431 0.228786
R26879 C9_P_btm.n156 C9_P_btm.n155 0.228786
R26880 C9_P_btm.n428 C9_P_btm.n161 0.228786
R26881 C9_P_btm.n163 C9_P_btm.n162 0.228786
R26882 C9_P_btm.n400 C9_P_btm.n179 0.228786
R26883 C9_P_btm.n401 C9_P_btm.n180 0.228786
R26884 C9_P_btm.n419 C9_P_btm.n182 0.228786
R26885 C9_P_btm.n418 C9_P_btm.n417 0.228786
R26886 C9_P_btm.n184 C9_P_btm.n183 0.228786
R26887 C9_P_btm.n205 C9_P_btm.n204 0.228786
R26888 C9_P_btm.n209 C9_P_btm.n208 0.228786
R26889 C9_P_btm.n210 C9_P_btm.n201 0.228786
R26890 C9_P_btm.n382 C9_P_btm.n381 0.228786
R26891 C9_P_btm.n245 C9_P_btm.n214 0.228786
R26892 C9_P_btm.n376 C9_P_btm.n212 0.228786
R26893 C9_P_btm.n378 C9_P_btm.n377 0.228786
R26894 C9_P_btm.n199 C9_P_btm.n198 0.228786
R26895 C9_P_btm.n384 C9_P_btm.n383 0.228786
R26896 C9_P_btm.n385 C9_P_btm.n197 0.228786
R26897 C9_P_btm.n207 C9_P_btm.n196 0.228786
R26898 C9_P_btm.n206 C9_P_btm.n189 0.228786
R26899 C9_P_btm.n414 C9_P_btm.n185 0.228786
R26900 C9_P_btm.n416 C9_P_btm.n415 0.228786
R26901 C9_P_btm.n187 C9_P_btm.n186 0.228786
R26902 C9_P_btm.n403 C9_P_btm.n402 0.228786
R26903 C9_P_btm.n399 C9_P_btm.n398 0.228786
R26904 C9_P_btm.n393 C9_P_btm.n160 0.228786
R26905 C9_P_btm.n397 C9_P_btm.n396 0.228786
R26906 C9_P_btm.n405 C9_P_btm.n404 0.228786
R26907 C9_P_btm.n406 C9_P_btm.n392 0.228786
R26908 C9_P_btm.n390 C9_P_btm.n188 0.228786
R26909 C9_P_btm.n413 C9_P_btm.n190 0.228786
R26910 C9_P_btm.n412 C9_P_btm.n411 0.228786
R26911 C9_P_btm.n192 C9_P_btm.n191 0.228786
R26912 C9_P_btm.n387 C9_P_btm.n386 0.228786
R26913 C9_P_btm.n195 C9_P_btm.n194 0.228786
R26914 C9_P_btm.n366 C9_P_btm.n363 0.228786
R26915 C9_P_btm.n365 C9_P_btm.n364 0.228786
R26916 C9_P_btm.n361 C9_P_btm.n215 0.228786
R26917 C9_P_btm.n373 C9_P_btm.n217 0.228786
R26918 C9_P_btm.n372 C9_P_btm.n371 0.228786
R26919 C9_P_btm.n250 C9_P_btm.n249 0.228786
R26920 C9_P_btm.n240 C9_P_btm.n239 0.228786
R26921 C9_P_btm.n243 C9_P_btm.n241 0.228786
R26922 C9_P_btm.n252 C9_P_btm.n251 0.228786
R26923 C9_P_btm.n254 C9_P_btm.n253 0.228786
R26924 C9_P_btm.n219 C9_P_btm.n218 0.228786
R26925 C9_P_btm.n255 C9_P_btm.n220 0.228786
R26926 C9_P_btm.n230 C9_P_btm.n224 0.228786
R26927 C9_P_btm.n256 C9_P_btm.n222 0.228786
R26928 C9_P_btm.n236 C9_P_btm.n235 0.228786
R26929 C9_P_btm.n267 C9_P_btm.n266 0.228786
R26930 C9_P_btm.n269 C9_P_btm.n268 0.228786
R26931 C9_P_btm.n232 C9_P_btm.n229 0.228786
R26932 C9_P_btm.n271 C9_P_btm.n270 0.228786
R26933 C9_P_btm.n273 C9_P_btm.n272 0.228786
R26934 C9_P_btm.n228 C9_P_btm.n226 0.228786
R26935 C9_P_btm.n360 C9_P_btm.n359 0.228786
R26936 C9_P_btm.n359 C9_P_btm.n221 0.228786
R26937 C9_P_btm.n357 C9_P_btm.n223 0.228786
R26938 C9_P_btm.n315 C9_P_btm.n221 0.228786
R26939 C9_P_btm.n318 C9_P_btm.n317 0.228786
R26940 C9_P_btm.n317 C9_P_btm.n316 0.228786
R26941 C9_P_btm.n316 C9_P_btm.n315 0.228786
R26942 C9_P_btm.n355 C9_P_btm.n225 0.228786
R26943 C9_P_btm.n314 C9_P_btm.n313 0.228786
R26944 C9_P_btm.n310 C9_P_btm.n309 0.228786
R26945 C9_P_btm.n311 C9_P_btm.n307 0.228786
R26946 C9_P_btm.n320 C9_P_btm.n319 0.228786
R26947 C9_P_btm.n318 C9_P_btm.n308 0.228786
R26948 C9_P_btm.n305 C9_P_btm.n304 0.228786
R26949 C9_P_btm.n306 C9_P_btm.n305 0.228786
R26950 C9_P_btm.n308 C9_P_btm.n306 0.228786
R26951 C9_P_btm.n322 C9_P_btm.n321 0.228786
R26952 C9_P_btm.n323 C9_P_btm.n301 0.228786
R26953 C9_P_btm.n283 C9_P_btm.n282 0.228786
R26954 C9_P_btm.n325 C9_P_btm.n324 0.228786
R26955 C9_P_btm.n300 C9_P_btm.n299 0.228786
R26956 C9_P_btm.n304 C9_P_btm.n303 0.228786
R26957 C9_P_btm.n294 C9_P_btm.n291 0.228786
R26958 C9_P_btm.n295 C9_P_btm.n294 0.228786
R26959 C9_P_btm.n302 C9_P_btm.n295 0.228786
R26960 C9_P_btm.n303 C9_P_btm.n302 0.228786
R26961 C9_P_btm.n329 C9_P_btm.n328 0.228786
R26962 C9_P_btm.n327 C9_P_btm.n326 0.228786
R26963 C9_P_btm.n288 C9_P_btm.n287 0.228786
R26964 C9_P_btm.n293 C9_P_btm.n292 0.228786
R26965 C9_P_btm.n331 C9_P_btm.n330 0.228786
R26966 C9_P_btm.n491 C9_P_btm.n490 0.228786
R26967 C9_P_btm.n493 C9_P_btm.n492 0.228786
R26968 C9_P_btm.n36 C9_P_btm.n33 0.228786
R26969 C9_P_btm.n495 C9_P_btm.n494 0.228786
R26970 C9_P_btm.n497 C9_P_btm.n496 0.228786
R26971 C9_P_btm.n32 C9_P_btm.n31 0.228786
R26972 C9_P_btm.n499 C9_P_btm.n498 0.228786
R26973 C9_P_btm.n501 C9_P_btm.n500 0.228786
R26974 C9_P_btm.n28 C9_P_btm.n25 0.228786
R26975 C9_P_btm.n503 C9_P_btm.n502 0.228786
R26976 C9_P_btm.n505 C9_P_btm.n504 0.228786
R26977 C9_P_btm.n24 C9_P_btm.n23 0.228786
R26978 C9_P_btm.n507 C9_P_btm.n506 0.228786
R26979 C9_P_btm.n509 C9_P_btm.n508 0.228786
R26980 C9_P_btm.n20 C9_P_btm.n17 0.228786
R26981 C9_P_btm.n511 C9_P_btm.n510 0.228786
R26982 C9_P_btm.n513 C9_P_btm.n512 0.228786
R26983 C9_P_btm.n203 C9_P_btm.n202 0.208893
R26984 C9_P_btm.n264 C9_P_btm.n263 0.208893
R26985 C9_P_btm.n334 C9_P_btm.n289 0.208893
R26986 C9_P_btm.n434 C9_P_btm.n433 0.208893
R26987 C9_P_btm.n107 C9_P_btm.n105 0.208893
R26988 C9_P_btm.n333 C9_P_btm.n332 0.208893
R26989 C9_P_btm.n407 C9_P_btm.n391 0.208893
R26990 C9_P_btm.n82 C9_P_btm.n81 0.208893
R26991 C9_P_btm.n475 C9_P_btm.n144 0.208893
R26992 C9_P_btm.n228 C9_P_btm.n224 0.09425
R26993 C9_P_btm.n230 C9_P_btm.n222 0.09425
R26994 C9_P_btm.n255 C9_P_btm.n219 0.09425
R26995 C9_P_btm.n397 C9_P_btm.n393 0.09425
R26996 C9_P_btm.n172 C9_P_btm.n158 0.09425
R26997 C9_P_btm.n174 C9_P_btm.n164 0.09425
R26998 C9_P_btm.n425 C9_P_btm.n165 0.09425
R26999 C9_P_btm.n84 C9_P_btm.n83 0.09425
R27000 C9_P_btm.n78 C9_P_btm.n77 0.09425
R27001 C9_P_btm.n81 C9_P_btm.n80 0.09425
R27002 C9_P_btm.n80 C9_P_btm.n51 0.09425
R27003 C9_P_btm.n137 C9_P_btm.n51 0.09425
R27004 C9_P_btm.n138 C9_P_btm.n137 0.09425
R27005 C9_P_btm.n482 C9_P_btm.n138 0.09425
R27006 C9_P_btm.n482 C9_P_btm.n481 0.09425
R27007 C9_P_btm.n481 C9_P_btm.n480 0.09425
R27008 C9_P_btm.n480 C9_P_btm.n479 0.09425
R27009 C9_P_btm.n479 C9_P_btm.n478 0.09425
R27010 C9_P_btm.n478 C9_P_btm.n477 0.09425
R27011 C9_P_btm.n477 C9_P_btm.n476 0.09425
R27012 C9_P_btm.n474 C9_P_btm.n145 0.09425
R27013 C9_P_btm.n168 C9_P_btm.n144 0.09425
R27014 C9_P_btm.n169 C9_P_btm.n167 0.09425
R27015 C9_P_btm.n169 C9_P_btm.n145 0.09425
R27016 C9_P_btm.n168 C9_P_btm.n166 0.09425
R27017 C9_P_btm.n176 C9_P_btm.n166 0.09425
R27018 C9_P_btm.n423 C9_P_btm.n178 0.09425
R27019 C9_P_btm.n178 C9_P_btm.n177 0.09425
R27020 C9_P_btm.n177 C9_P_btm.n176 0.09425
R27021 C9_P_btm.n175 C9_P_btm.n165 0.09425
R27022 C9_P_btm.n175 C9_P_btm.n167 0.09425
R27023 C9_P_btm.n174 C9_P_btm.n173 0.09425
R27024 C9_P_btm.n173 C9_P_btm.n170 0.09425
R27025 C9_P_btm.n172 C9_P_btm.n171 0.09425
R27026 C9_P_btm.n171 C9_P_btm.n147 0.09425
R27027 C9_P_btm.n170 C9_P_btm.n146 0.09425
R27028 C9_P_btm.n473 C9_P_btm.n146 0.09425
R27029 C9_P_btm.n472 C9_P_btm.n147 0.09425
R27030 C9_P_btm.n472 C9_P_btm.n148 0.09425
R27031 C9_P_btm.n473 C9_P_btm.n143 0.09425
R27032 C9_P_btm.n143 C9_P_btm.n142 0.09425
R27033 C9_P_btm.n458 C9_P_btm.n148 0.09425
R27034 C9_P_btm.n458 C9_P_btm.n457 0.09425
R27035 C9_P_btm.n142 C9_P_btm.n141 0.09425
R27036 C9_P_btm.n141 C9_P_btm.n140 0.09425
R27037 C9_P_btm.n457 C9_P_btm.n456 0.09425
R27038 C9_P_btm.n456 C9_P_btm.n439 0.09425
R27039 C9_P_btm.n140 C9_P_btm.n139 0.09425
R27040 C9_P_btm.n139 C9_P_btm.n49 0.09425
R27041 C9_P_btm.n439 C9_P_btm.n48 0.09425
R27042 C9_P_btm.n484 C9_P_btm.n48 0.09425
R27043 C9_P_btm.n483 C9_P_btm.n49 0.09425
R27044 C9_P_btm.n483 C9_P_btm.n50 0.09425
R27045 C9_P_btm.n484 C9_P_btm.n46 0.09425
R27046 C9_P_btm.n135 C9_P_btm.n46 0.09425
R27047 C9_P_btm.n136 C9_P_btm.n50 0.09425
R27048 C9_P_btm.n136 C9_P_btm.n52 0.09425
R27049 C9_P_btm.n135 C9_P_btm.n134 0.09425
R27050 C9_P_btm.n134 C9_P_btm.n53 0.09425
R27051 C9_P_btm.n79 C9_P_btm.n52 0.09425
R27052 C9_P_btm.n79 C9_P_btm.n78 0.09425
R27053 C9_P_btm.n133 C9_P_btm.n132 0.09425
R27054 C9_P_btm.n132 C9_P_btm.n54 0.09425
R27055 C9_P_btm.n76 C9_P_btm.n53 0.09425
R27056 C9_P_btm.n84 C9_P_btm.n76 0.09425
R27057 C9_P_btm.n131 C9_P_btm.n55 0.09425
R27058 C9_P_btm.n86 C9_P_btm.n55 0.09425
R27059 C9_P_btm.n85 C9_P_btm.n54 0.09425
R27060 C9_P_btm.n85 C9_P_btm.n75 0.09425
R27061 C9_P_btm.n86 C9_P_btm.n74 0.09425
R27062 C9_P_btm.n87 C9_P_btm.n56 0.09425
R27063 C9_P_btm.n88 C9_P_btm.n87 0.09425
R27064 C9_P_btm.n89 C9_P_btm.n57 0.09425
R27065 C9_P_btm.n127 C9_P_btm.n58 0.09425
R27066 C9_P_btm.n90 C9_P_btm.n58 0.09425
R27067 C9_P_btm.n91 C9_P_btm.n59 0.09425
R27068 C9_P_btm.n125 C9_P_btm.n60 0.09425
R27069 C9_P_btm.n92 C9_P_btm.n60 0.09425
R27070 C9_P_btm.n93 C9_P_btm.n61 0.09425
R27071 C9_P_btm.n123 C9_P_btm.n62 0.09425
R27072 C9_P_btm.n94 C9_P_btm.n62 0.09425
R27073 C9_P_btm.n95 C9_P_btm.n63 0.09425
R27074 C9_P_btm.n119 C9_P_btm.n64 0.09425
R27075 C9_P_btm.n96 C9_P_btm.n64 0.09425
R27076 C9_P_btm.n97 C9_P_btm.n65 0.09425
R27077 C9_P_btm.n117 C9_P_btm.n66 0.09425
R27078 C9_P_btm.n98 C9_P_btm.n66 0.09425
R27079 C9_P_btm.n99 C9_P_btm.n67 0.09425
R27080 C9_P_btm.n115 C9_P_btm.n68 0.09425
R27081 C9_P_btm.n100 C9_P_btm.n68 0.09425
R27082 C9_P_btm.n101 C9_P_btm.n69 0.09425
R27083 C9_P_btm.n111 C9_P_btm.n70 0.09425
R27084 C9_P_btm.n102 C9_P_btm.n70 0.09425
R27085 C9_P_btm.n103 C9_P_btm.n71 0.09425
R27086 C9_P_btm.n109 C9_P_btm.n72 0.09425
R27087 C9_P_btm.n104 C9_P_btm.n72 0.09425
R27088 C9_P_btm.n106 C9_P_btm.n16 0.09425
R27089 C9_P_btm.n107 C9_P_btm.n106 0.09425
R27090 C9_P_btm.n108 C9_P_btm.n18 0.09425
R27091 C9_P_btm.n108 C9_P_btm.n73 0.09425
R27092 C9_P_btm.n510 C9_P_btm.n19 0.09425
R27093 C9_P_btm.n109 C9_P_btm.n19 0.09425
R27094 C9_P_btm.n110 C9_P_btm.n21 0.09425
R27095 C9_P_btm.n110 C9_P_btm.n71 0.09425
R27096 C9_P_btm.n508 C9_P_btm.n22 0.09425
R27097 C9_P_btm.n111 C9_P_btm.n22 0.09425
R27098 C9_P_btm.n113 C9_P_btm.n112 0.09425
R27099 C9_P_btm.n112 C9_P_btm.n69 0.09425
R27100 C9_P_btm.n114 C9_P_btm.n24 0.09425
R27101 C9_P_btm.n115 C9_P_btm.n114 0.09425
R27102 C9_P_btm.n116 C9_P_btm.n26 0.09425
R27103 C9_P_btm.n116 C9_P_btm.n67 0.09425
R27104 C9_P_btm.n502 C9_P_btm.n27 0.09425
R27105 C9_P_btm.n117 C9_P_btm.n27 0.09425
R27106 C9_P_btm.n118 C9_P_btm.n29 0.09425
R27107 C9_P_btm.n118 C9_P_btm.n65 0.09425
R27108 C9_P_btm.n500 C9_P_btm.n30 0.09425
R27109 C9_P_btm.n119 C9_P_btm.n30 0.09425
R27110 C9_P_btm.n121 C9_P_btm.n120 0.09425
R27111 C9_P_btm.n120 C9_P_btm.n63 0.09425
R27112 C9_P_btm.n122 C9_P_btm.n32 0.09425
R27113 C9_P_btm.n123 C9_P_btm.n122 0.09425
R27114 C9_P_btm.n124 C9_P_btm.n34 0.09425
R27115 C9_P_btm.n124 C9_P_btm.n61 0.09425
R27116 C9_P_btm.n494 C9_P_btm.n35 0.09425
R27117 C9_P_btm.n125 C9_P_btm.n35 0.09425
R27118 C9_P_btm.n126 C9_P_btm.n37 0.09425
R27119 C9_P_btm.n126 C9_P_btm.n59 0.09425
R27120 C9_P_btm.n492 C9_P_btm.n38 0.09425
R27121 C9_P_btm.n127 C9_P_btm.n38 0.09425
R27122 C9_P_btm.n129 C9_P_btm.n128 0.09425
R27123 C9_P_btm.n128 C9_P_btm.n57 0.09425
R27124 C9_P_btm.n130 C9_P_btm.n42 0.09425
R27125 C9_P_btm.n130 C9_P_btm.n56 0.09425
R27126 C9_P_btm.n488 C9_P_btm.n43 0.09425
R27127 C9_P_btm.n131 C9_P_btm.n43 0.09425
R27128 C9_P_btm.n486 C9_P_btm.n44 0.09425
R27129 C9_P_btm.n133 C9_P_btm.n44 0.09425
R27130 C9_P_btm.n487 C9_P_btm.n45 0.09425
R27131 C9_P_btm.n488 C9_P_btm.n487 0.09425
R27132 C9_P_btm.n485 C9_P_btm.n47 0.09425
R27133 C9_P_btm.n486 C9_P_btm.n485 0.09425
R27134 C9_P_btm.n446 C9_P_btm.n441 0.09425
R27135 C9_P_btm.n446 C9_P_btm.n45 0.09425
R27136 C9_P_btm.n455 C9_P_btm.n440 0.09425
R27137 C9_P_btm.n440 C9_P_btm.n47 0.09425
R27138 C9_P_btm.n454 C9_P_btm.n437 0.09425
R27139 C9_P_btm.n454 C9_P_btm.n441 0.09425
R27140 C9_P_btm.n459 C9_P_btm.n438 0.09425
R27141 C9_P_btm.n455 C9_P_btm.n438 0.09425
R27142 C9_P_btm.n461 C9_P_btm.n460 0.09425
R27143 C9_P_btm.n460 C9_P_btm.n437 0.09425
R27144 C9_P_btm.n471 C9_P_btm.n149 0.09425
R27145 C9_P_btm.n459 C9_P_btm.n149 0.09425
R27146 C9_P_btm.n469 C9_P_btm.n150 0.09425
R27147 C9_P_btm.n461 C9_P_btm.n150 0.09425
R27148 C9_P_btm.n470 C9_P_btm.n151 0.09425
R27149 C9_P_btm.n471 C9_P_btm.n470 0.09425
R27150 C9_P_btm.n468 C9_P_btm.n153 0.09425
R27151 C9_P_btm.n469 C9_P_btm.n468 0.09425
R27152 C9_P_btm.n430 C9_P_btm.n157 0.09425
R27153 C9_P_btm.n157 C9_P_btm.n151 0.09425
R27154 C9_P_btm.n431 C9_P_btm.n156 0.09425
R27155 C9_P_btm.n431 C9_P_btm.n153 0.09425
R27156 C9_P_btm.n430 C9_P_btm.n429 0.09425
R27157 C9_P_btm.n428 C9_P_btm.n160 0.09425
R27158 C9_P_btm.n429 C9_P_btm.n428 0.09425
R27159 C9_P_btm.n427 C9_P_btm.n159 0.09425
R27160 C9_P_btm.n159 C9_P_btm.n158 0.09425
R27161 C9_P_btm.n426 C9_P_btm.n163 0.09425
R27162 C9_P_btm.n426 C9_P_btm.n164 0.09425
R27163 C9_P_btm.n424 C9_P_btm.n179 0.09425
R27164 C9_P_btm.n425 C9_P_btm.n424 0.09425
R27165 C9_P_btm.n422 C9_P_btm.n421 0.09425
R27166 C9_P_btm.n423 C9_P_btm.n422 0.09425
R27167 C9_P_btm.n419 C9_P_btm.n180 0.09425
R27168 C9_P_btm.n180 C9_P_btm.n179 0.09425
R27169 C9_P_btm.n420 C9_P_btm.n181 0.09425
R27170 C9_P_btm.n421 C9_P_btm.n420 0.09425
R27171 C9_P_btm.n418 C9_P_btm.n183 0.09425
R27172 C9_P_btm.n419 C9_P_btm.n418 0.09425
R27173 C9_P_btm.n202 C9_P_btm.n181 0.09425
R27174 C9_P_btm.n204 C9_P_btm.n183 0.09425
R27175 C9_P_btm.n210 C9_P_btm.n209 0.09425
R27176 C9_P_btm.n381 C9_P_btm.n210 0.09425
R27177 C9_P_btm.n247 C9_P_btm.n246 0.09425
R27178 C9_P_btm.n245 C9_P_btm.n244 0.09425
R27179 C9_P_btm.n245 C9_P_btm.n212 0.09425
R27180 C9_P_btm.n246 C9_P_btm.n211 0.09425
R27181 C9_P_btm.n379 C9_P_btm.n211 0.09425
R27182 C9_P_btm.n378 C9_P_btm.n212 0.09425
R27183 C9_P_btm.n378 C9_P_btm.n200 0.09425
R27184 C9_P_btm.n380 C9_P_btm.n379 0.09425
R27185 C9_P_btm.n381 C9_P_btm.n380 0.09425
R27186 C9_P_btm.n377 C9_P_btm.n199 0.09425
R27187 C9_P_btm.n383 C9_P_btm.n199 0.09425
R27188 C9_P_btm.n382 C9_P_btm.n200 0.09425
R27189 C9_P_btm.n382 C9_P_btm.n201 0.09425
R27190 C9_P_btm.n383 C9_P_btm.n197 0.09425
R27191 C9_P_btm.n207 C9_P_btm.n197 0.09425
R27192 C9_P_btm.n208 C9_P_btm.n201 0.09425
R27193 C9_P_btm.n208 C9_P_btm.n205 0.09425
R27194 C9_P_btm.n207 C9_P_btm.n206 0.09425
R27195 C9_P_btm.n206 C9_P_btm.n185 0.09425
R27196 C9_P_btm.n205 C9_P_btm.n184 0.09425
R27197 C9_P_btm.n417 C9_P_btm.n184 0.09425
R27198 C9_P_btm.n416 C9_P_btm.n185 0.09425
R27199 C9_P_btm.n416 C9_P_btm.n186 0.09425
R27200 C9_P_btm.n417 C9_P_btm.n182 0.09425
R27201 C9_P_btm.n401 C9_P_btm.n182 0.09425
R27202 C9_P_btm.n402 C9_P_btm.n186 0.09425
R27203 C9_P_btm.n402 C9_P_btm.n399 0.09425
R27204 C9_P_btm.n401 C9_P_btm.n400 0.09425
R27205 C9_P_btm.n400 C9_P_btm.n163 0.09425
R27206 C9_P_btm.n399 C9_P_btm.n162 0.09425
R27207 C9_P_btm.n427 C9_P_btm.n162 0.09425
R27208 C9_P_btm.n403 C9_P_btm.n398 0.09425
R27209 C9_P_btm.n398 C9_P_btm.n160 0.09425
R27210 C9_P_btm.n404 C9_P_btm.n392 0.09425
R27211 C9_P_btm.n404 C9_P_btm.n397 0.09425
R27212 C9_P_btm.n415 C9_P_btm.n187 0.09425
R27213 C9_P_btm.n403 C9_P_btm.n187 0.09425
R27214 C9_P_btm.n413 C9_P_btm.n188 0.09425
R27215 C9_P_btm.n392 C9_P_btm.n188 0.09425
R27216 C9_P_btm.n414 C9_P_btm.n189 0.09425
R27217 C9_P_btm.n415 C9_P_btm.n414 0.09425
R27218 C9_P_btm.n412 C9_P_btm.n191 0.09425
R27219 C9_P_btm.n413 C9_P_btm.n412 0.09425
R27220 C9_P_btm.n385 C9_P_btm.n196 0.09425
R27221 C9_P_btm.n196 C9_P_btm.n189 0.09425
R27222 C9_P_btm.n386 C9_P_btm.n195 0.09425
R27223 C9_P_btm.n386 C9_P_btm.n191 0.09425
R27224 C9_P_btm.n384 C9_P_btm.n198 0.09425
R27225 C9_P_btm.n385 C9_P_btm.n384 0.09425
R27226 C9_P_btm.n363 C9_P_btm.n215 0.09425
R27227 C9_P_btm.n364 C9_P_btm.n363 0.09425
R27228 C9_P_btm.n364 C9_P_btm.n195 0.09425
R27229 C9_P_btm.n375 C9_P_btm.n213 0.09425
R27230 C9_P_btm.n213 C9_P_btm.n198 0.09425
R27231 C9_P_btm.n376 C9_P_btm.n214 0.09425
R27232 C9_P_btm.n377 C9_P_btm.n376 0.09425
R27233 C9_P_btm.n373 C9_P_btm.n215 0.09425
R27234 C9_P_btm.n372 C9_P_btm.n218 0.09425
R27235 C9_P_btm.n373 C9_P_btm.n372 0.09425
R27236 C9_P_btm.n374 C9_P_btm.n216 0.09425
R27237 C9_P_btm.n375 C9_P_btm.n374 0.09425
R27238 C9_P_btm.n251 C9_P_btm.n242 0.09425
R27239 C9_P_btm.n242 C9_P_btm.n214 0.09425
R27240 C9_P_btm.n249 C9_P_btm.n247 0.09425
R27241 C9_P_btm.n263 C9_P_btm.n238 0.09425
R27242 C9_P_btm.n262 C9_P_btm.n239 0.09425
R27243 C9_P_btm.n243 C9_P_btm.n239 0.09425
R27244 C9_P_btm.n248 C9_P_btm.n238 0.09425
R27245 C9_P_btm.n249 C9_P_btm.n248 0.09425
R27246 C9_P_btm.n250 C9_P_btm.n243 0.09425
R27247 C9_P_btm.n250 C9_P_btm.n244 0.09425
R27248 C9_P_btm.n241 C9_P_btm.n240 0.09425
R27249 C9_P_btm.n251 C9_P_btm.n241 0.09425
R27250 C9_P_btm.n253 C9_P_btm.n252 0.09425
R27251 C9_P_btm.n252 C9_P_btm.n216 0.09425
R27252 C9_P_btm.n258 C9_P_btm.n254 0.09425
R27253 C9_P_btm.n254 C9_P_btm.n218 0.09425
R27254 C9_P_btm.n256 C9_P_btm.n220 0.09425
R27255 C9_P_btm.n270 C9_P_btm.n231 0.09425
R27256 C9_P_btm.n256 C9_P_btm.n231 0.09425
R27257 C9_P_btm.n257 C9_P_btm.n233 0.09425
R27258 C9_P_btm.n257 C9_P_btm.n255 0.09425
R27259 C9_P_btm.n268 C9_P_btm.n234 0.09425
R27260 C9_P_btm.n258 C9_P_btm.n234 0.09425
R27261 C9_P_btm.n260 C9_P_btm.n259 0.09425
R27262 C9_P_btm.n259 C9_P_btm.n253 0.09425
R27263 C9_P_btm.n261 C9_P_btm.n236 0.09425
R27264 C9_P_btm.n261 C9_P_btm.n240 0.09425
R27265 C9_P_btm.n262 C9_P_btm.n237 0.09425
R27266 C9_P_btm.n265 C9_P_btm.n236 0.09425
R27267 C9_P_btm.n266 C9_P_btm.n235 0.09425
R27268 C9_P_btm.n260 C9_P_btm.n235 0.09425
R27269 C9_P_btm.n268 C9_P_btm.n267 0.09425
R27270 C9_P_btm.n269 C9_P_btm.n232 0.09425
R27271 C9_P_btm.n269 C9_P_btm.n233 0.09425
R27272 C9_P_btm.n270 C9_P_btm.n229 0.09425
R27273 C9_P_btm.n272 C9_P_btm.n271 0.09425
R27274 C9_P_btm.n271 C9_P_btm.n230 0.09425
R27275 C9_P_btm.n273 C9_P_btm.n228 0.09425
R27276 C9_P_btm.n274 C9_P_btm.n226 0.09425
R27277 C9_P_btm.n330 C9_P_btm.n292 0.09425
R27278 C9_P_btm.n293 C9_P_btm.n287 0.09425
R27279 C9_P_btm.n297 C9_P_btm.n285 0.09425
R27280 C9_P_btm.n357 C9_P_btm.n221 0.09425
R27281 C9_P_btm.n316 C9_P_btm.n314 0.09425
R27282 C9_P_btm.n355 C9_P_btm.n223 0.09425
R27283 C9_P_btm.n315 C9_P_btm.n223 0.09425
R27284 C9_P_btm.n353 C9_P_btm.n225 0.09425
R27285 C9_P_btm.n314 C9_P_btm.n225 0.09425
R27286 C9_P_btm.n351 C9_P_btm.n227 0.09425
R27287 C9_P_btm.n312 C9_P_btm.n227 0.09425
R27288 C9_P_btm.n311 C9_P_btm.n310 0.09425
R27289 C9_P_btm.n319 C9_P_btm.n311 0.09425
R27290 C9_P_btm.n313 C9_P_btm.n312 0.09425
R27291 C9_P_btm.n317 C9_P_btm.n313 0.09425
R27292 C9_P_btm.n319 C9_P_btm.n318 0.09425
R27293 C9_P_btm.n321 C9_P_btm.n306 0.09425
R27294 C9_P_btm.n320 C9_P_btm.n307 0.09425
R27295 C9_P_btm.n320 C9_P_btm.n308 0.09425
R27296 C9_P_btm.n301 C9_P_btm.n279 0.09425
R27297 C9_P_btm.n321 C9_P_btm.n301 0.09425
R27298 C9_P_btm.n309 C9_P_btm.n277 0.09425
R27299 C9_P_btm.n309 C9_P_btm.n307 0.09425
R27300 C9_P_btm.n345 C9_P_btm.n280 0.09425
R27301 C9_P_btm.n323 C9_P_btm.n280 0.09425
R27302 C9_P_btm.n324 C9_P_btm.n282 0.09425
R27303 C9_P_btm.n324 C9_P_btm.n300 0.09425
R27304 C9_P_btm.n323 C9_P_btm.n322 0.09425
R27305 C9_P_btm.n322 C9_P_btm.n305 0.09425
R27306 C9_P_btm.n304 C9_P_btm.n300 0.09425
R27307 C9_P_btm.n328 C9_P_btm.n295 0.09425
R27308 C9_P_btm.n302 C9_P_btm.n296 0.09425
R27309 C9_P_btm.n325 C9_P_btm.n299 0.09425
R27310 C9_P_btm.n303 C9_P_btm.n299 0.09425
R27311 C9_P_btm.n326 C9_P_btm.n298 0.09425
R27312 C9_P_btm.n326 C9_P_btm.n296 0.09425
R27313 C9_P_btm.n343 C9_P_btm.n283 0.09425
R27314 C9_P_btm.n325 C9_P_btm.n283 0.09425
R27315 C9_P_btm.n327 C9_P_btm.n297 0.09425
R27316 C9_P_btm.n328 C9_P_btm.n327 0.09425
R27317 C9_P_btm.n329 C9_P_btm.n293 0.09425
R27318 C9_P_btm.n329 C9_P_btm.n294 0.09425
R27319 C9_P_btm.n330 C9_P_btm.n291 0.09425
R27320 C9_P_btm.n334 C9_P_btm.n333 0.09425
R27321 C9_P_btm.n335 C9_P_btm.n290 0.09425
R27322 C9_P_btm.n331 C9_P_btm.n290 0.09425
R27323 C9_P_btm.n337 C9_P_btm.n288 0.09425
R27324 C9_P_btm.n292 C9_P_btm.n288 0.09425
R27325 C9_P_btm.n336 C9_P_btm.n335 0.09425
R27326 C9_P_btm.n337 C9_P_btm.n286 0.09425
R27327 C9_P_btm.n339 C9_P_btm.n338 0.09425
R27328 C9_P_btm.n338 C9_P_btm.n287 0.09425
R27329 C9_P_btm.n340 C9_P_btm.n285 0.09425
R27330 C9_P_btm.n341 C9_P_btm.n284 0.09425
R27331 C9_P_btm.n298 C9_P_btm.n284 0.09425
R27332 C9_P_btm.n343 C9_P_btm.n342 0.09425
R27333 C9_P_btm.n344 C9_P_btm.n281 0.09425
R27334 C9_P_btm.n344 C9_P_btm.n282 0.09425
R27335 C9_P_btm.n345 C9_P_btm.n278 0.09425
R27336 C9_P_btm.n347 C9_P_btm.n346 0.09425
R27337 C9_P_btm.n346 C9_P_btm.n279 0.09425
R27338 C9_P_btm.n348 C9_P_btm.n277 0.09425
R27339 C9_P_btm.n349 C9_P_btm.n276 0.09425
R27340 C9_P_btm.n310 C9_P_btm.n276 0.09425
R27341 C9_P_btm.n351 C9_P_btm.n350 0.09425
R27342 C9_P_btm.n352 C9_P_btm.n275 0.09425
R27343 C9_P_btm.n353 C9_P_btm.n352 0.09425
R27344 C9_P_btm.n354 C9_P_btm.n226 0.09425
R27345 C9_P_btm.n355 C9_P_btm.n354 0.09425
R27346 C9_P_btm.n356 C9_P_btm.n224 0.09425
R27347 C9_P_btm.n357 C9_P_btm.n356 0.09425
R27348 C9_P_btm.n358 C9_P_btm.n222 0.09425
R27349 C9_P_btm.n359 C9_P_btm.n358 0.09425
R27350 C9_P_btm.n360 C9_P_btm.n220 0.09425
R27351 C9_P_btm.n370 C9_P_btm.n360 0.09425
R27352 C9_P_btm.n371 C9_P_btm.n219 0.09425
R27353 C9_P_btm.n371 C9_P_btm.n217 0.09425
R27354 C9_P_btm.n370 C9_P_btm.n369 0.09425
R27355 C9_P_btm.n369 C9_P_btm.n368 0.09425
R27356 C9_P_btm.n361 C9_P_btm.n217 0.09425
R27357 C9_P_btm.n366 C9_P_btm.n361 0.09425
R27358 C9_P_btm.n368 C9_P_btm.n367 0.09425
R27359 C9_P_btm.n367 C9_P_btm.n362 0.09425
R27360 C9_P_btm.n366 C9_P_btm.n365 0.09425
R27361 C9_P_btm.n365 C9_P_btm.n194 0.09425
R27362 C9_P_btm.n362 C9_P_btm.n193 0.09425
R27363 C9_P_btm.n388 C9_P_btm.n193 0.09425
R27364 C9_P_btm.n387 C9_P_btm.n194 0.09425
R27365 C9_P_btm.n387 C9_P_btm.n192 0.09425
R27366 C9_P_btm.n389 C9_P_btm.n388 0.09425
R27367 C9_P_btm.n410 C9_P_btm.n389 0.09425
R27368 C9_P_btm.n411 C9_P_btm.n192 0.09425
R27369 C9_P_btm.n411 C9_P_btm.n190 0.09425
R27370 C9_P_btm.n410 C9_P_btm.n409 0.09425
R27371 C9_P_btm.n409 C9_P_btm.n408 0.09425
R27372 C9_P_btm.n390 C9_P_btm.n190 0.09425
R27373 C9_P_btm.n406 C9_P_btm.n390 0.09425
R27374 C9_P_btm.n408 C9_P_btm.n407 0.09425
R27375 C9_P_btm.n406 C9_P_btm.n405 0.09425
R27376 C9_P_btm.n396 C9_P_btm.n395 0.09425
R27377 C9_P_btm.n395 C9_P_btm.n394 0.09425
R27378 C9_P_btm.n393 C9_P_btm.n161 0.09425
R27379 C9_P_btm.n161 C9_P_btm.n156 0.09425
R27380 C9_P_btm.n394 C9_P_btm.n155 0.09425
R27381 C9_P_btm.n432 C9_P_btm.n154 0.09425
R27382 C9_P_btm.n467 C9_P_btm.n154 0.09425
R27383 C9_P_btm.n466 C9_P_btm.n434 0.09425
R27384 C9_P_btm.n466 C9_P_btm.n465 0.09425
R27385 C9_P_btm.n467 C9_P_btm.n152 0.09425
R27386 C9_P_btm.n463 C9_P_btm.n152 0.09425
R27387 C9_P_btm.n465 C9_P_btm.n464 0.09425
R27388 C9_P_btm.n464 C9_P_btm.n435 0.09425
R27389 C9_P_btm.n463 C9_P_btm.n462 0.09425
R27390 C9_P_btm.n462 C9_P_btm.n436 0.09425
R27391 C9_P_btm.n443 C9_P_btm.n435 0.09425
R27392 C9_P_btm.n444 C9_P_btm.n443 0.09425
R27393 C9_P_btm.n442 C9_P_btm.n436 0.09425
R27394 C9_P_btm.n453 C9_P_btm.n442 0.09425
R27395 C9_P_btm.n445 C9_P_btm.n444 0.09425
R27396 C9_P_btm.n451 C9_P_btm.n445 0.09425
R27397 C9_P_btm.n453 C9_P_btm.n452 0.09425
R27398 C9_P_btm.n452 C9_P_btm.n447 0.09425
R27399 C9_P_btm.n451 C9_P_btm.n450 0.09425
R27400 C9_P_btm.n450 C9_P_btm.n449 0.09425
R27401 C9_P_btm.n448 C9_P_btm.n447 0.09425
R27402 C9_P_btm.n448 C9_P_btm.n41 0.09425
R27403 C9_P_btm.n449 C9_P_btm.n40 0.09425
R27404 C9_P_btm.n490 C9_P_btm.n40 0.09425
R27405 C9_P_btm.n489 C9_P_btm.n41 0.09425
R27406 C9_P_btm.n489 C9_P_btm.n42 0.09425
R27407 C9_P_btm.n490 C9_P_btm.n39 0.09425
R27408 C9_P_btm.n129 C9_P_btm.n39 0.09425
R27409 C9_P_btm.n492 C9_P_btm.n491 0.09425
R27410 C9_P_btm.n493 C9_P_btm.n36 0.09425
R27411 C9_P_btm.n493 C9_P_btm.n37 0.09425
R27412 C9_P_btm.n494 C9_P_btm.n33 0.09425
R27413 C9_P_btm.n496 C9_P_btm.n495 0.09425
R27414 C9_P_btm.n495 C9_P_btm.n34 0.09425
R27415 C9_P_btm.n497 C9_P_btm.n32 0.09425
R27416 C9_P_btm.n498 C9_P_btm.n31 0.09425
R27417 C9_P_btm.n121 C9_P_btm.n31 0.09425
R27418 C9_P_btm.n500 C9_P_btm.n499 0.09425
R27419 C9_P_btm.n501 C9_P_btm.n28 0.09425
R27420 C9_P_btm.n501 C9_P_btm.n29 0.09425
R27421 C9_P_btm.n502 C9_P_btm.n25 0.09425
R27422 C9_P_btm.n504 C9_P_btm.n503 0.09425
R27423 C9_P_btm.n503 C9_P_btm.n26 0.09425
R27424 C9_P_btm.n505 C9_P_btm.n24 0.09425
R27425 C9_P_btm.n506 C9_P_btm.n23 0.09425
R27426 C9_P_btm.n113 C9_P_btm.n23 0.09425
R27427 C9_P_btm.n508 C9_P_btm.n507 0.09425
R27428 C9_P_btm.n509 C9_P_btm.n20 0.09425
R27429 C9_P_btm.n509 C9_P_btm.n21 0.09425
R27430 C9_P_btm.n510 C9_P_btm.n17 0.09425
R27431 C9_P_btm.n512 C9_P_btm.n511 0.09425
R27432 C9_P_btm.n511 C9_P_btm.n18 0.09425
R27433 C9_P_btm.n513 C9_P_btm.n16 0.09425
R27434 C9_P_btm.n209 C9_P_btm.n203 0.047875
R27435 C9_P_btm.n396 C9_P_btm.n391 0.047875
R27436 C9_P_btm.n433 C9_P_btm.n155 0.047875
R27437 C9_P_btm.n476 C9_P_btm.n475 0.047875
R27438 C9_P_btm.n105 C9_P_btm.n73 0.0342289
R27439 C9_P_btm.n332 C9_P_btm.n331 0.0342289
R27440 C9_P_btm.n405 C9_P_btm.n391 0.0342289
R27441 C9_P_btm.n82 C9_P_btm.n77 0.0342289
R27442 C9_P_btm.n475 C9_P_btm.n474 0.0342289
R27443 C9_P_btm.n204 C9_P_btm.n203 0.0342289
R27444 C9_P_btm.n264 C9_P_btm.n237 0.0342289
R27445 C9_P_btm.n336 C9_P_btm.n289 0.0342289
R27446 C9_P_btm.n433 C9_P_btm.n432 0.0342289
R27447 a_n3565_39590.n4 a_n3565_39590.t9 756.547
R27448 a_n3565_39590.n6 a_n3565_39590.t13 756.226
R27449 a_n3565_39590.n5 a_n3565_39590.t10 756.226
R27450 a_n3565_39590.n4 a_n3565_39590.t12 756.226
R27451 a_n3565_39590.n11 a_n3565_39590.n10 340.637
R27452 a_n3565_39590.n3 a_n3565_39590.t11 241.536
R27453 a_n3565_39590.n10 a_n3565_39590.n9 195.577
R27454 a_n3565_39590.n3 a_n3565_39590.t8 169.237
R27455 a_n3565_39590.n7 a_n3565_39590.n3 168.505
R27456 a_n3565_39590.n2 a_n3565_39590.n0 137.189
R27457 a_n3565_39590.n2 a_n3565_39590.n1 98.788
R27458 a_n3565_39590.n7 a_n3565_39590.n6 75.687
R27459 a_n3565_39590.n10 a_n3565_39590.n8 39.0246
R27460 a_n3565_39590.n9 a_n3565_39590.t2 26.5955
R27461 a_n3565_39590.n9 a_n3565_39590.t1 26.5955
R27462 a_n3565_39590.n11 a_n3565_39590.t0 26.5955
R27463 a_n3565_39590.t3 a_n3565_39590.n11 26.5955
R27464 a_n3565_39590.n8 a_n3565_39590.n2 25.9824
R27465 a_n3565_39590.n0 a_n3565_39590.t5 24.9236
R27466 a_n3565_39590.n0 a_n3565_39590.t6 24.9236
R27467 a_n3565_39590.n1 a_n3565_39590.t4 24.9236
R27468 a_n3565_39590.n1 a_n3565_39590.t7 24.9236
R27469 a_n3565_39590.n8 a_n3565_39590.n7 9.38613
R27470 a_n3565_39590.n5 a_n3565_39590.n4 0.3205
R27471 a_n3565_39590.n6 a_n3565_39590.n5 0.304667
R27472 a_13661_43548.n10 a_13661_43548.t6 323.342
R27473 a_13661_43548.n7 a_13661_43548.t14 293.969
R27474 a_13661_43548.n22 a_13661_43548.n21 287.752
R27475 a_13661_43548.n21 a_13661_43548.n0 277.568
R27476 a_13661_43548.n16 a_13661_43548.t17 256.728
R27477 a_13661_43548.n6 a_13661_43548.t5 241.536
R27478 a_13661_43548.n9 a_13661_43548.t12 241.536
R27479 a_13661_43548.n4 a_13661_43548.t7 241.536
R27480 a_13661_43548.n8 a_13661_43548.t9 236.18
R27481 a_13661_43548.n5 a_13661_43548.n3 212.566
R27482 a_13661_43548.n2 a_13661_43548.t21 212.081
R27483 a_13661_43548.n3 a_13661_43548.t15 212.081
R27484 a_13661_43548.n5 a_13661_43548.n4 203.4
R27485 a_13661_43548.n10 a_13661_43548.t19 194.809
R27486 a_13661_43548.n11 a_13661_43548.n10 190.188
R27487 a_13661_43548.n14 a_13661_43548.n6 177.918
R27488 a_13661_43548.n11 a_13661_43548.n9 176.302
R27489 a_13661_43548.n20 a_13661_43548.n19 169.554
R27490 a_13661_43548.n6 a_13661_43548.t25 169.237
R27491 a_13661_43548.n9 a_13661_43548.t11 169.237
R27492 a_13661_43548.n4 a_13661_43548.t18 169.237
R27493 a_13661_43548.n18 a_13661_43548.n1 167.631
R27494 a_13661_43548.n17 a_13661_43548.n16 166.964
R27495 a_13661_43548.n13 a_13661_43548.n7 164.173
R27496 a_13661_43548.n8 a_13661_43548.t13 163.881
R27497 a_13661_43548.n12 a_13661_43548.n8 162.903
R27498 a_13661_43548.n16 a_13661_43548.t20 161.275
R27499 a_13661_43548.n2 a_13661_43548.t16 139.78
R27500 a_13661_43548.n3 a_13661_43548.t22 139.78
R27501 a_13661_43548.n7 a_13661_43548.t24 138.338
R27502 a_13661_43548.n19 a_13661_43548.t4 137.177
R27503 a_13661_43548.n1 a_13661_43548.t23 137.177
R27504 a_13661_43548.n19 a_13661_43548.t8 121.109
R27505 a_13661_43548.n1 a_13661_43548.t10 121.109
R27506 a_13661_43548.n3 a_13661_43548.n2 62.8066
R27507 a_13661_43548.n15 a_13661_43548.n14 27.2546
R27508 a_13661_43548.t1 a_13661_43548.n22 26.5955
R27509 a_13661_43548.n22 a_13661_43548.t0 26.5955
R27510 a_13661_43548.n21 a_13661_43548.n20 25.5469
R27511 a_13661_43548.n0 a_13661_43548.t3 24.9236
R27512 a_13661_43548.n0 a_13661_43548.t2 24.9236
R27513 a_13661_43548.n12 a_13661_43548.n11 21.8082
R27514 a_13661_43548.n14 a_13661_43548.n13 13.8439
R27515 a_13661_43548.n15 a_13661_43548.n5 7.51989
R27516 a_13661_43548.n20 a_13661_43548.n18 6.84528
R27517 a_13661_43548.n18 a_13661_43548.n17 4.72577
R27518 a_13661_43548.n13 a_13661_43548.n12 2.33292
R27519 a_13661_43548.n17 a_13661_43548.n15 0.779346
R27520 a_n4318_39768.n3 a_n4318_39768.n2 296.139
R27521 a_n4318_39768.n2 a_n4318_39768.n0 269.182
R27522 a_n4318_39768.n1 a_n4318_39768.t4 235.821
R27523 a_n4318_39768.n2 a_n4318_39768.n1 235.451
R27524 a_n4318_39768.n1 a_n4318_39768.t5 163.52
R27525 a_n4318_39768.t1 a_n4318_39768.n3 26.5955
R27526 a_n4318_39768.n3 a_n4318_39768.t0 26.5955
R27527 a_n4318_39768.n0 a_n4318_39768.t2 24.9236
R27528 a_n4318_39768.n0 a_n4318_39768.t3 24.9236
R27529 DATA[5].n6 DATA[5].n5 585
R27530 DATA[5].n2 DATA[5].n0 243.627
R27531 DATA[5].n2 DATA[5].n1 200.262
R27532 DATA[5].n4 DATA[5].n3 194.441
R27533 DATA[5].n6 DATA[5].n4 62.148
R27534 DATA[5].n4 DATA[5].n2 50.5705
R27535 DATA[5].n0 DATA[5].t6 40.0005
R27536 DATA[5].n0 DATA[5].t5 40.0005
R27537 DATA[5].n1 DATA[5].t4 40.0005
R27538 DATA[5].n1 DATA[5].t7 40.0005
R27539 DATA[5].n5 DATA[5].t2 27.5805
R27540 DATA[5].n5 DATA[5].t3 27.5805
R27541 DATA[5].n3 DATA[5].t1 27.5805
R27542 DATA[5].n3 DATA[5].t0 27.5805
R27543 DATA[5] DATA[5].n6 19.8133
R27544 a_8049_45260.n0 a_8049_45260.t3 276.464
R27545 a_8049_45260.n1 a_8049_45260.t5 230.155
R27546 a_8049_45260.n3 a_8049_45260.t1 199.456
R27547 a_8049_45260.n0 a_8049_45260.t4 196.131
R27548 a_8049_45260.n4 a_8049_45260.n3 190.911
R27549 a_8049_45260.n2 a_8049_45260.n0 182.242
R27550 a_8049_45260.n2 a_8049_45260.n1 175.762
R27551 a_8049_45260.n1 a_8049_45260.t6 157.856
R27552 a_8049_45260.n3 a_8049_45260.n2 27.5018
R27553 a_8049_45260.t0 a_8049_45260.n4 26.5955
R27554 a_8049_45260.n4 a_8049_45260.t2 26.5955
R27555 a_11691_44458.n2 a_11691_44458.t4 414.432
R27556 a_11691_44458.n2 a_11691_44458.t7 300.349
R27557 a_11691_44458.n4 a_11691_44458.t8 241.536
R27558 a_11691_44458.n1 a_11691_44458.t9 234.483
R27559 a_11691_44458.n7 a_11691_44458.n6 190.911
R27560 a_11691_44458.n3 a_11691_44458.n1 187.422
R27561 a_11691_44458.n5 a_11691_44458.n4 172.821
R27562 a_11691_44458.n4 a_11691_44458.t5 169.237
R27563 a_11691_44458.n1 a_11691_44458.t6 162.184
R27564 a_11691_44458.n6 a_11691_44458.n0 150.264
R27565 a_11691_44458.n6 a_11691_44458.n5 42.4857
R27566 a_11691_44458.n3 a_11691_44458.n2 37.7163
R27567 a_11691_44458.t1 a_11691_44458.n7 26.5955
R27568 a_11691_44458.n7 a_11691_44458.t0 26.5955
R27569 a_11691_44458.n0 a_11691_44458.t3 24.9236
R27570 a_11691_44458.n0 a_11691_44458.t2 24.9236
R27571 a_11691_44458.n5 a_11691_44458.n3 12.6927
R27572 a_n2442_46660.n3 a_n2442_46660.n2 287.752
R27573 a_n2442_46660.n2 a_n2442_46660.n0 277.568
R27574 a_n2442_46660.n2 a_n2442_46660.n1 273.709
R27575 a_n2442_46660.n1 a_n2442_46660.t4 228.649
R27576 a_n2442_46660.n1 a_n2442_46660.t5 156.35
R27577 a_n2442_46660.t1 a_n2442_46660.n3 26.5955
R27578 a_n2442_46660.n3 a_n2442_46660.t0 26.5955
R27579 a_n2442_46660.n0 a_n2442_46660.t2 24.9236
R27580 a_n2442_46660.n0 a_n2442_46660.t3 24.9236
R27581 a_4185_45028.n2 a_4185_45028.n0 293.272
R27582 a_4185_45028.n0 a_4185_45028.t3 276.464
R27583 a_4185_45028.n1 a_4185_45028.t4 230.155
R27584 a_4185_45028.n3 a_4185_45028.t1 199.456
R27585 a_4185_45028.n0 a_4185_45028.t5 196.131
R27586 a_4185_45028.n4 a_4185_45028.n3 190.911
R27587 a_4185_45028.n2 a_4185_45028.n1 178.535
R27588 a_4185_45028.n1 a_4185_45028.t6 157.856
R27589 a_4185_45028.t0 a_4185_45028.n4 26.5955
R27590 a_4185_45028.n4 a_4185_45028.t2 26.5955
R27591 a_4185_45028.n3 a_4185_45028.n2 18.9814
R27592 a_3537_45260.t22 a_3537_45260.t17 395.01
R27593 a_3537_45260.t26 a_3537_45260.t16 378.255
R27594 a_3537_45260.n20 a_3537_45260.t22 336.003
R27595 a_3537_45260.n21 a_3537_45260.t26 334.733
R27596 a_3537_45260.n23 a_3537_45260.n0 248.087
R27597 a_3537_45260.n17 a_3537_45260.t19 241.536
R27598 a_3537_45260.n15 a_3537_45260.t15 241.536
R27599 a_3537_45260.n12 a_3537_45260.t27 241.536
R27600 a_3537_45260.n5 a_3537_45260.t12 241.536
R27601 a_3537_45260.n8 a_3537_45260.t14 236.18
R27602 a_3537_45260.n6 a_3537_45260.t9 236.18
R27603 a_3537_45260.n4 a_3537_45260.t13 231.835
R27604 a_3537_45260.n10 a_3537_45260.t29 212.081
R27605 a_3537_45260.n11 a_3537_45260.t18 212.081
R27606 a_3537_45260.n24 a_3537_45260.n23 208.506
R27607 a_3537_45260.n13 a_3537_45260.n11 194.209
R27608 a_3537_45260.n9 a_3537_45260.n8 173.3
R27609 a_3537_45260.n18 a_3537_45260.n17 172.821
R27610 a_3537_45260.n13 a_3537_45260.n12 172.246
R27611 a_3537_45260.n7 a_3537_45260.n5 171.75
R27612 a_3537_45260.n19 a_3537_45260.n4 169.841
R27613 a_3537_45260.n17 a_3537_45260.t10 169.237
R27614 a_3537_45260.n15 a_3537_45260.t25 169.237
R27615 a_3537_45260.n12 a_3537_45260.t20 169.237
R27616 a_3537_45260.n5 a_3537_45260.t28 169.237
R27617 a_3537_45260.n7 a_3537_45260.n6 167.987
R27618 a_3537_45260.n16 a_3537_45260.n15 167.934
R27619 a_3537_45260.n8 a_3537_45260.t21 163.881
R27620 a_3537_45260.n6 a_3537_45260.t23 163.881
R27621 a_3537_45260.n4 a_3537_45260.t24 157.07
R27622 a_3537_45260.n10 a_3537_45260.t8 139.78
R27623 a_3537_45260.n11 a_3537_45260.t11 139.78
R27624 a_3537_45260.n3 a_3537_45260.n1 137.576
R27625 a_3537_45260.n3 a_3537_45260.n2 99.1759
R27626 a_3537_45260.n11 a_3537_45260.n10 61.346
R27627 a_3537_45260.n22 a_3537_45260.n3 36.0958
R27628 a_3537_45260.n0 a_3537_45260.t1 26.5955
R27629 a_3537_45260.n0 a_3537_45260.t2 26.5955
R27630 a_3537_45260.n24 a_3537_45260.t0 26.5955
R27631 a_3537_45260.t3 a_3537_45260.n24 26.5955
R27632 a_3537_45260.n1 a_3537_45260.t5 24.9236
R27633 a_3537_45260.n1 a_3537_45260.t4 24.9236
R27634 a_3537_45260.n2 a_3537_45260.t6 24.9236
R27635 a_3537_45260.n2 a_3537_45260.t7 24.9236
R27636 a_3537_45260.n18 a_3537_45260.n16 20.4274
R27637 a_3537_45260.n19 a_3537_45260.n18 17.7726
R27638 a_3537_45260.n23 a_3537_45260.n22 17.2539
R27639 a_3537_45260.n22 a_3537_45260.n21 15.3913
R27640 a_3537_45260.n20 a_3537_45260.n19 15.2725
R27641 a_3537_45260.n14 a_3537_45260.n9 8.92461
R27642 a_3537_45260.n14 a_3537_45260.n13 6.89885
R27643 a_3537_45260.n16 a_3537_45260.n14 5.02935
R27644 a_3537_45260.n21 a_3537_45260.n20 4.5005
R27645 a_3537_45260.n9 a_3537_45260.n7 0.1255
R27646 a_n1151_42308.n17 a_n1151_42308.n16 659.109
R27647 a_n1151_42308.n11 a_n1151_42308.t12 471.289
R27648 a_n1151_42308.n9 a_n1151_42308.t4 471.289
R27649 a_n1151_42308.n7 a_n1151_42308.t7 471.289
R27650 a_n1151_42308.n5 a_n1151_42308.t16 471.289
R27651 a_n1151_42308.n2 a_n1151_42308.t6 471.289
R27652 a_n1151_42308.n3 a_n1151_42308.t10 414.432
R27653 a_n1151_42308.n1 a_n1151_42308.t11 414.432
R27654 a_n1151_42308.n3 a_n1151_42308.t18 300.349
R27655 a_n1151_42308.n1 a_n1151_42308.t9 300.349
R27656 a_n1151_42308.n13 a_n1151_42308.t17 256.07
R27657 a_n1151_42308.n16 a_n1151_42308.n0 219.663
R27658 a_n1151_42308.n4 a_n1151_42308.n2 191.392
R27659 a_n1151_42308.n14 a_n1151_42308.n13 177.833
R27660 a_n1151_42308.n8 a_n1151_42308.n7 175.936
R27661 a_n1151_42308.n10 a_n1151_42308.n9 171.076
R27662 a_n1151_42308.n6 a_n1151_42308.n5 171.076
R27663 a_n1151_42308.n12 a_n1151_42308.n11 171.035
R27664 a_n1151_42308.n13 a_n1151_42308.t14 150.03
R27665 a_n1151_42308.n11 a_n1151_42308.t13 148.35
R27666 a_n1151_42308.n9 a_n1151_42308.t5 148.35
R27667 a_n1151_42308.n7 a_n1151_42308.t8 148.35
R27668 a_n1151_42308.n5 a_n1151_42308.t19 148.35
R27669 a_n1151_42308.n2 a_n1151_42308.t15 148.35
R27670 a_n1151_42308.n15 a_n1151_42308.n1 81.3745
R27671 a_n1151_42308.n0 a_n1151_42308.t2 38.5719
R27672 a_n1151_42308.n0 a_n1151_42308.t3 38.5719
R27673 a_n1151_42308.n4 a_n1151_42308.n3 33.2163
R27674 a_n1151_42308.n16 a_n1151_42308.n15 29.5163
R27675 a_n1151_42308.t1 a_n1151_42308.n17 26.5955
R27676 a_n1151_42308.n17 a_n1151_42308.t0 26.5955
R27677 a_n1151_42308.n15 a_n1151_42308.n14 16.0761
R27678 a_n1151_42308.n12 a_n1151_42308.n10 14.7159
R27679 a_n1151_42308.n6 a_n1151_42308.n4 14.7132
R27680 a_n1151_42308.n10 a_n1151_42308.n8 10.0982
R27681 a_n1151_42308.n14 a_n1151_42308.n12 8.84913
R27682 a_n1151_42308.n8 a_n1151_42308.n6 2.75891
R27683 a_17730_32519.n2 a_17730_32519.t4 1415.15
R27684 a_17730_32519.n1 a_17730_32519.t6 1330.32
R27685 a_17730_32519.n0 a_17730_32519.t5 1320.68
R27686 a_17730_32519.n2 a_17730_32519.t7 1320.68
R27687 a_17730_32519.n6 a_17730_32519.n5 380.32
R27688 a_17730_32519.n5 a_17730_32519.n4 185
R27689 a_17730_32519.n3 a_17730_32519.n0 161.764
R27690 a_17730_32519.n3 a_17730_32519.n2 161.3
R27691 a_17730_32519.n5 a_17730_32519.n3 117.606
R27692 a_17730_32519.n2 a_17730_32519.n1 84.8325
R27693 a_17730_32519.n1 a_17730_32519.n0 84.8325
R27694 a_17730_32519.n6 a_17730_32519.t0 26.5955
R27695 a_17730_32519.t1 a_17730_32519.n6 26.5955
R27696 a_17730_32519.n4 a_17730_32519.t3 24.9236
R27697 a_17730_32519.n4 a_17730_32519.t2 24.9236
R27698 EN_VIN_BSTR_N.n20 EN_VIN_BSTR_N.t18 1559.46
R27699 EN_VIN_BSTR_N.n19 EN_VIN_BSTR_N.t11 1415.15
R27700 EN_VIN_BSTR_N.n19 EN_VIN_BSTR_N.t15 1320.68
R27701 EN_VIN_BSTR_N.n4 EN_VIN_BSTR_N.t16 748.122
R27702 EN_VIN_BSTR_N.n4 EN_VIN_BSTR_N.t22 678.014
R27703 EN_VIN_BSTR_N.n11 EN_VIN_BSTR_N.t12 605.802
R27704 EN_VIN_BSTR_N.n10 EN_VIN_BSTR_N.t8 444.502
R27705 EN_VIN_BSTR_N.n5 EN_VIN_BSTR_N.t13 398.577
R27706 EN_VIN_BSTR_N.n9 EN_VIN_BSTR_N.t17 382.812
R27707 EN_VIN_BSTR_N.n17 EN_VIN_BSTR_N.t19 381.798
R27708 EN_VIN_BSTR_N.n9 EN_VIN_BSTR_N.t21 381.793
R27709 EN_VIN_BSTR_N.n16 EN_VIN_BSTR_N.t23 381.788
R27710 EN_VIN_BSTR_N.n15 EN_VIN_BSTR_N.t10 381.413
R27711 EN_VIN_BSTR_N.n14 EN_VIN_BSTR_N.t20 381.413
R27712 EN_VIN_BSTR_N.n13 EN_VIN_BSTR_N.t9 381.413
R27713 EN_VIN_BSTR_N.n12 EN_VIN_BSTR_N.t14 381.413
R27714 EN_VIN_BSTR_N.n10 EN_VIN_BSTR_N.t7 356.68
R27715 EN_VIN_BSTR_N.n5 EN_VIN_BSTR_N.n4 176.941
R27716 EN_VIN_BSTR_N.n11 EN_VIN_BSTR_N.n10 161.768
R27717 EN_VIN_BSTR_N.n20 EN_VIN_BSTR_N.n19 161.3
R27718 EN_VIN_BSTR_N.n7 EN_VIN_BSTR_N.n2 56.3527
R27719 EN_VIN_BSTR_N.n6 EN_VIN_BSTR_N.n3 56.3527
R27720 EN_VIN_BSTR_N.n21 EN_VIN_BSTR_N.n18 28.2777
R27721 EN_VIN_BSTR_N EN_VIN_BSTR_N.n21 26.0382
R27722 EN_VIN_BSTR_N.n0 EN_VIN_BSTR_N.t2 24.8342
R27723 EN_VIN_BSTR_N.n0 EN_VIN_BSTR_N.t1 24.1879
R27724 EN_VIN_BSTR_N.n1 EN_VIN_BSTR_N.t0 24.1612
R27725 EN_VIN_BSTR_N.n2 EN_VIN_BSTR_N.t4 8.12675
R27726 EN_VIN_BSTR_N.n2 EN_VIN_BSTR_N.t5 8.12675
R27727 EN_VIN_BSTR_N.n3 EN_VIN_BSTR_N.t6 8.12675
R27728 EN_VIN_BSTR_N.n3 EN_VIN_BSTR_N.t3 8.12675
R27729 EN_VIN_BSTR_N.n21 EN_VIN_BSTR_N.n20 4.51508
R27730 EN_VIN_BSTR_N EN_VIN_BSTR_N.n8 4.0544
R27731 EN_VIN_BSTR_N.n6 EN_VIN_BSTR_N.n5 2.39112
R27732 EN_VIN_BSTR_N.n8 EN_VIN_BSTR_N.n7 1.18584
R27733 EN_VIN_BSTR_N.n1 EN_VIN_BSTR_N.n0 0.989971
R27734 EN_VIN_BSTR_N.n17 EN_VIN_BSTR_N.n16 0.9005
R27735 EN_VIN_BSTR_N.n18 EN_VIN_BSTR_N.n17 0.7005
R27736 EN_VIN_BSTR_N.n13 EN_VIN_BSTR_N.n12 0.512318
R27737 EN_VIN_BSTR_N.n14 EN_VIN_BSTR_N.n13 0.512318
R27738 EN_VIN_BSTR_N.n15 EN_VIN_BSTR_N.n14 0.512318
R27739 EN_VIN_BSTR_N.n7 EN_VIN_BSTR_N.n6 0.462038
R27740 EN_VIN_BSTR_N.n18 EN_VIN_BSTR_N.n9 0.3755
R27741 EN_VIN_BSTR_N.n12 EN_VIN_BSTR_N.n11 0.267318
R27742 EN_VIN_BSTR_N.n16 EN_VIN_BSTR_N.n15 0.138909
R27743 EN_VIN_BSTR_N.n8 EN_VIN_BSTR_N.n1 0.018
R27744 a_10890_34112.n16 a_10890_34112.n15 21.0507
R27745 a_10890_34112.n17 a_10890_34112.n16 20.1816
R27746 a_10890_34112.t6 a_10890_34112.n1 9.23464
R27747 a_10890_34112.n12 a_10890_34112.t6 9.23464
R27748 a_10890_34112.n6 a_10890_34112.t7 9.23464
R27749 a_10890_34112.t7 a_10890_34112.n5 9.23464
R27750 a_10890_34112.t4 a_10890_34112.n6 9.23464
R27751 a_10890_34112.n7 a_10890_34112.t4 9.23464
R27752 a_10890_34112.n12 a_10890_34112.t5 9.23464
R27753 a_10890_34112.t5 a_10890_34112.n0 9.23464
R27754 a_10890_34112.n16 a_10890_34112.n14 8.608
R27755 a_10890_34112.n13 a_10890_34112.n1 7.21068
R27756 a_10890_34112.n5 a_10890_34112.n3 6.97192
R27757 a_10890_34112.n14 a_10890_34112.n0 6.82478
R27758 a_10890_34112.n10 a_10890_34112.n1 5.37812
R27759 a_10890_34112.n15 a_10890_34112.t2 4.9505
R27760 a_10890_34112.n15 a_10890_34112.t3 4.9505
R27761 a_10890_34112.n17 a_10890_34112.t1 4.9505
R27762 a_10890_34112.t0 a_10890_34112.n17 4.9505
R27763 a_10890_34112.n7 a_10890_34112.n4 4.27043
R27764 a_10890_34112.n5 a_10890_34112.n4 4.26906
R27765 a_10890_34112.n8 a_10890_34112.n7 3.68933
R27766 a_10890_34112.n13 a_10890_34112.n12 3.36562
R27767 a_10890_34112.n8 a_10890_34112.n3 3.27354
R27768 a_10890_34112.n10 a_10890_34112.n9 3.26815
R27769 a_10890_34112.n9 a_10890_34112.n8 3.08438
R27770 a_10890_34112.n6 a_10890_34112.n4 2.53415
R27771 a_10890_34112.n3 a_10890_34112.n2 2.24437
R27772 a_10890_34112.n11 a_10890_34112.n10 2.23841
R27773 a_10890_34112.n9 a_10890_34112.n0 2.1614
R27774 a_10890_34112.n6 a_10890_34112.n2 1.07306
R27775 a_10890_34112.n11 a_10890_34112.n2 0.911511
R27776 a_10890_34112.n12 a_10890_34112.n11 0.624254
R27777 a_10890_34112.n14 a_10890_34112.n13 0.34925
R27778 VIN_N.n2 VIN_N.t6 92.1604
R27779 VIN_N.n4 VIN_N.t8 91.0227
R27780 VIN_N.n8 VIN_N.t14 90.7102
R27781 VIN_N.n7 VIN_N.t9 90.7102
R27782 VIN_N.n6 VIN_N.t15 90.7102
R27783 VIN_N.n5 VIN_N.t11 90.7102
R27784 VIN_N.n2 VIN_N.t13 90.6265
R27785 VIN_N.n3 VIN_N.t10 90.6219
R27786 VIN_N.n11 VIN_N.t0 47.4586
R27787 VIN_N.n10 VIN_N.n9 37.5586
R27788 VIN_N.n14 VIN_N.n13 29.098
R27789 VIN_N.n0 VIN_N.t2 25.3459
R27790 VIN_N.n0 VIN_N.t3 25.1227
R27791 VIN_N.n14 VIN_N.n0 20.9238
R27792 VIN_N VIN_N.n14 20.705
R27793 VIN_N.n13 VIN_N.t4 16.5266
R27794 VIN_N.n12 VIN_N.n1 14.0516
R27795 VIN_N.n12 VIN_N.n11 11.2899
R27796 VIN_N.n9 VIN_N.t1 9.9005
R27797 VIN_N.n9 VIN_N.t12 9.9005
R27798 VIN_N.n1 VIN_N.t5 2.4755
R27799 VIN_N.n1 VIN_N.t7 2.4755
R27800 VIN_N.n3 VIN_N.n2 1.6255
R27801 VIN_N.n4 VIN_N.n3 1.2505
R27802 VIN_N.n10 VIN_N.n8 0.8755
R27803 VIN_N.n6 VIN_N.n5 0.563
R27804 VIN_N.n7 VIN_N.n6 0.563
R27805 VIN_N.n8 VIN_N.n7 0.563
R27806 VIN_N.n11 VIN_N.n10 0.453625
R27807 VIN_N.n13 VIN_N.n12 0.438
R27808 VIN_N.n5 VIN_N.n4 0.2505
R27809 a_4223_44672.t4 a_4223_44672.t8 378.255
R27810 a_4223_44672.n4 a_4223_44672.t4 368.628
R27811 a_4223_44672.n1 a_4223_44672.t7 241.536
R27812 a_4223_44672.n2 a_4223_44672.t5 231.835
R27813 a_4223_44672.n6 a_4223_44672.n5 190.911
R27814 a_4223_44672.n1 a_4223_44672.t6 169.237
R27815 a_4223_44672.n3 a_4223_44672.n1 169.059
R27816 a_4223_44672.n3 a_4223_44672.n2 167.75
R27817 a_4223_44672.n2 a_4223_44672.t9 157.07
R27818 a_4223_44672.n5 a_4223_44672.n0 150.263
R27819 a_4223_44672.t1 a_4223_44672.n6 26.5955
R27820 a_4223_44672.n6 a_4223_44672.t0 26.5955
R27821 a_4223_44672.n0 a_4223_44672.t3 24.9236
R27822 a_4223_44672.n0 a_4223_44672.t2 24.9236
R27823 a_4223_44672.n5 a_4223_44672.n4 23.3827
R27824 a_4223_44672.n4 a_4223_44672.n3 11.9043
R27825 a_3422_30871.n19 a_3422_30871.t15 1421.83
R27826 a_3422_30871.n9 a_3422_30871.t16 1421.83
R27827 a_3422_30871.n12 a_3422_30871.t17 1327.11
R27828 a_3422_30871.n16 a_3422_30871.t5 1327.11
R27829 a_3422_30871.n18 a_3422_30871.t10 1327.11
R27830 a_3422_30871.n8 a_3422_30871.t12 1327.11
R27831 a_3422_30871.n6 a_3422_30871.t6 1327.11
R27832 a_3422_30871.n2 a_3422_30871.t13 1327.11
R27833 a_3422_30871.n19 a_3422_30871.t9 1320.68
R27834 a_3422_30871.n17 a_3422_30871.t18 1320.68
R27835 a_3422_30871.n15 a_3422_30871.t19 1320.68
R27836 a_3422_30871.n13 a_3422_30871.t21 1320.68
R27837 a_3422_30871.n3 a_3422_30871.t8 1320.68
R27838 a_3422_30871.n5 a_3422_30871.t7 1320.68
R27839 a_3422_30871.n7 a_3422_30871.t20 1320.68
R27840 a_3422_30871.n9 a_3422_30871.t11 1320.68
R27841 a_3422_30871.n25 a_3422_30871.n24 296.139
R27842 a_3422_30871.n24 a_3422_30871.n0 269.182
R27843 a_3422_30871.n22 a_3422_30871.t14 260.322
R27844 a_3422_30871.n23 a_3422_30871.n22 185.969
R27845 a_3422_30871.n22 a_3422_30871.t4 175.169
R27846 a_3422_30871.n14 a_3422_30871.n13 161.701
R27847 a_3422_30871.n4 a_3422_30871.n3 161.701
R27848 a_3422_30871.n20 a_3422_30871.n19 161.3
R27849 a_3422_30871.n15 a_3422_30871.n14 161.3
R27850 a_3422_30871.n17 a_3422_30871.n11 161.3
R27851 a_3422_30871.n10 a_3422_30871.n9 161.3
R27852 a_3422_30871.n7 a_3422_30871.n1 161.3
R27853 a_3422_30871.n5 a_3422_30871.n4 161.3
R27854 a_3422_30871.n13 a_3422_30871.n12 94.7191
R27855 a_3422_30871.n15 a_3422_30871.n12 94.7191
R27856 a_3422_30871.n16 a_3422_30871.n15 94.7191
R27857 a_3422_30871.n17 a_3422_30871.n16 94.7191
R27858 a_3422_30871.n18 a_3422_30871.n17 94.7191
R27859 a_3422_30871.n19 a_3422_30871.n18 94.7191
R27860 a_3422_30871.n9 a_3422_30871.n8 94.7191
R27861 a_3422_30871.n8 a_3422_30871.n7 94.7191
R27862 a_3422_30871.n7 a_3422_30871.n6 94.7191
R27863 a_3422_30871.n6 a_3422_30871.n5 94.7191
R27864 a_3422_30871.n5 a_3422_30871.n2 94.7191
R27865 a_3422_30871.n3 a_3422_30871.n2 94.7191
R27866 a_3422_30871.n23 a_3422_30871.n21 88.0407
R27867 a_3422_30871.n21 a_3422_30871.n20 42.689
R27868 a_3422_30871.n21 a_3422_30871.n10 38.4682
R27869 a_3422_30871.n25 a_3422_30871.t0 26.5955
R27870 a_3422_30871.t1 a_3422_30871.n25 26.5955
R27871 a_3422_30871.n0 a_3422_30871.t2 24.9236
R27872 a_3422_30871.n0 a_3422_30871.t3 24.9236
R27873 a_3422_30871.n24 a_3422_30871.n23 24.5919
R27874 a_3422_30871.n14 a_3422_30871.n11 0.4005
R27875 a_3422_30871.n20 a_3422_30871.n11 0.4005
R27876 a_3422_30871.n10 a_3422_30871.n1 0.4005
R27877 a_3422_30871.n4 a_3422_30871.n1 0.4005
R27878 SMPL_ON_N.n7 SMPL_ON_N.t8 260.322
R27879 SMPL_ON_N.n5 SMPL_ON_N.n3 244.067
R27880 SMPL_ON_N.n2 SMPL_ON_N.n0 236.589
R27881 SMPL_ON_N.n5 SMPL_ON_N.n4 204.893
R27882 SMPL_ON_N.n2 SMPL_ON_N.n1 200.321
R27883 SMPL_ON_N SMPL_ON_N.n7 177.627
R27884 SMPL_ON_N.n7 SMPL_ON_N.t9 175.169
R27885 SMPL_ON_N SMPL_ON_N.n6 70.2992
R27886 SMPL_ON_N.n6 SMPL_ON_N.n5 27.3804
R27887 SMPL_ON_N.n4 SMPL_ON_N.t0 26.5955
R27888 SMPL_ON_N.n4 SMPL_ON_N.t2 26.5955
R27889 SMPL_ON_N.n3 SMPL_ON_N.t1 26.5955
R27890 SMPL_ON_N.n3 SMPL_ON_N.t3 26.5955
R27891 SMPL_ON_N.n0 SMPL_ON_N.t7 24.9236
R27892 SMPL_ON_N.n0 SMPL_ON_N.t5 24.9236
R27893 SMPL_ON_N.n1 SMPL_ON_N.t4 24.9236
R27894 SMPL_ON_N.n1 SMPL_ON_N.t6 24.9236
R27895 SMPL_ON_N.n6 SMPL_ON_N.n2 24.8775
R27896 a_4646_46812.n2 a_4646_46812.n0 333.392
R27897 a_4646_46812.n2 a_4646_46812.n1 301.392
R27898 a_4646_46812.n4 a_4646_46812.n3 301.392
R27899 a_4646_46812.n6 a_4646_46812.n5 301.392
R27900 a_4646_46812.n8 a_4646_46812.n7 301.392
R27901 a_4646_46812.n39 a_4646_46812.n38 301.392
R27902 a_4646_46812.n37 a_4646_46812.n21 297.863
R27903 a_4646_46812.n12 a_4646_46812.t40 294.557
R27904 a_4646_46812.n9 a_4646_46812.t34 294.557
R27905 a_4646_46812.n10 a_4646_46812.t41 294.557
R27906 a_4646_46812.n14 a_4646_46812.t32 294.557
R27907 a_4646_46812.n15 a_4646_46812.t39 294.557
R27908 a_4646_46812.n19 a_4646_46812.n18 287.303
R27909 a_4646_46812.n24 a_4646_46812.n22 248.638
R27910 a_4646_46812.n12 a_4646_46812.t36 211.01
R27911 a_4646_46812.n9 a_4646_46812.t37 211.01
R27912 a_4646_46812.n10 a_4646_46812.t33 211.01
R27913 a_4646_46812.n14 a_4646_46812.t35 211.01
R27914 a_4646_46812.n15 a_4646_46812.t38 211.01
R27915 a_4646_46812.n24 a_4646_46812.n23 203.463
R27916 a_4646_46812.n26 a_4646_46812.n25 203.463
R27917 a_4646_46812.n30 a_4646_46812.n29 203.463
R27918 a_4646_46812.n32 a_4646_46812.n31 203.463
R27919 a_4646_46812.n34 a_4646_46812.n33 203.463
R27920 a_4646_46812.n28 a_4646_46812.n27 202.456
R27921 a_4646_46812.n36 a_4646_46812.n35 200.212
R27922 a_4646_46812.n11 a_4646_46812.n10 187.215
R27923 a_4646_46812.n16 a_4646_46812.n14 181.066
R27924 a_4646_46812.n13 a_4646_46812.n12 180.447
R27925 a_4646_46812.n16 a_4646_46812.n15 176.706
R27926 a_4646_46812.n11 a_4646_46812.n9 162.398
R27927 a_4646_46812.n26 a_4646_46812.n24 45.177
R27928 a_4646_46812.n32 a_4646_46812.n30 45.177
R27929 a_4646_46812.n34 a_4646_46812.n32 45.177
R27930 a_4646_46812.n28 a_4646_46812.n26 44.0476
R27931 a_4646_46812.n30 a_4646_46812.n28 44.0476
R27932 a_4646_46812.n22 a_4646_46812.t26 40.0005
R27933 a_4646_46812.n22 a_4646_46812.t17 40.0005
R27934 a_4646_46812.n23 a_4646_46812.t19 40.0005
R27935 a_4646_46812.n23 a_4646_46812.t30 40.0005
R27936 a_4646_46812.n25 a_4646_46812.t25 40.0005
R27937 a_4646_46812.n25 a_4646_46812.t21 40.0005
R27938 a_4646_46812.n27 a_4646_46812.t27 40.0005
R27939 a_4646_46812.n27 a_4646_46812.t23 40.0005
R27940 a_4646_46812.n29 a_4646_46812.t16 40.0005
R27941 a_4646_46812.n29 a_4646_46812.t28 40.0005
R27942 a_4646_46812.n31 a_4646_46812.t29 40.0005
R27943 a_4646_46812.n31 a_4646_46812.t31 40.0005
R27944 a_4646_46812.n33 a_4646_46812.t18 40.0005
R27945 a_4646_46812.n33 a_4646_46812.t20 40.0005
R27946 a_4646_46812.n35 a_4646_46812.t24 40.0005
R27947 a_4646_46812.n35 a_4646_46812.t22 40.0005
R27948 a_4646_46812.n4 a_4646_46812.n2 32.0005
R27949 a_4646_46812.n6 a_4646_46812.n4 32.0005
R27950 a_4646_46812.n20 a_4646_46812.n8 32.0005
R27951 a_4646_46812.n38 a_4646_46812.n20 32.0005
R27952 a_4646_46812.n8 a_4646_46812.n6 31.2005
R27953 a_4646_46812.n19 a_4646_46812.n17 28.9224
R27954 a_4646_46812.n0 a_4646_46812.t4 27.5805
R27955 a_4646_46812.n0 a_4646_46812.t10 27.5805
R27956 a_4646_46812.n1 a_4646_46812.t9 27.5805
R27957 a_4646_46812.n1 a_4646_46812.t12 27.5805
R27958 a_4646_46812.n3 a_4646_46812.t7 27.5805
R27959 a_4646_46812.n3 a_4646_46812.t0 27.5805
R27960 a_4646_46812.n5 a_4646_46812.t2 27.5805
R27961 a_4646_46812.n5 a_4646_46812.t6 27.5805
R27962 a_4646_46812.n7 a_4646_46812.t11 27.5805
R27963 a_4646_46812.n7 a_4646_46812.t5 27.5805
R27964 a_4646_46812.n18 a_4646_46812.t13 27.5805
R27965 a_4646_46812.n18 a_4646_46812.t14 27.5805
R27966 a_4646_46812.n21 a_4646_46812.t3 27.5805
R27967 a_4646_46812.n21 a_4646_46812.t1 27.5805
R27968 a_4646_46812.t15 a_4646_46812.n39 27.5805
R27969 a_4646_46812.n39 a_4646_46812.t8 27.5805
R27970 a_4646_46812.n20 a_4646_46812.n19 14.0898
R27971 a_4646_46812.n36 a_4646_46812.n34 13.177
R27972 a_4646_46812.n38 a_4646_46812.n37 10.4484
R27973 a_4646_46812.n17 a_4646_46812.n16 9.52935
R27974 a_4646_46812.n13 a_4646_46812.n11 8.9222
R27975 a_4646_46812.n37 a_4646_46812.n36 8.62539
R27976 a_4646_46812.n17 a_4646_46812.n13 4.11863
R27977 a_18114_32519.n9 a_18114_32519.t11 1415.15
R27978 a_18114_32519.n8 a_18114_32519.t5 1330.32
R27979 a_18114_32519.n6 a_18114_32519.t9 1330.32
R27980 a_18114_32519.n2 a_18114_32519.t7 1330.32
R27981 a_18114_32519.n3 a_18114_32519.t10 1320.68
R27982 a_18114_32519.n5 a_18114_32519.t4 1320.68
R27983 a_18114_32519.n7 a_18114_32519.t6 1320.68
R27984 a_18114_32519.n9 a_18114_32519.t8 1320.68
R27985 a_18114_32519.n12 a_18114_32519.n11 287.752
R27986 a_18114_32519.n11 a_18114_32519.n0 277.568
R27987 a_18114_32519.n4 a_18114_32519.n3 161.78
R27988 a_18114_32519.n5 a_18114_32519.n4 161.3
R27989 a_18114_32519.n7 a_18114_32519.n1 161.3
R27990 a_18114_32519.n10 a_18114_32519.n9 161.3
R27991 a_18114_32519.n11 a_18114_32519.n10 125.153
R27992 a_18114_32519.n9 a_18114_32519.n8 84.8325
R27993 a_18114_32519.n8 a_18114_32519.n7 84.8325
R27994 a_18114_32519.n7 a_18114_32519.n6 84.8325
R27995 a_18114_32519.n6 a_18114_32519.n5 84.8325
R27996 a_18114_32519.n5 a_18114_32519.n2 84.8325
R27997 a_18114_32519.n3 a_18114_32519.n2 84.8325
R27998 a_18114_32519.n12 a_18114_32519.t0 26.5955
R27999 a_18114_32519.t1 a_18114_32519.n12 26.5955
R28000 a_18114_32519.n0 a_18114_32519.t2 24.9236
R28001 a_18114_32519.n0 a_18114_32519.t3 24.9236
R28002 a_18114_32519.n4 a_18114_32519.n1 0.4805
R28003 a_18114_32519.n10 a_18114_32519.n1 0.4655
R28004 VREF_GND VREF_GND.n43 56.7552
R28005 VREF_GND VREF_GND.n21 56.5923
R28006 VREF_GND.n0 VREF_GND.t21 47.7249
R28007 VREF_GND.n22 VREF_GND.t45 47.7249
R28008 VREF_GND.n6 VREF_GND.t20 47.1624
R28009 VREF_GND.n3 VREF_GND.t32 47.1624
R28010 VREF_GND.n2 VREF_GND.t33 47.1624
R28011 VREF_GND.n1 VREF_GND.t18 47.1624
R28012 VREF_GND.n0 VREF_GND.t44 47.1624
R28013 VREF_GND.n28 VREF_GND.t4 47.1624
R28014 VREF_GND.n25 VREF_GND.t24 47.1624
R28015 VREF_GND.n24 VREF_GND.t43 47.1624
R28016 VREF_GND.n23 VREF_GND.t27 47.1624
R28017 VREF_GND.n22 VREF_GND.t25 47.1624
R28018 VREF_GND.n5 VREF_GND.n4 37.2624
R28019 VREF_GND.n27 VREF_GND.n26 37.2624
R28020 VREF_GND.n8 VREF_GND.n6 23.1134
R28021 VREF_GND.n30 VREF_GND.n28 23.1134
R28022 VREF_GND.n21 VREF_GND.t17 16.1734
R28023 VREF_GND.n43 VREF_GND.t38 16.1734
R28024 VREF_GND.n20 VREF_GND.n19 13.6984
R28025 VREF_GND.n18 VREF_GND.n17 13.6984
R28026 VREF_GND.n16 VREF_GND.n15 13.6984
R28027 VREF_GND.n14 VREF_GND.n13 13.6984
R28028 VREF_GND.n12 VREF_GND.n11 13.6984
R28029 VREF_GND.n10 VREF_GND.n9 13.6984
R28030 VREF_GND.n8 VREF_GND.n7 13.6984
R28031 VREF_GND.n42 VREF_GND.n41 13.6984
R28032 VREF_GND.n40 VREF_GND.n39 13.6984
R28033 VREF_GND.n38 VREF_GND.n37 13.6984
R28034 VREF_GND.n36 VREF_GND.n35 13.6984
R28035 VREF_GND.n34 VREF_GND.n33 13.6984
R28036 VREF_GND.n32 VREF_GND.n31 13.6984
R28037 VREF_GND.n30 VREF_GND.n29 13.6984
R28038 VREF_GND.n4 VREF_GND.t19 9.9005
R28039 VREF_GND.n4 VREF_GND.t23 9.9005
R28040 VREF_GND.n26 VREF_GND.t26 9.9005
R28041 VREF_GND.n26 VREF_GND.t5 9.9005
R28042 VREF_GND.n19 VREF_GND.t11 2.4755
R28043 VREF_GND.n19 VREF_GND.t10 2.4755
R28044 VREF_GND.n17 VREF_GND.t15 2.4755
R28045 VREF_GND.n17 VREF_GND.t14 2.4755
R28046 VREF_GND.n15 VREF_GND.t16 2.4755
R28047 VREF_GND.n15 VREF_GND.t13 2.4755
R28048 VREF_GND.n13 VREF_GND.t12 2.4755
R28049 VREF_GND.n13 VREF_GND.t6 2.4755
R28050 VREF_GND.n11 VREF_GND.t9 2.4755
R28051 VREF_GND.n11 VREF_GND.t7 2.4755
R28052 VREF_GND.n9 VREF_GND.t8 2.4755
R28053 VREF_GND.n9 VREF_GND.t30 2.4755
R28054 VREF_GND.n7 VREF_GND.t31 2.4755
R28055 VREF_GND.n7 VREF_GND.t22 2.4755
R28056 VREF_GND.n41 VREF_GND.t41 2.4755
R28057 VREF_GND.n41 VREF_GND.t36 2.4755
R28058 VREF_GND.n39 VREF_GND.t37 2.4755
R28059 VREF_GND.n39 VREF_GND.t35 2.4755
R28060 VREF_GND.n37 VREF_GND.t34 2.4755
R28061 VREF_GND.n37 VREF_GND.t39 2.4755
R28062 VREF_GND.n35 VREF_GND.t1 2.4755
R28063 VREF_GND.n35 VREF_GND.t40 2.4755
R28064 VREF_GND.n33 VREF_GND.t0 2.4755
R28065 VREF_GND.n33 VREF_GND.t2 2.4755
R28066 VREF_GND.n31 VREF_GND.t29 2.4755
R28067 VREF_GND.n31 VREF_GND.t3 2.4755
R28068 VREF_GND.n29 VREF_GND.t42 2.4755
R28069 VREF_GND.n29 VREF_GND.t28 2.4755
R28070 VREF_GND.n1 VREF_GND.n0 0.563
R28071 VREF_GND.n2 VREF_GND.n1 0.563
R28072 VREF_GND.n3 VREF_GND.n2 0.563
R28073 VREF_GND.n5 VREF_GND.n3 0.563
R28074 VREF_GND.n23 VREF_GND.n22 0.563
R28075 VREF_GND.n24 VREF_GND.n23 0.563
R28076 VREF_GND.n25 VREF_GND.n24 0.563
R28077 VREF_GND.n27 VREF_GND.n25 0.563
R28078 VREF_GND.n18 VREF_GND.n16 0.53175
R28079 VREF_GND.n40 VREF_GND.n38 0.53175
R28080 VREF_GND.n6 VREF_GND.n5 0.507196
R28081 VREF_GND.n28 VREF_GND.n27 0.507196
R28082 VREF_GND.n10 VREF_GND.n8 0.5005
R28083 VREF_GND.n12 VREF_GND.n10 0.5005
R28084 VREF_GND.n14 VREF_GND.n12 0.5005
R28085 VREF_GND.n16 VREF_GND.n14 0.5005
R28086 VREF_GND.n20 VREF_GND.n18 0.5005
R28087 VREF_GND.n21 VREF_GND.n20 0.5005
R28088 VREF_GND.n32 VREF_GND.n30 0.5005
R28089 VREF_GND.n34 VREF_GND.n32 0.5005
R28090 VREF_GND.n36 VREF_GND.n34 0.5005
R28091 VREF_GND.n38 VREF_GND.n36 0.5005
R28092 VREF_GND.n42 VREF_GND.n40 0.5005
R28093 VREF_GND.n43 VREF_GND.n42 0.5005
R28094 a_n4209_38216.n4 a_n4209_38216.t10 553.458
R28095 a_n4209_38216.n8 a_n4209_38216.n7 340.637
R28096 a_n4209_38216.n3 a_n4209_38216.t8 241.536
R28097 a_n4209_38216.n7 a_n4209_38216.n6 195.577
R28098 a_n4209_38216.n4 a_n4209_38216.n3 174.202
R28099 a_n4209_38216.n3 a_n4209_38216.t9 169.237
R28100 a_n4209_38216.n2 a_n4209_38216.n0 137.189
R28101 a_n4209_38216.n2 a_n4209_38216.n1 98.787
R28102 a_n4209_38216.n5 a_n4209_38216.n2 38.9679
R28103 a_n4209_38216.n6 a_n4209_38216.t1 26.5955
R28104 a_n4209_38216.n6 a_n4209_38216.t0 26.5955
R28105 a_n4209_38216.n8 a_n4209_38216.t2 26.5955
R28106 a_n4209_38216.t3 a_n4209_38216.n8 26.5955
R28107 a_n4209_38216.n7 a_n4209_38216.n5 26.0391
R28108 a_n4209_38216.n0 a_n4209_38216.t6 24.9236
R28109 a_n4209_38216.n0 a_n4209_38216.t4 24.9236
R28110 a_n4209_38216.n1 a_n4209_38216.t5 24.9236
R28111 a_n4209_38216.n1 a_n4209_38216.t7 24.9236
R28112 a_n4209_38216.n5 a_n4209_38216.n4 9.30997
R28113 a_13747_46662.n9 a_13747_46662.n8 335.983
R28114 a_13747_46662.n8 a_13747_46662.t1 328.421
R28115 a_13747_46662.n5 a_13747_46662.t9 261.887
R28116 a_13747_46662.n0 a_13747_46662.t10 230.363
R28117 a_13747_46662.n4 a_13747_46662.t6 224.984
R28118 a_13747_46662.n3 a_13747_46662.n2 219.293
R28119 a_13747_46662.n1 a_13747_46662.t3 212.081
R28120 a_13747_46662.n2 a_13747_46662.t4 212.081
R28121 a_13747_46662.n4 a_13747_46662.t12 187.714
R28122 a_13747_46662.n6 a_13747_46662.n5 179.061
R28123 a_13747_46662.n3 a_13747_46662.n0 168.323
R28124 a_13747_46662.n6 a_13747_46662.n4 165.323
R28125 a_13747_46662.n0 a_13747_46662.t8 158.064
R28126 a_13747_46662.n5 a_13747_46662.t7 155.847
R28127 a_13747_46662.n1 a_13747_46662.t11 139.78
R28128 a_13747_46662.n2 a_13747_46662.t5 139.78
R28129 a_13747_46662.n2 a_13747_46662.n1 61.346
R28130 a_13747_46662.n9 a_13747_46662.t2 26.5955
R28131 a_13747_46662.t0 a_13747_46662.n9 26.5955
R28132 a_13747_46662.n8 a_13747_46662.n7 24.5342
R28133 a_13747_46662.n7 a_13747_46662.n6 20.6489
R28134 a_13747_46662.n7 a_13747_46662.n3 10.3618
R28135 a_n2956_39768.n3 a_n2956_39768.n2 287.752
R28136 a_n2956_39768.n2 a_n2956_39768.n0 277.568
R28137 a_n2956_39768.n2 a_n2956_39768.n1 261.014
R28138 a_n2956_39768.n1 a_n2956_39768.t5 228.649
R28139 a_n2956_39768.n1 a_n2956_39768.t4 156.35
R28140 a_n2956_39768.n3 a_n2956_39768.t0 26.5955
R28141 a_n2956_39768.t1 a_n2956_39768.n3 26.5955
R28142 a_n2956_39768.n0 a_n2956_39768.t3 24.9236
R28143 a_n2956_39768.n0 a_n2956_39768.t2 24.9236
R28144 DATA[3].n3 DATA[3].n2 647.148
R28145 DATA[3].n5 DATA[3].n4 200.262
R28146 DATA[3].n3 DATA[3].n1 194.441
R28147 DATA[3].n6 DATA[3].n0 185
R28148 DATA[3].n6 DATA[3].n5 58.6278
R28149 DATA[3].n5 DATA[3].n3 50.5705
R28150 DATA[3].n0 DATA[3].t7 40.0005
R28151 DATA[3].n0 DATA[3].t5 40.0005
R28152 DATA[3].n4 DATA[3].t6 40.0005
R28153 DATA[3].n4 DATA[3].t4 40.0005
R28154 DATA[3].n1 DATA[3].t2 27.5805
R28155 DATA[3].n1 DATA[3].t3 27.5805
R28156 DATA[3].n2 DATA[3].t0 27.5805
R28157 DATA[3].n2 DATA[3].t1 27.5805
R28158 DATA[3] DATA[3].n6 18.6693
R28159 a_n97_42460.n21 a_n97_42460.n20 380.32
R28160 a_n97_42460.n15 a_n97_42460.t23 239.505
R28161 a_n97_42460.n12 a_n97_42460.t8 239.505
R28162 a_n97_42460.n10 a_n97_42460.t5 239.505
R28163 a_n97_42460.n1 a_n97_42460.t10 239.505
R28164 a_n97_42460.n7 a_n97_42460.t18 239.505
R28165 a_n97_42460.n5 a_n97_42460.t21 239.505
R28166 a_n97_42460.n2 a_n97_42460.t22 239.505
R28167 a_n97_42460.n0 a_n97_42460.t7 239.505
R28168 a_n97_42460.n16 a_n97_42460.t17 231.017
R28169 a_n97_42460.n3 a_n97_42460.t20 231.017
R28170 a_n97_42460.n13 a_n97_42460.n12 196.069
R28171 a_n97_42460.n11 a_n97_42460.n10 196.069
R28172 a_n97_42460.n14 a_n97_42460.n0 186.174
R28173 a_n97_42460.n6 a_n97_42460.n5 185.987
R28174 a_n97_42460.n20 a_n97_42460.n19 185
R28175 a_n97_42460.n4 a_n97_42460.n2 182.804
R28176 a_n97_42460.n9 a_n97_42460.n1 174.34
R28177 a_n97_42460.n4 a_n97_42460.n3 174.03
R28178 a_n97_42460.n17 a_n97_42460.n15 173.066
R28179 a_n97_42460.n8 a_n97_42460.n7 169.514
R28180 a_n97_42460.n15 a_n97_42460.t4 167.204
R28181 a_n97_42460.n12 a_n97_42460.t16 167.204
R28182 a_n97_42460.n10 a_n97_42460.t9 167.204
R28183 a_n97_42460.n1 a_n97_42460.t6 167.204
R28184 a_n97_42460.n7 a_n97_42460.t19 167.204
R28185 a_n97_42460.n5 a_n97_42460.t15 167.204
R28186 a_n97_42460.n2 a_n97_42460.t13 167.204
R28187 a_n97_42460.n0 a_n97_42460.t14 167.204
R28188 a_n97_42460.n17 a_n97_42460.n16 163.046
R28189 a_n97_42460.n16 a_n97_42460.t12 158.716
R28190 a_n97_42460.n3 a_n97_42460.t11 158.716
R28191 a_n97_42460.n8 a_n97_42460.n6 47.2723
R28192 a_n97_42460.t1 a_n97_42460.n21 26.5955
R28193 a_n97_42460.n21 a_n97_42460.t0 26.5955
R28194 a_n97_42460.n20 a_n97_42460.n18 25.8732
R28195 a_n97_42460.n19 a_n97_42460.t2 24.9236
R28196 a_n97_42460.n19 a_n97_42460.t3 24.9236
R28197 a_n97_42460.n11 a_n97_42460.n9 19.5348
R28198 a_n97_42460.n14 a_n97_42460.n13 18.6173
R28199 a_n97_42460.n18 a_n97_42460.n14 17.8329
R28200 a_n97_42460.n9 a_n97_42460.n8 11.1185
R28201 a_n97_42460.n13 a_n97_42460.n11 7.6722
R28202 a_n97_42460.n18 a_n97_42460.n17 4.79462
R28203 a_n97_42460.n6 a_n97_42460.n4 1.11605
R28204 a_13258_32519.n1 a_13258_32519.t4 694.745
R28205 a_13258_32519.n2 a_13258_32519.n1 287.752
R28206 a_13258_32519.n1 a_13258_32519.n0 277.568
R28207 a_13258_32519.t1 a_13258_32519.n2 26.5955
R28208 a_13258_32519.n2 a_13258_32519.t0 26.5955
R28209 a_13258_32519.n0 a_13258_32519.t2 24.9236
R28210 a_13258_32519.n0 a_13258_32519.t3 24.9236
R28211 a_6171_45002.t0 a_6171_45002.n4 728.274
R28212 a_6171_45002.t0 a_6171_45002.n0 685.292
R28213 a_6171_45002.n0 a_6171_45002.t1 289.469
R28214 a_6171_45002.n1 a_6171_45002.t2 241.536
R28215 a_6171_45002.n2 a_6171_45002.t3 229.369
R28216 a_6171_45002.n3 a_6171_45002.n1 186.169
R28217 a_6171_45002.n3 a_6171_45002.n2 173.899
R28218 a_6171_45002.n1 a_6171_45002.t4 169.237
R28219 a_6171_45002.n2 a_6171_45002.t5 157.07
R28220 a_6171_45002.n4 a_6171_45002.n3 23.0309
R28221 a_6171_45002.n4 a_6171_45002.n0 15.826
R28222 a_n2017_45002.n1 a_n2017_45002.t4 260.322
R28223 a_n2017_45002.n2 a_n2017_45002.n0 238.784
R28224 a_n2017_45002.n2 a_n2017_45002.n1 235.232
R28225 a_n2017_45002.n3 a_n2017_45002.n2 191.194
R28226 a_n2017_45002.n1 a_n2017_45002.t5 175.169
R28227 a_n2017_45002.n3 a_n2017_45002.t0 26.5955
R28228 a_n2017_45002.t1 a_n2017_45002.n3 26.5955
R28229 a_n2017_45002.n0 a_n2017_45002.t2 24.9236
R28230 a_n2017_45002.n0 a_n2017_45002.t3 24.9236
R28231 a_n3674_37592.n3 a_n3674_37592.n2 380.32
R28232 a_n3674_37592.n0 a_n3674_37592.t4 235.821
R28233 a_n3674_37592.n2 a_n3674_37592.n0 235.3
R28234 a_n3674_37592.n2 a_n3674_37592.n1 185
R28235 a_n3674_37592.n0 a_n3674_37592.t5 163.52
R28236 a_n3674_37592.t1 a_n3674_37592.n3 26.5955
R28237 a_n3674_37592.n3 a_n3674_37592.t0 26.5955
R28238 a_n3674_37592.n1 a_n3674_37592.t3 24.9236
R28239 a_n3674_37592.n1 a_n3674_37592.t2 24.9236
R28240 a_n4064_39072.n4 a_n4064_39072.t9 1645.77
R28241 a_n4064_39072.n7 a_n4064_39072.n6 360.399
R28242 a_n4064_39072.n3 a_n4064_39072.t8 241.536
R28243 a_n4064_39072.n2 a_n4064_39072.n1 232.862
R28244 a_n4064_39072.n8 a_n4064_39072.n7 203.161
R28245 a_n4064_39072.n4 a_n4064_39072.n3 172.035
R28246 a_n4064_39072.n3 a_n4064_39072.t10 169.237
R28247 a_n4064_39072.n2 a_n4064_39072.n0 95.6721
R28248 a_n4064_39072.n5 a_n4064_39072.n2 60.5918
R28249 a_n4064_39072.n6 a_n4064_39072.t2 27.5805
R28250 a_n4064_39072.n6 a_n4064_39072.t0 27.5805
R28251 a_n4064_39072.n8 a_n4064_39072.t1 27.5805
R28252 a_n4064_39072.t3 a_n4064_39072.n8 27.5805
R28253 a_n4064_39072.n1 a_n4064_39072.t7 25.8467
R28254 a_n4064_39072.n1 a_n4064_39072.t6 25.8467
R28255 a_n4064_39072.n0 a_n4064_39072.t5 25.8467
R28256 a_n4064_39072.n0 a_n4064_39072.t4 25.8467
R28257 a_n4064_39072.n7 a_n4064_39072.n5 22.6489
R28258 a_n4064_39072.n5 a_n4064_39072.n4 9.40917
R28259 a_n3565_39304.n4 a_n3565_39304.t8 833.053
R28260 a_n3565_39304.n8 a_n3565_39304.n7 340.637
R28261 a_n3565_39304.n3 a_n3565_39304.t10 241.536
R28262 a_n3565_39304.n7 a_n3565_39304.n6 195.577
R28263 a_n3565_39304.n3 a_n3565_39304.t9 169.237
R28264 a_n3565_39304.n4 a_n3565_39304.n3 168.845
R28265 a_n3565_39304.n2 a_n3565_39304.n0 137.189
R28266 a_n3565_39304.n2 a_n3565_39304.n1 98.787
R28267 a_n3565_39304.n7 a_n3565_39304.n5 39.0246
R28268 a_n3565_39304.n6 a_n3565_39304.t2 26.5955
R28269 a_n3565_39304.n6 a_n3565_39304.t0 26.5955
R28270 a_n3565_39304.n8 a_n3565_39304.t1 26.5955
R28271 a_n3565_39304.t3 a_n3565_39304.n8 26.5955
R28272 a_n3565_39304.n5 a_n3565_39304.n2 25.9824
R28273 a_n3565_39304.n0 a_n3565_39304.t4 24.9236
R28274 a_n3565_39304.n0 a_n3565_39304.t7 24.9236
R28275 a_n3565_39304.n1 a_n3565_39304.t5 24.9236
R28276 a_n3565_39304.n1 a_n3565_39304.t6 24.9236
R28277 a_n3565_39304.n5 a_n3565_39304.n4 9.3005
R28278 C6_P_btm.n4 C6_P_btm.t5 97.811
R28279 C6_P_btm.n3 C6_P_btm.t2 68.0518
R28280 C6_P_btm C6_P_btm.n4 57.9172
R28281 C6_P_btm.n2 C6_P_btm.n1 45.0311
R28282 C6_P_btm.n2 C6_P_btm.n0 37.4635
R28283 C6_P_btm.n0 C6_P_btm.t3 9.9005
R28284 C6_P_btm.n0 C6_P_btm.t4 9.9005
R28285 C6_P_btm.n1 C6_P_btm.t1 9.9005
R28286 C6_P_btm.n1 C6_P_btm.t0 9.9005
R28287 C6_P_btm.n4 C6_P_btm.n3 8.0005
R28288 C6_P_btm.n3 C6_P_btm.n2 6.58904
R28289 a_10227_46804.n23 a_10227_46804.t24 408.63
R28290 a_10227_46804.n12 a_10227_46804.t14 408.63
R28291 a_10227_46804.n15 a_10227_46804.t23 408.63
R28292 a_10227_46804.n18 a_10227_46804.t26 408.63
R28293 a_10227_46804.n5 a_10227_46804.t16 408.63
R28294 a_10227_46804.n8 a_10227_46804.t32 408.63
R28295 a_10227_46804.n1 a_10227_46804.t12 408.63
R28296 a_10227_46804.n31 a_10227_46804.n30 380.32
R28297 a_10227_46804.n24 a_10227_46804.t18 347.577
R28298 a_10227_46804.n13 a_10227_46804.t6 347.577
R28299 a_10227_46804.n19 a_10227_46804.t31 347.577
R28300 a_10227_46804.n16 a_10227_46804.t5 347.577
R28301 a_10227_46804.n6 a_10227_46804.t27 347.577
R28302 a_10227_46804.n9 a_10227_46804.t8 347.577
R28303 a_10227_46804.n0 a_10227_46804.t28 347.577
R28304 a_10227_46804.n3 a_10227_46804.t29 238.59
R28305 a_10227_46804.n3 a_10227_46804.t21 203.244
R28306 a_10227_46804.n24 a_10227_46804.t4 193.337
R28307 a_10227_46804.n13 a_10227_46804.t20 193.337
R28308 a_10227_46804.n19 a_10227_46804.t15 193.337
R28309 a_10227_46804.n16 a_10227_46804.t10 193.337
R28310 a_10227_46804.n6 a_10227_46804.t11 193.337
R28311 a_10227_46804.n9 a_10227_46804.t33 193.337
R28312 a_10227_46804.n0 a_10227_46804.t30 193.337
R28313 a_10227_46804.n30 a_10227_46804.n29 185
R28314 a_10227_46804.n14 a_10227_46804.n12 167.808
R28315 a_10227_46804.n25 a_10227_46804.n23 167.666
R28316 a_10227_46804.n7 a_10227_46804.n5 167.666
R28317 a_10227_46804.n10 a_10227_46804.n8 167.663
R28318 a_10227_46804.n20 a_10227_46804.n18 167.603
R28319 a_10227_46804.n4 a_10227_46804.n3 165.343
R28320 a_10227_46804.n2 a_10227_46804.n1 165.077
R28321 a_10227_46804.n17 a_10227_46804.n15 165.049
R28322 a_10227_46804.n17 a_10227_46804.n16 163.196
R28323 a_10227_46804.n2 a_10227_46804.n0 163
R28324 a_10227_46804.n20 a_10227_46804.n19 160.476
R28325 a_10227_46804.n14 a_10227_46804.n13 160.448
R28326 a_10227_46804.n25 a_10227_46804.n24 160.415
R28327 a_10227_46804.n7 a_10227_46804.n6 160.415
R28328 a_10227_46804.n10 a_10227_46804.n9 160.415
R28329 a_10227_46804.n23 a_10227_46804.t13 132.282
R28330 a_10227_46804.n12 a_10227_46804.t9 132.282
R28331 a_10227_46804.n15 a_10227_46804.t17 132.282
R28332 a_10227_46804.n18 a_10227_46804.t25 132.282
R28333 a_10227_46804.n5 a_10227_46804.t19 132.282
R28334 a_10227_46804.n8 a_10227_46804.t22 132.282
R28335 a_10227_46804.n1 a_10227_46804.t7 132.282
R28336 a_10227_46804.n21 a_10227_46804.n20 36.8876
R28337 a_10227_46804.n11 a_10227_46804.n7 31.1142
R28338 a_10227_46804.n31 a_10227_46804.t0 26.5955
R28339 a_10227_46804.t1 a_10227_46804.n31 26.5955
R28340 a_10227_46804.n4 a_10227_46804.n2 24.9964
R28341 a_10227_46804.n29 a_10227_46804.t3 24.9236
R28342 a_10227_46804.n29 a_10227_46804.t2 24.9236
R28343 a_10227_46804.n27 a_10227_46804.n11 18.8555
R28344 a_10227_46804.n26 a_10227_46804.n22 18.6705
R28345 a_10227_46804.n28 a_10227_46804.n4 12.7475
R28346 a_10227_46804.n22 a_10227_46804.n21 10.8576
R28347 a_10227_46804.n30 a_10227_46804.n28 10.3044
R28348 a_10227_46804.n11 a_10227_46804.n10 10.1077
R28349 a_10227_46804.n28 a_10227_46804.n27 9.83292
R28350 a_10227_46804.n27 a_10227_46804.n26 4.503
R28351 a_10227_46804.n22 a_10227_46804.n14 1.61506
R28352 a_10227_46804.n21 a_10227_46804.n17 1.04321
R28353 a_10227_46804.n26 a_10227_46804.n25 0.0476225
R28354 a_7754_40130.n4 a_7754_40130.t12 578.173
R28355 a_7754_40130.t12 a_7754_40130.n3 578.173
R28356 a_7754_40130.n18 a_7754_40130.t11 578.173
R28357 a_7754_40130.n16 a_7754_40130.t11 577.779
R28358 a_7754_40130.n18 a_7754_40130.t9 577.749
R28359 a_7754_40130.t9 a_7754_40130.n17 577.749
R28360 a_7754_40130.n19 a_7754_40130.t13 577.749
R28361 a_7754_40130.t13 a_7754_40130.n14 577.749
R28362 a_7754_40130.t4 a_7754_40130.n20 577.749
R28363 a_7754_40130.n21 a_7754_40130.t4 577.749
R28364 a_7754_40130.t14 a_7754_40130.n13 577.749
R28365 a_7754_40130.n22 a_7754_40130.t14 577.749
R28366 a_7754_40130.n24 a_7754_40130.t8 577.749
R28367 a_7754_40130.t8 a_7754_40130.n23 577.749
R28368 a_7754_40130.n12 a_7754_40130.t0 577.749
R28369 a_7754_40130.t0 a_7754_40130.n11 577.749
R28370 a_7754_40130.t10 a_7754_40130.n1 577.749
R28371 a_7754_40130.n10 a_7754_40130.t10 577.749
R28372 a_7754_40130.t15 a_7754_40130.n8 577.749
R28373 a_7754_40130.n9 a_7754_40130.t15 577.749
R28374 a_7754_40130.n7 a_7754_40130.t5 577.749
R28375 a_7754_40130.t5 a_7754_40130.n2 577.749
R28376 a_7754_40130.n6 a_7754_40130.t7 577.749
R28377 a_7754_40130.t7 a_7754_40130.n5 577.749
R28378 a_7754_40130.t6 a_7754_40130.n3 577.749
R28379 a_7754_40130.n4 a_7754_40130.t6 577.749
R28380 a_7754_40130.n15 a_7754_40130.t2 233.501
R28381 a_7754_40130.n15 a_7754_40130.t3 48.461
R28382 a_7754_40130.t1 a_7754_40130.n26 29.4286
R28383 a_7754_40130.n16 a_7754_40130.n15 9.38245
R28384 a_7754_40130.n26 a_7754_40130.n25 2.29004
R28385 a_7754_40130.n26 a_7754_40130.n0 2.27754
R28386 a_7754_40130.n5 a_7754_40130.n4 0.4255
R28387 a_7754_40130.n5 a_7754_40130.n2 0.4255
R28388 a_7754_40130.n9 a_7754_40130.n2 0.4255
R28389 a_7754_40130.n10 a_7754_40130.n9 0.4255
R28390 a_7754_40130.n11 a_7754_40130.n10 0.4255
R28391 a_7754_40130.n23 a_7754_40130.n22 0.4255
R28392 a_7754_40130.n22 a_7754_40130.n21 0.4255
R28393 a_7754_40130.n21 a_7754_40130.n14 0.4255
R28394 a_7754_40130.n17 a_7754_40130.n14 0.4255
R28395 a_7754_40130.n6 a_7754_40130.n3 0.4255
R28396 a_7754_40130.n7 a_7754_40130.n6 0.4255
R28397 a_7754_40130.n8 a_7754_40130.n7 0.4255
R28398 a_7754_40130.n8 a_7754_40130.n1 0.4255
R28399 a_7754_40130.n12 a_7754_40130.n1 0.4255
R28400 a_7754_40130.n24 a_7754_40130.n13 0.4255
R28401 a_7754_40130.n20 a_7754_40130.n13 0.4255
R28402 a_7754_40130.n20 a_7754_40130.n19 0.4255
R28403 a_7754_40130.n19 a_7754_40130.n18 0.4255
R28404 a_7754_40130.n17 a_7754_40130.n16 0.395812
R28405 a_7754_40130.n23 a_7754_40130.n0 0.303625
R28406 a_7754_40130.n25 a_7754_40130.n24 0.303625
R28407 a_7754_40130.n11 a_7754_40130.n0 0.122375
R28408 a_7754_40130.n25 a_7754_40130.n12 0.122375
R28409 a_11206_38545.n2 a_11206_38545.n1 225.84
R28410 a_11206_38545.n0 a_11206_38545.t3 39.2429
R28411 a_11206_38545.n0 a_11206_38545.t2 34.125
R28412 a_11206_38545.n1 a_11206_38545.t1 34.125
R28413 a_11206_38545.n2 a_11206_38545.t4 28.5655
R28414 a_11206_38545.t0 a_11206_38545.n2 28.5655
R28415 a_11206_38545.n1 a_11206_38545.n0 0.563
R28416 a_3090_45724.n18 a_3090_45724.n0 311.288
R28417 a_3090_45724.n14 a_3090_45724.t20 241.536
R28418 a_3090_45724.n4 a_3090_45724.t19 236.18
R28419 a_3090_45724.n19 a_3090_45724.n18 234.267
R28420 a_3090_45724.n5 a_3090_45724.t15 231.718
R28421 a_3090_45724.n3 a_3090_45724.t18 230.793
R28422 a_3090_45724.n10 a_3090_45724.t14 230.793
R28423 a_3090_45724.n6 a_3090_45724.t11 230.793
R28424 a_3090_45724.n7 a_3090_45724.t21 230.363
R28425 a_3090_45724.n2 a_3090_45724.t10 206.19
R28426 a_3090_45724.n12 a_3090_45724.n4 193.694
R28427 a_3090_45724.n16 a_3090_45724.n2 191.525
R28428 a_3090_45724.n17 a_3090_45724.n1 190.839
R28429 a_3090_45724.n8 a_3090_45724.n6 179.93
R28430 a_3090_45724.n13 a_3090_45724.n3 173.03
R28431 a_3090_45724.n11 a_3090_45724.n10 172.69
R28432 a_3090_45724.n15 a_3090_45724.n14 170.581
R28433 a_3090_45724.n9 a_3090_45724.n5 170.536
R28434 a_3090_45724.n14 a_3090_45724.t6 169.237
R28435 a_3090_45724.n8 a_3090_45724.n7 168.618
R28436 a_3090_45724.n4 a_3090_45724.t7 163.881
R28437 a_3090_45724.n5 a_3090_45724.t16 159.417
R28438 a_3090_45724.n3 a_3090_45724.t13 158.494
R28439 a_3090_45724.n10 a_3090_45724.t8 158.494
R28440 a_3090_45724.n6 a_3090_45724.t9 158.494
R28441 a_3090_45724.n7 a_3090_45724.t12 158.064
R28442 a_3090_45724.n2 a_3090_45724.t17 148.35
R28443 a_3090_45724.n18 a_3090_45724.n17 48.8466
R28444 a_3090_45724.n13 a_3090_45724.n12 35.1042
R28445 a_3090_45724.n0 a_3090_45724.t3 32.5055
R28446 a_3090_45724.n0 a_3090_45724.t2 32.5055
R28447 a_3090_45724.t1 a_3090_45724.n19 26.5955
R28448 a_3090_45724.n19 a_3090_45724.t0 26.5955
R28449 a_3090_45724.n1 a_3090_45724.t4 24.9236
R28450 a_3090_45724.n1 a_3090_45724.t5 24.9236
R28451 a_3090_45724.n16 a_3090_45724.n15 16.5405
R28452 a_3090_45724.n15 a_3090_45724.n13 13.5684
R28453 a_3090_45724.n9 a_3090_45724.n8 12.1543
R28454 a_3090_45724.n17 a_3090_45724.n16 9.3005
R28455 a_3090_45724.n11 a_3090_45724.n9 9.06979
R28456 a_3090_45724.n12 a_3090_45724.n11 5.85607
R28457 a_n2438_43548.n42 a_n2438_43548.n41 333.392
R28458 a_n2438_43548.n18 a_n2438_43548.n0 301.392
R28459 a_n2438_43548.n36 a_n2438_43548.n35 301.392
R28460 a_n2438_43548.n38 a_n2438_43548.n37 301.392
R28461 a_n2438_43548.n40 a_n2438_43548.n39 301.392
R28462 a_n2438_43548.n43 a_n2438_43548.n42 301.392
R28463 a_n2438_43548.n17 a_n2438_43548.n1 297.863
R28464 a_n2438_43548.n29 a_n2438_43548.t33 294.557
R28465 a_n2438_43548.n27 a_n2438_43548.t40 294.557
R28466 a_n2438_43548.n25 a_n2438_43548.t44 294.557
R28467 a_n2438_43548.n23 a_n2438_43548.t42 294.557
R28468 a_n2438_43548.n21 a_n2438_43548.t38 294.557
R28469 a_n2438_43548.n20 a_n2438_43548.t43 294.557
R28470 a_n2438_43548.n19 a_n2438_43548.t34 294.557
R28471 a_n2438_43548.n33 a_n2438_43548.n32 287.303
R28472 a_n2438_43548.n4 a_n2438_43548.n2 248.638
R28473 a_n2438_43548.n29 a_n2438_43548.t37 211.01
R28474 a_n2438_43548.n27 a_n2438_43548.t36 211.01
R28475 a_n2438_43548.n25 a_n2438_43548.t41 211.01
R28476 a_n2438_43548.n23 a_n2438_43548.t39 211.01
R28477 a_n2438_43548.n21 a_n2438_43548.t45 211.01
R28478 a_n2438_43548.n20 a_n2438_43548.t35 211.01
R28479 a_n2438_43548.n19 a_n2438_43548.t32 211.01
R28480 a_n2438_43548.n4 a_n2438_43548.n3 203.463
R28481 a_n2438_43548.n6 a_n2438_43548.n5 203.463
R28482 a_n2438_43548.n10 a_n2438_43548.n9 203.463
R28483 a_n2438_43548.n12 a_n2438_43548.n11 203.463
R28484 a_n2438_43548.n14 a_n2438_43548.n13 203.463
R28485 a_n2438_43548.n8 a_n2438_43548.n7 202.456
R28486 a_n2438_43548.n16 a_n2438_43548.n15 200.212
R28487 a_n2438_43548.n26 a_n2438_43548.n25 180.447
R28488 a_n2438_43548.n22 a_n2438_43548.n21 180.447
R28489 a_n2438_43548.n31 a_n2438_43548.n19 179.643
R28490 a_n2438_43548.n30 a_n2438_43548.n29 174.832
R28491 a_n2438_43548.n22 a_n2438_43548.n20 169.195
R28492 a_n2438_43548.n24 a_n2438_43548.n23 167.191
R28493 a_n2438_43548.n28 a_n2438_43548.n27 166.898
R28494 a_n2438_43548.n6 a_n2438_43548.n4 45.177
R28495 a_n2438_43548.n12 a_n2438_43548.n10 45.177
R28496 a_n2438_43548.n14 a_n2438_43548.n12 45.177
R28497 a_n2438_43548.n8 a_n2438_43548.n6 44.0476
R28498 a_n2438_43548.n10 a_n2438_43548.n8 44.0476
R28499 a_n2438_43548.n33 a_n2438_43548.n31 42.1036
R28500 a_n2438_43548.n2 a_n2438_43548.t20 40.0005
R28501 a_n2438_43548.n2 a_n2438_43548.t18 40.0005
R28502 a_n2438_43548.n3 a_n2438_43548.t30 40.0005
R28503 a_n2438_43548.n3 a_n2438_43548.t28 40.0005
R28504 a_n2438_43548.n5 a_n2438_43548.t24 40.0005
R28505 a_n2438_43548.n5 a_n2438_43548.t29 40.0005
R28506 a_n2438_43548.n7 a_n2438_43548.t26 40.0005
R28507 a_n2438_43548.n7 a_n2438_43548.t21 40.0005
R28508 a_n2438_43548.n9 a_n2438_43548.t19 40.0005
R28509 a_n2438_43548.n9 a_n2438_43548.t31 40.0005
R28510 a_n2438_43548.n11 a_n2438_43548.t25 40.0005
R28511 a_n2438_43548.n11 a_n2438_43548.t27 40.0005
R28512 a_n2438_43548.n13 a_n2438_43548.t22 40.0005
R28513 a_n2438_43548.n13 a_n2438_43548.t17 40.0005
R28514 a_n2438_43548.n15 a_n2438_43548.t16 40.0005
R28515 a_n2438_43548.n15 a_n2438_43548.t23 40.0005
R28516 a_n2438_43548.n34 a_n2438_43548.n18 32.0005
R28517 a_n2438_43548.n36 a_n2438_43548.n34 32.0005
R28518 a_n2438_43548.n40 a_n2438_43548.n38 32.0005
R28519 a_n2438_43548.n42 a_n2438_43548.n40 32.0005
R28520 a_n2438_43548.n38 a_n2438_43548.n36 31.2005
R28521 a_n2438_43548.n41 a_n2438_43548.t11 27.5805
R28522 a_n2438_43548.n41 a_n2438_43548.t13 27.5805
R28523 a_n2438_43548.n0 a_n2438_43548.t2 27.5805
R28524 a_n2438_43548.n0 a_n2438_43548.t7 27.5805
R28525 a_n2438_43548.n1 a_n2438_43548.t5 27.5805
R28526 a_n2438_43548.n1 a_n2438_43548.t0 27.5805
R28527 a_n2438_43548.n32 a_n2438_43548.t1 27.5805
R28528 a_n2438_43548.n32 a_n2438_43548.t4 27.5805
R28529 a_n2438_43548.n35 a_n2438_43548.t12 27.5805
R28530 a_n2438_43548.n35 a_n2438_43548.t8 27.5805
R28531 a_n2438_43548.n37 a_n2438_43548.t3 27.5805
R28532 a_n2438_43548.n37 a_n2438_43548.t10 27.5805
R28533 a_n2438_43548.n39 a_n2438_43548.t14 27.5805
R28534 a_n2438_43548.n39 a_n2438_43548.t6 27.5805
R28535 a_n2438_43548.t15 a_n2438_43548.n43 27.5805
R28536 a_n2438_43548.n43 a_n2438_43548.t9 27.5805
R28537 a_n2438_43548.n30 a_n2438_43548.n28 15.7163
R28538 a_n2438_43548.n34 a_n2438_43548.n33 14.0898
R28539 a_n2438_43548.n16 a_n2438_43548.n14 13.177
R28540 a_n2438_43548.n18 a_n2438_43548.n17 10.4484
R28541 a_n2438_43548.n17 a_n2438_43548.n16 8.62539
R28542 a_n2438_43548.n28 a_n2438_43548.n26 7.15435
R28543 a_n2438_43548.n31 a_n2438_43548.n30 6.45533
R28544 a_n2438_43548.n24 a_n2438_43548.n22 2.2972
R28545 a_n2438_43548.n26 a_n2438_43548.n24 2.2972
R28546 a_15493_43396.t0 a_15493_43396.n1 223.757
R28547 a_15493_43396.n1 a_15493_43396.n0 206.781
R28548 a_15493_43396.n0 a_15493_43396.t2 206.19
R28549 a_15493_43396.n1 a_15493_43396.t1 186.736
R28550 a_15493_43396.n0 a_15493_43396.t3 142.344
R28551 a_5891_43370.n7 a_5891_43370.t15 256.728
R28552 a_5891_43370.n23 a_5891_43370.n22 248.087
R28553 a_5891_43370.n9 a_5891_43370.t11 241.536
R28554 a_5891_43370.n3 a_5891_43370.t18 236.18
R28555 a_5891_43370.n5 a_5891_43370.t16 231.835
R28556 a_5891_43370.n6 a_5891_43370.t23 229.369
R28557 a_5891_43370.n22 a_5891_43370.n21 208.508
R28558 a_5891_43370.n17 a_5891_43370.t21 201.369
R28559 a_5891_43370.n15 a_5891_43370.t22 183.505
R28560 a_5891_43370.n18 a_5891_43370.n17 182.165
R28561 a_5891_43370.n19 a_5891_43370.n3 178.9
R28562 a_5891_43370.n8 a_5891_43370.n7 178.311
R28563 a_5891_43370.n8 a_5891_43370.n6 173.828
R28564 a_5891_43370.n10 a_5891_43370.n9 172.821
R28565 a_5891_43370.n12 a_5891_43370.n4 171.267
R28566 a_5891_43370.n11 a_5891_43370.n5 169.833
R28567 a_5891_43370.n9 a_5891_43370.t8 169.237
R28568 a_5891_43370.n14 a_5891_43370.n13 168.282
R28569 a_5891_43370.n3 a_5891_43370.t9 163.881
R28570 a_5891_43370.n16 a_5891_43370.n15 163.162
R28571 a_5891_43370.n7 a_5891_43370.t12 161.275
R28572 a_5891_43370.n6 a_5891_43370.t10 157.07
R28573 a_5891_43370.n5 a_5891_43370.t13 157.07
R28574 a_5891_43370.n13 a_5891_43370.t20 142.994
R28575 a_5891_43370.n2 a_5891_43370.n0 137.575
R28576 a_5891_43370.n4 a_5891_43370.t14 137.177
R28577 a_5891_43370.n17 a_5891_43370.t19 132.282
R28578 a_5891_43370.n13 a_5891_43370.t24 126.927
R28579 a_5891_43370.n4 a_5891_43370.t25 121.109
R28580 a_5891_43370.n15 a_5891_43370.t17 114.532
R28581 a_5891_43370.n2 a_5891_43370.n1 99.1749
R28582 a_5891_43370.n22 a_5891_43370.n20 38.4831
R28583 a_5891_43370.n21 a_5891_43370.t1 26.5955
R28584 a_5891_43370.n21 a_5891_43370.t2 26.5955
R28585 a_5891_43370.n23 a_5891_43370.t0 26.5955
R28586 a_5891_43370.t3 a_5891_43370.n23 26.5955
R28587 a_5891_43370.n0 a_5891_43370.t7 24.9236
R28588 a_5891_43370.n0 a_5891_43370.t5 24.9236
R28589 a_5891_43370.n1 a_5891_43370.t6 24.9236
R28590 a_5891_43370.n1 a_5891_43370.t4 24.9236
R28591 a_5891_43370.n16 a_5891_43370.n14 15.1928
R28592 a_5891_43370.n20 a_5891_43370.n2 14.8665
R28593 a_5891_43370.n20 a_5891_43370.n19 9.3005
R28594 a_5891_43370.n11 a_5891_43370.n10 9.27676
R28595 a_5891_43370.n18 a_5891_43370.n16 8.39198
R28596 a_5891_43370.n19 a_5891_43370.n18 6.43748
R28597 a_5891_43370.n12 a_5891_43370.n11 5.63649
R28598 a_5891_43370.n10 a_5891_43370.n8 5.42752
R28599 a_5891_43370.n14 a_5891_43370.n12 4.5005
R28600 a_18184_42460.n0 a_18184_42460.t5 241.536
R28601 a_18184_42460.n1 a_18184_42460.t7 241.536
R28602 a_18184_42460.n2 a_18184_42460.t6 231.835
R28603 a_18184_42460.n5 a_18184_42460.t1 223.441
R28604 a_18184_42460.n4 a_18184_42460.n0 193.537
R28605 a_18184_42460.n3 a_18184_42460.n1 185.968
R28606 a_18184_42460.n3 a_18184_42460.n2 182.538
R28607 a_18184_42460.n6 a_18184_42460.n5 175.648
R28608 a_18184_42460.n0 a_18184_42460.t3 169.237
R28609 a_18184_42460.n1 a_18184_42460.t8 169.237
R28610 a_18184_42460.n2 a_18184_42460.t4 157.07
R28611 a_18184_42460.n6 a_18184_42460.t2 24.9236
R28612 a_18184_42460.t0 a_18184_42460.n6 24.9236
R28613 a_18184_42460.n5 a_18184_42460.n4 22.9867
R28614 a_18184_42460.n4 a_18184_42460.n3 0.705335
R28615 a_10903_43370.n21 a_10903_43370.n20 589.152
R28616 a_10903_43370.n15 a_10903_43370.t18 334.723
R28617 a_10903_43370.n17 a_10903_43370.t13 334.723
R28618 a_10903_43370.n9 a_10903_43370.t11 327.99
R28619 a_10903_43370.n20 a_10903_43370.n0 289.462
R28620 a_10903_43370.n14 a_10903_43370.t6 241.536
R28621 a_10903_43370.n6 a_10903_43370.t8 241.536
R28622 a_10903_43370.n2 a_10903_43370.t4 241.536
R28623 a_10903_43370.n3 a_10903_43370.t19 236.18
R28624 a_10903_43370.n11 a_10903_43370.t16 230.576
R28625 a_10903_43370.n1 a_10903_43370.t15 230.155
R28626 a_10903_43370.n15 a_10903_43370.t21 206.19
R28627 a_10903_43370.n17 a_10903_43370.t22 206.19
R28628 a_10903_43370.n9 a_10903_43370.t10 199.457
R28629 a_10903_43370.n4 a_10903_43370.n2 194.036
R28630 a_10903_43370.n16 a_10903_43370.n15 192.115
R28631 a_10903_43370.n12 a_10903_43370.n11 185.613
R28632 a_10903_43370.n10 a_10903_43370.n9 181.588
R28633 a_10903_43370.n7 a_10903_43370.n6 179.196
R28634 a_10903_43370.n4 a_10903_43370.n3 177.173
R28635 a_10903_43370.n18 a_10903_43370.n17 176.702
R28636 a_10903_43370.n16 a_10903_43370.n14 175.984
R28637 a_10903_43370.n14 a_10903_43370.t14 169.237
R28638 a_10903_43370.n6 a_10903_43370.t12 169.237
R28639 a_10903_43370.n2 a_10903_43370.t20 169.237
R28640 a_10903_43370.n13 a_10903_43370.n1 169.178
R28641 a_10903_43370.n7 a_10903_43370.n5 163.888
R28642 a_10903_43370.n3 a_10903_43370.t17 163.881
R28643 a_10903_43370.n11 a_10903_43370.t5 158.275
R28644 a_10903_43370.n1 a_10903_43370.t23 157.856
R28645 a_10903_43370.n5 a_10903_43370.t9 137.177
R28646 a_10903_43370.n5 a_10903_43370.t7 121.109
R28647 a_10903_43370.n0 a_10903_43370.t2 38.5719
R28648 a_10903_43370.n0 a_10903_43370.t3 38.5719
R28649 a_10903_43370.t1 a_10903_43370.n21 26.5955
R28650 a_10903_43370.n21 a_10903_43370.t0 26.5955
R28651 a_10903_43370.n20 a_10903_43370.n19 11.6482
R28652 a_10903_43370.n19 a_10903_43370.n18 10.9936
R28653 a_10903_43370.n10 a_10903_43370.n8 8.90435
R28654 a_10903_43370.n19 a_10903_43370.n13 7.24363
R28655 a_10903_43370.n12 a_10903_43370.n10 2.90435
R28656 a_10903_43370.n18 a_10903_43370.n16 2.53913
R28657 a_10903_43370.n8 a_10903_43370.n4 2.34819
R28658 a_10903_43370.n13 a_10903_43370.n12 1.08292
R28659 a_10903_43370.n8 a_10903_43370.n7 0.34528
R28660 a_3483_46348.n7 a_3483_46348.t18 722.096
R28661 a_3483_46348.n5 a_3483_46348.t22 722.096
R28662 a_3483_46348.n4 a_3483_46348.t16 722.096
R28663 a_3483_46348.n21 a_3483_46348.n20 380.32
R28664 a_3483_46348.n3 a_3483_46348.t11 241.536
R28665 a_3483_46348.n2 a_3483_46348.t20 241.536
R28666 a_3483_46348.n13 a_3483_46348.t7 241.536
R28667 a_3483_46348.n1 a_3483_46348.t9 239.505
R28668 a_3483_46348.n0 a_3483_46348.t6 238.59
R28669 a_3483_46348.n15 a_3483_46348.t8 230.923
R28670 a_3483_46348.n10 a_3483_46348.t19 230.923
R28671 a_3483_46348.n0 a_3483_46348.t23 203.244
R28672 a_3483_46348.n12 a_3483_46348.n2 191.306
R28673 a_3483_46348.n6 a_3483_46348.n4 187.928
R28674 a_3483_46348.n9 a_3483_46348.n3 187.328
R28675 a_3483_46348.n20 a_3483_46348.n19 185
R28676 a_3483_46348.n18 a_3483_46348.n0 184.639
R28677 a_3483_46348.n11 a_3483_46348.n10 179.589
R28678 a_3483_46348.n16 a_3483_46348.n15 177.131
R28679 a_3483_46348.n14 a_3483_46348.n13 171.482
R28680 a_3483_46348.n3 a_3483_46348.t12 169.237
R28681 a_3483_46348.n2 a_3483_46348.t21 169.237
R28682 a_3483_46348.n13 a_3483_46348.t15 169.237
R28683 a_3483_46348.n8 a_3483_46348.n7 168.016
R28684 a_3483_46348.n6 a_3483_46348.n5 168.016
R28685 a_3483_46348.n17 a_3483_46348.n1 167.879
R28686 a_3483_46348.n1 a_3483_46348.t10 167.204
R28687 a_3483_46348.n15 a_3483_46348.t14 163.881
R28688 a_3483_46348.n10 a_3483_46348.t4 163.881
R28689 a_3483_46348.n7 a_3483_46348.t17 162.963
R28690 a_3483_46348.n5 a_3483_46348.t5 162.963
R28691 a_3483_46348.n4 a_3483_46348.t13 162.963
R28692 a_3483_46348.n21 a_3483_46348.t0 26.5955
R28693 a_3483_46348.t1 a_3483_46348.n21 26.5955
R28694 a_3483_46348.n19 a_3483_46348.t2 24.9236
R28695 a_3483_46348.n19 a_3483_46348.t3 24.9236
R28696 a_3483_46348.n11 a_3483_46348.n9 17.9222
R28697 a_3483_46348.n18 a_3483_46348.n17 17.5257
R28698 a_3483_46348.n20 a_3483_46348.n18 15.0985
R28699 a_3483_46348.n17 a_3483_46348.n16 14.7674
R28700 a_3483_46348.n16 a_3483_46348.n14 10.1186
R28701 a_3483_46348.n9 a_3483_46348.n8 9.83292
R28702 a_3483_46348.n12 a_3483_46348.n11 8.88649
R28703 a_3483_46348.n8 a_3483_46348.n6 7.29462
R28704 a_3483_46348.n14 a_3483_46348.n12 0.779346
R28705 a_9290_44172.n4 a_9290_44172.t29 330.12
R28706 a_9290_44172.n15 a_9290_44172.t8 293.969
R28707 a_9290_44172.n11 a_9290_44172.t11 256.716
R28708 a_9290_44172.n25 a_9290_44172.n0 248.088
R28709 a_9290_44172.n8 a_9290_44172.t21 241.536
R28710 a_9290_44172.n9 a_9290_44172.t17 241.536
R28711 a_9290_44172.n7 a_9290_44172.t19 241.536
R28712 a_9290_44172.n5 a_9290_44172.t28 236.18
R28713 a_9290_44172.n6 a_9290_44172.t10 231.835
R28714 a_9290_44172.n16 a_9290_44172.n14 219.542
R28715 a_9290_44172.n14 a_9290_44172.t22 212.081
R28716 a_9290_44172.n13 a_9290_44172.t25 212.081
R28717 a_9290_44172.n26 a_9290_44172.n25 208.507
R28718 a_9290_44172.n4 a_9290_44172.t20 201.587
R28719 a_9290_44172.n19 a_9290_44172.t24 201.369
R28720 a_9290_44172.n23 a_9290_44172.n4 191.014
R28721 a_9290_44172.n20 a_9290_44172.n19 180.903
R28722 a_9290_44172.n18 a_9290_44172.n7 180.822
R28723 a_9290_44172.n10 a_9290_44172.n8 178.106
R28724 a_9290_44172.n22 a_9290_44172.n5 177.312
R28725 a_9290_44172.n10 a_9290_44172.n9 173.597
R28726 a_9290_44172.n12 a_9290_44172.n11 169.565
R28727 a_9290_44172.n8 a_9290_44172.t16 169.237
R28728 a_9290_44172.n9 a_9290_44172.t15 169.237
R28729 a_9290_44172.n7 a_9290_44172.t14 169.237
R28730 a_9290_44172.n16 a_9290_44172.n15 164.994
R28731 a_9290_44172.n5 a_9290_44172.t23 163.881
R28732 a_9290_44172.n21 a_9290_44172.n6 163.536
R28733 a_9290_44172.n11 a_9290_44172.t9 161.275
R28734 a_9290_44172.n6 a_9290_44172.t26 157.07
R28735 a_9290_44172.n14 a_9290_44172.t27 139.78
R28736 a_9290_44172.n13 a_9290_44172.t12 139.78
R28737 a_9290_44172.n15 a_9290_44172.t13 138.338
R28738 a_9290_44172.n3 a_9290_44172.n1 137.575
R28739 a_9290_44172.n19 a_9290_44172.t18 132.282
R28740 a_9290_44172.n3 a_9290_44172.n2 99.1749
R28741 a_9290_44172.n14 a_9290_44172.n13 61.346
R28742 a_9290_44172.n24 a_9290_44172.n3 36.0958
R28743 a_9290_44172.n0 a_9290_44172.t2 26.5955
R28744 a_9290_44172.n0 a_9290_44172.t0 26.5955
R28745 a_9290_44172.n26 a_9290_44172.t1 26.5955
R28746 a_9290_44172.t3 a_9290_44172.n26 26.5955
R28747 a_9290_44172.n1 a_9290_44172.t7 24.9236
R28748 a_9290_44172.n1 a_9290_44172.t4 24.9236
R28749 a_9290_44172.n2 a_9290_44172.t6 24.9236
R28750 a_9290_44172.n2 a_9290_44172.t5 24.9236
R28751 a_9290_44172.n24 a_9290_44172.n23 21.5163
R28752 a_9290_44172.n17 a_9290_44172.n16 17.6543
R28753 a_9290_44172.n25 a_9290_44172.n24 17.2539
R28754 a_9290_44172.n17 a_9290_44172.n12 9.36863
R28755 a_9290_44172.n12 a_9290_44172.n10 9.31227
R28756 a_9290_44172.n20 a_9290_44172.n18 7.09391
R28757 a_9290_44172.n18 a_9290_44172.n17 6.83292
R28758 a_9290_44172.n23 a_9290_44172.n22 6.22028
R28759 a_9290_44172.n22 a_9290_44172.n21 1.98814
R28760 a_9290_44172.n21 a_9290_44172.n20 0.755995
R28761 a_11823_42460.t17 a_11823_42460.t16 378.255
R28762 a_11823_42460.n4 a_11823_42460.t17 363.978
R28763 a_11823_42460.n17 a_11823_42460.t9 334.723
R28764 a_11823_42460.n5 a_11823_42460.t22 334.723
R28765 a_11823_42460.n6 a_11823_42460.t25 293.969
R28766 a_11823_42460.n13 a_11823_42460.t24 256.716
R28767 a_11823_42460.n24 a_11823_42460.n23 248.087
R28768 a_11823_42460.n3 a_11823_42460.t10 241.536
R28769 a_11823_42460.n12 a_11823_42460.t11 241.536
R28770 a_11823_42460.n20 a_11823_42460.t13 231.835
R28771 a_11823_42460.n9 a_11823_42460.t14 212.081
R28772 a_11823_42460.n8 a_11823_42460.t26 212.081
R28773 a_11823_42460.n25 a_11823_42460.n24 208.506
R28774 a_11823_42460.n17 a_11823_42460.t28 206.19
R28775 a_11823_42460.n5 a_11823_42460.t23 206.19
R28776 a_11823_42460.n16 a_11823_42460.t18 201.369
R28777 a_11823_42460.n10 a_11823_42460.n9 194.022
R28778 a_11823_42460.n14 a_11823_42460.n12 185.038
R28779 a_11823_42460.n7 a_11823_42460.n5 179.22
R28780 a_11823_42460.n4 a_11823_42460.n3 178.106
R28781 a_11823_42460.n18 a_11823_42460.n17 174.528
R28782 a_11823_42460.n7 a_11823_42460.n6 172.155
R28783 a_11823_42460.n3 a_11823_42460.t19 169.237
R28784 a_11823_42460.n12 a_11823_42460.t29 169.237
R28785 a_11823_42460.n14 a_11823_42460.n13 167.819
R28786 a_11823_42460.n18 a_11823_42460.n16 164.242
R28787 a_11823_42460.n21 a_11823_42460.n20 163.349
R28788 a_11823_42460.n13 a_11823_42460.t27 161.275
R28789 a_11823_42460.n20 a_11823_42460.t20 157.07
R28790 a_11823_42460.n9 a_11823_42460.t15 139.78
R28791 a_11823_42460.n8 a_11823_42460.t12 139.78
R28792 a_11823_42460.n6 a_11823_42460.t8 138.338
R28793 a_11823_42460.n2 a_11823_42460.n0 137.576
R28794 a_11823_42460.n16 a_11823_42460.t21 132.282
R28795 a_11823_42460.n2 a_11823_42460.n1 99.1759
R28796 a_11823_42460.n9 a_11823_42460.n8 61.346
R28797 a_11823_42460.n22 a_11823_42460.n2 36.0958
R28798 a_11823_42460.n23 a_11823_42460.t0 26.5955
R28799 a_11823_42460.n23 a_11823_42460.t1 26.5955
R28800 a_11823_42460.n25 a_11823_42460.t2 26.5955
R28801 a_11823_42460.t3 a_11823_42460.n25 26.5955
R28802 a_11823_42460.n0 a_11823_42460.t6 24.9236
R28803 a_11823_42460.n0 a_11823_42460.t4 24.9236
R28804 a_11823_42460.n1 a_11823_42460.t5 24.9236
R28805 a_11823_42460.n1 a_11823_42460.t7 24.9236
R28806 a_11823_42460.n22 a_11823_42460.n21 20.5972
R28807 a_11823_42460.n24 a_11823_42460.n22 17.2539
R28808 a_11823_42460.n19 a_11823_42460.n15 15.2546
R28809 a_11823_42460.n11 a_11823_42460.n4 11.9991
R28810 a_11823_42460.n21 a_11823_42460.n19 10.5142
R28811 a_11823_42460.n15 a_11823_42460.n14 10.4401
R28812 a_11823_42460.n11 a_11823_42460.n10 6.01149
R28813 a_11823_42460.n15 a_11823_42460.n11 5.63649
R28814 a_11823_42460.n10 a_11823_42460.n7 4.5005
R28815 a_11823_42460.n19 a_11823_42460.n18 4.5005
R28816 a_n2312_40392.n3 a_n2312_40392.n2 380.32
R28817 a_n2312_40392.n2 a_n2312_40392.n0 263.784
R28818 a_n2312_40392.n0 a_n2312_40392.t5 228.649
R28819 a_n2312_40392.n2 a_n2312_40392.n1 185
R28820 a_n2312_40392.n0 a_n2312_40392.t4 156.35
R28821 a_n2312_40392.t1 a_n2312_40392.n3 26.5955
R28822 a_n2312_40392.n3 a_n2312_40392.t0 26.5955
R28823 a_n2312_40392.n1 a_n2312_40392.t2 24.9236
R28824 a_n2312_40392.n1 a_n2312_40392.t3 24.9236
R28825 a_2063_45854.n9 a_2063_45854.t10 471.289
R28826 a_2063_45854.n10 a_2063_45854.t14 471.289
R28827 a_2063_45854.n15 a_2063_45854.n14 288.212
R28828 a_2063_45854.n14 a_2063_45854.n0 261.81
R28829 a_2063_45854.n1 a_2063_45854.t15 256.07
R28830 a_2063_45854.n5 a_2063_45854.t16 236.18
R28831 a_2063_45854.n2 a_2063_45854.t7 230.363
R28832 a_2063_45854.n3 a_2063_45854.t4 230.155
R28833 a_2063_45854.n7 a_2063_45854.t8 229.369
R28834 a_2063_45854.n11 a_2063_45854.n10 190.51
R28835 a_2063_45854.n6 a_2063_45854.n5 189.482
R28836 a_2063_45854.n13 a_2063_45854.n1 188.681
R28837 a_2063_45854.n11 a_2063_45854.n9 181.641
R28838 a_2063_45854.n8 a_2063_45854.n7 171.438
R28839 a_2063_45854.n4 a_2063_45854.n2 168.891
R28840 a_2063_45854.n4 a_2063_45854.n3 168.81
R28841 a_2063_45854.n5 a_2063_45854.t5 163.881
R28842 a_2063_45854.n2 a_2063_45854.t11 158.064
R28843 a_2063_45854.n3 a_2063_45854.t12 157.856
R28844 a_2063_45854.n7 a_2063_45854.t9 157.07
R28845 a_2063_45854.n1 a_2063_45854.t6 150.03
R28846 a_2063_45854.n9 a_2063_45854.t17 148.35
R28847 a_2063_45854.n10 a_2063_45854.t13 148.35
R28848 a_2063_45854.n12 a_2063_45854.n11 39.613
R28849 a_2063_45854.n15 a_2063_45854.t0 26.5955
R28850 a_2063_45854.t1 a_2063_45854.n15 26.5955
R28851 a_2063_45854.n14 a_2063_45854.n13 25.0133
R28852 a_2063_45854.n0 a_2063_45854.t2 24.9236
R28853 a_2063_45854.n0 a_2063_45854.t3 24.9236
R28854 a_2063_45854.n12 a_2063_45854.n8 7.30536
R28855 a_2063_45854.n6 a_2063_45854.n4 5.32742
R28856 a_2063_45854.n13 a_2063_45854.n12 3.4105
R28857 a_2063_45854.n8 a_2063_45854.n6 2.45242
R28858 a_n3565_38502.n4 a_n3565_38502.t10 557.081
R28859 a_n3565_38502.n8 a_n3565_38502.n7 340.637
R28860 a_n3565_38502.n3 a_n3565_38502.t8 241.536
R28861 a_n3565_38502.n7 a_n3565_38502.n6 195.577
R28862 a_n3565_38502.n3 a_n3565_38502.t9 169.237
R28863 a_n3565_38502.n4 a_n3565_38502.n3 168.505
R28864 a_n3565_38502.n2 a_n3565_38502.n0 137.189
R28865 a_n3565_38502.n2 a_n3565_38502.n1 98.788
R28866 a_n3565_38502.n7 a_n3565_38502.n5 39.0246
R28867 a_n3565_38502.n6 a_n3565_38502.t0 26.5955
R28868 a_n3565_38502.n6 a_n3565_38502.t2 26.5955
R28869 a_n3565_38502.t3 a_n3565_38502.n8 26.5955
R28870 a_n3565_38502.n8 a_n3565_38502.t1 26.5955
R28871 a_n3565_38502.n5 a_n3565_38502.n2 25.9824
R28872 a_n3565_38502.n0 a_n3565_38502.t4 24.9236
R28873 a_n3565_38502.n0 a_n3565_38502.t6 24.9236
R28874 a_n3565_38502.n1 a_n3565_38502.t5 24.9236
R28875 a_n3565_38502.n1 a_n3565_38502.t7 24.9236
R28876 a_n3565_38502.n5 a_n3565_38502.n4 9.38613
R28877 a_4883_46098.t0 a_4883_46098.n7 427.791
R28878 a_4883_46098.n0 a_4883_46098.t6 323.55
R28879 a_4883_46098.n2 a_4883_46098.t5 276.464
R28880 a_4883_46098.n1 a_4883_46098.t4 276.464
R28881 a_4883_46098.n4 a_4883_46098.t7 224.984
R28882 a_4883_46098.n7 a_4883_46098.t1 209.923
R28883 a_4883_46098.n2 a_4883_46098.t3 196.131
R28884 a_4883_46098.n1 a_4883_46098.t8 196.131
R28885 a_4883_46098.n0 a_4883_46098.t2 195.017
R28886 a_4883_46098.n3 a_4883_46098.n2 193.362
R28887 a_4883_46098.n4 a_4883_46098.t9 187.714
R28888 a_4883_46098.n6 a_4883_46098.n0 179.174
R28889 a_4883_46098.n3 a_4883_46098.n1 175.321
R28890 a_4883_46098.n5 a_4883_46098.n4 172.817
R28891 a_4883_46098.n7 a_4883_46098.n6 19.824
R28892 a_4883_46098.n6 a_4883_46098.n5 13.5596
R28893 a_4883_46098.n5 a_4883_46098.n3 0.356133
R28894 a_n784_42308.n0 a_n784_42308.t4 585.907
R28895 a_n784_42308.n0 a_n784_42308.t6 585.436
R28896 a_n784_42308.n5 a_n784_42308.n4 380.32
R28897 a_n784_42308.n1 a_n784_42308.t5 260.322
R28898 a_n784_42308.n2 a_n784_42308.n1 186.899
R28899 a_n784_42308.n4 a_n784_42308.n3 185
R28900 a_n784_42308.n1 a_n784_42308.t7 175.169
R28901 a_n784_42308.n2 a_n784_42308.n0 129.095
R28902 a_n784_42308.n5 a_n784_42308.t0 26.5955
R28903 a_n784_42308.t1 a_n784_42308.n5 26.5955
R28904 a_n784_42308.n3 a_n784_42308.t2 24.9236
R28905 a_n784_42308.n3 a_n784_42308.t3 24.9236
R28906 a_n784_42308.n4 a_n784_42308.n2 22.9371
R28907 C0_P_btm.n1 C0_P_btm.t0 101.944
R28908 C0_P_btm.n2 C0_P_btm.t3 99.4985
R28909 C0_P_btm.n0 C0_P_btm.t2 54.9098
R28910 C0_P_btm C0_P_btm.n2 47.6359
R28911 C0_P_btm.n0 C0_P_btm.t1 47.3635
R28912 C0_P_btm.n1 C0_P_btm.n0 8.27654
R28913 C0_P_btm.n2 C0_P_btm.n1 6.33383
R28914 a_n237_47217.n4 a_n237_47217.t13 471.289
R28915 a_n237_47217.n5 a_n237_47217.t12 414.432
R28916 a_n237_47217.n12 a_n237_47217.n11 365.022
R28917 a_n237_47217.n5 a_n237_47217.t11 300.349
R28918 a_n237_47217.n3 a_n237_47217.t8 256.07
R28919 a_n237_47217.n2 a_n237_47217.t15 230.155
R28920 a_n237_47217.n0 a_n237_47217.t6 212.081
R28921 a_n237_47217.n1 a_n237_47217.t5 212.081
R28922 a_n237_47217.n6 a_n237_47217.n4 202.714
R28923 a_n237_47217.n9 a_n237_47217.n1 200.113
R28924 a_n237_47217.n7 a_n237_47217.n3 190.47
R28925 a_n237_47217.n11 a_n237_47217.n10 185
R28926 a_n237_47217.n8 a_n237_47217.n2 164.554
R28927 a_n237_47217.n2 a_n237_47217.t7 157.856
R28928 a_n237_47217.n3 a_n237_47217.t4 150.03
R28929 a_n237_47217.n4 a_n237_47217.t10 148.35
R28930 a_n237_47217.n0 a_n237_47217.t9 139.78
R28931 a_n237_47217.n1 a_n237_47217.t14 139.78
R28932 a_n237_47217.n6 a_n237_47217.n5 64.1409
R28933 a_n237_47217.n1 a_n237_47217.n0 61.346
R28934 a_n237_47217.n7 a_n237_47217.n6 37.0081
R28935 a_n237_47217.n12 a_n237_47217.t0 26.5955
R28936 a_n237_47217.t1 a_n237_47217.n12 26.5955
R28937 a_n237_47217.n10 a_n237_47217.t3 24.9236
R28938 a_n237_47217.n10 a_n237_47217.t2 24.9236
R28939 a_n237_47217.n11 a_n237_47217.n9 20.2386
R28940 a_n237_47217.n8 a_n237_47217.n7 9.29785
R28941 a_n237_47217.n9 a_n237_47217.n8 5.9277
R28942 a_6123_31319.n0 a_6123_31319.t7 581.852
R28943 a_6123_31319.n0 a_6123_31319.t4 578.573
R28944 a_6123_31319.n5 a_6123_31319.n4 380.32
R28945 a_6123_31319.n1 a_6123_31319.t5 260.322
R28946 a_6123_31319.n4 a_6123_31319.n3 185
R28947 a_6123_31319.n1 a_6123_31319.t6 175.169
R28948 a_6123_31319.n2 a_6123_31319.n1 173.462
R28949 a_6123_31319.n2 a_6123_31319.n0 116.695
R28950 a_6123_31319.t1 a_6123_31319.n5 26.5955
R28951 a_6123_31319.n5 a_6123_31319.t0 26.5955
R28952 a_6123_31319.n3 a_6123_31319.t2 24.9236
R28953 a_6123_31319.n3 a_6123_31319.t3 24.9236
R28954 a_6123_31319.n4 a_6123_31319.n2 18.0103
R28955 a_5534_30871.n1 a_5534_30871.t4 1614.4
R28956 a_5534_30871.n1 a_5534_30871.t5 1613.18
R28957 a_5534_30871.n5 a_5534_30871.n4 380.32
R28958 a_5534_30871.n0 a_5534_30871.t6 260.322
R28959 a_5534_30871.n4 a_5534_30871.n3 185
R28960 a_5534_30871.n2 a_5534_30871.n0 179.272
R28961 a_5534_30871.n0 a_5534_30871.t7 175.169
R28962 a_5534_30871.n2 a_5534_30871.n1 74.8947
R28963 a_5534_30871.n5 a_5534_30871.t0 26.5955
R28964 a_5534_30871.t1 a_5534_30871.n5 26.5955
R28965 a_5534_30871.n3 a_5534_30871.t3 24.9236
R28966 a_5534_30871.n3 a_5534_30871.t2 24.9236
R28967 a_5534_30871.n4 a_5534_30871.n2 23.017
R28968 C7_P_btm C7_P_btm.n3 60.563
R28969 C7_P_btm.n3 C7_P_btm.t4 53.6613
R28970 C7_P_btm.n1 C7_P_btm.n0 52.9499
R28971 C7_P_btm.n1 C7_P_btm.t0 23.6451
R28972 C7_P_btm.n2 C7_P_btm.t1 23.6328
R28973 C7_P_btm.n2 C7_P_btm.n1 11.2505
R28974 C7_P_btm.n3 C7_P_btm.n2 8.41717
R28975 C7_P_btm.n0 C7_P_btm.t3 3.57113
R28976 C7_P_btm.n0 C7_P_btm.t2 3.57113
R28977 a_22612_30879.n0 a_22612_30879.t10 756.547
R28978 a_22612_30879.n14 a_22612_30879.t6 756.226
R28979 a_22612_30879.n0 a_22612_30879.t8 756.226
R28980 a_22612_30879.n1 a_22612_30879.t16 756.226
R28981 a_22612_30879.n2 a_22612_30879.t14 756.226
R28982 a_22612_30879.n3 a_22612_30879.t4 756.226
R28983 a_22612_30879.n4 a_22612_30879.t11 756.226
R28984 a_22612_30879.n5 a_22612_30879.t17 756.226
R28985 a_22612_30879.n6 a_22612_30879.t7 756.226
R28986 a_22612_30879.n7 a_22612_30879.t15 756.226
R28987 a_22612_30879.n8 a_22612_30879.t19 756.226
R28988 a_22612_30879.n9 a_22612_30879.t12 756.226
R28989 a_22612_30879.n10 a_22612_30879.t9 756.226
R28990 a_22612_30879.n11 a_22612_30879.t13 756.226
R28991 a_22612_30879.n12 a_22612_30879.t18 756.226
R28992 a_22612_30879.n13 a_22612_30879.t5 756.226
R28993 a_22612_30879.n17 a_22612_30879.n16 380.32
R28994 a_22612_30879.n16 a_22612_30879.n15 185
R28995 a_22612_30879.n16 a_22612_30879.n14 98.9943
R28996 a_22612_30879.t1 a_22612_30879.n17 26.5955
R28997 a_22612_30879.n17 a_22612_30879.t0 26.5955
R28998 a_22612_30879.n15 a_22612_30879.t3 24.9236
R28999 a_22612_30879.n15 a_22612_30879.t2 24.9236
R29000 a_22612_30879.n13 a_22612_30879.n12 0.3205
R29001 a_22612_30879.n12 a_22612_30879.n11 0.3205
R29002 a_22612_30879.n11 a_22612_30879.n10 0.3205
R29003 a_22612_30879.n10 a_22612_30879.n9 0.3205
R29004 a_22612_30879.n9 a_22612_30879.n8 0.3205
R29005 a_22612_30879.n8 a_22612_30879.n7 0.3205
R29006 a_22612_30879.n7 a_22612_30879.n6 0.3205
R29007 a_22612_30879.n6 a_22612_30879.n5 0.3205
R29008 a_22612_30879.n5 a_22612_30879.n4 0.3205
R29009 a_22612_30879.n4 a_22612_30879.n3 0.3205
R29010 a_22612_30879.n3 a_22612_30879.n2 0.3205
R29011 a_22612_30879.n2 a_22612_30879.n1 0.3205
R29012 a_22612_30879.n1 a_22612_30879.n0 0.3205
R29013 a_22612_30879.n14 a_22612_30879.n13 0.303833
R29014 a_n4064_37984.n5 a_n4064_37984.t9 634.832
R29015 a_n4064_37984.n8 a_n4064_37984.n7 360.399
R29016 a_n4064_37984.n4 a_n4064_37984.t10 241.536
R29017 a_n4064_37984.n3 a_n4064_37984.n2 232.862
R29018 a_n4064_37984.n7 a_n4064_37984.n0 203.161
R29019 a_n4064_37984.n5 a_n4064_37984.n4 172.035
R29020 a_n4064_37984.n4 a_n4064_37984.t8 169.237
R29021 a_n4064_37984.n3 a_n4064_37984.n1 95.6721
R29022 a_n4064_37984.n6 a_n4064_37984.n3 60.5918
R29023 a_n4064_37984.n0 a_n4064_37984.t0 27.5805
R29024 a_n4064_37984.n0 a_n4064_37984.t2 27.5805
R29025 a_n4064_37984.n8 a_n4064_37984.t1 27.5805
R29026 a_n4064_37984.t3 a_n4064_37984.n8 27.5805
R29027 a_n4064_37984.n2 a_n4064_37984.t5 25.8467
R29028 a_n4064_37984.n2 a_n4064_37984.t4 25.8467
R29029 a_n4064_37984.n1 a_n4064_37984.t7 25.8467
R29030 a_n4064_37984.n1 a_n4064_37984.t6 25.8467
R29031 a_n4064_37984.n7 a_n4064_37984.n6 22.6489
R29032 a_n4064_37984.n6 a_n4064_37984.n5 9.40917
R29033 a_n3674_38680.n3 a_n3674_38680.n2 287.752
R29034 a_n3674_38680.n2 a_n3674_38680.n0 277.568
R29035 a_n3674_38680.n2 a_n3674_38680.n1 238.288
R29036 a_n3674_38680.n1 a_n3674_38680.t4 235.821
R29037 a_n3674_38680.n1 a_n3674_38680.t5 163.52
R29038 a_n3674_38680.n3 a_n3674_38680.t0 26.5955
R29039 a_n3674_38680.t1 a_n3674_38680.n3 26.5955
R29040 a_n3674_38680.n0 a_n3674_38680.t3 24.9236
R29041 a_n3674_38680.n0 a_n3674_38680.t2 24.9236
R29042 a_13467_32519.n1 a_13467_32519.t4 677.61
R29043 a_13467_32519.n2 a_13467_32519.n1 380.32
R29044 a_13467_32519.n1 a_13467_32519.n0 185
R29045 a_13467_32519.n2 a_13467_32519.t0 26.5955
R29046 a_13467_32519.t1 a_13467_32519.n2 26.5955
R29047 a_13467_32519.n0 a_13467_32519.t2 24.9236
R29048 a_13467_32519.n0 a_13467_32519.t3 24.9236
R29049 a_n4064_40160.n13 a_n4064_40160.t13 1415.15
R29050 a_n4064_40160.n12 a_n4064_40160.t17 1330.32
R29051 a_n4064_40160.n6 a_n4064_40160.t8 1330.32
R29052 a_n4064_40160.n10 a_n4064_40160.t11 1330.32
R29053 a_n4064_40160.n11 a_n4064_40160.t9 1320.68
R29054 a_n4064_40160.n13 a_n4064_40160.t10 1320.68
R29055 a_n4064_40160.n9 a_n4064_40160.t15 1320.68
R29056 a_n4064_40160.n7 a_n4064_40160.t16 1320.68
R29057 a_n4064_40160.n18 a_n4064_40160.n17 360.399
R29058 a_n4064_40160.n4 a_n4064_40160.t12 241.536
R29059 a_n4064_40160.n3 a_n4064_40160.n2 232.862
R29060 a_n4064_40160.n17 a_n4064_40160.n0 203.161
R29061 a_n4064_40160.n15 a_n4064_40160.n4 172.035
R29062 a_n4064_40160.n4 a_n4064_40160.t14 169.237
R29063 a_n4064_40160.n8 a_n4064_40160.n7 161.78
R29064 a_n4064_40160.n11 a_n4064_40160.n5 161.3
R29065 a_n4064_40160.n9 a_n4064_40160.n8 161.3
R29066 a_n4064_40160.n14 a_n4064_40160.n13 161.3
R29067 a_n4064_40160.n3 a_n4064_40160.n1 95.6721
R29068 a_n4064_40160.n13 a_n4064_40160.n12 84.8325
R29069 a_n4064_40160.n12 a_n4064_40160.n11 84.8325
R29070 a_n4064_40160.n7 a_n4064_40160.n6 84.8325
R29071 a_n4064_40160.n9 a_n4064_40160.n6 84.8325
R29072 a_n4064_40160.n10 a_n4064_40160.n9 84.8325
R29073 a_n4064_40160.n11 a_n4064_40160.n10 84.8325
R29074 a_n4064_40160.n15 a_n4064_40160.n14 77.6708
R29075 a_n4064_40160.n16 a_n4064_40160.n3 60.5918
R29076 a_n4064_40160.n0 a_n4064_40160.t0 27.5805
R29077 a_n4064_40160.n0 a_n4064_40160.t1 27.5805
R29078 a_n4064_40160.n18 a_n4064_40160.t2 27.5805
R29079 a_n4064_40160.t3 a_n4064_40160.n18 27.5805
R29080 a_n4064_40160.n2 a_n4064_40160.t4 25.8467
R29081 a_n4064_40160.n2 a_n4064_40160.t6 25.8467
R29082 a_n4064_40160.n1 a_n4064_40160.t5 25.8467
R29083 a_n4064_40160.n1 a_n4064_40160.t7 25.8467
R29084 a_n4064_40160.n17 a_n4064_40160.n16 22.6489
R29085 a_n4064_40160.n16 a_n4064_40160.n15 9.40917
R29086 a_n4064_40160.n8 a_n4064_40160.n5 0.4805
R29087 a_n4064_40160.n14 a_n4064_40160.n5 0.4655
R29088 C10_P_btm C10_P_btm.n32 90.4588
R29089 C10_P_btm.n2 C10_P_btm.n0 33.0802
R29090 C10_P_btm.n14 C10_P_btm.n13 32.3614
R29091 C10_P_btm.n12 C10_P_btm.n11 32.3614
R29092 C10_P_btm.n10 C10_P_btm.n9 32.3614
R29093 C10_P_btm.n8 C10_P_btm.n7 32.3614
R29094 C10_P_btm.n6 C10_P_btm.n5 32.3614
R29095 C10_P_btm.n4 C10_P_btm.n3 32.3614
R29096 C10_P_btm.n2 C10_P_btm.n1 32.3614
R29097 C10_P_btm.n22 C10_P_btm.n14 29.1203
R29098 C10_P_btm.n24 C10_P_btm.n23 20.3263
R29099 C10_P_btm.n27 C10_P_btm.n25 15.4755
R29100 C10_P_btm.n17 C10_P_btm.n15 15.394
R29101 C10_P_btm.n29 C10_P_btm.n28 14.9755
R29102 C10_P_btm.n27 C10_P_btm.n26 14.9755
R29103 C10_P_btm.n31 C10_P_btm.n30 14.9755
R29104 C10_P_btm.n21 C10_P_btm.n20 14.894
R29105 C10_P_btm.n19 C10_P_btm.n18 14.894
R29106 C10_P_btm.n17 C10_P_btm.n16 14.894
R29107 C10_P_btm.n24 C10_P_btm.n22 6.29217
R29108 C10_P_btm.n22 C10_P_btm.n21 5.43279
R29109 C10_P_btm C10_P_btm.n1044 5.41222
R29110 C10_P_btm.n32 C10_P_btm.n31 5.33904
R29111 C10_P_btm.n32 C10_P_btm.n24 4.7505
R29112 C10_P_btm.n13 C10_P_btm.t26 3.57113
R29113 C10_P_btm.n13 C10_P_btm.t16 3.57113
R29114 C10_P_btm.n11 C10_P_btm.t24 3.57113
R29115 C10_P_btm.n11 C10_P_btm.t28 3.57113
R29116 C10_P_btm.n9 C10_P_btm.t25 3.57113
R29117 C10_P_btm.n9 C10_P_btm.t18 3.57113
R29118 C10_P_btm.n7 C10_P_btm.t23 3.57113
R29119 C10_P_btm.n7 C10_P_btm.t29 3.57113
R29120 C10_P_btm.n5 C10_P_btm.t31 3.57113
R29121 C10_P_btm.n5 C10_P_btm.t27 3.57113
R29122 C10_P_btm.n3 C10_P_btm.t30 3.57113
R29123 C10_P_btm.n3 C10_P_btm.t19 3.57113
R29124 C10_P_btm.n1 C10_P_btm.t22 3.57113
R29125 C10_P_btm.n1 C10_P_btm.t17 3.57113
R29126 C10_P_btm.n0 C10_P_btm.t20 3.57113
R29127 C10_P_btm.n0 C10_P_btm.t21 3.57113
R29128 C10_P_btm.n28 C10_P_btm.t1 2.4755
R29129 C10_P_btm.n28 C10_P_btm.t4 2.4755
R29130 C10_P_btm.n26 C10_P_btm.t0 2.4755
R29131 C10_P_btm.n26 C10_P_btm.t3 2.4755
R29132 C10_P_btm.n25 C10_P_btm.t5 2.4755
R29133 C10_P_btm.n25 C10_P_btm.t2 2.4755
R29134 C10_P_btm.n23 C10_P_btm.t32 2.4755
R29135 C10_P_btm.n23 C10_P_btm.t33 2.4755
R29136 C10_P_btm.n20 C10_P_btm.t10 2.4755
R29137 C10_P_btm.n20 C10_P_btm.t15 2.4755
R29138 C10_P_btm.n18 C10_P_btm.t9 2.4755
R29139 C10_P_btm.n18 C10_P_btm.t8 2.4755
R29140 C10_P_btm.n16 C10_P_btm.t12 2.4755
R29141 C10_P_btm.n16 C10_P_btm.t14 2.4755
R29142 C10_P_btm.n15 C10_P_btm.t11 2.4755
R29143 C10_P_btm.n15 C10_P_btm.t13 2.4755
R29144 C10_P_btm.n30 C10_P_btm.t7 2.4755
R29145 C10_P_btm.n30 C10_P_btm.t6 2.4755
R29146 C10_P_btm.n4 C10_P_btm.n2 0.71925
R29147 C10_P_btm.n8 C10_P_btm.n6 0.71925
R29148 C10_P_btm.n12 C10_P_btm.n10 0.71925
R29149 C10_P_btm.n6 C10_P_btm.n4 0.688
R29150 C10_P_btm.n10 C10_P_btm.n8 0.688
R29151 C10_P_btm.n14 C10_P_btm.n12 0.672375
R29152 C10_P_btm.n29 C10_P_btm.n27 0.5005
R29153 C10_P_btm.n19 C10_P_btm.n17 0.5005
R29154 C10_P_btm.n31 C10_P_btm.n29 0.484875
R29155 C10_P_btm.n21 C10_P_btm.n19 0.453625
R29156 C10_P_btm.n519 C10_P_btm.n518 0.276161
R29157 C10_P_btm.n768 C10_P_btm.n553 0.276161
R29158 C10_P_btm.n268 C10_P_btm.n174 0.276161
R29159 C10_P_btm.n130 C10_P_btm.n126 0.276161
R29160 C10_P_btm.n654 C10_P_btm.n653 0.276161
R29161 C10_P_btm.n265 C10_P_btm.n264 0.228786
R29162 C10_P_btm.n263 C10_P_btm.n176 0.228786
R29163 C10_P_btm.n261 C10_P_btm.n260 0.228786
R29164 C10_P_btm.n180 C10_P_btm.n177 0.228786
R29165 C10_P_btm.n195 C10_P_btm.n193 0.228786
R29166 C10_P_btm.n194 C10_P_btm.n175 0.228786
R29167 C10_P_btm.n267 C10_P_btm.n173 0.228786
R29168 C10_P_btm.n273 C10_P_btm.n171 0.228786
R29169 C10_P_btm.n172 C10_P_btm.n171 0.228786
R29170 C10_P_btm.n192 C10_P_btm.n191 0.228786
R29171 C10_P_btm.n191 C10_P_btm.n168 0.228786
R29172 C10_P_btm.n201 C10_P_btm.n190 0.228786
R29173 C10_P_btm.n200 C10_P_btm.n199 0.228786
R29174 C10_P_btm.n199 C10_P_btm.n198 0.228786
R29175 C10_P_btm.n197 C10_P_btm.n190 0.228786
R29176 C10_P_btm.n197 C10_P_btm.n196 0.228786
R29177 C10_P_btm.n188 C10_P_btm.n181 0.228786
R29178 C10_P_btm.n259 C10_P_btm.n181 0.228786
R29179 C10_P_btm.n258 C10_P_btm.n257 0.228786
R29180 C10_P_btm.n258 C10_P_btm.n179 0.228786
R29181 C10_P_btm.n187 C10_P_btm.n186 0.228786
R29182 C10_P_btm.n186 C10_P_btm.n185 0.228786
R29183 C10_P_btm.n184 C10_P_btm.n183 0.228786
R29184 C10_P_btm.n79 C10_P_btm.n78 0.228786
R29185 C10_P_btm.n355 C10_P_btm.n354 0.228786
R29186 C10_P_btm.n356 C10_P_btm.n77 0.228786
R29187 C10_P_btm.n1004 C10_P_btm.n357 0.228786
R29188 C10_P_btm.n1003 C10_P_btm.n1002 0.228786
R29189 C10_P_btm.n1001 C10_P_btm.n358 0.228786
R29190 C10_P_btm.n1000 C10_P_btm.n359 0.228786
R29191 C10_P_btm.n999 C10_P_btm.n998 0.228786
R29192 C10_P_btm.n997 C10_P_btm.n360 0.228786
R29193 C10_P_btm.n385 C10_P_btm.n362 0.228786
R29194 C10_P_btm.n387 C10_P_btm.n386 0.228786
R29195 C10_P_btm.n384 C10_P_btm.n383 0.228786
R29196 C10_P_btm.n425 C10_P_btm.n421 0.228786
R29197 C10_P_btm.n424 C10_P_btm.n423 0.228786
R29198 C10_P_btm.n406 C10_P_btm.n405 0.228786
R29199 C10_P_btm.n945 C10_P_btm.n944 0.228786
R29200 C10_P_btm.n944 C10_P_btm.n943 0.228786
R29201 C10_P_btm.n408 C10_P_btm.n404 0.228786
R29202 C10_P_btm.n927 C10_P_btm.n403 0.228786
R29203 C10_P_btm.n928 C10_P_btm.n402 0.228786
R29204 C10_P_btm.n923 C10_P_btm.n401 0.228786
R29205 C10_P_btm.n922 C10_P_btm.n400 0.228786
R29206 C10_P_btm.n921 C10_P_btm.n399 0.228786
R29207 C10_P_btm.n896 C10_P_btm.n398 0.228786
R29208 C10_P_btm.n905 C10_P_btm.n397 0.228786
R29209 C10_P_btm.n904 C10_P_btm.n396 0.228786
R29210 C10_P_btm.n381 C10_P_btm.n380 0.228786
R29211 C10_P_btm.n958 C10_P_btm.n957 0.228786
R29212 C10_P_btm.n382 C10_P_btm.n378 0.228786
R29213 C10_P_btm.n393 C10_P_btm.n392 0.228786
R29214 C10_P_btm.n392 C10_P_btm.n376 0.228786
R29215 C10_P_btm.n391 C10_P_btm.n390 0.228786
R29216 C10_P_btm.n389 C10_P_btm.n388 0.228786
R29217 C10_P_btm.n364 C10_P_btm.n363 0.228786
R29218 C10_P_btm.n996 C10_P_btm.n995 0.228786
R29219 C10_P_btm.n365 C10_P_btm.n361 0.228786
R29220 C10_P_btm.n981 C10_P_btm.n980 0.228786
R29221 C10_P_btm.n979 C10_P_btm.n978 0.228786
R29222 C10_P_btm.n75 C10_P_btm.n74 0.228786
R29223 C10_P_btm.n1006 C10_P_btm.n1005 0.228786
R29224 C10_P_btm.n76 C10_P_btm.n72 0.228786
R29225 C10_P_btm.n353 C10_P_btm.n352 0.228786
R29226 C10_P_btm.n351 C10_P_btm.n80 0.228786
R29227 C10_P_btm.n182 C10_P_btm.n81 0.228786
R29228 C10_P_btm.n82 C10_P_btm.n81 0.228786
R29229 C10_P_btm.n256 C10_P_btm.n255 0.228786
R29230 C10_P_btm.n255 C10_P_btm.n83 0.228786
R29231 C10_P_btm.n254 C10_P_btm.n253 0.228786
R29232 C10_P_btm.n252 C10_P_btm.n251 0.228786
R29233 C10_P_btm.n189 C10_P_btm.n86 0.228786
R29234 C10_P_btm.n343 C10_P_btm.n86 0.228786
R29235 C10_P_btm.n250 C10_P_btm.n88 0.228786
R29236 C10_P_btm.n249 C10_P_btm.n248 0.228786
R29237 C10_P_btm.n167 C10_P_btm.n166 0.228786
R29238 C10_P_btm.n276 C10_P_btm.n275 0.228786
R29239 C10_P_btm.n274 C10_P_btm.n164 0.228786
R29240 C10_P_btm.n279 C10_P_btm.n278 0.228786
R29241 C10_P_btm.n277 C10_P_btm.n159 0.228786
R29242 C10_P_btm.n202 C10_P_btm.n165 0.228786
R29243 C10_P_btm.n247 C10_P_btm.n246 0.228786
R29244 C10_P_btm.n90 C10_P_btm.n89 0.228786
R29245 C10_P_btm.n342 C10_P_btm.n341 0.228786
R29246 C10_P_btm.n341 C10_P_btm.n91 0.228786
R29247 C10_P_btm.n92 C10_P_btm.n91 0.228786
R29248 C10_P_btm.n204 C10_P_btm.n203 0.228786
R29249 C10_P_btm.n245 C10_P_btm.n244 0.228786
R29250 C10_P_btm.n158 C10_P_btm.n157 0.228786
R29251 C10_P_btm.n282 C10_P_btm.n281 0.228786
R29252 C10_P_btm.n280 C10_P_btm.n155 0.228786
R29253 C10_P_btm.n285 C10_P_btm.n284 0.228786
R29254 C10_P_btm.n283 C10_P_btm.n150 0.228786
R29255 C10_P_btm.n206 C10_P_btm.n156 0.228786
R29256 C10_P_btm.n243 C10_P_btm.n242 0.228786
R29257 C10_P_btm.n241 C10_P_btm.n205 0.228786
R29258 C10_P_btm.n94 C10_P_btm.n93 0.228786
R29259 C10_P_btm.n95 C10_P_btm.n94 0.228786
R29260 C10_P_btm.n96 C10_P_btm.n95 0.228786
R29261 C10_P_btm.n240 C10_P_btm.n239 0.228786
R29262 C10_P_btm.n238 C10_P_btm.n207 0.228786
R29263 C10_P_btm.n149 C10_P_btm.n148 0.228786
R29264 C10_P_btm.n288 C10_P_btm.n287 0.228786
R29265 C10_P_btm.n286 C10_P_btm.n146 0.228786
R29266 C10_P_btm.n291 C10_P_btm.n290 0.228786
R29267 C10_P_btm.n289 C10_P_btm.n144 0.228786
R29268 C10_P_btm.n209 C10_P_btm.n147 0.228786
R29269 C10_P_btm.n237 C10_P_btm.n236 0.228786
R29270 C10_P_btm.n235 C10_P_btm.n208 0.228786
R29271 C10_P_btm.n98 C10_P_btm.n97 0.228786
R29272 C10_P_btm.n99 C10_P_btm.n98 0.228786
R29273 C10_P_btm.n100 C10_P_btm.n99 0.228786
R29274 C10_P_btm.n234 C10_P_btm.n233 0.228786
R29275 C10_P_btm.n232 C10_P_btm.n210 0.228786
R29276 C10_P_btm.n213 C10_P_btm.n212 0.228786
R29277 C10_P_btm.n215 C10_P_btm.n143 0.228786
R29278 C10_P_btm.n292 C10_P_btm.n141 0.228786
R29279 C10_P_btm.n298 C10_P_btm.n139 0.228786
R29280 C10_P_btm.n140 C10_P_btm.n139 0.228786
R29281 C10_P_btm.n217 C10_P_btm.n216 0.228786
R29282 C10_P_btm.n218 C10_P_btm.n214 0.228786
R29283 C10_P_btm.n231 C10_P_btm.n230 0.228786
R29284 C10_P_btm.n229 C10_P_btm.n211 0.228786
R29285 C10_P_btm.n102 C10_P_btm.n101 0.228786
R29286 C10_P_btm.n103 C10_P_btm.n102 0.228786
R29287 C10_P_btm.n104 C10_P_btm.n103 0.228786
R29288 C10_P_btm.n228 C10_P_btm.n227 0.228786
R29289 C10_P_btm.n221 C10_P_btm.n220 0.228786
R29290 C10_P_btm.n219 C10_P_btm.n124 0.228786
R29291 C10_P_btm.n300 C10_P_btm.n125 0.228786
R29292 C10_P_btm.n301 C10_P_btm.n300 0.228786
R29293 C10_P_btm.n299 C10_P_btm.n123 0.228786
R29294 C10_P_btm.n121 C10_P_btm.n120 0.228786
R29295 C10_P_btm.n303 C10_P_btm.n302 0.228786
R29296 C10_P_btm.n304 C10_P_btm.n119 0.228786
R29297 C10_P_btm.n122 C10_P_btm.n119 0.228786
R29298 C10_P_btm.n223 C10_P_btm.n222 0.228786
R29299 C10_P_btm.n226 C10_P_btm.n225 0.228786
R29300 C10_P_btm.n106 C10_P_btm.n105 0.228786
R29301 C10_P_btm.n107 C10_P_btm.n106 0.228786
R29302 C10_P_btm.n108 C10_P_btm.n107 0.228786
R29303 C10_P_btm.n224 C10_P_btm.n116 0.228786
R29304 C10_P_btm.n306 C10_P_btm.n117 0.228786
R29305 C10_P_btm.n307 C10_P_btm.n306 0.228786
R29306 C10_P_btm.n305 C10_P_btm.n115 0.228786
R29307 C10_P_btm.n127 C10_P_btm.n118 0.228786
R29308 C10_P_btm.n133 C10_P_btm.n132 0.228786
R29309 C10_P_btm.n129 C10_P_btm.n128 0.228786
R29310 C10_P_btm.n113 C10_P_btm.n112 0.228786
R29311 C10_P_btm.n309 C10_P_btm.n308 0.228786
R29312 C10_P_btm.n310 C10_P_btm.n111 0.228786
R29313 C10_P_btm.n114 C10_P_btm.n111 0.228786
R29314 C10_P_btm.n110 C10_P_btm.n109 0.228786
R29315 C10_P_btm.n311 C10_P_btm.n110 0.228786
R29316 C10_P_btm.n312 C10_P_btm.n35 0.228786
R29317 C10_P_btm.n314 C10_P_btm.n313 0.228786
R29318 C10_P_btm.n315 C10_P_btm.n314 0.228786
R29319 C10_P_btm.n36 C10_P_btm.n35 0.228786
R29320 C10_P_btm.n38 C10_P_btm.n36 0.228786
R29321 C10_P_btm.n316 C10_P_btm.n315 0.228786
R29322 C10_P_btm.n317 C10_P_btm.n316 0.228786
R29323 C10_P_btm.n39 C10_P_btm.n38 0.228786
R29324 C10_P_btm.n319 C10_P_btm.n39 0.228786
R29325 C10_P_btm.n318 C10_P_btm.n317 0.228786
R29326 C10_P_btm.n321 C10_P_btm.n318 0.228786
R29327 C10_P_btm.n320 C10_P_btm.n319 0.228786
R29328 C10_P_btm.n320 C10_P_btm.n43 0.228786
R29329 C10_P_btm.n322 C10_P_btm.n321 0.228786
R29330 C10_P_btm.n323 C10_P_btm.n322 0.228786
R29331 C10_P_btm.n44 C10_P_btm.n43 0.228786
R29332 C10_P_btm.n46 C10_P_btm.n44 0.228786
R29333 C10_P_btm.n324 C10_P_btm.n323 0.228786
R29334 C10_P_btm.n325 C10_P_btm.n324 0.228786
R29335 C10_P_btm.n47 C10_P_btm.n46 0.228786
R29336 C10_P_btm.n327 C10_P_btm.n47 0.228786
R29337 C10_P_btm.n326 C10_P_btm.n325 0.228786
R29338 C10_P_btm.n329 C10_P_btm.n326 0.228786
R29339 C10_P_btm.n328 C10_P_btm.n327 0.228786
R29340 C10_P_btm.n328 C10_P_btm.n51 0.228786
R29341 C10_P_btm.n330 C10_P_btm.n329 0.228786
R29342 C10_P_btm.n331 C10_P_btm.n330 0.228786
R29343 C10_P_btm.n52 C10_P_btm.n51 0.228786
R29344 C10_P_btm.n54 C10_P_btm.n52 0.228786
R29345 C10_P_btm.n332 C10_P_btm.n331 0.228786
R29346 C10_P_btm.n333 C10_P_btm.n332 0.228786
R29347 C10_P_btm.n55 C10_P_btm.n54 0.228786
R29348 C10_P_btm.n335 C10_P_btm.n55 0.228786
R29349 C10_P_btm.n334 C10_P_btm.n333 0.228786
R29350 C10_P_btm.n337 C10_P_btm.n334 0.228786
R29351 C10_P_btm.n336 C10_P_btm.n335 0.228786
R29352 C10_P_btm.n336 C10_P_btm.n59 0.228786
R29353 C10_P_btm.n338 C10_P_btm.n337 0.228786
R29354 C10_P_btm.n339 C10_P_btm.n338 0.228786
R29355 C10_P_btm.n60 C10_P_btm.n59 0.228786
R29356 C10_P_btm.n62 C10_P_btm.n60 0.228786
R29357 C10_P_btm.n340 C10_P_btm.n339 0.228786
R29358 C10_P_btm.n340 C10_P_btm.n87 0.228786
R29359 C10_P_btm.n63 C10_P_btm.n62 0.228786
R29360 C10_P_btm.n85 C10_P_btm.n63 0.228786
R29361 C10_P_btm.n346 C10_P_btm.n85 0.228786
R29362 C10_P_btm.n345 C10_P_btm.n344 0.228786
R29363 C10_P_btm.n345 C10_P_btm.n84 0.228786
R29364 C10_P_btm.n67 C10_P_btm.n66 0.228786
R29365 C10_P_btm.n347 C10_P_btm.n346 0.228786
R29366 C10_P_btm.n348 C10_P_btm.n347 0.228786
R29367 C10_P_btm.n349 C10_P_btm.n67 0.228786
R29368 C10_P_btm.n350 C10_P_btm.n349 0.228786
R29369 C10_P_btm.n71 C10_P_btm.n68 0.228786
R29370 C10_P_btm.n1011 C10_P_btm.n68 0.228786
R29371 C10_P_btm.n1009 C10_P_btm.n1008 0.228786
R29372 C10_P_btm.n1007 C10_P_btm.n70 0.228786
R29373 C10_P_btm.n975 C10_P_btm.n73 0.228786
R29374 C10_P_btm.n977 C10_P_btm.n976 0.228786
R29375 C10_P_btm.n983 C10_P_btm.n982 0.228786
R29376 C10_P_btm.n969 C10_P_btm.n366 0.228786
R29377 C10_P_btm.n994 C10_P_btm.n367 0.228786
R29378 C10_P_btm.n993 C10_P_btm.n992 0.228786
R29379 C10_P_btm.n991 C10_P_btm.n368 0.228786
R29380 C10_P_btm.n375 C10_P_btm.n370 0.228786
R29381 C10_P_btm.n963 C10_P_btm.n962 0.228786
R29382 C10_P_btm.n961 C10_P_btm.n374 0.228786
R29383 C10_P_btm.n961 C10_P_btm.n960 0.228786
R29384 C10_P_btm.n959 C10_P_btm.n377 0.228786
R29385 C10_P_btm.n910 C10_P_btm.n377 0.228786
R29386 C10_P_btm.n911 C10_P_btm.n379 0.228786
R29387 C10_P_btm.n908 C10_P_btm.n903 0.228786
R29388 C10_P_btm.n907 C10_P_btm.n906 0.228786
R29389 C10_P_btm.n898 C10_P_btm.n897 0.228786
R29390 C10_P_btm.n920 C10_P_btm.n919 0.228786
R29391 C10_P_btm.n895 C10_P_btm.n894 0.228786
R29392 C10_P_btm.n931 C10_P_btm.n930 0.228786
R29393 C10_P_btm.n929 C10_P_btm.n892 0.228786
R29394 C10_P_btm.n926 C10_P_btm.n925 0.228786
R29395 C10_P_btm.n924 C10_P_btm.n409 0.228786
R29396 C10_P_btm.n942 C10_P_btm.n410 0.228786
R29397 C10_P_btm.n941 C10_P_btm.n940 0.228786
R29398 C10_P_btm.n941 C10_P_btm.n407 0.228786
R29399 C10_P_btm.n422 C10_P_btm.n411 0.228786
R29400 C10_P_btm.n412 C10_P_btm.n411 0.228786
R29401 C10_P_btm.n883 C10_P_btm.n882 0.228786
R29402 C10_P_btm.n884 C10_P_btm.n416 0.228786
R29403 C10_P_btm.n420 C10_P_btm.n416 0.228786
R29404 C10_P_btm.n882 C10_P_btm.n881 0.228786
R29405 C10_P_btm.n881 C10_P_btm.n880 0.228786
R29406 C10_P_btm.n879 C10_P_btm.n419 0.228786
R29407 C10_P_btm.n879 C10_P_btm.n878 0.228786
R29408 C10_P_btm.n877 C10_P_btm.n427 0.228786
R29409 C10_P_btm.n876 C10_P_btm.n428 0.228786
R29410 C10_P_btm.n875 C10_P_btm.n874 0.228786
R29411 C10_P_btm.n873 C10_P_btm.n429 0.228786
R29412 C10_P_btm.n451 C10_P_btm.n431 0.228786
R29413 C10_P_btm.n453 C10_P_btm.n452 0.228786
R29414 C10_P_btm.n459 C10_P_btm.n458 0.228786
R29415 C10_P_btm.n460 C10_P_btm.n450 0.228786
R29416 C10_P_btm.n837 C10_P_btm.n461 0.228786
R29417 C10_P_btm.n833 C10_P_btm.n832 0.228786
R29418 C10_P_btm.n832 C10_P_btm.n831 0.228786
R29419 C10_P_btm.n830 C10_P_btm.n462 0.228786
R29420 C10_P_btm.n836 C10_P_btm.n448 0.228786
R29421 C10_P_btm.n448 C10_P_btm.n447 0.228786
R29422 C10_P_btm.n839 C10_P_btm.n838 0.228786
R29423 C10_P_btm.n449 C10_P_btm.n445 0.228786
R29424 C10_P_btm.n457 C10_P_btm.n456 0.228786
R29425 C10_P_btm.n455 C10_P_btm.n454 0.228786
R29426 C10_P_btm.n433 C10_P_btm.n432 0.228786
R29427 C10_P_btm.n872 C10_P_btm.n871 0.228786
R29428 C10_P_btm.n434 C10_P_btm.n430 0.228786
R29429 C10_P_btm.n857 C10_P_btm.n856 0.228786
R29430 C10_P_btm.n855 C10_P_btm.n854 0.228786
R29431 C10_P_btm.n418 C10_P_btm.n417 0.228786
R29432 C10_P_btm.n853 C10_P_btm.n852 0.228786
R29433 C10_P_btm.n859 C10_P_btm.n858 0.228786
R29434 C10_P_btm.n848 C10_P_btm.n435 0.228786
R29435 C10_P_btm.n870 C10_P_btm.n436 0.228786
R29436 C10_P_btm.n869 C10_P_btm.n868 0.228786
R29437 C10_P_btm.n867 C10_P_btm.n437 0.228786
R29438 C10_P_btm.n444 C10_P_btm.n439 0.228786
R29439 C10_P_btm.n842 C10_P_btm.n841 0.228786
R29440 C10_P_btm.n840 C10_P_btm.n443 0.228786
R29441 C10_P_btm.n826 C10_P_btm.n446 0.228786
R29442 C10_P_btm.n828 C10_P_btm.n827 0.228786
R29443 C10_P_btm.n829 C10_P_btm.n828 0.228786
R29444 C10_P_btm.n467 C10_P_btm.n465 0.228786
R29445 C10_P_btm.n468 C10_P_btm.n467 0.228786
R29446 C10_P_btm.n818 C10_P_btm.n471 0.228786
R29447 C10_P_btm.n818 C10_P_btm.n817 0.228786
R29448 C10_P_btm.n819 C10_P_btm.n472 0.228786
R29449 C10_P_btm.n476 C10_P_btm.n472 0.228786
R29450 C10_P_btm.n817 C10_P_btm.n816 0.228786
R29451 C10_P_btm.n816 C10_P_btm.n815 0.228786
R29452 C10_P_btm.n476 C10_P_btm.n466 0.228786
R29453 C10_P_btm.n466 C10_P_btm.n464 0.228786
R29454 C10_P_btm.n815 C10_P_btm.n814 0.228786
R29455 C10_P_btm.n814 C10_P_btm.n813 0.228786
R29456 C10_P_btm.n812 C10_P_btm.n478 0.228786
R29457 C10_P_btm.n810 C10_P_btm.n809 0.228786
R29458 C10_P_btm.n477 C10_P_btm.n475 0.228786
R29459 C10_P_btm.n721 C10_P_btm.n481 0.228786
R29460 C10_P_btm.n474 C10_P_btm.n473 0.228786
R29461 C10_P_btm.n723 C10_P_btm.n722 0.228786
R29462 C10_P_btm.n725 C10_P_btm.n685 0.228786
R29463 C10_P_btm.n724 C10_P_btm.n683 0.228786
R29464 C10_P_btm.n690 C10_P_btm.n688 0.228786
R29465 C10_P_btm.n716 C10_P_btm.n688 0.228786
R29466 C10_P_btm.n715 C10_P_btm.n714 0.228786
R29467 C10_P_btm.n715 C10_P_btm.n686 0.228786
R29468 C10_P_btm.n717 C10_P_btm.n716 0.228786
R29469 C10_P_btm.n718 C10_P_btm.n717 0.228786
R29470 C10_P_btm.n719 C10_P_btm.n686 0.228786
R29471 C10_P_btm.n720 C10_P_btm.n719 0.228786
R29472 C10_P_btm.n718 C10_P_btm.n485 0.228786
R29473 C10_P_btm.n805 C10_P_btm.n485 0.228786
R29474 C10_P_btm.n720 C10_P_btm.n483 0.228786
R29475 C10_P_btm.n807 C10_P_btm.n483 0.228786
R29476 C10_P_btm.n806 C10_P_btm.n805 0.228786
R29477 C10_P_btm.n806 C10_P_btm.n482 0.228786
R29478 C10_P_btm.n808 C10_P_btm.n807 0.228786
R29479 C10_P_btm.n808 C10_P_btm.n480 0.228786
R29480 C10_P_btm.n504 C10_P_btm.n482 0.228786
R29481 C10_P_btm.n506 C10_P_btm.n504 0.228786
R29482 C10_P_btm.n508 C10_P_btm.n507 0.228786
R29483 C10_P_btm.n510 C10_P_btm.n503 0.228786
R29484 C10_P_btm.n509 C10_P_btm.n484 0.228786
R29485 C10_P_btm.n511 C10_P_btm.n486 0.228786
R29486 C10_P_btm.n804 C10_P_btm.n803 0.228786
R29487 C10_P_btm.n802 C10_P_btm.n801 0.228786
R29488 C10_P_btm.n687 C10_P_btm.n487 0.228786
R29489 C10_P_btm.n705 C10_P_btm.n489 0.228786
R29490 C10_P_btm.n704 C10_P_btm.n689 0.228786
R29491 C10_P_btm.n707 C10_P_btm.n706 0.228786
R29492 C10_P_btm.n709 C10_P_btm.n692 0.228786
R29493 C10_P_btm.n708 C10_P_btm.n699 0.228786
R29494 C10_P_btm.n534 C10_P_btm.n532 0.228786
R29495 C10_P_btm.n532 C10_P_btm.n531 0.228786
R29496 C10_P_btm.n698 C10_P_btm.n697 0.228786
R29497 C10_P_btm.n698 C10_P_btm.n693 0.228786
R29498 C10_P_btm.n700 C10_P_btm.n531 0.228786
R29499 C10_P_btm.n701 C10_P_btm.n700 0.228786
R29500 C10_P_btm.n702 C10_P_btm.n693 0.228786
R29501 C10_P_btm.n703 C10_P_btm.n702 0.228786
R29502 C10_P_btm.n701 C10_P_btm.n493 0.228786
R29503 C10_P_btm.n797 C10_P_btm.n493 0.228786
R29504 C10_P_btm.n703 C10_P_btm.n491 0.228786
R29505 C10_P_btm.n799 C10_P_btm.n491 0.228786
R29506 C10_P_btm.n798 C10_P_btm.n797 0.228786
R29507 C10_P_btm.n798 C10_P_btm.n490 0.228786
R29508 C10_P_btm.n800 C10_P_btm.n799 0.228786
R29509 C10_P_btm.n800 C10_P_btm.n488 0.228786
R29510 C10_P_btm.n495 C10_P_btm.n490 0.228786
R29511 C10_P_btm.n497 C10_P_btm.n495 0.228786
R29512 C10_P_btm.n512 C10_P_btm.n488 0.228786
R29513 C10_P_btm.n513 C10_P_btm.n512 0.228786
R29514 C10_P_btm.n498 C10_P_btm.n497 0.228786
R29515 C10_P_btm.n515 C10_P_btm.n498 0.228786
R29516 C10_P_btm.n514 C10_P_btm.n513 0.228786
R29517 C10_P_btm.n514 C10_P_btm.n502 0.228786
R29518 C10_P_btm.n516 C10_P_btm.n515 0.228786
R29519 C10_P_btm.n517 C10_P_btm.n516 0.228786
R29520 C10_P_btm.n521 C10_P_btm.n499 0.228786
R29521 C10_P_btm.n520 C10_P_btm.n496 0.228786
R29522 C10_P_btm.n523 C10_P_btm.n522 0.228786
R29523 C10_P_btm.n525 C10_P_btm.n494 0.228786
R29524 C10_P_btm.n524 C10_P_btm.n492 0.228786
R29525 C10_P_btm.n527 C10_P_btm.n526 0.228786
R29526 C10_P_btm.n796 C10_P_btm.n795 0.228786
R29527 C10_P_btm.n794 C10_P_btm.n793 0.228786
R29528 C10_P_btm.n529 C10_P_btm.n528 0.228786
R29529 C10_P_btm.n792 C10_P_btm.n791 0.228786
R29530 C10_P_btm.n790 C10_P_btm.n789 0.228786
R29531 C10_P_btm.n533 C10_P_btm.n530 0.228786
R29532 C10_P_btm.n788 C10_P_btm.n787 0.228786
R29533 C10_P_btm.n786 C10_P_btm.n785 0.228786
R29534 C10_P_btm.n785 C10_P_btm.n784 0.228786
R29535 C10_P_btm.n731 C10_P_btm.n680 0.228786
R29536 C10_P_btm.n733 C10_P_btm.n603 0.228786
R29537 C10_P_btm.n735 C10_P_btm.n600 0.228786
R29538 C10_P_btm.n734 C10_P_btm.n733 0.228786
R29539 C10_P_btm.n732 C10_P_btm.n601 0.228786
R29540 C10_P_btm.n675 C10_P_btm.n604 0.228786
R29541 C10_P_btm.n606 C10_P_btm.n602 0.228786
R29542 C10_P_btm.n633 C10_P_btm.n598 0.228786
R29543 C10_P_btm.n737 C10_P_btm.n595 0.228786
R29544 C10_P_btm.n740 C10_P_btm.n739 0.228786
R29545 C10_P_btm.n741 C10_P_btm.n593 0.228786
R29546 C10_P_btm.n592 C10_P_btm.n590 0.228786
R29547 C10_P_btm.n742 C10_P_btm.n741 0.228786
R29548 C10_P_btm.n740 C10_P_btm.n587 0.228786
R29549 C10_P_btm.n632 C10_P_btm.n594 0.228786
R29550 C10_P_btm.n635 C10_P_btm.n634 0.228786
R29551 C10_P_btm.n608 C10_P_btm.n607 0.228786
R29552 C10_P_btm.n674 C10_P_btm.n673 0.228786
R29553 C10_P_btm.n669 C10_P_btm.n609 0.228786
R29554 C10_P_btm.n631 C10_P_btm.n611 0.228786
R29555 C10_P_btm.n637 C10_P_btm.n636 0.228786
R29556 C10_P_btm.n586 C10_P_btm.n585 0.228786
R29557 C10_P_btm.n745 C10_P_btm.n744 0.228786
R29558 C10_P_btm.n743 C10_P_btm.n583 0.228786
R29559 C10_P_btm.n589 C10_P_btm.n588 0.228786
R29560 C10_P_btm.n541 C10_P_btm.n539 0.228786
R29561 C10_P_btm.n542 C10_P_btm.n541 0.228786
R29562 C10_P_btm.n580 C10_P_btm.n542 0.228786
R29563 C10_P_btm.n582 C10_P_btm.n581 0.228786
R29564 C10_P_btm.n748 C10_P_btm.n747 0.228786
R29565 C10_P_btm.n746 C10_P_btm.n576 0.228786
R29566 C10_P_btm.n630 C10_P_btm.n584 0.228786
R29567 C10_P_btm.n639 C10_P_btm.n638 0.228786
R29568 C10_P_btm.n613 C10_P_btm.n612 0.228786
R29569 C10_P_btm.n668 C10_P_btm.n667 0.228786
R29570 C10_P_btm.n663 C10_P_btm.n614 0.228786
R29571 C10_P_btm.n629 C10_P_btm.n616 0.228786
R29572 C10_P_btm.n641 C10_P_btm.n640 0.228786
R29573 C10_P_btm.n575 C10_P_btm.n574 0.228786
R29574 C10_P_btm.n751 C10_P_btm.n750 0.228786
R29575 C10_P_btm.n749 C10_P_btm.n572 0.228786
R29576 C10_P_btm.n578 C10_P_btm.n577 0.228786
R29577 C10_P_btm.n579 C10_P_btm.n546 0.228786
R29578 C10_P_btm.n547 C10_P_btm.n546 0.228786
R29579 C10_P_btm.n549 C10_P_btm.n547 0.228786
R29580 C10_P_btm.n571 C10_P_btm.n570 0.228786
R29581 C10_P_btm.n754 C10_P_btm.n753 0.228786
R29582 C10_P_btm.n752 C10_P_btm.n565 0.228786
R29583 C10_P_btm.n628 C10_P_btm.n573 0.228786
R29584 C10_P_btm.n643 C10_P_btm.n642 0.228786
R29585 C10_P_btm.n618 C10_P_btm.n617 0.228786
R29586 C10_P_btm.n662 C10_P_btm.n661 0.228786
R29587 C10_P_btm.n657 C10_P_btm.n619 0.228786
R29588 C10_P_btm.n627 C10_P_btm.n621 0.228786
R29589 C10_P_btm.n645 C10_P_btm.n644 0.228786
R29590 C10_P_btm.n564 C10_P_btm.n563 0.228786
R29591 C10_P_btm.n757 C10_P_btm.n756 0.228786
R29592 C10_P_btm.n755 C10_P_btm.n561 0.228786
R29593 C10_P_btm.n569 C10_P_btm.n568 0.228786
R29594 C10_P_btm.n567 C10_P_btm.n550 0.228786
R29595 C10_P_btm.n567 C10_P_btm.n566 0.228786
R29596 C10_P_btm.n566 C10_P_btm.n554 0.228786
R29597 C10_P_btm.n560 C10_P_btm.n558 0.228786
R29598 C10_P_btm.n760 C10_P_btm.n759 0.228786
R29599 C10_P_btm.n758 C10_P_btm.n559 0.228786
R29600 C10_P_btm.n648 C10_P_btm.n562 0.228786
R29601 C10_P_btm.n647 C10_P_btm.n646 0.228786
R29602 C10_P_btm.n623 C10_P_btm.n622 0.228786
R29603 C10_P_btm.n656 C10_P_btm.n655 0.228786
R29604 C10_P_btm.n652 C10_P_btm.n625 0.228786
R29605 C10_P_btm.n651 C10_P_btm.n650 0.228786
R29606 C10_P_btm.n649 C10_P_btm.n626 0.228786
R29607 C10_P_btm.n557 C10_P_btm.n556 0.228786
R29608 C10_P_btm.n762 C10_P_btm.n761 0.228786
R29609 C10_P_btm.n763 C10_P_btm.n555 0.228786
R29610 C10_P_btm.n765 C10_P_btm.n764 0.228786
R29611 C10_P_btm.n767 C10_P_btm.n766 0.228786
R29612 C10_P_btm.n767 C10_P_btm.n552 0.228786
R29613 C10_P_btm.n769 C10_P_btm.n768 0.228786
R29614 C10_P_btm.n770 C10_P_btm.n769 0.228786
R29615 C10_P_btm.n552 C10_P_btm.n551 0.228786
R29616 C10_P_btm.n772 C10_P_btm.n551 0.228786
R29617 C10_P_btm.n771 C10_P_btm.n770 0.228786
R29618 C10_P_btm.n771 C10_P_btm.n548 0.228786
R29619 C10_P_btm.n773 C10_P_btm.n772 0.228786
R29620 C10_P_btm.n774 C10_P_btm.n773 0.228786
R29621 C10_P_btm.n548 C10_P_btm.n545 0.228786
R29622 C10_P_btm.n776 C10_P_btm.n545 0.228786
R29623 C10_P_btm.n775 C10_P_btm.n774 0.228786
R29624 C10_P_btm.n775 C10_P_btm.n544 0.228786
R29625 C10_P_btm.n777 C10_P_btm.n776 0.228786
R29626 C10_P_btm.n778 C10_P_btm.n777 0.228786
R29627 C10_P_btm.n544 C10_P_btm.n543 0.228786
R29628 C10_P_btm.n780 C10_P_btm.n543 0.228786
R29629 C10_P_btm.n779 C10_P_btm.n778 0.228786
R29630 C10_P_btm.n779 C10_P_btm.n540 0.228786
R29631 C10_P_btm.n781 C10_P_btm.n780 0.228786
R29632 C10_P_btm.n782 C10_P_btm.n781 0.228786
R29633 C10_P_btm.n540 C10_P_btm.n537 0.228786
R29634 C10_P_btm.n784 C10_P_btm.n537 0.228786
R29635 C10_P_btm.n783 C10_P_btm.n782 0.228786
R29636 C10_P_btm.n783 C10_P_btm.n536 0.228786
R29637 C10_P_btm.n591 C10_P_btm.n538 0.228786
R29638 C10_P_btm.n591 C10_P_btm.n535 0.228786
R29639 C10_P_btm.n695 C10_P_btm.n592 0.228786
R29640 C10_P_btm.n696 C10_P_btm.n695 0.228786
R29641 C10_P_btm.n596 C10_P_btm.n593 0.228786
R29642 C10_P_btm.n694 C10_P_btm.n596 0.228786
R29643 C10_P_btm.n738 C10_P_btm.n597 0.228786
R29644 C10_P_btm.n691 C10_P_btm.n597 0.228786
R29645 C10_P_btm.n736 C10_P_btm.n599 0.228786
R29646 C10_P_btm.n710 C10_P_btm.n599 0.228786
R29647 C10_P_btm.n711 C10_P_btm.n600 0.228786
R29648 C10_P_btm.n713 C10_P_btm.n711 0.228786
R29649 C10_P_btm.n712 C10_P_btm.n603 0.228786
R29650 C10_P_btm.n712 C10_P_btm.n682 0.228786
R29651 C10_P_btm.n727 C10_P_btm.n680 0.228786
R29652 C10_P_btm.n727 C10_P_btm.n726 0.228786
R29653 C10_P_btm.n820 C10_P_btm.n470 0.228786
R29654 C10_P_btm.n822 C10_P_btm.n821 0.228786
R29655 C10_P_btm.n823 C10_P_btm.n469 0.228786
R29656 C10_P_btm.n825 C10_P_btm.n824 0.228786
R29657 C10_P_btm.n442 C10_P_btm.n441 0.228786
R29658 C10_P_btm.n844 C10_P_btm.n843 0.228786
R29659 C10_P_btm.n845 C10_P_btm.n440 0.228786
R29660 C10_P_btm.n866 C10_P_btm.n865 0.228786
R29661 C10_P_btm.n864 C10_P_btm.n438 0.228786
R29662 C10_P_btm.n863 C10_P_btm.n846 0.228786
R29663 C10_P_btm.n862 C10_P_btm.n861 0.228786
R29664 C10_P_btm.n850 C10_P_btm.n849 0.228786
R29665 C10_P_btm.n415 C10_P_btm.n414 0.228786
R29666 C10_P_btm.n886 C10_P_btm.n885 0.228786
R29667 C10_P_btm.n887 C10_P_btm.n413 0.228786
R29668 C10_P_btm.n939 C10_P_btm.n888 0.228786
R29669 C10_P_btm.n938 C10_P_btm.n937 0.228786
R29670 C10_P_btm.n936 C10_P_btm.n889 0.228786
R29671 C10_P_btm.n935 C10_P_btm.n890 0.228786
R29672 C10_P_btm.n934 C10_P_btm.n933 0.228786
R29673 C10_P_btm.n932 C10_P_btm.n891 0.228786
R29674 C10_P_btm.n900 C10_P_btm.n893 0.228786
R29675 C10_P_btm.n918 C10_P_btm.n917 0.228786
R29676 C10_P_btm.n916 C10_P_btm.n899 0.228786
R29677 C10_P_btm.n915 C10_P_btm.n901 0.228786
R29678 C10_P_btm.n914 C10_P_btm.n913 0.228786
R29679 C10_P_btm.n912 C10_P_btm.n902 0.228786
R29680 C10_P_btm.n965 C10_P_btm.n964 0.228786
R29681 C10_P_btm.n966 C10_P_btm.n371 0.228786
R29682 C10_P_btm.n990 C10_P_btm.n989 0.228786
R29683 C10_P_btm.n988 C10_P_btm.n369 0.228786
R29684 C10_P_btm.n987 C10_P_btm.n967 0.228786
R29685 C10_P_btm.n986 C10_P_btm.n985 0.228786
R29686 C10_P_btm.n984 C10_P_btm.n968 0.228786
R29687 C10_P_btm.n971 C10_P_btm.n970 0.228786
R29688 C10_P_btm.n974 C10_P_btm.n973 0.228786
R29689 C10_P_btm.n972 C10_P_btm.n69 0.228786
R29690 C10_P_btm.n1010 C10_P_btm.n65 0.228786
R29691 C10_P_btm.n1013 C10_P_btm.n1012 0.228786
R29692 C10_P_btm.n1015 C10_P_btm.n64 0.228786
R29693 C10_P_btm.n1014 C10_P_btm.n61 0.228786
R29694 C10_P_btm.n1017 C10_P_btm.n1016 0.228786
R29695 C10_P_btm.n1019 C10_P_btm.n58 0.228786
R29696 C10_P_btm.n1018 C10_P_btm.n57 0.228786
R29697 C10_P_btm.n1021 C10_P_btm.n1020 0.228786
R29698 C10_P_btm.n1023 C10_P_btm.n56 0.228786
R29699 C10_P_btm.n1022 C10_P_btm.n53 0.228786
R29700 C10_P_btm.n1025 C10_P_btm.n1024 0.228786
R29701 C10_P_btm.n1027 C10_P_btm.n50 0.228786
R29702 C10_P_btm.n1026 C10_P_btm.n49 0.228786
R29703 C10_P_btm.n1029 C10_P_btm.n1028 0.228786
R29704 C10_P_btm.n1031 C10_P_btm.n48 0.228786
R29705 C10_P_btm.n1030 C10_P_btm.n45 0.228786
R29706 C10_P_btm.n1033 C10_P_btm.n1032 0.228786
R29707 C10_P_btm.n1035 C10_P_btm.n42 0.228786
R29708 C10_P_btm.n1034 C10_P_btm.n41 0.228786
R29709 C10_P_btm.n1037 C10_P_btm.n1036 0.228786
R29710 C10_P_btm.n1039 C10_P_btm.n40 0.228786
R29711 C10_P_btm.n1038 C10_P_btm.n37 0.228786
R29712 C10_P_btm.n1041 C10_P_btm.n1040 0.228786
R29713 C10_P_btm.n1043 C10_P_btm.n34 0.228786
R29714 C10_P_btm.n1042 C10_P_btm.n33 0.228786
R29715 C10_P_btm.n684 C10_P_btm.n471 0.228786
R29716 C10_P_btm.n269 C10_P_btm.n268 0.228786
R29717 C10_P_btm.n267 C10_P_btm.n266 0.228786
R29718 C10_P_btm.n265 C10_P_btm.n175 0.228786
R29719 C10_P_btm.n193 C10_P_btm.n176 0.228786
R29720 C10_P_btm.n262 C10_P_btm.n177 0.228786
R29721 C10_P_btm.n179 C10_P_btm.n178 0.228786
R29722 C10_P_btm.n260 C10_P_btm.n259 0.228786
R29723 C10_P_btm.n196 C10_P_btm.n180 0.228786
R29724 C10_P_btm.n198 C10_P_btm.n195 0.228786
R29725 C10_P_btm.n194 C10_P_btm.n192 0.228786
R29726 C10_P_btm.n173 C10_P_btm.n172 0.228786
R29727 C10_P_btm.n270 C10_P_btm.n269 0.228786
R29728 C10_P_btm.n271 C10_P_btm.n270 0.228786
R29729 C10_P_btm.n170 C10_P_btm.n169 0.228786
R29730 C10_P_btm.n272 C10_P_btm.n170 0.228786
R29731 C10_P_btm.n274 C10_P_btm.n273 0.228786
R29732 C10_P_btm.n272 C10_P_btm.n271 0.228786
R29733 C10_P_btm.n275 C10_P_btm.n168 0.228786
R29734 C10_P_btm.n200 C10_P_btm.n167 0.228786
R29735 C10_P_btm.n249 C10_P_btm.n201 0.228786
R29736 C10_P_btm.n252 C10_P_btm.n188 0.228786
R29737 C10_P_btm.n257 C10_P_btm.n254 0.228786
R29738 C10_P_btm.n256 C10_P_btm.n187 0.228786
R29739 C10_P_btm.n183 C10_P_btm.n182 0.228786
R29740 C10_P_btm.n80 C10_P_btm.n79 0.228786
R29741 C10_P_btm.n354 C10_P_btm.n353 0.228786
R29742 C10_P_btm.n77 C10_P_btm.n76 0.228786
R29743 C10_P_btm.n1005 C10_P_btm.n1004 0.228786
R29744 C10_P_btm.n1003 C10_P_btm.n75 0.228786
R29745 C10_P_btm.n979 C10_P_btm.n358 0.228786
R29746 C10_P_btm.n980 C10_P_btm.n359 0.228786
R29747 C10_P_btm.n998 C10_P_btm.n361 0.228786
R29748 C10_P_btm.n997 C10_P_btm.n996 0.228786
R29749 C10_P_btm.n363 C10_P_btm.n362 0.228786
R29750 C10_P_btm.n388 C10_P_btm.n387 0.228786
R29751 C10_P_btm.n391 C10_P_btm.n384 0.228786
R29752 C10_P_btm.n394 C10_P_btm.n393 0.228786
R29753 C10_P_btm.n395 C10_P_btm.n382 0.228786
R29754 C10_P_btm.n957 C10_P_btm.n956 0.228786
R29755 C10_P_btm.n955 C10_P_btm.n381 0.228786
R29756 C10_P_btm.n954 C10_P_btm.n396 0.228786
R29757 C10_P_btm.n953 C10_P_btm.n397 0.228786
R29758 C10_P_btm.n952 C10_P_btm.n398 0.228786
R29759 C10_P_btm.n951 C10_P_btm.n399 0.228786
R29760 C10_P_btm.n950 C10_P_btm.n400 0.228786
R29761 C10_P_btm.n949 C10_P_btm.n401 0.228786
R29762 C10_P_btm.n948 C10_P_btm.n402 0.228786
R29763 C10_P_btm.n947 C10_P_btm.n403 0.228786
R29764 C10_P_btm.n946 C10_P_btm.n404 0.228786
R29765 C10_P_btm.n880 C10_P_btm.n426 0.228786
R29766 C10_P_btm.n421 C10_P_btm.n420 0.228786
R29767 C10_P_btm.n423 C10_P_btm.n422 0.228786
R29768 C10_P_btm.n407 C10_P_btm.n406 0.228786
R29769 C10_P_btm.n943 C10_P_btm.n942 0.228786
R29770 C10_P_btm.n409 C10_P_btm.n408 0.228786
R29771 C10_P_btm.n927 C10_P_btm.n926 0.228786
R29772 C10_P_btm.n929 C10_P_btm.n928 0.228786
R29773 C10_P_btm.n930 C10_P_btm.n923 0.228786
R29774 C10_P_btm.n922 C10_P_btm.n895 0.228786
R29775 C10_P_btm.n921 C10_P_btm.n920 0.228786
R29776 C10_P_btm.n897 C10_P_btm.n896 0.228786
R29777 C10_P_btm.n906 C10_P_btm.n905 0.228786
R29778 C10_P_btm.n904 C10_P_btm.n903 0.228786
R29779 C10_P_btm.n380 C10_P_btm.n379 0.228786
R29780 C10_P_btm.n959 C10_P_btm.n958 0.228786
R29781 C10_P_btm.n960 C10_P_btm.n378 0.228786
R29782 C10_P_btm.n962 C10_P_btm.n376 0.228786
R29783 C10_P_btm.n390 C10_P_btm.n375 0.228786
R29784 C10_P_btm.n389 C10_P_btm.n368 0.228786
R29785 C10_P_btm.n993 C10_P_btm.n364 0.228786
R29786 C10_P_btm.n995 C10_P_btm.n994 0.228786
R29787 C10_P_btm.n366 C10_P_btm.n365 0.228786
R29788 C10_P_btm.n982 C10_P_btm.n981 0.228786
R29789 C10_P_btm.n978 C10_P_btm.n977 0.228786
R29790 C10_P_btm.n74 C10_P_btm.n73 0.228786
R29791 C10_P_btm.n1007 C10_P_btm.n1006 0.228786
R29792 C10_P_btm.n1008 C10_P_btm.n72 0.228786
R29793 C10_P_btm.n352 C10_P_btm.n71 0.228786
R29794 C10_P_btm.n351 C10_P_btm.n350 0.228786
R29795 C10_P_btm.n348 C10_P_btm.n82 0.228786
R29796 C10_P_btm.n84 C10_P_btm.n83 0.228786
R29797 C10_P_btm.n253 C10_P_btm.n189 0.228786
R29798 C10_P_btm.n251 C10_P_btm.n250 0.228786
R29799 C10_P_btm.n344 C10_P_btm.n87 0.228786
R29800 C10_P_btm.n343 C10_P_btm.n342 0.228786
R29801 C10_P_btm.n89 C10_P_btm.n88 0.228786
R29802 C10_P_btm.n248 C10_P_btm.n247 0.228786
R29803 C10_P_btm.n166 C10_P_btm.n165 0.228786
R29804 C10_P_btm.n277 C10_P_btm.n276 0.228786
R29805 C10_P_btm.n278 C10_P_btm.n164 0.228786
R29806 C10_P_btm.n169 C10_P_btm.n163 0.228786
R29807 C10_P_btm.n163 C10_P_btm.n162 0.228786
R29808 C10_P_btm.n161 C10_P_btm.n160 0.228786
R29809 C10_P_btm.n162 C10_P_btm.n161 0.228786
R29810 C10_P_btm.n280 C10_P_btm.n279 0.228786
R29811 C10_P_btm.n281 C10_P_btm.n159 0.228786
R29812 C10_P_btm.n202 C10_P_btm.n158 0.228786
R29813 C10_P_btm.n246 C10_P_btm.n245 0.228786
R29814 C10_P_btm.n203 C10_P_btm.n90 0.228786
R29815 C10_P_btm.n93 C10_P_btm.n92 0.228786
R29816 C10_P_btm.n205 C10_P_btm.n204 0.228786
R29817 C10_P_btm.n244 C10_P_btm.n243 0.228786
R29818 C10_P_btm.n157 C10_P_btm.n156 0.228786
R29819 C10_P_btm.n283 C10_P_btm.n282 0.228786
R29820 C10_P_btm.n284 C10_P_btm.n155 0.228786
R29821 C10_P_btm.n160 C10_P_btm.n154 0.228786
R29822 C10_P_btm.n154 C10_P_btm.n153 0.228786
R29823 C10_P_btm.n152 C10_P_btm.n151 0.228786
R29824 C10_P_btm.n153 C10_P_btm.n152 0.228786
R29825 C10_P_btm.n286 C10_P_btm.n285 0.228786
R29826 C10_P_btm.n287 C10_P_btm.n150 0.228786
R29827 C10_P_btm.n206 C10_P_btm.n149 0.228786
R29828 C10_P_btm.n242 C10_P_btm.n207 0.228786
R29829 C10_P_btm.n241 C10_P_btm.n240 0.228786
R29830 C10_P_btm.n97 C10_P_btm.n96 0.228786
R29831 C10_P_btm.n239 C10_P_btm.n208 0.228786
R29832 C10_P_btm.n238 C10_P_btm.n237 0.228786
R29833 C10_P_btm.n148 C10_P_btm.n147 0.228786
R29834 C10_P_btm.n289 C10_P_btm.n288 0.228786
R29835 C10_P_btm.n290 C10_P_btm.n146 0.228786
R29836 C10_P_btm.n151 C10_P_btm.n145 0.228786
R29837 C10_P_btm.n145 C10_P_btm.n142 0.228786
R29838 C10_P_btm.n294 C10_P_btm.n293 0.228786
R29839 C10_P_btm.n293 C10_P_btm.n142 0.228786
R29840 C10_P_btm.n292 C10_P_btm.n291 0.228786
R29841 C10_P_btm.n144 C10_P_btm.n143 0.228786
R29842 C10_P_btm.n212 C10_P_btm.n209 0.228786
R29843 C10_P_btm.n236 C10_P_btm.n210 0.228786
R29844 C10_P_btm.n235 C10_P_btm.n234 0.228786
R29845 C10_P_btm.n101 C10_P_btm.n100 0.228786
R29846 C10_P_btm.n233 C10_P_btm.n211 0.228786
R29847 C10_P_btm.n232 C10_P_btm.n231 0.228786
R29848 C10_P_btm.n214 C10_P_btm.n213 0.228786
R29849 C10_P_btm.n216 C10_P_btm.n215 0.228786
R29850 C10_P_btm.n141 C10_P_btm.n140 0.228786
R29851 C10_P_btm.n295 C10_P_btm.n294 0.228786
R29852 C10_P_btm.n296 C10_P_btm.n295 0.228786
R29853 C10_P_btm.n138 C10_P_btm.n137 0.228786
R29854 C10_P_btm.n297 C10_P_btm.n138 0.228786
R29855 C10_P_btm.n299 C10_P_btm.n298 0.228786
R29856 C10_P_btm.n297 C10_P_btm.n296 0.228786
R29857 C10_P_btm.n217 C10_P_btm.n125 0.228786
R29858 C10_P_btm.n219 C10_P_btm.n218 0.228786
R29859 C10_P_btm.n230 C10_P_btm.n220 0.228786
R29860 C10_P_btm.n229 C10_P_btm.n228 0.228786
R29861 C10_P_btm.n105 C10_P_btm.n104 0.228786
R29862 C10_P_btm.n227 C10_P_btm.n226 0.228786
R29863 C10_P_btm.n222 C10_P_btm.n221 0.228786
R29864 C10_P_btm.n124 C10_P_btm.n122 0.228786
R29865 C10_P_btm.n302 C10_P_btm.n301 0.228786
R29866 C10_P_btm.n123 C10_P_btm.n121 0.228786
R29867 C10_P_btm.n137 C10_P_btm.n136 0.228786
R29868 C10_P_btm.n134 C10_P_btm.n126 0.228786
R29869 C10_P_btm.n135 C10_P_btm.n134 0.228786
R29870 C10_P_btm.n136 C10_P_btm.n135 0.228786
R29871 C10_P_btm.n133 C10_P_btm.n120 0.228786
R29872 C10_P_btm.n305 C10_P_btm.n304 0.228786
R29873 C10_P_btm.n303 C10_P_btm.n118 0.228786
R29874 C10_P_btm.n223 C10_P_btm.n117 0.228786
R29875 C10_P_btm.n225 C10_P_btm.n224 0.228786
R29876 C10_P_btm.n109 C10_P_btm.n108 0.228786
R29877 C10_P_btm.n116 C10_P_btm.n114 0.228786
R29878 C10_P_btm.n308 C10_P_btm.n307 0.228786
R29879 C10_P_btm.n115 C10_P_btm.n113 0.228786
R29880 C10_P_btm.n128 C10_P_btm.n127 0.228786
R29881 C10_P_btm.n132 C10_P_btm.n131 0.228786
R29882 C10_P_btm.n66 C10_P_btm.n64 0.228786
R29883 C10_P_btm.n1012 C10_P_btm.n1011 0.228786
R29884 C10_P_btm.n1010 C10_P_btm.n1009 0.228786
R29885 C10_P_btm.n70 C10_P_btm.n69 0.228786
R29886 C10_P_btm.n975 C10_P_btm.n974 0.228786
R29887 C10_P_btm.n976 C10_P_btm.n970 0.228786
R29888 C10_P_btm.n984 C10_P_btm.n983 0.228786
R29889 C10_P_btm.n985 C10_P_btm.n969 0.228786
R29890 C10_P_btm.n967 C10_P_btm.n367 0.228786
R29891 C10_P_btm.n992 C10_P_btm.n369 0.228786
R29892 C10_P_btm.n991 C10_P_btm.n990 0.228786
R29893 C10_P_btm.n371 C10_P_btm.n370 0.228786
R29894 C10_P_btm.n374 C10_P_btm.n373 0.228786
R29895 C10_P_btm.n964 C10_P_btm.n963 0.228786
R29896 C10_P_btm.n910 C10_P_btm.n909 0.228786
R29897 C10_P_btm.n912 C10_P_btm.n911 0.228786
R29898 C10_P_btm.n913 C10_P_btm.n908 0.228786
R29899 C10_P_btm.n907 C10_P_btm.n901 0.228786
R29900 C10_P_btm.n899 C10_P_btm.n898 0.228786
R29901 C10_P_btm.n919 C10_P_btm.n918 0.228786
R29902 C10_P_btm.n894 C10_P_btm.n893 0.228786
R29903 C10_P_btm.n932 C10_P_btm.n931 0.228786
R29904 C10_P_btm.n933 C10_P_btm.n892 0.228786
R29905 C10_P_btm.n925 C10_P_btm.n890 0.228786
R29906 C10_P_btm.n924 C10_P_btm.n889 0.228786
R29907 C10_P_btm.n940 C10_P_btm.n939 0.228786
R29908 C10_P_btm.n938 C10_P_btm.n410 0.228786
R29909 C10_P_btm.n413 C10_P_btm.n412 0.228786
R29910 C10_P_btm.n885 C10_P_btm.n884 0.228786
R29911 C10_P_btm.n883 C10_P_btm.n415 0.228786
R29912 C10_P_btm.n419 C10_P_btm.n418 0.228786
R29913 C10_P_btm.n855 C10_P_btm.n427 0.228786
R29914 C10_P_btm.n856 C10_P_btm.n428 0.228786
R29915 C10_P_btm.n874 C10_P_btm.n430 0.228786
R29916 C10_P_btm.n873 C10_P_btm.n872 0.228786
R29917 C10_P_btm.n432 C10_P_btm.n431 0.228786
R29918 C10_P_btm.n454 C10_P_btm.n453 0.228786
R29919 C10_P_btm.n458 C10_P_btm.n457 0.228786
R29920 C10_P_btm.n450 C10_P_btm.n449 0.228786
R29921 C10_P_btm.n838 C10_P_btm.n837 0.228786
R29922 C10_P_btm.n836 C10_P_btm.n835 0.228786
R29923 C10_P_btm.n834 C10_P_btm.n462 0.228786
R29924 C10_P_btm.n464 C10_P_btm.n463 0.228786
R29925 C10_P_btm.n831 C10_P_btm.n465 0.228786
R29926 C10_P_btm.n830 C10_P_btm.n829 0.228786
R29927 C10_P_btm.n447 C10_P_btm.n446 0.228786
R29928 C10_P_btm.n840 C10_P_btm.n839 0.228786
R29929 C10_P_btm.n841 C10_P_btm.n445 0.228786
R29930 C10_P_btm.n456 C10_P_btm.n444 0.228786
R29931 C10_P_btm.n455 C10_P_btm.n437 0.228786
R29932 C10_P_btm.n869 C10_P_btm.n433 0.228786
R29933 C10_P_btm.n871 C10_P_btm.n870 0.228786
R29934 C10_P_btm.n435 C10_P_btm.n434 0.228786
R29935 C10_P_btm.n858 C10_P_btm.n857 0.228786
R29936 C10_P_btm.n854 C10_P_btm.n853 0.228786
R29937 C10_P_btm.n849 C10_P_btm.n417 0.228786
R29938 C10_P_btm.n852 C10_P_btm.n851 0.228786
R29939 C10_P_btm.n860 C10_P_btm.n859 0.228786
R29940 C10_P_btm.n861 C10_P_btm.n848 0.228786
R29941 C10_P_btm.n846 C10_P_btm.n436 0.228786
R29942 C10_P_btm.n868 C10_P_btm.n438 0.228786
R29943 C10_P_btm.n867 C10_P_btm.n866 0.228786
R29944 C10_P_btm.n440 C10_P_btm.n439 0.228786
R29945 C10_P_btm.n843 C10_P_btm.n842 0.228786
R29946 C10_P_btm.n443 C10_P_btm.n442 0.228786
R29947 C10_P_btm.n827 C10_P_btm.n469 0.228786
R29948 C10_P_btm.n826 C10_P_btm.n825 0.228786
R29949 C10_P_btm.n821 C10_P_btm.n468 0.228786
R29950 C10_P_btm.n820 C10_P_btm.n819 0.228786
R29951 C10_P_btm.n480 C10_P_btm.n479 0.228786
R29952 C10_P_btm.n811 C10_P_btm.n810 0.228786
R29953 C10_P_btm.n478 C10_P_btm.n477 0.228786
R29954 C10_P_btm.n809 C10_P_btm.n481 0.228786
R29955 C10_P_btm.n475 C10_P_btm.n474 0.228786
R29956 C10_P_btm.n722 C10_P_btm.n721 0.228786
R29957 C10_P_btm.n685 C10_P_btm.n473 0.228786
R29958 C10_P_btm.n724 C10_P_btm.n723 0.228786
R29959 C10_P_btm.n726 C10_P_btm.n725 0.228786
R29960 C10_P_btm.n683 C10_P_btm.n682 0.228786
R29961 C10_P_btm.n710 C10_P_btm.n690 0.228786
R29962 C10_P_btm.n714 C10_P_btm.n713 0.228786
R29963 C10_P_btm.n502 C10_P_btm.n501 0.228786
R29964 C10_P_btm.n505 C10_P_btm.n503 0.228786
R29965 C10_P_btm.n509 C10_P_btm.n508 0.228786
R29966 C10_P_btm.n511 C10_P_btm.n510 0.228786
R29967 C10_P_btm.n804 C10_P_btm.n484 0.228786
R29968 C10_P_btm.n802 C10_P_btm.n486 0.228786
R29969 C10_P_btm.n803 C10_P_btm.n487 0.228786
R29970 C10_P_btm.n801 C10_P_btm.n489 0.228786
R29971 C10_P_btm.n689 C10_P_btm.n687 0.228786
R29972 C10_P_btm.n706 C10_P_btm.n705 0.228786
R29973 C10_P_btm.n704 C10_P_btm.n692 0.228786
R29974 C10_P_btm.n708 C10_P_btm.n707 0.228786
R29975 C10_P_btm.n709 C10_P_btm.n691 0.228786
R29976 C10_P_btm.n699 C10_P_btm.n694 0.228786
R29977 C10_P_btm.n535 C10_P_btm.n534 0.228786
R29978 C10_P_btm.n697 C10_P_btm.n696 0.228786
R29979 C10_P_btm.n500 C10_P_btm.n499 0.228786
R29980 C10_P_btm.n520 C10_P_btm.n519 0.228786
R29981 C10_P_btm.n522 C10_P_btm.n521 0.228786
R29982 C10_P_btm.n496 C10_P_btm.n494 0.228786
R29983 C10_P_btm.n524 C10_P_btm.n523 0.228786
R29984 C10_P_btm.n526 C10_P_btm.n525 0.228786
R29985 C10_P_btm.n796 C10_P_btm.n492 0.228786
R29986 C10_P_btm.n794 C10_P_btm.n527 0.228786
R29987 C10_P_btm.n795 C10_P_btm.n528 0.228786
R29988 C10_P_btm.n793 C10_P_btm.n792 0.228786
R29989 C10_P_btm.n790 C10_P_btm.n529 0.228786
R29990 C10_P_btm.n791 C10_P_btm.n530 0.228786
R29991 C10_P_btm.n789 C10_P_btm.n788 0.228786
R29992 C10_P_btm.n786 C10_P_btm.n533 0.228786
R29993 C10_P_btm.n787 C10_P_btm.n536 0.228786
R29994 C10_P_btm.n728 C10_P_btm.n681 0.228786
R29995 C10_P_btm.n729 C10_P_btm.n728 0.228786
R29996 C10_P_btm.n730 C10_P_btm.n729 0.228786
R29997 C10_P_btm.n732 C10_P_btm.n731 0.228786
R29998 C10_P_btm.n730 C10_P_btm.n679 0.228786
R29999 C10_P_btm.n679 C10_P_btm.n678 0.228786
R30000 C10_P_btm.n737 C10_P_btm.n736 0.228786
R30001 C10_P_btm.n735 C10_P_btm.n598 0.228786
R30002 C10_P_btm.n734 C10_P_btm.n602 0.228786
R30003 C10_P_btm.n604 C10_P_btm.n601 0.228786
R30004 C10_P_btm.n678 C10_P_btm.n677 0.228786
R30005 C10_P_btm.n677 C10_P_btm.n676 0.228786
R30006 C10_P_btm.n672 C10_P_btm.n605 0.228786
R30007 C10_P_btm.n676 C10_P_btm.n605 0.228786
R30008 C10_P_btm.n675 C10_P_btm.n674 0.228786
R30009 C10_P_btm.n607 C10_P_btm.n606 0.228786
R30010 C10_P_btm.n634 C10_P_btm.n633 0.228786
R30011 C10_P_btm.n739 C10_P_btm.n738 0.228786
R30012 C10_P_btm.n595 C10_P_btm.n594 0.228786
R30013 C10_P_btm.n539 C10_P_btm.n538 0.228786
R30014 C10_P_btm.n590 C10_P_btm.n589 0.228786
R30015 C10_P_btm.n743 C10_P_btm.n742 0.228786
R30016 C10_P_btm.n744 C10_P_btm.n587 0.228786
R30017 C10_P_btm.n632 C10_P_btm.n586 0.228786
R30018 C10_P_btm.n636 C10_P_btm.n635 0.228786
R30019 C10_P_btm.n631 C10_P_btm.n608 0.228786
R30020 C10_P_btm.n673 C10_P_btm.n609 0.228786
R30021 C10_P_btm.n672 C10_P_btm.n671 0.228786
R30022 C10_P_btm.n671 C10_P_btm.n670 0.228786
R30023 C10_P_btm.n666 C10_P_btm.n610 0.228786
R30024 C10_P_btm.n670 C10_P_btm.n610 0.228786
R30025 C10_P_btm.n669 C10_P_btm.n668 0.228786
R30026 C10_P_btm.n612 C10_P_btm.n611 0.228786
R30027 C10_P_btm.n638 C10_P_btm.n637 0.228786
R30028 C10_P_btm.n585 C10_P_btm.n584 0.228786
R30029 C10_P_btm.n746 C10_P_btm.n745 0.228786
R30030 C10_P_btm.n747 C10_P_btm.n583 0.228786
R30031 C10_P_btm.n588 C10_P_btm.n582 0.228786
R30032 C10_P_btm.n580 C10_P_btm.n579 0.228786
R30033 C10_P_btm.n581 C10_P_btm.n578 0.228786
R30034 C10_P_btm.n749 C10_P_btm.n748 0.228786
R30035 C10_P_btm.n750 C10_P_btm.n576 0.228786
R30036 C10_P_btm.n630 C10_P_btm.n575 0.228786
R30037 C10_P_btm.n640 C10_P_btm.n639 0.228786
R30038 C10_P_btm.n629 C10_P_btm.n613 0.228786
R30039 C10_P_btm.n667 C10_P_btm.n614 0.228786
R30040 C10_P_btm.n666 C10_P_btm.n665 0.228786
R30041 C10_P_btm.n665 C10_P_btm.n664 0.228786
R30042 C10_P_btm.n660 C10_P_btm.n615 0.228786
R30043 C10_P_btm.n664 C10_P_btm.n615 0.228786
R30044 C10_P_btm.n663 C10_P_btm.n662 0.228786
R30045 C10_P_btm.n617 C10_P_btm.n616 0.228786
R30046 C10_P_btm.n642 C10_P_btm.n641 0.228786
R30047 C10_P_btm.n574 C10_P_btm.n573 0.228786
R30048 C10_P_btm.n752 C10_P_btm.n751 0.228786
R30049 C10_P_btm.n753 C10_P_btm.n572 0.228786
R30050 C10_P_btm.n577 C10_P_btm.n571 0.228786
R30051 C10_P_btm.n550 C10_P_btm.n549 0.228786
R30052 C10_P_btm.n570 C10_P_btm.n569 0.228786
R30053 C10_P_btm.n755 C10_P_btm.n754 0.228786
R30054 C10_P_btm.n756 C10_P_btm.n565 0.228786
R30055 C10_P_btm.n628 C10_P_btm.n564 0.228786
R30056 C10_P_btm.n644 C10_P_btm.n643 0.228786
R30057 C10_P_btm.n627 C10_P_btm.n618 0.228786
R30058 C10_P_btm.n661 C10_P_btm.n619 0.228786
R30059 C10_P_btm.n660 C10_P_btm.n659 0.228786
R30060 C10_P_btm.n659 C10_P_btm.n658 0.228786
R30061 C10_P_btm.n654 C10_P_btm.n620 0.228786
R30062 C10_P_btm.n658 C10_P_btm.n620 0.228786
R30063 C10_P_btm.n657 C10_P_btm.n656 0.228786
R30064 C10_P_btm.n622 C10_P_btm.n621 0.228786
R30065 C10_P_btm.n646 C10_P_btm.n645 0.228786
R30066 C10_P_btm.n563 C10_P_btm.n562 0.228786
R30067 C10_P_btm.n758 C10_P_btm.n757 0.228786
R30068 C10_P_btm.n759 C10_P_btm.n561 0.228786
R30069 C10_P_btm.n568 C10_P_btm.n560 0.228786
R30070 C10_P_btm.n765 C10_P_btm.n554 0.228786
R30071 C10_P_btm.n558 C10_P_btm.n555 0.228786
R30072 C10_P_btm.n761 C10_P_btm.n760 0.228786
R30073 C10_P_btm.n559 C10_P_btm.n557 0.228786
R30074 C10_P_btm.n649 C10_P_btm.n648 0.228786
R30075 C10_P_btm.n650 C10_P_btm.n647 0.228786
R30076 C10_P_btm.n625 C10_P_btm.n623 0.228786
R30077 C10_P_btm.n655 C10_P_btm.n624 0.228786
R30078 C10_P_btm.n684 C10_P_btm.n681 0.228786
R30079 C10_P_btm.n1014 C10_P_btm.n1013 0.228786
R30080 C10_P_btm.n1016 C10_P_btm.n1015 0.228786
R30081 C10_P_btm.n61 C10_P_btm.n58 0.228786
R30082 C10_P_btm.n1018 C10_P_btm.n1017 0.228786
R30083 C10_P_btm.n1020 C10_P_btm.n1019 0.228786
R30084 C10_P_btm.n57 C10_P_btm.n56 0.228786
R30085 C10_P_btm.n1022 C10_P_btm.n1021 0.228786
R30086 C10_P_btm.n1024 C10_P_btm.n1023 0.228786
R30087 C10_P_btm.n53 C10_P_btm.n50 0.228786
R30088 C10_P_btm.n1026 C10_P_btm.n1025 0.228786
R30089 C10_P_btm.n1028 C10_P_btm.n1027 0.228786
R30090 C10_P_btm.n49 C10_P_btm.n48 0.228786
R30091 C10_P_btm.n1030 C10_P_btm.n1029 0.228786
R30092 C10_P_btm.n1032 C10_P_btm.n1031 0.228786
R30093 C10_P_btm.n45 C10_P_btm.n42 0.228786
R30094 C10_P_btm.n1034 C10_P_btm.n1033 0.228786
R30095 C10_P_btm.n1036 C10_P_btm.n1035 0.228786
R30096 C10_P_btm.n41 C10_P_btm.n40 0.228786
R30097 C10_P_btm.n1038 C10_P_btm.n1037 0.228786
R30098 C10_P_btm.n1040 C10_P_btm.n1039 0.228786
R30099 C10_P_btm.n37 C10_P_btm.n34 0.228786
R30100 C10_P_btm.n1042 C10_P_btm.n1041 0.228786
R30101 C10_P_btm.n1044 C10_P_btm.n1043 0.228786
R30102 C10_P_btm.n764 C10_P_btm.n553 0.208893
R30103 C10_P_btm.n965 C10_P_btm.n372 0.208893
R30104 C10_P_btm.n130 C10_P_btm.n129 0.208893
R30105 C10_P_btm.n518 C10_P_btm.n517 0.208893
R30106 C10_P_btm.n653 C10_P_btm.n652 0.208893
R30107 C10_P_btm.n862 C10_P_btm.n847 0.208893
R30108 C10_P_btm.n264 C10_P_btm.n174 0.208893
R30109 C10_P_btm.n787 C10_P_btm.n535 0.09425
R30110 C10_P_btm.n696 C10_P_btm.n534 0.09425
R30111 C10_P_btm.n699 C10_P_btm.n691 0.09425
R30112 C10_P_btm.n710 C10_P_btm.n709 0.09425
R30113 C10_P_btm.n713 C10_P_btm.n690 0.09425
R30114 C10_P_btm.n726 C10_P_btm.n683 0.09425
R30115 C10_P_btm.n725 C10_P_btm.n684 0.09425
R30116 C10_P_btm.n820 C10_P_btm.n471 0.09425
R30117 C10_P_btm.n852 C10_P_btm.n849 0.09425
R30118 C10_P_btm.n346 C10_P_btm.n66 0.09425
R30119 C10_P_btm.n233 C10_P_btm.n100 0.09425
R30120 C10_P_btm.n329 C10_P_btm.n99 0.09425
R30121 C10_P_btm.n239 C10_P_btm.n96 0.09425
R30122 C10_P_btm.n333 C10_P_btm.n95 0.09425
R30123 C10_P_btm.n204 C10_P_btm.n92 0.09425
R30124 C10_P_btm.n339 C10_P_btm.n91 0.09425
R30125 C10_P_btm.n196 C10_P_btm.n195 0.09425
R30126 C10_P_btm.n259 C10_P_btm.n180 0.09425
R30127 C10_P_btm.n260 C10_P_btm.n179 0.09425
R30128 C10_P_btm.n265 C10_P_btm.n176 0.09425
R30129 C10_P_btm.n266 C10_P_btm.n265 0.09425
R30130 C10_P_btm.n264 C10_P_btm.n263 0.09425
R30131 C10_P_btm.n263 C10_P_btm.n262 0.09425
R30132 C10_P_btm.n185 C10_P_btm.n178 0.09425
R30133 C10_P_btm.n261 C10_P_btm.n178 0.09425
R30134 C10_P_btm.n262 C10_P_btm.n261 0.09425
R30135 C10_P_btm.n260 C10_P_btm.n177 0.09425
R30136 C10_P_btm.n177 C10_P_btm.n176 0.09425
R30137 C10_P_btm.n193 C10_P_btm.n180 0.09425
R30138 C10_P_btm.n193 C10_P_btm.n175 0.09425
R30139 C10_P_btm.n195 C10_P_btm.n194 0.09425
R30140 C10_P_btm.n194 C10_P_btm.n173 0.09425
R30141 C10_P_btm.n267 C10_P_btm.n175 0.09425
R30142 C10_P_btm.n268 C10_P_btm.n267 0.09425
R30143 C10_P_btm.n269 C10_P_btm.n173 0.09425
R30144 C10_P_btm.n270 C10_P_btm.n172 0.09425
R30145 C10_P_btm.n273 C10_P_btm.n168 0.09425
R30146 C10_P_btm.n273 C10_P_btm.n272 0.09425
R30147 C10_P_btm.n191 C10_P_btm.n171 0.09425
R30148 C10_P_btm.n271 C10_P_btm.n171 0.09425
R30149 C10_P_btm.n198 C10_P_btm.n192 0.09425
R30150 C10_P_btm.n192 C10_P_btm.n172 0.09425
R30151 C10_P_btm.n200 C10_P_btm.n168 0.09425
R30152 C10_P_btm.n251 C10_P_btm.n201 0.09425
R30153 C10_P_btm.n201 C10_P_btm.n200 0.09425
R30154 C10_P_btm.n199 C10_P_btm.n190 0.09425
R30155 C10_P_btm.n199 C10_P_btm.n191 0.09425
R30156 C10_P_btm.n197 C10_P_btm.n188 0.09425
R30157 C10_P_btm.n198 C10_P_btm.n197 0.09425
R30158 C10_P_btm.n257 C10_P_btm.n181 0.09425
R30159 C10_P_btm.n196 C10_P_btm.n181 0.09425
R30160 C10_P_btm.n258 C10_P_btm.n187 0.09425
R30161 C10_P_btm.n259 C10_P_btm.n258 0.09425
R30162 C10_P_btm.n186 C10_P_btm.n183 0.09425
R30163 C10_P_btm.n186 C10_P_btm.n179 0.09425
R30164 C10_P_btm.n184 C10_P_btm.n78 0.09425
R30165 C10_P_btm.n185 C10_P_btm.n184 0.09425
R30166 C10_P_btm.n354 C10_P_btm.n79 0.09425
R30167 C10_P_btm.n183 C10_P_btm.n79 0.09425
R30168 C10_P_btm.n356 C10_P_btm.n355 0.09425
R30169 C10_P_btm.n355 C10_P_btm.n78 0.09425
R30170 C10_P_btm.n1004 C10_P_btm.n77 0.09425
R30171 C10_P_btm.n354 C10_P_btm.n77 0.09425
R30172 C10_P_btm.n1002 C10_P_btm.n357 0.09425
R30173 C10_P_btm.n357 C10_P_btm.n356 0.09425
R30174 C10_P_btm.n1003 C10_P_btm.n358 0.09425
R30175 C10_P_btm.n1004 C10_P_btm.n1003 0.09425
R30176 C10_P_btm.n1001 C10_P_btm.n1000 0.09425
R30177 C10_P_btm.n1002 C10_P_btm.n1001 0.09425
R30178 C10_P_btm.n998 C10_P_btm.n359 0.09425
R30179 C10_P_btm.n359 C10_P_btm.n358 0.09425
R30180 C10_P_btm.n999 C10_P_btm.n360 0.09425
R30181 C10_P_btm.n1000 C10_P_btm.n999 0.09425
R30182 C10_P_btm.n997 C10_P_btm.n362 0.09425
R30183 C10_P_btm.n998 C10_P_btm.n997 0.09425
R30184 C10_P_btm.n386 C10_P_btm.n385 0.09425
R30185 C10_P_btm.n385 C10_P_btm.n360 0.09425
R30186 C10_P_btm.n387 C10_P_btm.n384 0.09425
R30187 C10_P_btm.n387 C10_P_btm.n362 0.09425
R30188 C10_P_btm.n386 C10_P_btm.n383 0.09425
R30189 C10_P_btm.n394 C10_P_btm.n383 0.09425
R30190 C10_P_btm.n395 C10_P_btm.n394 0.09425
R30191 C10_P_btm.n956 C10_P_btm.n395 0.09425
R30192 C10_P_btm.n956 C10_P_btm.n955 0.09425
R30193 C10_P_btm.n955 C10_P_btm.n954 0.09425
R30194 C10_P_btm.n954 C10_P_btm.n953 0.09425
R30195 C10_P_btm.n953 C10_P_btm.n952 0.09425
R30196 C10_P_btm.n952 C10_P_btm.n951 0.09425
R30197 C10_P_btm.n951 C10_P_btm.n950 0.09425
R30198 C10_P_btm.n950 C10_P_btm.n949 0.09425
R30199 C10_P_btm.n949 C10_P_btm.n948 0.09425
R30200 C10_P_btm.n948 C10_P_btm.n947 0.09425
R30201 C10_P_btm.n947 C10_P_btm.n946 0.09425
R30202 C10_P_btm.n878 C10_P_btm.n426 0.09425
R30203 C10_P_btm.n426 C10_P_btm.n425 0.09425
R30204 C10_P_btm.n880 C10_P_btm.n421 0.09425
R30205 C10_P_btm.n423 C10_P_btm.n421 0.09425
R30206 C10_P_btm.n425 C10_P_btm.n424 0.09425
R30207 C10_P_btm.n424 C10_P_btm.n405 0.09425
R30208 C10_P_btm.n423 C10_P_btm.n406 0.09425
R30209 C10_P_btm.n944 C10_P_btm.n406 0.09425
R30210 C10_P_btm.n945 C10_P_btm.n405 0.09425
R30211 C10_P_btm.n946 C10_P_btm.n945 0.09425
R30212 C10_P_btm.n943 C10_P_btm.n407 0.09425
R30213 C10_P_btm.n943 C10_P_btm.n408 0.09425
R30214 C10_P_btm.n944 C10_P_btm.n404 0.09425
R30215 C10_P_btm.n404 C10_P_btm.n403 0.09425
R30216 C10_P_btm.n927 C10_P_btm.n408 0.09425
R30217 C10_P_btm.n928 C10_P_btm.n927 0.09425
R30218 C10_P_btm.n403 C10_P_btm.n402 0.09425
R30219 C10_P_btm.n402 C10_P_btm.n401 0.09425
R30220 C10_P_btm.n928 C10_P_btm.n923 0.09425
R30221 C10_P_btm.n923 C10_P_btm.n922 0.09425
R30222 C10_P_btm.n401 C10_P_btm.n400 0.09425
R30223 C10_P_btm.n400 C10_P_btm.n399 0.09425
R30224 C10_P_btm.n922 C10_P_btm.n921 0.09425
R30225 C10_P_btm.n921 C10_P_btm.n896 0.09425
R30226 C10_P_btm.n399 C10_P_btm.n398 0.09425
R30227 C10_P_btm.n398 C10_P_btm.n397 0.09425
R30228 C10_P_btm.n905 C10_P_btm.n896 0.09425
R30229 C10_P_btm.n905 C10_P_btm.n904 0.09425
R30230 C10_P_btm.n397 C10_P_btm.n396 0.09425
R30231 C10_P_btm.n396 C10_P_btm.n381 0.09425
R30232 C10_P_btm.n904 C10_P_btm.n380 0.09425
R30233 C10_P_btm.n958 C10_P_btm.n380 0.09425
R30234 C10_P_btm.n957 C10_P_btm.n381 0.09425
R30235 C10_P_btm.n957 C10_P_btm.n382 0.09425
R30236 C10_P_btm.n958 C10_P_btm.n378 0.09425
R30237 C10_P_btm.n392 C10_P_btm.n378 0.09425
R30238 C10_P_btm.n393 C10_P_btm.n382 0.09425
R30239 C10_P_btm.n393 C10_P_btm.n384 0.09425
R30240 C10_P_btm.n960 C10_P_btm.n376 0.09425
R30241 C10_P_btm.n390 C10_P_btm.n376 0.09425
R30242 C10_P_btm.n392 C10_P_btm.n391 0.09425
R30243 C10_P_btm.n391 C10_P_btm.n388 0.09425
R30244 C10_P_btm.n390 C10_P_btm.n389 0.09425
R30245 C10_P_btm.n389 C10_P_btm.n364 0.09425
R30246 C10_P_btm.n388 C10_P_btm.n363 0.09425
R30247 C10_P_btm.n996 C10_P_btm.n363 0.09425
R30248 C10_P_btm.n995 C10_P_btm.n364 0.09425
R30249 C10_P_btm.n995 C10_P_btm.n365 0.09425
R30250 C10_P_btm.n996 C10_P_btm.n361 0.09425
R30251 C10_P_btm.n980 C10_P_btm.n361 0.09425
R30252 C10_P_btm.n981 C10_P_btm.n365 0.09425
R30253 C10_P_btm.n981 C10_P_btm.n978 0.09425
R30254 C10_P_btm.n980 C10_P_btm.n979 0.09425
R30255 C10_P_btm.n979 C10_P_btm.n75 0.09425
R30256 C10_P_btm.n978 C10_P_btm.n74 0.09425
R30257 C10_P_btm.n1006 C10_P_btm.n74 0.09425
R30258 C10_P_btm.n1005 C10_P_btm.n75 0.09425
R30259 C10_P_btm.n1005 C10_P_btm.n76 0.09425
R30260 C10_P_btm.n1006 C10_P_btm.n72 0.09425
R30261 C10_P_btm.n352 C10_P_btm.n72 0.09425
R30262 C10_P_btm.n353 C10_P_btm.n76 0.09425
R30263 C10_P_btm.n353 C10_P_btm.n80 0.09425
R30264 C10_P_btm.n352 C10_P_btm.n351 0.09425
R30265 C10_P_btm.n351 C10_P_btm.n81 0.09425
R30266 C10_P_btm.n182 C10_P_btm.n80 0.09425
R30267 C10_P_btm.n187 C10_P_btm.n182 0.09425
R30268 C10_P_btm.n350 C10_P_btm.n82 0.09425
R30269 C10_P_btm.n255 C10_P_btm.n82 0.09425
R30270 C10_P_btm.n256 C10_P_btm.n81 0.09425
R30271 C10_P_btm.n257 C10_P_btm.n256 0.09425
R30272 C10_P_btm.n348 C10_P_btm.n83 0.09425
R30273 C10_P_btm.n253 C10_P_btm.n83 0.09425
R30274 C10_P_btm.n255 C10_P_btm.n254 0.09425
R30275 C10_P_btm.n254 C10_P_btm.n188 0.09425
R30276 C10_P_btm.n253 C10_P_btm.n252 0.09425
R30277 C10_P_btm.n252 C10_P_btm.n190 0.09425
R30278 C10_P_btm.n189 C10_P_btm.n84 0.09425
R30279 C10_P_btm.n251 C10_P_btm.n189 0.09425
R30280 C10_P_btm.n344 C10_P_btm.n85 0.09425
R30281 C10_P_btm.n344 C10_P_btm.n343 0.09425
R30282 C10_P_btm.n343 C10_P_btm.n88 0.09425
R30283 C10_P_btm.n250 C10_P_btm.n86 0.09425
R30284 C10_P_btm.n250 C10_P_btm.n249 0.09425
R30285 C10_P_btm.n248 C10_P_btm.n88 0.09425
R30286 C10_P_btm.n248 C10_P_btm.n166 0.09425
R30287 C10_P_btm.n249 C10_P_btm.n167 0.09425
R30288 C10_P_btm.n275 C10_P_btm.n167 0.09425
R30289 C10_P_btm.n276 C10_P_btm.n166 0.09425
R30290 C10_P_btm.n276 C10_P_btm.n164 0.09425
R30291 C10_P_btm.n275 C10_P_btm.n274 0.09425
R30292 C10_P_btm.n274 C10_P_btm.n170 0.09425
R30293 C10_P_btm.n169 C10_P_btm.n164 0.09425
R30294 C10_P_btm.n278 C10_P_btm.n163 0.09425
R30295 C10_P_btm.n279 C10_P_btm.n159 0.09425
R30296 C10_P_btm.n279 C10_P_btm.n162 0.09425
R30297 C10_P_btm.n277 C10_P_btm.n165 0.09425
R30298 C10_P_btm.n278 C10_P_btm.n277 0.09425
R30299 C10_P_btm.n246 C10_P_btm.n202 0.09425
R30300 C10_P_btm.n202 C10_P_btm.n159 0.09425
R30301 C10_P_btm.n247 C10_P_btm.n89 0.09425
R30302 C10_P_btm.n247 C10_P_btm.n165 0.09425
R30303 C10_P_btm.n341 C10_P_btm.n90 0.09425
R30304 C10_P_btm.n246 C10_P_btm.n90 0.09425
R30305 C10_P_btm.n342 C10_P_btm.n87 0.09425
R30306 C10_P_btm.n342 C10_P_btm.n89 0.09425
R30307 C10_P_btm.n203 C10_P_btm.n91 0.09425
R30308 C10_P_btm.n245 C10_P_btm.n203 0.09425
R30309 C10_P_btm.n244 C10_P_btm.n204 0.09425
R30310 C10_P_btm.n244 C10_P_btm.n157 0.09425
R30311 C10_P_btm.n245 C10_P_btm.n158 0.09425
R30312 C10_P_btm.n281 C10_P_btm.n158 0.09425
R30313 C10_P_btm.n282 C10_P_btm.n157 0.09425
R30314 C10_P_btm.n282 C10_P_btm.n155 0.09425
R30315 C10_P_btm.n281 C10_P_btm.n280 0.09425
R30316 C10_P_btm.n280 C10_P_btm.n161 0.09425
R30317 C10_P_btm.n160 C10_P_btm.n155 0.09425
R30318 C10_P_btm.n284 C10_P_btm.n154 0.09425
R30319 C10_P_btm.n285 C10_P_btm.n150 0.09425
R30320 C10_P_btm.n285 C10_P_btm.n153 0.09425
R30321 C10_P_btm.n283 C10_P_btm.n156 0.09425
R30322 C10_P_btm.n284 C10_P_btm.n283 0.09425
R30323 C10_P_btm.n242 C10_P_btm.n206 0.09425
R30324 C10_P_btm.n206 C10_P_btm.n150 0.09425
R30325 C10_P_btm.n243 C10_P_btm.n205 0.09425
R30326 C10_P_btm.n243 C10_P_btm.n156 0.09425
R30327 C10_P_btm.n241 C10_P_btm.n94 0.09425
R30328 C10_P_btm.n242 C10_P_btm.n241 0.09425
R30329 C10_P_btm.n337 C10_P_btm.n93 0.09425
R30330 C10_P_btm.n205 C10_P_btm.n93 0.09425
R30331 C10_P_btm.n240 C10_P_btm.n95 0.09425
R30332 C10_P_btm.n240 C10_P_btm.n207 0.09425
R30333 C10_P_btm.n239 C10_P_btm.n238 0.09425
R30334 C10_P_btm.n238 C10_P_btm.n148 0.09425
R30335 C10_P_btm.n207 C10_P_btm.n149 0.09425
R30336 C10_P_btm.n287 C10_P_btm.n149 0.09425
R30337 C10_P_btm.n288 C10_P_btm.n148 0.09425
R30338 C10_P_btm.n288 C10_P_btm.n146 0.09425
R30339 C10_P_btm.n287 C10_P_btm.n286 0.09425
R30340 C10_P_btm.n286 C10_P_btm.n152 0.09425
R30341 C10_P_btm.n151 C10_P_btm.n146 0.09425
R30342 C10_P_btm.n290 C10_P_btm.n145 0.09425
R30343 C10_P_btm.n291 C10_P_btm.n144 0.09425
R30344 C10_P_btm.n291 C10_P_btm.n142 0.09425
R30345 C10_P_btm.n289 C10_P_btm.n147 0.09425
R30346 C10_P_btm.n290 C10_P_btm.n289 0.09425
R30347 C10_P_btm.n236 C10_P_btm.n209 0.09425
R30348 C10_P_btm.n209 C10_P_btm.n144 0.09425
R30349 C10_P_btm.n237 C10_P_btm.n208 0.09425
R30350 C10_P_btm.n237 C10_P_btm.n147 0.09425
R30351 C10_P_btm.n235 C10_P_btm.n98 0.09425
R30352 C10_P_btm.n236 C10_P_btm.n235 0.09425
R30353 C10_P_btm.n331 C10_P_btm.n97 0.09425
R30354 C10_P_btm.n208 C10_P_btm.n97 0.09425
R30355 C10_P_btm.n234 C10_P_btm.n99 0.09425
R30356 C10_P_btm.n234 C10_P_btm.n210 0.09425
R30357 C10_P_btm.n233 C10_P_btm.n232 0.09425
R30358 C10_P_btm.n232 C10_P_btm.n213 0.09425
R30359 C10_P_btm.n212 C10_P_btm.n210 0.09425
R30360 C10_P_btm.n212 C10_P_btm.n143 0.09425
R30361 C10_P_btm.n215 C10_P_btm.n213 0.09425
R30362 C10_P_btm.n215 C10_P_btm.n141 0.09425
R30363 C10_P_btm.n292 C10_P_btm.n143 0.09425
R30364 C10_P_btm.n293 C10_P_btm.n292 0.09425
R30365 C10_P_btm.n294 C10_P_btm.n141 0.09425
R30366 C10_P_btm.n295 C10_P_btm.n140 0.09425
R30367 C10_P_btm.n298 C10_P_btm.n297 0.09425
R30368 C10_P_btm.n217 C10_P_btm.n139 0.09425
R30369 C10_P_btm.n296 C10_P_btm.n139 0.09425
R30370 C10_P_btm.n216 C10_P_btm.n214 0.09425
R30371 C10_P_btm.n216 C10_P_btm.n140 0.09425
R30372 C10_P_btm.n230 C10_P_btm.n218 0.09425
R30373 C10_P_btm.n218 C10_P_btm.n217 0.09425
R30374 C10_P_btm.n231 C10_P_btm.n211 0.09425
R30375 C10_P_btm.n231 C10_P_btm.n214 0.09425
R30376 C10_P_btm.n229 C10_P_btm.n102 0.09425
R30377 C10_P_btm.n230 C10_P_btm.n229 0.09425
R30378 C10_P_btm.n325 C10_P_btm.n101 0.09425
R30379 C10_P_btm.n211 C10_P_btm.n101 0.09425
R30380 C10_P_btm.n323 C10_P_btm.n103 0.09425
R30381 C10_P_btm.n228 C10_P_btm.n103 0.09425
R30382 C10_P_btm.n227 C10_P_btm.n104 0.09425
R30383 C10_P_btm.n227 C10_P_btm.n221 0.09425
R30384 C10_P_btm.n228 C10_P_btm.n220 0.09425
R30385 C10_P_btm.n220 C10_P_btm.n219 0.09425
R30386 C10_P_btm.n221 C10_P_btm.n124 0.09425
R30387 C10_P_btm.n300 C10_P_btm.n124 0.09425
R30388 C10_P_btm.n219 C10_P_btm.n125 0.09425
R30389 C10_P_btm.n298 C10_P_btm.n125 0.09425
R30390 C10_P_btm.n301 C10_P_btm.n122 0.09425
R30391 C10_P_btm.n301 C10_P_btm.n123 0.09425
R30392 C10_P_btm.n300 C10_P_btm.n299 0.09425
R30393 C10_P_btm.n299 C10_P_btm.n138 0.09425
R30394 C10_P_btm.n137 C10_P_btm.n123 0.09425
R30395 C10_P_btm.n135 C10_P_btm.n120 0.09425
R30396 C10_P_btm.n302 C10_P_btm.n121 0.09425
R30397 C10_P_btm.n136 C10_P_btm.n121 0.09425
R30398 C10_P_btm.n304 C10_P_btm.n303 0.09425
R30399 C10_P_btm.n303 C10_P_btm.n120 0.09425
R30400 C10_P_btm.n223 C10_P_btm.n119 0.09425
R30401 C10_P_btm.n302 C10_P_btm.n119 0.09425
R30402 C10_P_btm.n226 C10_P_btm.n222 0.09425
R30403 C10_P_btm.n222 C10_P_btm.n122 0.09425
R30404 C10_P_btm.n225 C10_P_btm.n106 0.09425
R30405 C10_P_btm.n225 C10_P_btm.n223 0.09425
R30406 C10_P_btm.n321 C10_P_btm.n105 0.09425
R30407 C10_P_btm.n226 C10_P_btm.n105 0.09425
R30408 C10_P_btm.n317 C10_P_btm.n107 0.09425
R30409 C10_P_btm.n224 C10_P_btm.n107 0.09425
R30410 C10_P_btm.n116 C10_P_btm.n108 0.09425
R30411 C10_P_btm.n306 C10_P_btm.n116 0.09425
R30412 C10_P_btm.n224 C10_P_btm.n117 0.09425
R30413 C10_P_btm.n304 C10_P_btm.n117 0.09425
R30414 C10_P_btm.n307 C10_P_btm.n114 0.09425
R30415 C10_P_btm.n307 C10_P_btm.n115 0.09425
R30416 C10_P_btm.n306 C10_P_btm.n305 0.09425
R30417 C10_P_btm.n305 C10_P_btm.n118 0.09425
R30418 C10_P_btm.n127 C10_P_btm.n115 0.09425
R30419 C10_P_btm.n132 C10_P_btm.n127 0.09425
R30420 C10_P_btm.n133 C10_P_btm.n118 0.09425
R30421 C10_P_btm.n134 C10_P_btm.n133 0.09425
R30422 C10_P_btm.n132 C10_P_btm.n126 0.09425
R30423 C10_P_btm.n131 C10_P_btm.n128 0.09425
R30424 C10_P_btm.n129 C10_P_btm.n112 0.09425
R30425 C10_P_btm.n308 C10_P_btm.n113 0.09425
R30426 C10_P_btm.n128 C10_P_btm.n113 0.09425
R30427 C10_P_btm.n311 C10_P_btm.n310 0.09425
R30428 C10_P_btm.n310 C10_P_btm.n309 0.09425
R30429 C10_P_btm.n309 C10_P_btm.n112 0.09425
R30430 C10_P_btm.n111 C10_P_btm.n110 0.09425
R30431 C10_P_btm.n308 C10_P_btm.n111 0.09425
R30432 C10_P_btm.n315 C10_P_btm.n109 0.09425
R30433 C10_P_btm.n114 C10_P_btm.n109 0.09425
R30434 C10_P_btm.n313 C10_P_btm.n311 0.09425
R30435 C10_P_btm.n312 C10_P_btm.n33 0.09425
R30436 C10_P_btm.n313 C10_P_btm.n312 0.09425
R30437 C10_P_btm.n314 C10_P_btm.n35 0.09425
R30438 C10_P_btm.n314 C10_P_btm.n110 0.09425
R30439 C10_P_btm.n1041 C10_P_btm.n36 0.09425
R30440 C10_P_btm.n315 C10_P_btm.n36 0.09425
R30441 C10_P_btm.n316 C10_P_btm.n38 0.09425
R30442 C10_P_btm.n316 C10_P_btm.n108 0.09425
R30443 C10_P_btm.n1039 C10_P_btm.n39 0.09425
R30444 C10_P_btm.n317 C10_P_btm.n39 0.09425
R30445 C10_P_btm.n319 C10_P_btm.n318 0.09425
R30446 C10_P_btm.n318 C10_P_btm.n106 0.09425
R30447 C10_P_btm.n320 C10_P_btm.n41 0.09425
R30448 C10_P_btm.n321 C10_P_btm.n320 0.09425
R30449 C10_P_btm.n322 C10_P_btm.n43 0.09425
R30450 C10_P_btm.n322 C10_P_btm.n104 0.09425
R30451 C10_P_btm.n1033 C10_P_btm.n44 0.09425
R30452 C10_P_btm.n323 C10_P_btm.n44 0.09425
R30453 C10_P_btm.n324 C10_P_btm.n46 0.09425
R30454 C10_P_btm.n324 C10_P_btm.n102 0.09425
R30455 C10_P_btm.n1031 C10_P_btm.n47 0.09425
R30456 C10_P_btm.n325 C10_P_btm.n47 0.09425
R30457 C10_P_btm.n327 C10_P_btm.n326 0.09425
R30458 C10_P_btm.n326 C10_P_btm.n100 0.09425
R30459 C10_P_btm.n328 C10_P_btm.n49 0.09425
R30460 C10_P_btm.n329 C10_P_btm.n328 0.09425
R30461 C10_P_btm.n330 C10_P_btm.n51 0.09425
R30462 C10_P_btm.n330 C10_P_btm.n98 0.09425
R30463 C10_P_btm.n1025 C10_P_btm.n52 0.09425
R30464 C10_P_btm.n331 C10_P_btm.n52 0.09425
R30465 C10_P_btm.n332 C10_P_btm.n54 0.09425
R30466 C10_P_btm.n332 C10_P_btm.n96 0.09425
R30467 C10_P_btm.n1023 C10_P_btm.n55 0.09425
R30468 C10_P_btm.n333 C10_P_btm.n55 0.09425
R30469 C10_P_btm.n335 C10_P_btm.n334 0.09425
R30470 C10_P_btm.n334 C10_P_btm.n94 0.09425
R30471 C10_P_btm.n336 C10_P_btm.n57 0.09425
R30472 C10_P_btm.n337 C10_P_btm.n336 0.09425
R30473 C10_P_btm.n338 C10_P_btm.n59 0.09425
R30474 C10_P_btm.n338 C10_P_btm.n92 0.09425
R30475 C10_P_btm.n1017 C10_P_btm.n60 0.09425
R30476 C10_P_btm.n339 C10_P_btm.n60 0.09425
R30477 C10_P_btm.n340 C10_P_btm.n62 0.09425
R30478 C10_P_btm.n341 C10_P_btm.n340 0.09425
R30479 C10_P_btm.n1015 C10_P_btm.n63 0.09425
R30480 C10_P_btm.n87 C10_P_btm.n63 0.09425
R30481 C10_P_btm.n346 C10_P_btm.n345 0.09425
R30482 C10_P_btm.n345 C10_P_btm.n86 0.09425
R30483 C10_P_btm.n1011 C10_P_btm.n67 0.09425
R30484 C10_P_btm.n347 C10_P_btm.n67 0.09425
R30485 C10_P_btm.n347 C10_P_btm.n84 0.09425
R30486 C10_P_btm.n349 C10_P_btm.n68 0.09425
R30487 C10_P_btm.n349 C10_P_btm.n348 0.09425
R30488 C10_P_btm.n1008 C10_P_btm.n71 0.09425
R30489 C10_P_btm.n350 C10_P_btm.n71 0.09425
R30490 C10_P_btm.n1009 C10_P_btm.n70 0.09425
R30491 C10_P_btm.n1009 C10_P_btm.n68 0.09425
R30492 C10_P_btm.n1007 C10_P_btm.n73 0.09425
R30493 C10_P_btm.n1008 C10_P_btm.n1007 0.09425
R30494 C10_P_btm.n976 C10_P_btm.n975 0.09425
R30495 C10_P_btm.n975 C10_P_btm.n70 0.09425
R30496 C10_P_btm.n982 C10_P_btm.n977 0.09425
R30497 C10_P_btm.n977 C10_P_btm.n73 0.09425
R30498 C10_P_btm.n983 C10_P_btm.n969 0.09425
R30499 C10_P_btm.n983 C10_P_btm.n976 0.09425
R30500 C10_P_btm.n994 C10_P_btm.n366 0.09425
R30501 C10_P_btm.n982 C10_P_btm.n366 0.09425
R30502 C10_P_btm.n992 C10_P_btm.n367 0.09425
R30503 C10_P_btm.n969 C10_P_btm.n367 0.09425
R30504 C10_P_btm.n993 C10_P_btm.n368 0.09425
R30505 C10_P_btm.n994 C10_P_btm.n993 0.09425
R30506 C10_P_btm.n991 C10_P_btm.n370 0.09425
R30507 C10_P_btm.n992 C10_P_btm.n991 0.09425
R30508 C10_P_btm.n962 C10_P_btm.n375 0.09425
R30509 C10_P_btm.n375 C10_P_btm.n368 0.09425
R30510 C10_P_btm.n910 C10_P_btm.n374 0.09425
R30511 C10_P_btm.n963 C10_P_btm.n374 0.09425
R30512 C10_P_btm.n963 C10_P_btm.n370 0.09425
R30513 C10_P_btm.n961 C10_P_btm.n377 0.09425
R30514 C10_P_btm.n962 C10_P_btm.n961 0.09425
R30515 C10_P_btm.n959 C10_P_btm.n379 0.09425
R30516 C10_P_btm.n960 C10_P_btm.n959 0.09425
R30517 C10_P_btm.n911 C10_P_btm.n908 0.09425
R30518 C10_P_btm.n911 C10_P_btm.n377 0.09425
R30519 C10_P_btm.n906 C10_P_btm.n903 0.09425
R30520 C10_P_btm.n903 C10_P_btm.n379 0.09425
R30521 C10_P_btm.n907 C10_P_btm.n898 0.09425
R30522 C10_P_btm.n908 C10_P_btm.n907 0.09425
R30523 C10_P_btm.n920 C10_P_btm.n897 0.09425
R30524 C10_P_btm.n906 C10_P_btm.n897 0.09425
R30525 C10_P_btm.n919 C10_P_btm.n894 0.09425
R30526 C10_P_btm.n919 C10_P_btm.n898 0.09425
R30527 C10_P_btm.n930 C10_P_btm.n895 0.09425
R30528 C10_P_btm.n920 C10_P_btm.n895 0.09425
R30529 C10_P_btm.n931 C10_P_btm.n892 0.09425
R30530 C10_P_btm.n931 C10_P_btm.n894 0.09425
R30531 C10_P_btm.n929 C10_P_btm.n926 0.09425
R30532 C10_P_btm.n930 C10_P_btm.n929 0.09425
R30533 C10_P_btm.n925 C10_P_btm.n924 0.09425
R30534 C10_P_btm.n925 C10_P_btm.n892 0.09425
R30535 C10_P_btm.n942 C10_P_btm.n409 0.09425
R30536 C10_P_btm.n926 C10_P_btm.n409 0.09425
R30537 C10_P_btm.n940 C10_P_btm.n412 0.09425
R30538 C10_P_btm.n940 C10_P_btm.n410 0.09425
R30539 C10_P_btm.n924 C10_P_btm.n410 0.09425
R30540 C10_P_btm.n941 C10_P_btm.n411 0.09425
R30541 C10_P_btm.n942 C10_P_btm.n941 0.09425
R30542 C10_P_btm.n422 C10_P_btm.n420 0.09425
R30543 C10_P_btm.n422 C10_P_btm.n407 0.09425
R30544 C10_P_btm.n884 C10_P_btm.n412 0.09425
R30545 C10_P_btm.n883 C10_P_btm.n417 0.09425
R30546 C10_P_btm.n884 C10_P_btm.n883 0.09425
R30547 C10_P_btm.n882 C10_P_btm.n416 0.09425
R30548 C10_P_btm.n416 C10_P_btm.n411 0.09425
R30549 C10_P_btm.n881 C10_P_btm.n419 0.09425
R30550 C10_P_btm.n881 C10_P_btm.n420 0.09425
R30551 C10_P_btm.n879 C10_P_btm.n427 0.09425
R30552 C10_P_btm.n880 C10_P_btm.n879 0.09425
R30553 C10_P_btm.n877 C10_P_btm.n876 0.09425
R30554 C10_P_btm.n878 C10_P_btm.n877 0.09425
R30555 C10_P_btm.n874 C10_P_btm.n428 0.09425
R30556 C10_P_btm.n428 C10_P_btm.n427 0.09425
R30557 C10_P_btm.n875 C10_P_btm.n429 0.09425
R30558 C10_P_btm.n876 C10_P_btm.n875 0.09425
R30559 C10_P_btm.n873 C10_P_btm.n431 0.09425
R30560 C10_P_btm.n874 C10_P_btm.n873 0.09425
R30561 C10_P_btm.n452 C10_P_btm.n451 0.09425
R30562 C10_P_btm.n451 C10_P_btm.n429 0.09425
R30563 C10_P_btm.n458 C10_P_btm.n453 0.09425
R30564 C10_P_btm.n453 C10_P_btm.n431 0.09425
R30565 C10_P_btm.n460 C10_P_btm.n459 0.09425
R30566 C10_P_btm.n459 C10_P_btm.n452 0.09425
R30567 C10_P_btm.n837 C10_P_btm.n450 0.09425
R30568 C10_P_btm.n458 C10_P_btm.n450 0.09425
R30569 C10_P_btm.n461 C10_P_btm.n460 0.09425
R30570 C10_P_btm.n835 C10_P_btm.n461 0.09425
R30571 C10_P_btm.n835 C10_P_btm.n834 0.09425
R30572 C10_P_btm.n813 C10_P_btm.n463 0.09425
R30573 C10_P_btm.n833 C10_P_btm.n463 0.09425
R30574 C10_P_btm.n834 C10_P_btm.n833 0.09425
R30575 C10_P_btm.n832 C10_P_btm.n464 0.09425
R30576 C10_P_btm.n832 C10_P_btm.n462 0.09425
R30577 C10_P_btm.n831 C10_P_btm.n830 0.09425
R30578 C10_P_btm.n830 C10_P_btm.n448 0.09425
R30579 C10_P_btm.n836 C10_P_btm.n462 0.09425
R30580 C10_P_btm.n837 C10_P_btm.n836 0.09425
R30581 C10_P_btm.n829 C10_P_btm.n447 0.09425
R30582 C10_P_btm.n839 C10_P_btm.n447 0.09425
R30583 C10_P_btm.n838 C10_P_btm.n448 0.09425
R30584 C10_P_btm.n838 C10_P_btm.n449 0.09425
R30585 C10_P_btm.n839 C10_P_btm.n445 0.09425
R30586 C10_P_btm.n456 C10_P_btm.n445 0.09425
R30587 C10_P_btm.n457 C10_P_btm.n449 0.09425
R30588 C10_P_btm.n457 C10_P_btm.n454 0.09425
R30589 C10_P_btm.n456 C10_P_btm.n455 0.09425
R30590 C10_P_btm.n455 C10_P_btm.n433 0.09425
R30591 C10_P_btm.n454 C10_P_btm.n432 0.09425
R30592 C10_P_btm.n872 C10_P_btm.n432 0.09425
R30593 C10_P_btm.n871 C10_P_btm.n433 0.09425
R30594 C10_P_btm.n871 C10_P_btm.n434 0.09425
R30595 C10_P_btm.n872 C10_P_btm.n430 0.09425
R30596 C10_P_btm.n856 C10_P_btm.n430 0.09425
R30597 C10_P_btm.n857 C10_P_btm.n434 0.09425
R30598 C10_P_btm.n857 C10_P_btm.n854 0.09425
R30599 C10_P_btm.n856 C10_P_btm.n855 0.09425
R30600 C10_P_btm.n855 C10_P_btm.n419 0.09425
R30601 C10_P_btm.n854 C10_P_btm.n418 0.09425
R30602 C10_P_btm.n882 C10_P_btm.n418 0.09425
R30603 C10_P_btm.n858 C10_P_btm.n853 0.09425
R30604 C10_P_btm.n853 C10_P_btm.n417 0.09425
R30605 C10_P_btm.n859 C10_P_btm.n848 0.09425
R30606 C10_P_btm.n859 C10_P_btm.n852 0.09425
R30607 C10_P_btm.n870 C10_P_btm.n435 0.09425
R30608 C10_P_btm.n858 C10_P_btm.n435 0.09425
R30609 C10_P_btm.n868 C10_P_btm.n436 0.09425
R30610 C10_P_btm.n848 C10_P_btm.n436 0.09425
R30611 C10_P_btm.n869 C10_P_btm.n437 0.09425
R30612 C10_P_btm.n870 C10_P_btm.n869 0.09425
R30613 C10_P_btm.n867 C10_P_btm.n439 0.09425
R30614 C10_P_btm.n868 C10_P_btm.n867 0.09425
R30615 C10_P_btm.n841 C10_P_btm.n444 0.09425
R30616 C10_P_btm.n444 C10_P_btm.n437 0.09425
R30617 C10_P_btm.n842 C10_P_btm.n443 0.09425
R30618 C10_P_btm.n842 C10_P_btm.n439 0.09425
R30619 C10_P_btm.n840 C10_P_btm.n446 0.09425
R30620 C10_P_btm.n841 C10_P_btm.n840 0.09425
R30621 C10_P_btm.n827 C10_P_btm.n468 0.09425
R30622 C10_P_btm.n827 C10_P_btm.n826 0.09425
R30623 C10_P_btm.n826 C10_P_btm.n443 0.09425
R30624 C10_P_btm.n828 C10_P_btm.n467 0.09425
R30625 C10_P_btm.n828 C10_P_btm.n446 0.09425
R30626 C10_P_btm.n476 C10_P_btm.n465 0.09425
R30627 C10_P_btm.n829 C10_P_btm.n465 0.09425
R30628 C10_P_btm.n819 C10_P_btm.n468 0.09425
R30629 C10_P_btm.n818 C10_P_btm.n473 0.09425
R30630 C10_P_btm.n819 C10_P_btm.n818 0.09425
R30631 C10_P_btm.n817 C10_P_btm.n472 0.09425
R30632 C10_P_btm.n472 C10_P_btm.n467 0.09425
R30633 C10_P_btm.n816 C10_P_btm.n475 0.09425
R30634 C10_P_btm.n816 C10_P_btm.n476 0.09425
R30635 C10_P_btm.n815 C10_P_btm.n466 0.09425
R30636 C10_P_btm.n831 C10_P_btm.n466 0.09425
R30637 C10_P_btm.n814 C10_P_btm.n478 0.09425
R30638 C10_P_btm.n814 C10_P_btm.n464 0.09425
R30639 C10_P_btm.n506 C10_P_btm.n479 0.09425
R30640 C10_P_btm.n811 C10_P_btm.n479 0.09425
R30641 C10_P_btm.n812 C10_P_btm.n811 0.09425
R30642 C10_P_btm.n813 C10_P_btm.n812 0.09425
R30643 C10_P_btm.n810 C10_P_btm.n480 0.09425
R30644 C10_P_btm.n810 C10_P_btm.n478 0.09425
R30645 C10_P_btm.n809 C10_P_btm.n477 0.09425
R30646 C10_P_btm.n815 C10_P_btm.n477 0.09425
R30647 C10_P_btm.n807 C10_P_btm.n481 0.09425
R30648 C10_P_btm.n481 C10_P_btm.n475 0.09425
R30649 C10_P_btm.n721 C10_P_btm.n474 0.09425
R30650 C10_P_btm.n817 C10_P_btm.n474 0.09425
R30651 C10_P_btm.n722 C10_P_btm.n720 0.09425
R30652 C10_P_btm.n722 C10_P_btm.n473 0.09425
R30653 C10_P_btm.n723 C10_P_btm.n685 0.09425
R30654 C10_P_btm.n685 C10_P_btm.n471 0.09425
R30655 C10_P_btm.n724 C10_P_btm.n686 0.09425
R30656 C10_P_btm.n725 C10_P_btm.n724 0.09425
R30657 C10_P_btm.n714 C10_P_btm.n682 0.09425
R30658 C10_P_btm.n704 C10_P_btm.n688 0.09425
R30659 C10_P_btm.n714 C10_P_btm.n688 0.09425
R30660 C10_P_btm.n716 C10_P_btm.n715 0.09425
R30661 C10_P_btm.n715 C10_P_btm.n683 0.09425
R30662 C10_P_btm.n717 C10_P_btm.n687 0.09425
R30663 C10_P_btm.n717 C10_P_btm.n686 0.09425
R30664 C10_P_btm.n719 C10_P_btm.n718 0.09425
R30665 C10_P_btm.n723 C10_P_btm.n719 0.09425
R30666 C10_P_btm.n803 C10_P_btm.n485 0.09425
R30667 C10_P_btm.n720 C10_P_btm.n485 0.09425
R30668 C10_P_btm.n805 C10_P_btm.n483 0.09425
R30669 C10_P_btm.n721 C10_P_btm.n483 0.09425
R30670 C10_P_btm.n806 C10_P_btm.n484 0.09425
R30671 C10_P_btm.n807 C10_P_btm.n806 0.09425
R30672 C10_P_btm.n808 C10_P_btm.n482 0.09425
R30673 C10_P_btm.n809 C10_P_btm.n808 0.09425
R30674 C10_P_btm.n508 C10_P_btm.n504 0.09425
R30675 C10_P_btm.n504 C10_P_btm.n480 0.09425
R30676 C10_P_btm.n517 C10_P_btm.n501 0.09425
R30677 C10_P_btm.n505 C10_P_btm.n501 0.09425
R30678 C10_P_btm.n507 C10_P_btm.n505 0.09425
R30679 C10_P_btm.n507 C10_P_btm.n506 0.09425
R30680 C10_P_btm.n503 C10_P_btm.n502 0.09425
R30681 C10_P_btm.n508 C10_P_btm.n503 0.09425
R30682 C10_P_btm.n510 C10_P_btm.n509 0.09425
R30683 C10_P_btm.n509 C10_P_btm.n482 0.09425
R30684 C10_P_btm.n513 C10_P_btm.n511 0.09425
R30685 C10_P_btm.n511 C10_P_btm.n484 0.09425
R30686 C10_P_btm.n804 C10_P_btm.n486 0.09425
R30687 C10_P_btm.n805 C10_P_btm.n804 0.09425
R30688 C10_P_btm.n802 C10_P_btm.n488 0.09425
R30689 C10_P_btm.n803 C10_P_btm.n802 0.09425
R30690 C10_P_btm.n801 C10_P_btm.n487 0.09425
R30691 C10_P_btm.n718 C10_P_btm.n487 0.09425
R30692 C10_P_btm.n799 C10_P_btm.n489 0.09425
R30693 C10_P_btm.n687 C10_P_btm.n489 0.09425
R30694 C10_P_btm.n705 C10_P_btm.n689 0.09425
R30695 C10_P_btm.n716 C10_P_btm.n689 0.09425
R30696 C10_P_btm.n706 C10_P_btm.n703 0.09425
R30697 C10_P_btm.n706 C10_P_btm.n704 0.09425
R30698 C10_P_btm.n707 C10_P_btm.n692 0.09425
R30699 C10_P_btm.n692 C10_P_btm.n690 0.09425
R30700 C10_P_btm.n708 C10_P_btm.n693 0.09425
R30701 C10_P_btm.n709 C10_P_btm.n708 0.09425
R30702 C10_P_btm.n697 C10_P_btm.n694 0.09425
R30703 C10_P_btm.n789 C10_P_btm.n532 0.09425
R30704 C10_P_btm.n697 C10_P_btm.n532 0.09425
R30705 C10_P_btm.n698 C10_P_btm.n531 0.09425
R30706 C10_P_btm.n699 C10_P_btm.n698 0.09425
R30707 C10_P_btm.n700 C10_P_btm.n529 0.09425
R30708 C10_P_btm.n700 C10_P_btm.n693 0.09425
R30709 C10_P_btm.n702 C10_P_btm.n701 0.09425
R30710 C10_P_btm.n707 C10_P_btm.n702 0.09425
R30711 C10_P_btm.n795 C10_P_btm.n493 0.09425
R30712 C10_P_btm.n703 C10_P_btm.n493 0.09425
R30713 C10_P_btm.n797 C10_P_btm.n491 0.09425
R30714 C10_P_btm.n705 C10_P_btm.n491 0.09425
R30715 C10_P_btm.n798 C10_P_btm.n492 0.09425
R30716 C10_P_btm.n799 C10_P_btm.n798 0.09425
R30717 C10_P_btm.n800 C10_P_btm.n490 0.09425
R30718 C10_P_btm.n801 C10_P_btm.n800 0.09425
R30719 C10_P_btm.n523 C10_P_btm.n495 0.09425
R30720 C10_P_btm.n495 C10_P_btm.n488 0.09425
R30721 C10_P_btm.n512 C10_P_btm.n497 0.09425
R30722 C10_P_btm.n512 C10_P_btm.n486 0.09425
R30723 C10_P_btm.n521 C10_P_btm.n498 0.09425
R30724 C10_P_btm.n513 C10_P_btm.n498 0.09425
R30725 C10_P_btm.n515 C10_P_btm.n514 0.09425
R30726 C10_P_btm.n514 C10_P_btm.n510 0.09425
R30727 C10_P_btm.n516 C10_P_btm.n500 0.09425
R30728 C10_P_btm.n516 C10_P_btm.n502 0.09425
R30729 C10_P_btm.n519 C10_P_btm.n499 0.09425
R30730 C10_P_btm.n515 C10_P_btm.n499 0.09425
R30731 C10_P_btm.n521 C10_P_btm.n520 0.09425
R30732 C10_P_btm.n522 C10_P_btm.n496 0.09425
R30733 C10_P_btm.n522 C10_P_btm.n497 0.09425
R30734 C10_P_btm.n523 C10_P_btm.n494 0.09425
R30735 C10_P_btm.n525 C10_P_btm.n524 0.09425
R30736 C10_P_btm.n524 C10_P_btm.n490 0.09425
R30737 C10_P_btm.n526 C10_P_btm.n492 0.09425
R30738 C10_P_btm.n796 C10_P_btm.n527 0.09425
R30739 C10_P_btm.n797 C10_P_btm.n796 0.09425
R30740 C10_P_btm.n795 C10_P_btm.n794 0.09425
R30741 C10_P_btm.n793 C10_P_btm.n528 0.09425
R30742 C10_P_btm.n701 C10_P_btm.n528 0.09425
R30743 C10_P_btm.n792 C10_P_btm.n529 0.09425
R30744 C10_P_btm.n791 C10_P_btm.n790 0.09425
R30745 C10_P_btm.n790 C10_P_btm.n531 0.09425
R30746 C10_P_btm.n789 C10_P_btm.n530 0.09425
R30747 C10_P_btm.n788 C10_P_btm.n533 0.09425
R30748 C10_P_btm.n788 C10_P_btm.n534 0.09425
R30749 C10_P_btm.n787 C10_P_btm.n786 0.09425
R30750 C10_P_btm.n785 C10_P_btm.n536 0.09425
R30751 C10_P_btm.n558 C10_P_btm.n554 0.09425
R30752 C10_P_btm.n566 C10_P_btm.n552 0.09425
R30753 C10_P_btm.n570 C10_P_btm.n549 0.09425
R30754 C10_P_btm.n774 C10_P_btm.n547 0.09425
R30755 C10_P_btm.n581 C10_P_btm.n580 0.09425
R30756 C10_P_btm.n780 C10_P_btm.n542 0.09425
R30757 C10_P_btm.n729 C10_P_btm.n680 0.09425
R30758 C10_P_btm.n731 C10_P_btm.n603 0.09425
R30759 C10_P_btm.n731 C10_P_btm.n730 0.09425
R30760 C10_P_btm.n733 C10_P_btm.n600 0.09425
R30761 C10_P_btm.n736 C10_P_btm.n735 0.09425
R30762 C10_P_btm.n735 C10_P_btm.n734 0.09425
R30763 C10_P_btm.n734 C10_P_btm.n601 0.09425
R30764 C10_P_btm.n733 C10_P_btm.n732 0.09425
R30765 C10_P_btm.n732 C10_P_btm.n679 0.09425
R30766 C10_P_btm.n678 C10_P_btm.n601 0.09425
R30767 C10_P_btm.n677 C10_P_btm.n604 0.09425
R30768 C10_P_btm.n675 C10_P_btm.n606 0.09425
R30769 C10_P_btm.n676 C10_P_btm.n675 0.09425
R30770 C10_P_btm.n602 C10_P_btm.n598 0.09425
R30771 C10_P_btm.n604 C10_P_btm.n602 0.09425
R30772 C10_P_btm.n633 C10_P_btm.n595 0.09425
R30773 C10_P_btm.n633 C10_P_btm.n606 0.09425
R30774 C10_P_btm.n738 C10_P_btm.n737 0.09425
R30775 C10_P_btm.n737 C10_P_btm.n598 0.09425
R30776 C10_P_btm.n739 C10_P_btm.n593 0.09425
R30777 C10_P_btm.n739 C10_P_btm.n595 0.09425
R30778 C10_P_btm.n741 C10_P_btm.n592 0.09425
R30779 C10_P_btm.n590 C10_P_btm.n538 0.09425
R30780 C10_P_btm.n742 C10_P_btm.n590 0.09425
R30781 C10_P_btm.n742 C10_P_btm.n587 0.09425
R30782 C10_P_btm.n741 C10_P_btm.n740 0.09425
R30783 C10_P_btm.n740 C10_P_btm.n594 0.09425
R30784 C10_P_btm.n632 C10_P_btm.n587 0.09425
R30785 C10_P_btm.n635 C10_P_btm.n632 0.09425
R30786 C10_P_btm.n634 C10_P_btm.n594 0.09425
R30787 C10_P_btm.n634 C10_P_btm.n607 0.09425
R30788 C10_P_btm.n635 C10_P_btm.n608 0.09425
R30789 C10_P_btm.n673 C10_P_btm.n608 0.09425
R30790 C10_P_btm.n674 C10_P_btm.n607 0.09425
R30791 C10_P_btm.n674 C10_P_btm.n605 0.09425
R30792 C10_P_btm.n673 C10_P_btm.n672 0.09425
R30793 C10_P_btm.n671 C10_P_btm.n609 0.09425
R30794 C10_P_btm.n669 C10_P_btm.n611 0.09425
R30795 C10_P_btm.n670 C10_P_btm.n669 0.09425
R30796 C10_P_btm.n636 C10_P_btm.n631 0.09425
R30797 C10_P_btm.n631 C10_P_btm.n609 0.09425
R30798 C10_P_btm.n637 C10_P_btm.n585 0.09425
R30799 C10_P_btm.n637 C10_P_btm.n611 0.09425
R30800 C10_P_btm.n744 C10_P_btm.n586 0.09425
R30801 C10_P_btm.n636 C10_P_btm.n586 0.09425
R30802 C10_P_btm.n745 C10_P_btm.n583 0.09425
R30803 C10_P_btm.n745 C10_P_btm.n585 0.09425
R30804 C10_P_btm.n743 C10_P_btm.n589 0.09425
R30805 C10_P_btm.n744 C10_P_btm.n743 0.09425
R30806 C10_P_btm.n588 C10_P_btm.n541 0.09425
R30807 C10_P_btm.n588 C10_P_btm.n583 0.09425
R30808 C10_P_btm.n782 C10_P_btm.n539 0.09425
R30809 C10_P_btm.n589 C10_P_btm.n539 0.09425
R30810 C10_P_btm.n582 C10_P_btm.n542 0.09425
R30811 C10_P_btm.n747 C10_P_btm.n582 0.09425
R30812 C10_P_btm.n748 C10_P_btm.n581 0.09425
R30813 C10_P_btm.n748 C10_P_btm.n576 0.09425
R30814 C10_P_btm.n747 C10_P_btm.n746 0.09425
R30815 C10_P_btm.n746 C10_P_btm.n584 0.09425
R30816 C10_P_btm.n630 C10_P_btm.n576 0.09425
R30817 C10_P_btm.n639 C10_P_btm.n630 0.09425
R30818 C10_P_btm.n638 C10_P_btm.n584 0.09425
R30819 C10_P_btm.n638 C10_P_btm.n612 0.09425
R30820 C10_P_btm.n639 C10_P_btm.n613 0.09425
R30821 C10_P_btm.n667 C10_P_btm.n613 0.09425
R30822 C10_P_btm.n668 C10_P_btm.n612 0.09425
R30823 C10_P_btm.n668 C10_P_btm.n610 0.09425
R30824 C10_P_btm.n667 C10_P_btm.n666 0.09425
R30825 C10_P_btm.n665 C10_P_btm.n614 0.09425
R30826 C10_P_btm.n663 C10_P_btm.n616 0.09425
R30827 C10_P_btm.n664 C10_P_btm.n663 0.09425
R30828 C10_P_btm.n640 C10_P_btm.n629 0.09425
R30829 C10_P_btm.n629 C10_P_btm.n614 0.09425
R30830 C10_P_btm.n641 C10_P_btm.n574 0.09425
R30831 C10_P_btm.n641 C10_P_btm.n616 0.09425
R30832 C10_P_btm.n750 C10_P_btm.n575 0.09425
R30833 C10_P_btm.n640 C10_P_btm.n575 0.09425
R30834 C10_P_btm.n751 C10_P_btm.n572 0.09425
R30835 C10_P_btm.n751 C10_P_btm.n574 0.09425
R30836 C10_P_btm.n749 C10_P_btm.n578 0.09425
R30837 C10_P_btm.n750 C10_P_btm.n749 0.09425
R30838 C10_P_btm.n577 C10_P_btm.n546 0.09425
R30839 C10_P_btm.n577 C10_P_btm.n572 0.09425
R30840 C10_P_btm.n579 C10_P_btm.n544 0.09425
R30841 C10_P_btm.n579 C10_P_btm.n578 0.09425
R30842 C10_P_btm.n571 C10_P_btm.n547 0.09425
R30843 C10_P_btm.n753 C10_P_btm.n571 0.09425
R30844 C10_P_btm.n754 C10_P_btm.n570 0.09425
R30845 C10_P_btm.n754 C10_P_btm.n565 0.09425
R30846 C10_P_btm.n753 C10_P_btm.n752 0.09425
R30847 C10_P_btm.n752 C10_P_btm.n573 0.09425
R30848 C10_P_btm.n628 C10_P_btm.n565 0.09425
R30849 C10_P_btm.n643 C10_P_btm.n628 0.09425
R30850 C10_P_btm.n642 C10_P_btm.n573 0.09425
R30851 C10_P_btm.n642 C10_P_btm.n617 0.09425
R30852 C10_P_btm.n643 C10_P_btm.n618 0.09425
R30853 C10_P_btm.n661 C10_P_btm.n618 0.09425
R30854 C10_P_btm.n662 C10_P_btm.n617 0.09425
R30855 C10_P_btm.n662 C10_P_btm.n615 0.09425
R30856 C10_P_btm.n661 C10_P_btm.n660 0.09425
R30857 C10_P_btm.n659 C10_P_btm.n619 0.09425
R30858 C10_P_btm.n657 C10_P_btm.n621 0.09425
R30859 C10_P_btm.n658 C10_P_btm.n657 0.09425
R30860 C10_P_btm.n644 C10_P_btm.n627 0.09425
R30861 C10_P_btm.n627 C10_P_btm.n619 0.09425
R30862 C10_P_btm.n645 C10_P_btm.n563 0.09425
R30863 C10_P_btm.n645 C10_P_btm.n621 0.09425
R30864 C10_P_btm.n756 C10_P_btm.n564 0.09425
R30865 C10_P_btm.n644 C10_P_btm.n564 0.09425
R30866 C10_P_btm.n757 C10_P_btm.n561 0.09425
R30867 C10_P_btm.n757 C10_P_btm.n563 0.09425
R30868 C10_P_btm.n755 C10_P_btm.n569 0.09425
R30869 C10_P_btm.n756 C10_P_btm.n755 0.09425
R30870 C10_P_btm.n568 C10_P_btm.n567 0.09425
R30871 C10_P_btm.n568 C10_P_btm.n561 0.09425
R30872 C10_P_btm.n772 C10_P_btm.n550 0.09425
R30873 C10_P_btm.n569 C10_P_btm.n550 0.09425
R30874 C10_P_btm.n566 C10_P_btm.n560 0.09425
R30875 C10_P_btm.n759 C10_P_btm.n560 0.09425
R30876 C10_P_btm.n760 C10_P_btm.n558 0.09425
R30877 C10_P_btm.n760 C10_P_btm.n559 0.09425
R30878 C10_P_btm.n759 C10_P_btm.n758 0.09425
R30879 C10_P_btm.n758 C10_P_btm.n562 0.09425
R30880 C10_P_btm.n648 C10_P_btm.n559 0.09425
R30881 C10_P_btm.n648 C10_P_btm.n647 0.09425
R30882 C10_P_btm.n646 C10_P_btm.n562 0.09425
R30883 C10_P_btm.n646 C10_P_btm.n622 0.09425
R30884 C10_P_btm.n647 C10_P_btm.n623 0.09425
R30885 C10_P_btm.n655 C10_P_btm.n623 0.09425
R30886 C10_P_btm.n656 C10_P_btm.n622 0.09425
R30887 C10_P_btm.n656 C10_P_btm.n620 0.09425
R30888 C10_P_btm.n655 C10_P_btm.n654 0.09425
R30889 C10_P_btm.n650 C10_P_btm.n625 0.09425
R30890 C10_P_btm.n625 C10_P_btm.n624 0.09425
R30891 C10_P_btm.n651 C10_P_btm.n626 0.09425
R30892 C10_P_btm.n652 C10_P_btm.n651 0.09425
R30893 C10_P_btm.n649 C10_P_btm.n557 0.09425
R30894 C10_P_btm.n650 C10_P_btm.n649 0.09425
R30895 C10_P_btm.n762 C10_P_btm.n556 0.09425
R30896 C10_P_btm.n626 C10_P_btm.n556 0.09425
R30897 C10_P_btm.n761 C10_P_btm.n555 0.09425
R30898 C10_P_btm.n761 C10_P_btm.n557 0.09425
R30899 C10_P_btm.n764 C10_P_btm.n763 0.09425
R30900 C10_P_btm.n763 C10_P_btm.n762 0.09425
R30901 C10_P_btm.n766 C10_P_btm.n765 0.09425
R30902 C10_P_btm.n765 C10_P_btm.n555 0.09425
R30903 C10_P_btm.n768 C10_P_btm.n767 0.09425
R30904 C10_P_btm.n767 C10_P_btm.n554 0.09425
R30905 C10_P_btm.n769 C10_P_btm.n552 0.09425
R30906 C10_P_btm.n770 C10_P_btm.n551 0.09425
R30907 C10_P_btm.n567 C10_P_btm.n551 0.09425
R30908 C10_P_btm.n772 C10_P_btm.n771 0.09425
R30909 C10_P_btm.n773 C10_P_btm.n548 0.09425
R30910 C10_P_btm.n773 C10_P_btm.n549 0.09425
R30911 C10_P_btm.n774 C10_P_btm.n545 0.09425
R30912 C10_P_btm.n776 C10_P_btm.n775 0.09425
R30913 C10_P_btm.n775 C10_P_btm.n546 0.09425
R30914 C10_P_btm.n777 C10_P_btm.n544 0.09425
R30915 C10_P_btm.n778 C10_P_btm.n543 0.09425
R30916 C10_P_btm.n580 C10_P_btm.n543 0.09425
R30917 C10_P_btm.n780 C10_P_btm.n779 0.09425
R30918 C10_P_btm.n781 C10_P_btm.n540 0.09425
R30919 C10_P_btm.n781 C10_P_btm.n541 0.09425
R30920 C10_P_btm.n782 C10_P_btm.n537 0.09425
R30921 C10_P_btm.n784 C10_P_btm.n783 0.09425
R30922 C10_P_btm.n783 C10_P_btm.n538 0.09425
R30923 C10_P_btm.n591 C10_P_btm.n536 0.09425
R30924 C10_P_btm.n592 C10_P_btm.n591 0.09425
R30925 C10_P_btm.n695 C10_P_btm.n535 0.09425
R30926 C10_P_btm.n695 C10_P_btm.n593 0.09425
R30927 C10_P_btm.n696 C10_P_btm.n596 0.09425
R30928 C10_P_btm.n738 C10_P_btm.n596 0.09425
R30929 C10_P_btm.n694 C10_P_btm.n597 0.09425
R30930 C10_P_btm.n736 C10_P_btm.n597 0.09425
R30931 C10_P_btm.n691 C10_P_btm.n599 0.09425
R30932 C10_P_btm.n600 C10_P_btm.n599 0.09425
R30933 C10_P_btm.n711 C10_P_btm.n710 0.09425
R30934 C10_P_btm.n711 C10_P_btm.n603 0.09425
R30935 C10_P_btm.n713 C10_P_btm.n712 0.09425
R30936 C10_P_btm.n712 C10_P_btm.n680 0.09425
R30937 C10_P_btm.n727 C10_P_btm.n682 0.09425
R30938 C10_P_btm.n728 C10_P_btm.n727 0.09425
R30939 C10_P_btm.n726 C10_P_btm.n681 0.09425
R30940 C10_P_btm.n684 C10_P_btm.n470 0.09425
R30941 C10_P_btm.n822 C10_P_btm.n470 0.09425
R30942 C10_P_btm.n821 C10_P_btm.n820 0.09425
R30943 C10_P_btm.n821 C10_P_btm.n469 0.09425
R30944 C10_P_btm.n823 C10_P_btm.n822 0.09425
R30945 C10_P_btm.n824 C10_P_btm.n823 0.09425
R30946 C10_P_btm.n825 C10_P_btm.n469 0.09425
R30947 C10_P_btm.n825 C10_P_btm.n442 0.09425
R30948 C10_P_btm.n824 C10_P_btm.n441 0.09425
R30949 C10_P_btm.n844 C10_P_btm.n441 0.09425
R30950 C10_P_btm.n843 C10_P_btm.n442 0.09425
R30951 C10_P_btm.n843 C10_P_btm.n440 0.09425
R30952 C10_P_btm.n845 C10_P_btm.n844 0.09425
R30953 C10_P_btm.n865 C10_P_btm.n845 0.09425
R30954 C10_P_btm.n866 C10_P_btm.n440 0.09425
R30955 C10_P_btm.n866 C10_P_btm.n438 0.09425
R30956 C10_P_btm.n865 C10_P_btm.n864 0.09425
R30957 C10_P_btm.n864 C10_P_btm.n863 0.09425
R30958 C10_P_btm.n846 C10_P_btm.n438 0.09425
R30959 C10_P_btm.n861 C10_P_btm.n846 0.09425
R30960 C10_P_btm.n863 C10_P_btm.n862 0.09425
R30961 C10_P_btm.n861 C10_P_btm.n860 0.09425
R30962 C10_P_btm.n851 C10_P_btm.n850 0.09425
R30963 C10_P_btm.n850 C10_P_btm.n414 0.09425
R30964 C10_P_btm.n849 C10_P_btm.n415 0.09425
R30965 C10_P_btm.n885 C10_P_btm.n415 0.09425
R30966 C10_P_btm.n886 C10_P_btm.n414 0.09425
R30967 C10_P_btm.n887 C10_P_btm.n886 0.09425
R30968 C10_P_btm.n885 C10_P_btm.n413 0.09425
R30969 C10_P_btm.n939 C10_P_btm.n413 0.09425
R30970 C10_P_btm.n888 C10_P_btm.n887 0.09425
R30971 C10_P_btm.n937 C10_P_btm.n888 0.09425
R30972 C10_P_btm.n939 C10_P_btm.n938 0.09425
R30973 C10_P_btm.n938 C10_P_btm.n889 0.09425
R30974 C10_P_btm.n937 C10_P_btm.n936 0.09425
R30975 C10_P_btm.n936 C10_P_btm.n935 0.09425
R30976 C10_P_btm.n890 C10_P_btm.n889 0.09425
R30977 C10_P_btm.n933 C10_P_btm.n890 0.09425
R30978 C10_P_btm.n935 C10_P_btm.n934 0.09425
R30979 C10_P_btm.n934 C10_P_btm.n891 0.09425
R30980 C10_P_btm.n933 C10_P_btm.n932 0.09425
R30981 C10_P_btm.n932 C10_P_btm.n893 0.09425
R30982 C10_P_btm.n900 C10_P_btm.n891 0.09425
R30983 C10_P_btm.n917 C10_P_btm.n900 0.09425
R30984 C10_P_btm.n918 C10_P_btm.n893 0.09425
R30985 C10_P_btm.n918 C10_P_btm.n899 0.09425
R30986 C10_P_btm.n917 C10_P_btm.n916 0.09425
R30987 C10_P_btm.n916 C10_P_btm.n915 0.09425
R30988 C10_P_btm.n901 C10_P_btm.n899 0.09425
R30989 C10_P_btm.n913 C10_P_btm.n901 0.09425
R30990 C10_P_btm.n915 C10_P_btm.n914 0.09425
R30991 C10_P_btm.n914 C10_P_btm.n902 0.09425
R30992 C10_P_btm.n913 C10_P_btm.n912 0.09425
R30993 C10_P_btm.n912 C10_P_btm.n910 0.09425
R30994 C10_P_btm.n909 C10_P_btm.n902 0.09425
R30995 C10_P_btm.n964 C10_P_btm.n373 0.09425
R30996 C10_P_btm.n964 C10_P_btm.n371 0.09425
R30997 C10_P_btm.n966 C10_P_btm.n965 0.09425
R30998 C10_P_btm.n989 C10_P_btm.n966 0.09425
R30999 C10_P_btm.n990 C10_P_btm.n371 0.09425
R31000 C10_P_btm.n990 C10_P_btm.n369 0.09425
R31001 C10_P_btm.n989 C10_P_btm.n988 0.09425
R31002 C10_P_btm.n988 C10_P_btm.n987 0.09425
R31003 C10_P_btm.n967 C10_P_btm.n369 0.09425
R31004 C10_P_btm.n985 C10_P_btm.n967 0.09425
R31005 C10_P_btm.n987 C10_P_btm.n986 0.09425
R31006 C10_P_btm.n986 C10_P_btm.n968 0.09425
R31007 C10_P_btm.n985 C10_P_btm.n984 0.09425
R31008 C10_P_btm.n984 C10_P_btm.n970 0.09425
R31009 C10_P_btm.n971 C10_P_btm.n968 0.09425
R31010 C10_P_btm.n973 C10_P_btm.n971 0.09425
R31011 C10_P_btm.n974 C10_P_btm.n970 0.09425
R31012 C10_P_btm.n974 C10_P_btm.n69 0.09425
R31013 C10_P_btm.n973 C10_P_btm.n972 0.09425
R31014 C10_P_btm.n972 C10_P_btm.n65 0.09425
R31015 C10_P_btm.n1010 C10_P_btm.n69 0.09425
R31016 C10_P_btm.n1011 C10_P_btm.n1010 0.09425
R31017 C10_P_btm.n1012 C10_P_btm.n65 0.09425
R31018 C10_P_btm.n1012 C10_P_btm.n66 0.09425
R31019 C10_P_btm.n1013 C10_P_btm.n64 0.09425
R31020 C10_P_btm.n85 C10_P_btm.n64 0.09425
R31021 C10_P_btm.n1015 C10_P_btm.n1014 0.09425
R31022 C10_P_btm.n1016 C10_P_btm.n61 0.09425
R31023 C10_P_btm.n1016 C10_P_btm.n62 0.09425
R31024 C10_P_btm.n1017 C10_P_btm.n58 0.09425
R31025 C10_P_btm.n1019 C10_P_btm.n1018 0.09425
R31026 C10_P_btm.n1018 C10_P_btm.n59 0.09425
R31027 C10_P_btm.n1020 C10_P_btm.n57 0.09425
R31028 C10_P_btm.n1021 C10_P_btm.n56 0.09425
R31029 C10_P_btm.n335 C10_P_btm.n56 0.09425
R31030 C10_P_btm.n1023 C10_P_btm.n1022 0.09425
R31031 C10_P_btm.n1024 C10_P_btm.n53 0.09425
R31032 C10_P_btm.n1024 C10_P_btm.n54 0.09425
R31033 C10_P_btm.n1025 C10_P_btm.n50 0.09425
R31034 C10_P_btm.n1027 C10_P_btm.n1026 0.09425
R31035 C10_P_btm.n1026 C10_P_btm.n51 0.09425
R31036 C10_P_btm.n1028 C10_P_btm.n49 0.09425
R31037 C10_P_btm.n1029 C10_P_btm.n48 0.09425
R31038 C10_P_btm.n327 C10_P_btm.n48 0.09425
R31039 C10_P_btm.n1031 C10_P_btm.n1030 0.09425
R31040 C10_P_btm.n1032 C10_P_btm.n45 0.09425
R31041 C10_P_btm.n1032 C10_P_btm.n46 0.09425
R31042 C10_P_btm.n1033 C10_P_btm.n42 0.09425
R31043 C10_P_btm.n1035 C10_P_btm.n1034 0.09425
R31044 C10_P_btm.n1034 C10_P_btm.n43 0.09425
R31045 C10_P_btm.n1036 C10_P_btm.n41 0.09425
R31046 C10_P_btm.n1037 C10_P_btm.n40 0.09425
R31047 C10_P_btm.n319 C10_P_btm.n40 0.09425
R31048 C10_P_btm.n1039 C10_P_btm.n1038 0.09425
R31049 C10_P_btm.n1040 C10_P_btm.n37 0.09425
R31050 C10_P_btm.n1040 C10_P_btm.n38 0.09425
R31051 C10_P_btm.n1041 C10_P_btm.n34 0.09425
R31052 C10_P_btm.n1043 C10_P_btm.n1042 0.09425
R31053 C10_P_btm.n1042 C10_P_btm.n35 0.09425
R31054 C10_P_btm.n1044 C10_P_btm.n33 0.09425
R31055 C10_P_btm.n851 C10_P_btm.n847 0.047875
R31056 C10_P_btm.n909 C10_P_btm.n372 0.047875
R31057 C10_P_btm.n131 C10_P_btm.n130 0.0342289
R31058 C10_P_btm.n518 C10_P_btm.n500 0.0342289
R31059 C10_P_btm.n653 C10_P_btm.n624 0.0342289
R31060 C10_P_btm.n860 C10_P_btm.n847 0.0342289
R31061 C10_P_btm.n266 C10_P_btm.n174 0.0342289
R31062 C10_P_btm.n766 C10_P_btm.n553 0.0342289
R31063 C10_P_btm.n373 C10_P_btm.n372 0.0342289
R31064 EN_VIN_BSTR_P.n20 EN_VIN_BSTR_P.t11 1559.46
R31065 EN_VIN_BSTR_P.n19 EN_VIN_BSTR_P.t18 1415.15
R31066 EN_VIN_BSTR_P.n19 EN_VIN_BSTR_P.t9 1320.68
R31067 EN_VIN_BSTR_P.n2 EN_VIN_BSTR_P.t16 748.122
R31068 EN_VIN_BSTR_P.n2 EN_VIN_BSTR_P.t7 678.014
R31069 EN_VIN_BSTR_P.n11 EN_VIN_BSTR_P.t12 605.802
R31070 EN_VIN_BSTR_P.n10 EN_VIN_BSTR_P.t8 444.502
R31071 EN_VIN_BSTR_P.n3 EN_VIN_BSTR_P.t10 398.575
R31072 EN_VIN_BSTR_P.n9 EN_VIN_BSTR_P.t17 382.812
R31073 EN_VIN_BSTR_P.n17 EN_VIN_BSTR_P.t20 381.798
R31074 EN_VIN_BSTR_P.n9 EN_VIN_BSTR_P.t21 381.793
R31075 EN_VIN_BSTR_P.n16 EN_VIN_BSTR_P.t23 381.788
R31076 EN_VIN_BSTR_P.n15 EN_VIN_BSTR_P.t14 381.413
R31077 EN_VIN_BSTR_P.n14 EN_VIN_BSTR_P.t22 381.413
R31078 EN_VIN_BSTR_P.n13 EN_VIN_BSTR_P.t13 381.413
R31079 EN_VIN_BSTR_P.n12 EN_VIN_BSTR_P.t19 381.413
R31080 EN_VIN_BSTR_P.n10 EN_VIN_BSTR_P.t15 356.68
R31081 EN_VIN_BSTR_P.n3 EN_VIN_BSTR_P.n2 176.945
R31082 EN_VIN_BSTR_P.n11 EN_VIN_BSTR_P.n10 161.768
R31083 EN_VIN_BSTR_P.n20 EN_VIN_BSTR_P.n19 161.3
R31084 EN_VIN_BSTR_P.n4 EN_VIN_BSTR_P.n1 56.3527
R31085 EN_VIN_BSTR_P.n5 EN_VIN_BSTR_P.n0 56.3527
R31086 EN_VIN_BSTR_P.n21 EN_VIN_BSTR_P.n18 28.2777
R31087 EN_VIN_BSTR_P EN_VIN_BSTR_P.n21 26.0445
R31088 EN_VIN_BSTR_P.n6 EN_VIN_BSTR_P.t0 24.8352
R31089 EN_VIN_BSTR_P.n6 EN_VIN_BSTR_P.t1 24.1869
R31090 EN_VIN_BSTR_P.n7 EN_VIN_BSTR_P.t2 24.1612
R31091 EN_VIN_BSTR_P.n1 EN_VIN_BSTR_P.t3 8.12675
R31092 EN_VIN_BSTR_P.n1 EN_VIN_BSTR_P.t4 8.12675
R31093 EN_VIN_BSTR_P.n0 EN_VIN_BSTR_P.t6 8.12675
R31094 EN_VIN_BSTR_P.n0 EN_VIN_BSTR_P.t5 8.12675
R31095 EN_VIN_BSTR_P.n21 EN_VIN_BSTR_P.n20 4.51508
R31096 EN_VIN_BSTR_P EN_VIN_BSTR_P.n8 4.04813
R31097 EN_VIN_BSTR_P.n4 EN_VIN_BSTR_P.n3 2.39112
R31098 EN_VIN_BSTR_P.n8 EN_VIN_BSTR_P.n5 1.18584
R31099 EN_VIN_BSTR_P.n7 EN_VIN_BSTR_P.n6 0.989971
R31100 EN_VIN_BSTR_P.n17 EN_VIN_BSTR_P.n16 0.9005
R31101 EN_VIN_BSTR_P.n18 EN_VIN_BSTR_P.n17 0.7005
R31102 EN_VIN_BSTR_P.n13 EN_VIN_BSTR_P.n12 0.512318
R31103 EN_VIN_BSTR_P.n14 EN_VIN_BSTR_P.n13 0.512318
R31104 EN_VIN_BSTR_P.n15 EN_VIN_BSTR_P.n14 0.512318
R31105 EN_VIN_BSTR_P.n5 EN_VIN_BSTR_P.n4 0.462038
R31106 EN_VIN_BSTR_P.n18 EN_VIN_BSTR_P.n9 0.3755
R31107 EN_VIN_BSTR_P.n12 EN_VIN_BSTR_P.n11 0.267318
R31108 EN_VIN_BSTR_P.n16 EN_VIN_BSTR_P.n15 0.138909
R31109 EN_VIN_BSTR_P.n8 EN_VIN_BSTR_P.n7 0.018
R31110 w_1575_34786.n57 w_1575_34786.n10 15667.1
R31111 w_1575_34786.n43 w_1575_34786.n10 15667.1
R31112 w_1575_34786.n43 w_1575_34786.n41 15667.1
R31113 w_1575_34786.n41 w_1575_34786.n40 12324.7
R31114 w_1575_34786.n8 w_1575_34786.n6 3017.65
R31115 w_1575_34786.n61 w_1575_34786.n5 3017.65
R31116 w_1575_34786.n61 w_1575_34786.n6 3017.65
R31117 w_1575_34786.n40 w_1575_34786.n9 1757.65
R31118 w_1575_34786.n33 w_1575_34786.n26 1757.65
R31119 w_1575_34786.n44 w_1575_34786.n12 1671.15
R31120 w_1575_34786.n45 w_1575_34786.n25 1494.32
R31121 w_1575_34786.n57 w_1575_34786.n9 1464.71
R31122 w_1575_34786.n26 w_1575_34786.n5 1080
R31123 w_1575_34786.n56 w_1575_34786.n55 965.508
R31124 w_1575_34786.n39 w_1575_34786.t8 905.04
R31125 w_1575_34786.n43 w_1575_34786.t13 849.226
R31126 w_1575_34786.n58 w_1575_34786.t10 842.11
R31127 w_1575_34786.t8 w_1575_34786.n7 812.54
R31128 w_1575_34786.t13 w_1575_34786.n42 788.865
R31129 w_1575_34786.n42 w_1575_34786.t10 788.865
R31130 w_1575_34786.n27 w_1575_34786.n25 693.082
R31131 w_1575_34786.n55 w_1575_34786.n12 673.732
R31132 w_1575_34786.n28 w_1575_34786.n27 621.553
R31133 w_1575_34786.n34 w_1575_34786.n9 557.648
R31134 w_1575_34786.n34 w_1575_34786.n33 557.648
R31135 w_1575_34786.n40 w_1575_34786.n39 557.648
R31136 w_1575_34786.n39 w_1575_34786.n26 557.648
R31137 w_1575_34786.n32 w_1575_34786.n3 298.877
R31138 w_1575_34786.n30 w_1575_34786.n4 280.202
R31139 w_1575_34786.n63 w_1575_34786.n62 277.776
R31140 w_1575_34786.n17 w_1575_34786.t9 228.215
R31141 w_1575_34786.n28 w_1575_34786.n11 187.482
R31142 w_1575_34786.n37 w_1575_34786.n36 187.482
R31143 w_1575_34786.n45 w_1575_34786.n44 169.53
R31144 w_1575_34786.n56 w_1575_34786.n11 156.236
R31145 w_1575_34786.n61 w_1575_34786.t4 137.529
R31146 w_1575_34786.n37 w_1575_34786.n31 115.201
R31147 w_1575_34786.n59 w_1575_34786.n7 103.859
R31148 w_1575_34786.n39 w_1575_34786.n38 92.5005
R31149 w_1575_34786.n35 w_1575_34786.n34 92.5005
R31150 w_1575_34786.n34 w_1575_34786.n7 92.5005
R31151 w_1575_34786.t0 w_1575_34786.n59 75.2024
R31152 w_1575_34786.t2 w_1575_34786.t0 73.6677
R31153 w_1575_34786.t4 w_1575_34786.t6 73.6677
R31154 w_1575_34786.n52 w_1575_34786.t12 67.9353
R31155 w_1575_34786.t15 w_1575_34786.n49 67.9353
R31156 w_1575_34786.n21 w_1575_34786.t17 67.9353
R31157 w_1575_34786.n24 w_1575_34786.t14 67.9353
R31158 w_1575_34786.n68 w_1575_34786.t5 65.4041
R31159 w_1575_34786.n66 w_1575_34786.t1 62.5643
R31160 w_1575_34786.n33 w_1575_34786.n8 60.0005
R31161 w_1575_34786.n51 w_1575_34786.n50 59.5338
R31162 w_1575_34786.n23 w_1575_34786.n22 59.5338
R31163 w_1575_34786.n38 w_1575_34786.n28 59.4829
R31164 w_1575_34786.n38 w_1575_34786.n37 59.4829
R31165 w_1575_34786.n35 w_1575_34786.n11 59.4829
R31166 w_1575_34786.n36 w_1575_34786.n35 59.4829
R31167 w_1575_34786.n69 w_1575_34786.n68 56.8163
R31168 w_1575_34786.n60 w_1575_34786.t2 36.8341
R31169 w_1575_34786.t6 w_1575_34786.n60 36.8341
R31170 w_1575_34786.n59 w_1575_34786.n58 35.2823
R31171 w_1575_34786.n6 w_1575_34786.n3 26.4291
R31172 w_1575_34786.n60 w_1575_34786.n6 26.4291
R31173 w_1575_34786.n31 w_1575_34786.n5 26.4291
R31174 w_1575_34786.n60 w_1575_34786.n5 26.4291
R31175 w_1575_34786.n62 w_1575_34786.n4 20.4805
R31176 w_1575_34786.n31 w_1575_34786.n30 16.9417
R31177 w_1575_34786.n19 w_1575_34786.n18 15.2505
R31178 w_1575_34786.n62 w_1575_34786.n61 13.2148
R31179 w_1575_34786.n32 w_1575_34786.n8 13.2148
R31180 w_1575_34786.n59 w_1575_34786.n8 13.2148
R31181 w_1575_34786.n50 w_1575_34786.t15 8.40197
R31182 w_1575_34786.n50 w_1575_34786.t11 8.40197
R31183 w_1575_34786.t14 w_1575_34786.n23 8.40197
R31184 w_1575_34786.n23 w_1575_34786.t16 8.40197
R31185 w_1575_34786.n63 w_1575_34786.n3 8.2968
R31186 w_1575_34786.n69 w_1575_34786.t3 8.12675
R31187 w_1575_34786.t7 w_1575_34786.n69 8.12675
R31188 w_1575_34786.n47 w_1575_34786.n13 7.19895
R31189 w_1575_34786.n57 w_1575_34786.n56 7.11588
R31190 w_1575_34786.n58 w_1575_34786.n57 7.11588
R31191 w_1575_34786.n44 w_1575_34786.n43 7.11588
R31192 w_1575_34786.n54 w_1575_34786.n48 7.06493
R31193 w_1575_34786.n36 w_1575_34786.n32 6.4005
R31194 w_1575_34786.n68 w_1575_34786.n67 2.72081
R31195 w_1575_34786.n54 w_1575_34786.n53 2.33582
R31196 w_1575_34786.n14 w_1575_34786.n13 2.12421
R31197 w_1575_34786.n41 w_1575_34786.n25 1.8505
R31198 w_1575_34786.n42 w_1575_34786.n41 1.8505
R31199 w_1575_34786.n12 w_1575_34786.n10 1.8505
R31200 w_1575_34786.n42 w_1575_34786.n10 1.8505
R31201 w_1575_34786.n64 w_1575_34786.n63 1.5505
R31202 w_1575_34786.n30 w_1575_34786.n29 1.5505
R31203 w_1575_34786.n64 w_1575_34786.n2 1.26141
R31204 w_1575_34786.n4 w_1575_34786.n2 1.03383
R31205 w_1575_34786.n46 w_1575_34786.n45 1.03383
R31206 w_1575_34786.n16 w_1575_34786.n11 1.03383
R31207 w_1575_34786.n66 w_1575_34786.n65 1.00774
R31208 w_1575_34786.n24 w_1575_34786.n22 0.984766
R31209 w_1575_34786.n22 w_1575_34786.n21 0.984766
R31210 w_1575_34786.n51 w_1575_34786.n49 0.984766
R31211 w_1575_34786.n52 w_1575_34786.n51 0.984766
R31212 w_1575_34786.n29 w_1575_34786.n2 0.938644
R31213 w_1575_34786.n48 w_1575_34786.n47 0.741479
R31214 w_1575_34786.n65 w_1575_34786.n64 0.542875
R31215 w_1575_34786.n14 w_1575_34786.n0 0.494823
R31216 w_1575_34786.n29 w_1575_34786.n0 0.441222
R31217 w_1575_34786.n67 w_1575_34786.n0 0.428803
R31218 w_1575_34786.n19 w_1575_34786.n1 0.286876
R31219 w_1575_34786.n53 w_1575_34786.n1 0.260002
R31220 w_1575_34786.n15 w_1575_34786.n14 0.253077
R31221 w_1575_34786.n27 w_1575_34786.n13 0.227329
R31222 w_1575_34786.n55 w_1575_34786.n54 0.227329
R31223 w_1575_34786.n65 w_1575_34786.n1 0.19304
R31224 w_1575_34786.n20 w_1575_34786.n19 0.178335
R31225 w_1575_34786.n18 w_1575_34786.n17 0.0711522
R31226 w_1575_34786.n20 w_1575_34786.n15 0.0700876
R31227 w_1575_34786.n67 w_1575_34786.n66 0.057539
R31228 w_1575_34786.n49 w_1575_34786.n48 0.0345909
R31229 w_1575_34786.n46 w_1575_34786.n24 0.0334254
R31230 w_1575_34786.n53 w_1575_34786.n52 0.0333453
R31231 w_1575_34786.n21 w_1575_34786.n20 0.0328427
R31232 w_1575_34786.n17 w_1575_34786.n15 0.0303913
R31233 w_1575_34786.n18 w_1575_34786.n16 0.0136119
R31234 w_1575_34786.n47 w_1575_34786.n46 0.0016655
R31235 w_1575_34786.n20 w_1575_34786.n16 0.00137413
R31236 a_10341_43396.t0 a_10341_43396.n1 463.529
R31237 a_10341_43396.n0 a_10341_43396.t3 276.464
R31238 a_10341_43396.n1 a_10341_43396.t1 254.047
R31239 a_10341_43396.n1 a_10341_43396.n0 197.768
R31240 a_10341_43396.n0 a_10341_43396.t2 196.131
R31241 a_n4209_38502.n4 a_n4209_38502.t9 553.635
R31242 a_n4209_38502.n7 a_n4209_38502.n6 340.637
R31243 a_n4209_38502.n3 a_n4209_38502.t8 241.536
R31244 a_n4209_38502.n8 a_n4209_38502.n7 195.577
R31245 a_n4209_38502.n4 a_n4209_38502.n3 173.952
R31246 a_n4209_38502.n3 a_n4209_38502.t10 169.237
R31247 a_n4209_38502.n2 a_n4209_38502.n0 137.189
R31248 a_n4209_38502.n2 a_n4209_38502.n1 98.788
R31249 a_n4209_38502.n7 a_n4209_38502.n5 37.1695
R31250 a_n4209_38502.n5 a_n4209_38502.n2 27.8375
R31251 a_n4209_38502.n6 a_n4209_38502.t2 26.5955
R31252 a_n4209_38502.n6 a_n4209_38502.t1 26.5955
R31253 a_n4209_38502.t3 a_n4209_38502.n8 26.5955
R31254 a_n4209_38502.n8 a_n4209_38502.t0 26.5955
R31255 a_n4209_38502.n0 a_n4209_38502.t7 24.9236
R31256 a_n4209_38502.n0 a_n4209_38502.t4 24.9236
R31257 a_n4209_38502.n1 a_n4209_38502.t6 24.9236
R31258 a_n4209_38502.n1 a_n4209_38502.t5 24.9236
R31259 a_n4209_38502.n5 a_n4209_38502.n4 9.30997
R31260 a_13887_32519.n1 a_13887_32519.t4 676.072
R31261 a_13887_32519.n2 a_13887_32519.n1 380.32
R31262 a_13887_32519.n1 a_13887_32519.n0 185
R31263 a_13887_32519.n2 a_13887_32519.t0 26.5955
R31264 a_13887_32519.t1 a_13887_32519.n2 26.5955
R31265 a_13887_32519.n0 a_13887_32519.t2 24.9236
R31266 a_13887_32519.n0 a_13887_32519.t3 24.9236
R31267 a_n881_46662.n21 a_n881_46662.n20 659.109
R31268 a_n881_46662.n2 a_n881_46662.t16 261.887
R31269 a_n881_46662.n16 a_n881_46662.t22 261.887
R31270 a_n881_46662.n14 a_n881_46662.t6 261.887
R31271 a_n881_46662.n11 a_n881_46662.t14 261.887
R31272 a_n881_46662.n4 a_n881_46662.t5 261.887
R31273 a_n881_46662.n6 a_n881_46662.t20 261.887
R31274 a_n881_46662.n5 a_n881_46662.t13 261.887
R31275 a_n881_46662.n3 a_n881_46662.t18 261.887
R31276 a_n881_46662.n8 a_n881_46662.t21 241.536
R31277 a_n881_46662.n1 a_n881_46662.t19 239.505
R31278 a_n881_46662.n20 a_n881_46662.n0 219.663
R31279 a_n881_46662.n9 a_n881_46662.n8 179.173
R31280 a_n881_46662.n19 a_n881_46662.n1 175.8
R31281 a_n881_46662.n7 a_n881_46662.n6 175.201
R31282 a_n881_46662.n7 a_n881_46662.n5 172.376
R31283 a_n881_46662.n13 a_n881_46662.n3 169.52
R31284 a_n881_46662.n8 a_n881_46662.t23 169.237
R31285 a_n881_46662.n1 a_n881_46662.t7 167.204
R31286 a_n881_46662.n18 a_n881_46662.n2 162.429
R31287 a_n881_46662.n17 a_n881_46662.n16 162.429
R31288 a_n881_46662.n15 a_n881_46662.n14 162.429
R31289 a_n881_46662.n12 a_n881_46662.n11 162.429
R31290 a_n881_46662.n10 a_n881_46662.n4 162.429
R31291 a_n881_46662.n2 a_n881_46662.t11 155.847
R31292 a_n881_46662.n16 a_n881_46662.t9 155.847
R31293 a_n881_46662.n14 a_n881_46662.t12 155.847
R31294 a_n881_46662.n11 a_n881_46662.t4 155.847
R31295 a_n881_46662.n4 a_n881_46662.t8 155.847
R31296 a_n881_46662.n6 a_n881_46662.t15 155.847
R31297 a_n881_46662.n5 a_n881_46662.t10 155.847
R31298 a_n881_46662.n3 a_n881_46662.t17 155.847
R31299 a_n881_46662.n0 a_n881_46662.t3 38.5719
R31300 a_n881_46662.n0 a_n881_46662.t2 38.5719
R31301 a_n881_46662.n19 a_n881_46662.n18 33.6375
R31302 a_n881_46662.n12 a_n881_46662.n10 28.8638
R31303 a_n881_46662.n21 a_n881_46662.t0 26.5955
R31304 a_n881_46662.t1 a_n881_46662.n21 26.5955
R31305 a_n881_46662.n15 a_n881_46662.n13 26.5513
R31306 a_n881_46662.n10 a_n881_46662.n9 10.3151
R31307 a_n881_46662.n13 a_n881_46662.n12 10.2972
R31308 a_n881_46662.n9 a_n881_46662.n7 9.87017
R31309 a_n881_46662.n20 a_n881_46662.n19 9.3005
R31310 a_n881_46662.n17 a_n881_46662.n15 8.50891
R31311 a_n881_46662.n18 a_n881_46662.n17 5.23847
R31312 a_4791_45118.n19 a_4791_45118.n18 620.708
R31313 a_4791_45118.n8 a_4791_45118.n6 459.668
R31314 a_4791_45118.n3 a_4791_45118.n1 459.668
R31315 a_4791_45118.n9 a_4791_45118.t5 382.425
R31316 a_4791_45118.t5 a_4791_45118.t14 378.255
R31317 a_4791_45118.n7 a_4791_45118.t9 329.902
R31318 a_4791_45118.n2 a_4791_45118.t17 329.902
R31319 a_4791_45118.n6 a_4791_45118.t8 272.062
R31320 a_4791_45118.n1 a_4791_45118.t20 272.062
R31321 a_4791_45118.n18 a_4791_45118.n0 258.063
R31322 a_4791_45118.n15 a_4791_45118.t11 231.835
R31323 a_4791_45118.n5 a_4791_45118.t12 212.081
R31324 a_4791_45118.n4 a_4791_45118.t16 212.081
R31325 a_4791_45118.n6 a_4791_45118.t22 206.19
R31326 a_4791_45118.n1 a_4791_45118.t21 206.19
R31327 a_4791_45118.n14 a_4791_45118.t7 201.369
R31328 a_4791_45118.n10 a_4791_45118.n5 194.209
R31329 a_4791_45118.n16 a_4791_45118.n14 180.572
R31330 a_4791_45118.n13 a_4791_45118.n12 171.97
R31331 a_4791_45118.n16 a_4791_45118.n15 170.369
R31332 a_4791_45118.n15 a_4791_45118.t15 157.07
R31333 a_4791_45118.n8 a_4791_45118.n7 152
R31334 a_4791_45118.n3 a_4791_45118.n2 152
R31335 a_4791_45118.n7 a_4791_45118.t4 148.35
R31336 a_4791_45118.n2 a_4791_45118.t10 148.35
R31337 a_4791_45118.n5 a_4791_45118.t13 139.78
R31338 a_4791_45118.n4 a_4791_45118.t23 139.78
R31339 a_4791_45118.n12 a_4791_45118.t19 137.177
R31340 a_4791_45118.n14 a_4791_45118.t6 132.282
R31341 a_4791_45118.n12 a_4791_45118.t18 121.109
R31342 a_4791_45118.n5 a_4791_45118.n4 61.346
R31343 a_4791_45118.n0 a_4791_45118.t2 38.5719
R31344 a_4791_45118.n0 a_4791_45118.t3 38.5719
R31345 a_4791_45118.n19 a_4791_45118.t0 26.5955
R31346 a_4791_45118.t1 a_4791_45118.n19 26.5955
R31347 a_4791_45118.n9 a_4791_45118.n8 23.4916
R31348 a_4791_45118.n11 a_4791_45118.n3 23.3393
R31349 a_4791_45118.n18 a_4791_45118.n17 14.5053
R31350 a_4791_45118.n17 a_4791_45118.n16 11.1935
R31351 a_4791_45118.n13 a_4791_45118.n11 8.4824
R31352 a_4791_45118.n11 a_4791_45118.n10 6.89885
R31353 a_4791_45118.n17 a_4791_45118.n13 5.53876
R31354 a_4791_45118.n10 a_4791_45118.n9 0.755995
R31355 a_n3674_39768.n3 a_n3674_39768.n2 296.139
R31356 a_n3674_39768.n2 a_n3674_39768.n0 269.182
R31357 a_n3674_39768.n1 a_n3674_39768.t5 235.821
R31358 a_n3674_39768.n2 a_n3674_39768.n1 227.056
R31359 a_n3674_39768.n1 a_n3674_39768.t4 163.52
R31360 a_n3674_39768.n3 a_n3674_39768.t0 26.5955
R31361 a_n3674_39768.t1 a_n3674_39768.n3 26.5955
R31362 a_n3674_39768.n0 a_n3674_39768.t2 24.9236
R31363 a_n3674_39768.n0 a_n3674_39768.t3 24.9236
R31364 a_10809_44734.n0 a_10809_44734.t4 276.464
R31365 a_10809_44734.n1 a_10809_44734.t5 230.155
R31366 a_10809_44734.n4 a_10809_44734.n3 207.219
R31367 a_10809_44734.n2 a_10809_44734.n0 200.749
R31368 a_10809_44734.n0 a_10809_44734.t6 196.131
R31369 a_10809_44734.n3 a_10809_44734.t2 183.06
R31370 a_10809_44734.n2 a_10809_44734.n1 163.605
R31371 a_10809_44734.n1 a_10809_44734.t3 157.856
R31372 a_10809_44734.n3 a_10809_44734.n2 36.5845
R31373 a_10809_44734.n4 a_10809_44734.t1 26.5955
R31374 a_10809_44734.t0 a_10809_44734.n4 26.5955
R31375 a_n2661_42834.n0 a_n2661_42834.t3 276.464
R31376 a_n2661_42834.n2 a_n2661_42834.n1 259.06
R31377 a_n2661_42834.n1 a_n2661_42834.n0 206.895
R31378 a_n2661_42834.n0 a_n2661_42834.t4 196.131
R31379 a_n2661_42834.n1 a_n2661_42834.t1 131.308
R31380 a_n2661_42834.t0 a_n2661_42834.n2 26.5955
R31381 a_n2661_42834.n2 a_n2661_42834.t2 26.5955
R31382 a_n743_46660.n6 a_n743_46660.t4 471.289
R31383 a_n743_46660.n5 a_n743_46660.t3 471.289
R31384 a_n743_46660.n0 a_n743_46660.t8 471.289
R31385 a_n743_46660.t0 a_n743_46660.n9 414.534
R31386 a_n743_46660.n3 a_n743_46660.t5 414.432
R31387 a_n743_46660.n3 a_n743_46660.t7 300.349
R31388 a_n743_46660.n9 a_n743_46660.t1 273.178
R31389 a_n743_46660.n1 a_n743_46660.t9 230.155
R31390 a_n743_46660.n2 a_n743_46660.n0 189.501
R31391 a_n743_46660.n7 a_n743_46660.n5 186.798
R31392 a_n743_46660.n7 a_n743_46660.n6 183.177
R31393 a_n743_46660.n2 a_n743_46660.n1 171.56
R31394 a_n743_46660.n1 a_n743_46660.t11 157.856
R31395 a_n743_46660.n6 a_n743_46660.t6 148.35
R31396 a_n743_46660.n5 a_n743_46660.t10 148.35
R31397 a_n743_46660.n0 a_n743_46660.t2 148.35
R31398 a_n743_46660.n9 a_n743_46660.n8 23.9092
R31399 a_n743_46660.n4 a_n743_46660.n3 18.2969
R31400 a_n743_46660.n8 a_n743_46660.n4 10.8778
R31401 a_n743_46660.n4 a_n743_46660.n2 8.73873
R31402 a_n743_46660.n8 a_n743_46660.n7 7.65435
R31403 a_1606_42308.n2 a_1606_42308.t7 579.59
R31404 a_1606_42308.n2 a_1606_42308.t5 579.311
R31405 a_1606_42308.n5 a_1606_42308.n4 287.752
R31406 a_1606_42308.n4 a_1606_42308.n0 277.568
R31407 a_1606_42308.n1 a_1606_42308.t4 260.322
R31408 a_1606_42308.n1 a_1606_42308.t6 175.169
R31409 a_1606_42308.n3 a_1606_42308.n1 169.016
R31410 a_1606_42308.n3 a_1606_42308.n2 123.073
R31411 a_1606_42308.n4 a_1606_42308.n3 31.8043
R31412 a_1606_42308.t1 a_1606_42308.n5 26.5955
R31413 a_1606_42308.n5 a_1606_42308.t0 26.5955
R31414 a_1606_42308.n0 a_1606_42308.t3 24.9236
R31415 a_1606_42308.n0 a_1606_42308.t2 24.9236
R31416 C0_N_btm.n1 C0_N_btm.t0 101.944
R31417 C0_N_btm.n2 C0_N_btm.t1 99.4985
R31418 C0_N_btm.n0 C0_N_btm.t2 54.9098
R31419 C0_N_btm C0_N_btm.n2 47.6047
R31420 C0_N_btm.n0 C0_N_btm.t3 47.3635
R31421 C0_N_btm.n1 C0_N_btm.n0 8.27654
R31422 C0_N_btm.n2 C0_N_btm.n1 6.33383
R31423 a_18194_34908.n3 a_18194_34908.t11 749.612
R31424 a_18194_34908.n9 a_18194_34908.t9 748.122
R31425 a_18194_34908.n7 a_18194_34908.t12 748.122
R31426 a_18194_34908.n5 a_18194_34908.t13 684.441
R31427 a_18194_34908.n3 a_18194_34908.t15 684.441
R31428 a_18194_34908.n4 a_18194_34908.t14 684.441
R31429 a_18194_34908.n9 a_18194_34908.t8 678.014
R31430 a_18194_34908.n7 a_18194_34908.t10 678.014
R31431 a_18194_34908.n13 a_18194_34908.n12 244.069
R31432 a_18194_34908.n2 a_18194_34908.n0 236.589
R31433 a_18194_34908.n14 a_18194_34908.n13 204.893
R31434 a_18194_34908.n2 a_18194_34908.n1 200.321
R31435 a_18194_34908.n8 a_18194_34908.n7 163.538
R31436 a_18194_34908.n10 a_18194_34908.n9 163.538
R31437 a_18194_34908.n6 a_18194_34908.n5 161.513
R31438 a_18194_34908.n6 a_18194_34908.n3 161.487
R31439 a_18194_34908.n5 a_18194_34908.n4 65.1723
R31440 a_18194_34908.n4 a_18194_34908.n3 65.1723
R31441 a_18194_34908.n11 a_18194_34908.n2 26.8022
R31442 a_18194_34908.n12 a_18194_34908.t1 26.5955
R31443 a_18194_34908.n12 a_18194_34908.t0 26.5955
R31444 a_18194_34908.t3 a_18194_34908.n14 26.5955
R31445 a_18194_34908.n14 a_18194_34908.t2 26.5955
R31446 a_18194_34908.n13 a_18194_34908.n11 25.4552
R31447 a_18194_34908.n0 a_18194_34908.t6 24.9236
R31448 a_18194_34908.n0 a_18194_34908.t4 24.9236
R31449 a_18194_34908.n1 a_18194_34908.t7 24.9236
R31450 a_18194_34908.n1 a_18194_34908.t5 24.9236
R31451 a_18194_34908.n8 a_18194_34908.n6 8.34106
R31452 a_18194_34908.n11 a_18194_34908.n10 6.0248
R31453 a_18194_34908.n10 a_18194_34908.n8 2.47042
R31454 a_1423_45028.n1 a_1423_45028.t7 323.55
R31455 a_1423_45028.n2 a_1423_45028.t4 238.59
R31456 a_1423_45028.n3 a_1423_45028.n1 204.679
R31457 a_1423_45028.n2 a_1423_45028.t6 203.244
R31458 a_1423_45028.n1 a_1423_45028.t5 195.017
R31459 a_1423_45028.n5 a_1423_45028.n4 190.911
R31460 a_1423_45028.n3 a_1423_45028.n2 175.121
R31461 a_1423_45028.n4 a_1423_45028.n0 150.264
R31462 a_1423_45028.n4 a_1423_45028.n3 36.0212
R31463 a_1423_45028.n5 a_1423_45028.t0 26.5955
R31464 a_1423_45028.t1 a_1423_45028.n5 26.5955
R31465 a_1423_45028.n0 a_1423_45028.t3 24.9236
R31466 a_1423_45028.n0 a_1423_45028.t2 24.9236
R31467 a_12741_44636.n0 a_12741_44636.t4 276.464
R31468 a_12741_44636.n1 a_12741_44636.t3 230.155
R31469 a_12741_44636.n2 a_12741_44636.n0 198.028
R31470 a_12741_44636.n4 a_12741_44636.n3 196.846
R31471 a_12741_44636.n0 a_12741_44636.t5 196.131
R31472 a_12741_44636.n3 a_12741_44636.t2 193.519
R31473 a_12741_44636.n2 a_12741_44636.n1 178.474
R31474 a_12741_44636.n1 a_12741_44636.t6 157.856
R31475 a_12741_44636.n4 a_12741_44636.t1 26.5955
R31476 a_12741_44636.t0 a_12741_44636.n4 26.5955
R31477 a_12741_44636.n3 a_12741_44636.n2 16.5418
R31478 a_n3565_38216.n4 a_n3565_38216.t10 557.019
R31479 a_n3565_38216.n8 a_n3565_38216.n7 340.637
R31480 a_n3565_38216.n3 a_n3565_38216.t8 241.536
R31481 a_n3565_38216.n7 a_n3565_38216.n6 195.577
R31482 a_n3565_38216.n3 a_n3565_38216.t9 169.237
R31483 a_n3565_38216.n4 a_n3565_38216.n3 168.845
R31484 a_n3565_38216.n2 a_n3565_38216.n0 137.189
R31485 a_n3565_38216.n2 a_n3565_38216.n1 98.787
R31486 a_n3565_38216.n7 a_n3565_38216.n5 39.0246
R31487 a_n3565_38216.n6 a_n3565_38216.t2 26.5955
R31488 a_n3565_38216.n6 a_n3565_38216.t0 26.5955
R31489 a_n3565_38216.t3 a_n3565_38216.n8 26.5955
R31490 a_n3565_38216.n8 a_n3565_38216.t1 26.5955
R31491 a_n3565_38216.n5 a_n3565_38216.n2 25.9824
R31492 a_n3565_38216.n0 a_n3565_38216.t4 24.9236
R31493 a_n3565_38216.n0 a_n3565_38216.t7 24.9236
R31494 a_n3565_38216.n1 a_n3565_38216.t5 24.9236
R31495 a_n3565_38216.n1 a_n3565_38216.t6 24.9236
R31496 a_n3565_38216.n5 a_n3565_38216.n4 9.3005
R31497 a_765_45546.n9 a_765_45546.n8 680.03
R31498 a_765_45546.n6 a_765_45546.t4 325.774
R31499 a_765_45546.n8 a_765_45546.n0 290.231
R31500 a_765_45546.n2 a_765_45546.t8 241.536
R31501 a_765_45546.n1 a_765_45546.t6 241.536
R31502 a_765_45546.n4 a_765_45546.t9 241.536
R31503 a_765_45546.n3 a_765_45546.n1 190.942
R31504 a_765_45546.n5 a_765_45546.n4 189.668
R31505 a_765_45546.n2 a_765_45546.t7 169.237
R31506 a_765_45546.n1 a_765_45546.t11 169.237
R31507 a_765_45546.n4 a_765_45546.t10 169.237
R31508 a_765_45546.n3 a_765_45546.n2 167.159
R31509 a_765_45546.n6 a_765_45546.t5 129
R31510 a_765_45546.n9 a_765_45546.t0 33.4905
R31511 a_765_45546.n7 a_765_45546.n6 31.393
R31512 a_765_45546.n0 a_765_45546.t2 26.5955
R31513 a_765_45546.n0 a_765_45546.t3 26.5955
R31514 a_765_45546.t1 a_765_45546.n9 26.5955
R31515 a_765_45546.n8 a_765_45546.n7 24.4794
R31516 a_765_45546.n5 a_765_45546.n3 24.147
R31517 a_765_45546.n7 a_765_45546.n5 14.1287
R31518 a_17517_44484.n1 a_17517_44484.t1 352.276
R31519 a_17517_44484.t0 a_17517_44484.n1 327.652
R31520 a_17517_44484.n0 a_17517_44484.t2 276.464
R31521 a_17517_44484.n0 a_17517_44484.t3 196.131
R31522 a_17517_44484.n1 a_17517_44484.n0 195.496
R31523 a_4915_47217.t0 a_4915_47217.n8 717.596
R31524 a_4915_47217.t0 a_4915_47217.n9 710.019
R31525 a_4915_47217.n0 a_4915_47217.t4 471.289
R31526 a_4915_47217.n9 a_4915_47217.t1 276.649
R31527 a_4915_47217.n1 a_4915_47217.t2 256.07
R31528 a_4915_47217.n6 a_4915_47217.t10 230.155
R31529 a_4915_47217.n4 a_4915_47217.t5 212.081
R31530 a_4915_47217.n3 a_4915_47217.t6 212.081
R31531 a_4915_47217.n2 a_4915_47217.n0 203.351
R31532 a_4915_47217.n5 a_4915_47217.n4 194.022
R31533 a_4915_47217.n7 a_4915_47217.n6 188.001
R31534 a_4915_47217.n2 a_4915_47217.n1 186.349
R31535 a_4915_47217.n6 a_4915_47217.t9 157.856
R31536 a_4915_47217.n1 a_4915_47217.t7 150.03
R31537 a_4915_47217.n0 a_4915_47217.t11 148.35
R31538 a_4915_47217.n4 a_4915_47217.t3 139.78
R31539 a_4915_47217.n3 a_4915_47217.t8 139.78
R31540 a_4915_47217.n4 a_4915_47217.n3 61.346
R31541 a_4915_47217.n9 a_4915_47217.n8 17.0672
R31542 a_4915_47217.n5 a_4915_47217.n2 15.5125
R31543 a_4915_47217.n8 a_4915_47217.n7 11.8103
R31544 a_4915_47217.n7 a_4915_47217.n5 11.8056
R31545 a_20820_30879.n0 a_20820_30879.t4 756.514
R31546 a_20820_30879.n0 a_20820_30879.t5 756.239
R31547 a_20820_30879.n3 a_20820_30879.n2 380.32
R31548 a_20820_30879.n2 a_20820_30879.n1 185
R31549 a_20820_30879.n2 a_20820_30879.n0 110.659
R31550 a_20820_30879.t1 a_20820_30879.n3 26.5955
R31551 a_20820_30879.n3 a_20820_30879.t0 26.5955
R31552 a_20820_30879.n1 a_20820_30879.t3 24.9236
R31553 a_20820_30879.n1 a_20820_30879.t2 24.9236
R31554 a_n4209_37414.n4 a_n4209_37414.t9 553.064
R31555 a_n4209_37414.n7 a_n4209_37414.n6 340.637
R31556 a_n4209_37414.n3 a_n4209_37414.t8 241.536
R31557 a_n4209_37414.n8 a_n4209_37414.n7 195.577
R31558 a_n4209_37414.n4 a_n4209_37414.n3 173.952
R31559 a_n4209_37414.n3 a_n4209_37414.t10 169.237
R31560 a_n4209_37414.n2 a_n4209_37414.n0 137.189
R31561 a_n4209_37414.n2 a_n4209_37414.n1 98.788
R31562 a_n4209_37414.n7 a_n4209_37414.n5 37.1695
R31563 a_n4209_37414.n5 a_n4209_37414.n2 27.8375
R31564 a_n4209_37414.n6 a_n4209_37414.t2 26.5955
R31565 a_n4209_37414.n6 a_n4209_37414.t0 26.5955
R31566 a_n4209_37414.t3 a_n4209_37414.n8 26.5955
R31567 a_n4209_37414.n8 a_n4209_37414.t1 26.5955
R31568 a_n4209_37414.n0 a_n4209_37414.t4 24.9236
R31569 a_n4209_37414.n0 a_n4209_37414.t6 24.9236
R31570 a_n4209_37414.n1 a_n4209_37414.t5 24.9236
R31571 a_n4209_37414.n1 a_n4209_37414.t7 24.9236
R31572 a_n4209_37414.n5 a_n4209_37414.n4 9.30997
R31573 a_768_44030.n4 a_768_44030.n0 252.931
R31574 a_768_44030.n19 a_768_44030.t19 241.536
R31575 a_768_44030.n5 a_768_44030.t8 241.536
R31576 a_768_44030.n16 a_768_44030.t16 241.536
R31577 a_768_44030.n12 a_768_44030.t14 241.536
R31578 a_768_44030.n3 a_768_44030.n1 238.163
R31579 a_768_44030.n9 a_768_44030.t13 212.081
R31580 a_768_44030.n10 a_768_44030.t23 212.081
R31581 a_768_44030.n11 a_768_44030.n10 210.942
R31582 a_768_44030.n14 a_768_44030.t11 206.19
R31583 a_768_44030.n6 a_768_44030.t15 206.19
R31584 a_768_44030.n22 a_768_44030.n21 188.983
R31585 a_768_44030.n7 a_768_44030.t20 185.376
R31586 a_768_44030.n17 a_768_44030.n16 177.773
R31587 a_768_44030.n13 a_768_44030.n12 176.047
R31588 a_768_44030.n18 a_768_44030.n5 174.227
R31589 a_768_44030.n20 a_768_44030.n19 173.752
R31590 a_768_44030.n8 a_768_44030.n6 172.607
R31591 a_768_44030.n8 a_768_44030.n7 171.845
R31592 a_768_44030.n15 a_768_44030.n14 171.078
R31593 a_768_44030.n19 a_768_44030.t9 169.237
R31594 a_768_44030.n5 a_768_44030.t22 169.237
R31595 a_768_44030.n16 a_768_44030.t18 169.237
R31596 a_768_44030.n12 a_768_44030.t25 169.237
R31597 a_768_44030.n14 a_768_44030.t12 148.35
R31598 a_768_44030.n6 a_768_44030.t10 148.35
R31599 a_768_44030.n9 a_768_44030.t17 139.78
R31600 a_768_44030.n10 a_768_44030.t24 139.78
R31601 a_768_44030.n7 a_768_44030.t21 137.177
R31602 a_768_44030.n3 a_768_44030.n2 98.981
R31603 a_768_44030.n4 a_768_44030.n3 70.96
R31604 a_768_44030.n10 a_768_44030.n9 61.346
R31605 a_768_44030.n21 a_768_44030.n20 39.2218
R31606 a_768_44030.n0 a_768_44030.t0 26.5955
R31607 a_768_44030.n0 a_768_44030.t2 26.5955
R31608 a_768_44030.t3 a_768_44030.n22 26.5955
R31609 a_768_44030.n22 a_768_44030.t1 26.5955
R31610 a_768_44030.n1 a_768_44030.t7 24.9236
R31611 a_768_44030.n1 a_768_44030.t6 24.9236
R31612 a_768_44030.n2 a_768_44030.t5 24.9236
R31613 a_768_44030.n2 a_768_44030.t4 24.9236
R31614 a_768_44030.n21 a_768_44030.n4 19.5257
R31615 a_768_44030.n20 a_768_44030.n18 12.2189
R31616 a_768_44030.n18 a_768_44030.n17 7.18714
R31617 a_768_44030.n15 a_768_44030.n13 5.63228
R31618 a_768_44030.n13 a_768_44030.n11 4.6495
R31619 a_768_44030.n17 a_768_44030.n15 3.16673
R31620 a_768_44030.n11 a_768_44030.n8 0.6444
R31621 a_n4209_39304.n4 a_n4209_39304.t11 756.514
R31622 a_n4209_39304.n4 a_n4209_39304.t8 756.239
R31623 a_n4209_39304.n9 a_n4209_39304.n8 340.637
R31624 a_n4209_39304.n3 a_n4209_39304.t10 241.536
R31625 a_n4209_39304.n8 a_n4209_39304.n7 195.577
R31626 a_n4209_39304.n5 a_n4209_39304.n3 174.202
R31627 a_n4209_39304.n3 a_n4209_39304.t9 169.237
R31628 a_n4209_39304.n2 a_n4209_39304.n0 137.189
R31629 a_n4209_39304.n2 a_n4209_39304.n1 98.787
R31630 a_n4209_39304.n5 a_n4209_39304.n4 73.3836
R31631 a_n4209_39304.n6 a_n4209_39304.n2 38.9679
R31632 a_n4209_39304.n7 a_n4209_39304.t2 26.5955
R31633 a_n4209_39304.n7 a_n4209_39304.t0 26.5955
R31634 a_n4209_39304.n9 a_n4209_39304.t1 26.5955
R31635 a_n4209_39304.t3 a_n4209_39304.n9 26.5955
R31636 a_n4209_39304.n8 a_n4209_39304.n6 26.0391
R31637 a_n4209_39304.n0 a_n4209_39304.t6 24.9236
R31638 a_n4209_39304.n0 a_n4209_39304.t7 24.9236
R31639 a_n4209_39304.n1 a_n4209_39304.t5 24.9236
R31640 a_n4209_39304.n1 a_n4209_39304.t4 24.9236
R31641 a_n4209_39304.n6 a_n4209_39304.n5 9.30997
R31642 a_n2956_38680.n3 a_n2956_38680.n2 296.139
R31643 a_n2956_38680.n2 a_n2956_38680.n0 269.182
R31644 a_n2956_38680.n2 a_n2956_38680.n1 254.305
R31645 a_n2956_38680.n1 a_n2956_38680.t4 228.649
R31646 a_n2956_38680.n1 a_n2956_38680.t5 156.35
R31647 a_n2956_38680.n3 a_n2956_38680.t0 26.5955
R31648 a_n2956_38680.t1 a_n2956_38680.n3 26.5955
R31649 a_n2956_38680.n0 a_n2956_38680.t2 24.9236
R31650 a_n2956_38680.n0 a_n2956_38680.t3 24.9236
R31651 a_14097_32519.n1 a_14097_32519.t4 672.947
R31652 a_14097_32519.n2 a_14097_32519.n1 380.32
R31653 a_14097_32519.n1 a_14097_32519.n0 185
R31654 a_14097_32519.n2 a_14097_32519.t0 26.5955
R31655 a_14097_32519.t1 a_14097_32519.n2 26.5955
R31656 a_14097_32519.n0 a_14097_32519.t3 24.9236
R31657 a_14097_32519.n0 a_14097_32519.t2 24.9236
R31658 C4_N_btm.n1 C4_N_btm.t3 101.361
R31659 C4_N_btm.n2 C4_N_btm.t0 98.3735
R31660 C4_N_btm.n0 C4_N_btm.t2 54.9311
R31661 C4_N_btm C4_N_btm.n2 52.9172
R31662 C4_N_btm.n0 C4_N_btm.t1 47.3635
R31663 C4_N_btm.n2 C4_N_btm.n1 8.08383
R31664 C4_N_btm.n1 C4_N_btm.n0 7.15154
R31665 a_20692_30879.n1 a_20692_30879.t4 866.769
R31666 a_20692_30879.n2 a_20692_30879.n1 380.32
R31667 a_20692_30879.n1 a_20692_30879.n0 185
R31668 a_20692_30879.t1 a_20692_30879.n2 26.5955
R31669 a_20692_30879.n2 a_20692_30879.t0 26.5955
R31670 a_20692_30879.n0 a_20692_30879.t3 24.9236
R31671 a_20692_30879.n0 a_20692_30879.t2 24.9236
R31672 C6_N_btm.n4 C6_N_btm.t0 97.811
R31673 C6_N_btm.n3 C6_N_btm.t1 68.0518
R31674 C6_N_btm C6_N_btm.n4 57.8859
R31675 C6_N_btm.n2 C6_N_btm.n0 45.0311
R31676 C6_N_btm.n2 C6_N_btm.n1 37.4635
R31677 C6_N_btm.n1 C6_N_btm.t5 9.9005
R31678 C6_N_btm.n1 C6_N_btm.t4 9.9005
R31679 C6_N_btm.n0 C6_N_btm.t3 9.9005
R31680 C6_N_btm.n0 C6_N_btm.t2 9.9005
R31681 C6_N_btm.n4 C6_N_btm.n3 8.0005
R31682 C6_N_btm.n3 C6_N_btm.n2 6.58904
R31683 a_n2293_42834.n0 a_n2293_42834.t3 276.464
R31684 a_n2293_42834.n2 a_n2293_42834.n1 254.679
R31685 a_n2293_42834.n1 a_n2293_42834.n0 207.022
R31686 a_n2293_42834.n0 a_n2293_42834.t4 196.131
R31687 a_n2293_42834.n1 a_n2293_42834.t1 135.579
R31688 a_n2293_42834.n2 a_n2293_42834.t2 26.5955
R31689 a_n2293_42834.t0 a_n2293_42834.n2 26.5955
R31690 a_21588_30879.n0 a_21588_30879.t8 756.547
R31691 a_21588_30879.n6 a_21588_30879.t6 756.231
R31692 a_21588_30879.n0 a_21588_30879.t4 756.226
R31693 a_21588_30879.n1 a_21588_30879.t11 756.226
R31694 a_21588_30879.n2 a_21588_30879.t7 756.226
R31695 a_21588_30879.n3 a_21588_30879.t9 756.226
R31696 a_21588_30879.n4 a_21588_30879.t10 756.226
R31697 a_21588_30879.n5 a_21588_30879.t5 756.226
R31698 a_21588_30879.n9 a_21588_30879.n8 380.32
R31699 a_21588_30879.n8 a_21588_30879.n7 185
R31700 a_21588_30879.n8 a_21588_30879.n6 104.999
R31701 a_21588_30879.n9 a_21588_30879.t0 26.5955
R31702 a_21588_30879.t1 a_21588_30879.n9 26.5955
R31703 a_21588_30879.n7 a_21588_30879.t3 24.9236
R31704 a_21588_30879.n7 a_21588_30879.t2 24.9236
R31705 a_21588_30879.n5 a_21588_30879.n4 0.3205
R31706 a_21588_30879.n4 a_21588_30879.n3 0.3205
R31707 a_21588_30879.n3 a_21588_30879.n2 0.3205
R31708 a_21588_30879.n2 a_21588_30879.n1 0.3205
R31709 a_21588_30879.n1 a_21588_30879.n0 0.3205
R31710 a_21588_30879.n6 a_21588_30879.n5 0.298833
R31711 C9_N_btm C9_N_btm.n15 80.4693
R31712 C9_N_btm.n2 C9_N_btm.n0 33.0802
R31713 C9_N_btm.n6 C9_N_btm.n5 32.3614
R31714 C9_N_btm.n4 C9_N_btm.n3 32.3614
R31715 C9_N_btm.n2 C9_N_btm.n1 32.3614
R31716 C9_N_btm.n10 C9_N_btm.n6 24.0265
R31717 C9_N_btm.n11 C9_N_btm.t8 23.0826
R31718 C9_N_btm.n14 C9_N_btm.n13 15.4287
R31719 C9_N_btm.n9 C9_N_btm.n7 15.3784
R31720 C9_N_btm.n14 C9_N_btm.n12 14.9755
R31721 C9_N_btm.n9 C9_N_btm.n8 14.894
R31722 C9_N_btm.n15 C9_N_btm.n11 7.16717
R31723 C9_N_btm.n10 C9_N_btm.n9 5.71404
R31724 C9_N_btm.n15 C9_N_btm.n14 5.62029
R31725 C9_N_btm C9_N_btm.n513 5.59972
R31726 C9_N_btm.n11 C9_N_btm.n10 3.91717
R31727 C9_N_btm.n5 C9_N_btm.t11 3.57113
R31728 C9_N_btm.n5 C9_N_btm.t12 3.57113
R31729 C9_N_btm.n3 C9_N_btm.t15 3.57113
R31730 C9_N_btm.n3 C9_N_btm.t13 3.57113
R31731 C9_N_btm.n1 C9_N_btm.t14 3.57113
R31732 C9_N_btm.n1 C9_N_btm.t16 3.57113
R31733 C9_N_btm.n0 C9_N_btm.t9 3.57113
R31734 C9_N_btm.n0 C9_N_btm.t10 3.57113
R31735 C9_N_btm.n12 C9_N_btm.t0 2.4755
R31736 C9_N_btm.n12 C9_N_btm.t2 2.4755
R31737 C9_N_btm.n8 C9_N_btm.t4 2.4755
R31738 C9_N_btm.n8 C9_N_btm.t7 2.4755
R31739 C9_N_btm.n7 C9_N_btm.t5 2.4755
R31740 C9_N_btm.n7 C9_N_btm.t6 2.4755
R31741 C9_N_btm.n13 C9_N_btm.t3 2.4755
R31742 C9_N_btm.n13 C9_N_btm.t1 2.4755
R31743 C9_N_btm.n4 C9_N_btm.n2 0.688
R31744 C9_N_btm.n6 C9_N_btm.n4 0.672375
R31745 C9_N_btm.n104 C9_N_btm.n100 0.276161
R31746 C9_N_btm.n68 C9_N_btm.n67 0.276161
R31747 C9_N_btm.n301 C9_N_btm.n298 0.276161
R31748 C9_N_btm.n331 C9_N_btm.n330 0.276161
R31749 C9_N_btm.n305 C9_N_btm.n304 0.276161
R31750 C9_N_btm.n98 C9_N_btm.n97 0.228786
R31751 C9_N_btm.n100 C9_N_btm.n98 0.228786
R31752 C9_N_btm.n97 C9_N_btm.n96 0.228786
R31753 C9_N_btm.n91 C9_N_btm.n90 0.228786
R31754 C9_N_btm.n95 C9_N_btm.n91 0.228786
R31755 C9_N_btm.n96 C9_N_btm.n95 0.228786
R31756 C9_N_btm.n90 C9_N_btm.n82 0.228786
R31757 C9_N_btm.n121 C9_N_btm.n120 0.228786
R31758 C9_N_btm.n120 C9_N_btm.n119 0.228786
R31759 C9_N_btm.n119 C9_N_btm.n82 0.228786
R31760 C9_N_btm.n122 C9_N_btm.n121 0.228786
R31761 C9_N_btm.n76 C9_N_btm.n75 0.228786
R31762 C9_N_btm.n78 C9_N_btm.n76 0.228786
R31763 C9_N_btm.n122 C9_N_btm.n78 0.228786
R31764 C9_N_btm.n75 C9_N_btm.n74 0.228786
R31765 C9_N_btm.n59 C9_N_btm.n58 0.228786
R31766 C9_N_btm.n73 C9_N_btm.n58 0.228786
R31767 C9_N_btm.n74 C9_N_btm.n73 0.228786
R31768 C9_N_btm.n68 C9_N_btm.n59 0.228786
R31769 C9_N_btm.n66 C9_N_btm.n65 0.228786
R31770 C9_N_btm.n64 C9_N_btm.n63 0.228786
R31771 C9_N_btm.n62 C9_N_btm.n51 0.228786
R31772 C9_N_btm.n136 C9_N_btm.n50 0.228786
R31773 C9_N_btm.n138 C9_N_btm.n137 0.228786
R31774 C9_N_btm.n139 C9_N_btm.n48 0.228786
R31775 C9_N_btm.n482 C9_N_btm.n140 0.228786
R31776 C9_N_btm.n298 C9_N_btm.n297 0.228786
R31777 C9_N_btm.n297 C9_N_btm.n296 0.228786
R31778 C9_N_btm.n296 C9_N_btm.n295 0.228786
R31779 C9_N_btm.n295 C9_N_btm.n294 0.228786
R31780 C9_N_btm.n294 C9_N_btm.n293 0.228786
R31781 C9_N_btm.n293 C9_N_btm.n290 0.228786
R31782 C9_N_btm.n290 C9_N_btm.n289 0.228786
R31783 C9_N_btm.n289 C9_N_btm.n288 0.228786
R31784 C9_N_btm.n288 C9_N_btm.n287 0.228786
R31785 C9_N_btm.n287 C9_N_btm.n286 0.228786
R31786 C9_N_btm.n286 C9_N_btm.n285 0.228786
R31787 C9_N_btm.n285 C9_N_btm.n282 0.228786
R31788 C9_N_btm.n281 C9_N_btm.n280 0.228786
R31789 C9_N_btm.n282 C9_N_btm.n281 0.228786
R31790 C9_N_btm.n237 C9_N_btm.n236 0.228786
R31791 C9_N_btm.n362 C9_N_btm.n361 0.228786
R31792 C9_N_btm.n363 C9_N_btm.n235 0.228786
R31793 C9_N_btm.n384 C9_N_btm.n364 0.228786
R31794 C9_N_btm.n383 C9_N_btm.n382 0.228786
R31795 C9_N_btm.n381 C9_N_btm.n365 0.228786
R31796 C9_N_btm.n380 C9_N_btm.n366 0.228786
R31797 C9_N_btm.n379 C9_N_btm.n378 0.228786
R31798 C9_N_btm.n377 C9_N_btm.n368 0.228786
R31799 C9_N_btm.n367 C9_N_btm.n202 0.228786
R31800 C9_N_btm.n401 C9_N_btm.n200 0.228786
R31801 C9_N_btm.n425 C9_N_btm.n424 0.228786
R31802 C9_N_btm.n423 C9_N_btm.n197 0.228786
R31803 C9_N_btm.n422 C9_N_btm.n405 0.228786
R31804 C9_N_btm.n421 C9_N_btm.n420 0.228786
R31805 C9_N_btm.n419 C9_N_btm.n406 0.228786
R31806 C9_N_btm.n409 C9_N_btm.n408 0.228786
R31807 C9_N_btm.n411 C9_N_btm.n410 0.228786
R31808 C9_N_btm.n167 C9_N_btm.n166 0.228786
R31809 C9_N_btm.n445 C9_N_btm.n444 0.228786
R31810 C9_N_btm.n446 C9_N_btm.n165 0.228786
R31811 C9_N_btm.n453 C9_N_btm.n452 0.228786
R31812 C9_N_btm.n451 C9_N_btm.n163 0.228786
R31813 C9_N_btm.n449 C9_N_btm.n448 0.228786
R31814 C9_N_btm.n143 C9_N_btm.n142 0.228786
R31815 C9_N_btm.n478 C9_N_btm.n477 0.228786
R31816 C9_N_btm.n479 C9_N_btm.n141 0.228786
R31817 C9_N_btm.n102 C9_N_btm.n18 0.228786
R31818 C9_N_btm.n103 C9_N_btm.n101 0.228786
R31819 C9_N_btm.n106 C9_N_btm.n105 0.228786
R31820 C9_N_btm.n107 C9_N_btm.n106 0.228786
R31821 C9_N_btm.n99 C9_N_btm.n94 0.228786
R31822 C9_N_btm.n101 C9_N_btm.n99 0.228786
R31823 C9_N_btm.n19 C9_N_btm.n18 0.228786
R31824 C9_N_btm.n21 C9_N_btm.n19 0.228786
R31825 C9_N_btm.n22 C9_N_btm.n21 0.228786
R31826 C9_N_btm.n111 C9_N_btm.n22 0.228786
R31827 C9_N_btm.n110 C9_N_btm.n109 0.228786
R31828 C9_N_btm.n109 C9_N_btm.n94 0.228786
R31829 C9_N_btm.n108 C9_N_btm.n107 0.228786
R31830 C9_N_btm.n108 C9_N_btm.n93 0.228786
R31831 C9_N_btm.n93 C9_N_btm.n92 0.228786
R31832 C9_N_btm.n115 C9_N_btm.n92 0.228786
R31833 C9_N_btm.n114 C9_N_btm.n113 0.228786
R31834 C9_N_btm.n113 C9_N_btm.n110 0.228786
R31835 C9_N_btm.n112 C9_N_btm.n111 0.228786
R31836 C9_N_btm.n112 C9_N_btm.n26 0.228786
R31837 C9_N_btm.n27 C9_N_btm.n26 0.228786
R31838 C9_N_btm.n29 C9_N_btm.n27 0.228786
R31839 C9_N_btm.n89 C9_N_btm.n88 0.228786
R31840 C9_N_btm.n114 C9_N_btm.n89 0.228786
R31841 C9_N_btm.n116 C9_N_btm.n115 0.228786
R31842 C9_N_btm.n117 C9_N_btm.n116 0.228786
R31843 C9_N_btm.n118 C9_N_btm.n117 0.228786
R31844 C9_N_btm.n118 C9_N_btm.n81 0.228786
R31845 C9_N_btm.n87 C9_N_btm.n86 0.228786
R31846 C9_N_btm.n88 C9_N_btm.n87 0.228786
R31847 C9_N_btm.n30 C9_N_btm.n29 0.228786
R31848 C9_N_btm.n83 C9_N_btm.n30 0.228786
R31849 C9_N_btm.n84 C9_N_btm.n83 0.228786
R31850 C9_N_btm.n84 C9_N_btm.n34 0.228786
R31851 C9_N_btm.n85 C9_N_btm.n79 0.228786
R31852 C9_N_btm.n86 C9_N_btm.n85 0.228786
R31853 C9_N_btm.n81 C9_N_btm.n80 0.228786
R31854 C9_N_btm.n123 C9_N_btm.n80 0.228786
R31855 C9_N_btm.n124 C9_N_btm.n123 0.228786
R31856 C9_N_btm.n125 C9_N_btm.n124 0.228786
R31857 C9_N_btm.n77 C9_N_btm.n57 0.228786
R31858 C9_N_btm.n79 C9_N_btm.n77 0.228786
R31859 C9_N_btm.n35 C9_N_btm.n34 0.228786
R31860 C9_N_btm.n37 C9_N_btm.n35 0.228786
R31861 C9_N_btm.n38 C9_N_btm.n37 0.228786
R31862 C9_N_btm.n129 C9_N_btm.n38 0.228786
R31863 C9_N_btm.n128 C9_N_btm.n127 0.228786
R31864 C9_N_btm.n127 C9_N_btm.n57 0.228786
R31865 C9_N_btm.n126 C9_N_btm.n125 0.228786
R31866 C9_N_btm.n126 C9_N_btm.n56 0.228786
R31867 C9_N_btm.n72 C9_N_btm.n56 0.228786
R31868 C9_N_btm.n72 C9_N_btm.n71 0.228786
R31869 C9_N_btm.n55 C9_N_btm.n54 0.228786
R31870 C9_N_btm.n128 C9_N_btm.n55 0.228786
R31871 C9_N_btm.n42 C9_N_btm.n39 0.228786
R31872 C9_N_btm.n130 C9_N_btm.n129 0.228786
R31873 C9_N_btm.n131 C9_N_btm.n130 0.228786
R31874 C9_N_btm.n43 C9_N_btm.n42 0.228786
R31875 C9_N_btm.n489 C9_N_btm.n488 0.228786
R31876 C9_N_btm.n485 C9_N_btm.n484 0.228786
R31877 C9_N_btm.n486 C9_N_btm.n46 0.228786
R31878 C9_N_btm.n487 C9_N_btm.n486 0.228786
R31879 C9_N_btm.n488 C9_N_btm.n44 0.228786
R31880 C9_N_btm.n135 C9_N_btm.n44 0.228786
R31881 C9_N_btm.n134 C9_N_btm.n133 0.228786
R31882 C9_N_btm.n133 C9_N_btm.n43 0.228786
R31883 C9_N_btm.n132 C9_N_btm.n131 0.228786
R31884 C9_N_btm.n132 C9_N_btm.n52 0.228786
R31885 C9_N_btm.n60 C9_N_btm.n53 0.228786
R31886 C9_N_btm.n54 C9_N_btm.n53 0.228786
R31887 C9_N_btm.n71 C9_N_btm.n70 0.228786
R31888 C9_N_btm.n70 C9_N_btm.n69 0.228786
R31889 C9_N_btm.n69 C9_N_btm.n61 0.228786
R31890 C9_N_btm.n65 C9_N_btm.n60 0.228786
R31891 C9_N_btm.n64 C9_N_btm.n52 0.228786
R31892 C9_N_btm.n134 C9_N_btm.n51 0.228786
R31893 C9_N_btm.n136 C9_N_btm.n135 0.228786
R31894 C9_N_btm.n137 C9_N_btm.n46 0.228786
R31895 C9_N_btm.n484 C9_N_btm.n48 0.228786
R31896 C9_N_btm.n483 C9_N_btm.n482 0.228786
R31897 C9_N_btm.n481 C9_N_btm.n480 0.228786
R31898 C9_N_btm.n466 C9_N_btm.n465 0.228786
R31899 C9_N_btm.n472 C9_N_btm.n471 0.228786
R31900 C9_N_btm.n470 C9_N_btm.n151 0.228786
R31901 C9_N_btm.n469 C9_N_btm.n468 0.228786
R31902 C9_N_btm.n468 C9_N_btm.n467 0.228786
R31903 C9_N_btm.n151 C9_N_btm.n149 0.228786
R31904 C9_N_btm.n149 C9_N_btm.n148 0.228786
R31905 C9_N_btm.n474 C9_N_btm.n145 0.228786
R31906 C9_N_btm.n476 C9_N_btm.n475 0.228786
R31907 C9_N_btm.n475 C9_N_btm.n147 0.228786
R31908 C9_N_btm.n474 C9_N_btm.n473 0.228786
R31909 C9_N_btm.n473 C9_N_btm.n472 0.228786
R31910 C9_N_btm.n154 C9_N_btm.n152 0.228786
R31911 C9_N_btm.n150 C9_N_btm.n147 0.228786
R31912 C9_N_btm.n464 C9_N_btm.n150 0.228786
R31913 C9_N_btm.n463 C9_N_btm.n152 0.228786
R31914 C9_N_btm.n462 C9_N_btm.n461 0.228786
R31915 C9_N_btm.n460 C9_N_btm.n153 0.228786
R31916 C9_N_btm.n176 C9_N_btm.n156 0.228786
R31917 C9_N_btm.n178 C9_N_btm.n177 0.228786
R31918 C9_N_btm.n184 C9_N_btm.n183 0.228786
R31919 C9_N_btm.n432 C9_N_btm.n188 0.228786
R31920 C9_N_btm.n212 C9_N_btm.n190 0.228786
R31921 C9_N_btm.n300 C9_N_btm.n299 0.228786
R31922 C9_N_btm.n299 C9_N_btm.n274 0.228786
R31923 C9_N_btm.n274 C9_N_btm.n273 0.228786
R31924 C9_N_btm.n273 C9_N_btm.n271 0.228786
R31925 C9_N_btm.n271 C9_N_btm.n270 0.228786
R31926 C9_N_btm.n292 C9_N_btm.n270 0.228786
R31927 C9_N_btm.n292 C9_N_btm.n291 0.228786
R31928 C9_N_btm.n291 C9_N_btm.n262 0.228786
R31929 C9_N_btm.n262 C9_N_btm.n261 0.228786
R31930 C9_N_btm.n261 C9_N_btm.n259 0.228786
R31931 C9_N_btm.n259 C9_N_btm.n258 0.228786
R31932 C9_N_btm.n284 C9_N_btm.n258 0.228786
R31933 C9_N_btm.n284 C9_N_btm.n283 0.228786
R31934 C9_N_btm.n283 C9_N_btm.n250 0.228786
R31935 C9_N_btm.n250 C9_N_btm.n249 0.228786
R31936 C9_N_btm.n249 C9_N_btm.n247 0.228786
R31937 C9_N_btm.n247 C9_N_btm.n246 0.228786
R31938 C9_N_btm.n228 C9_N_btm.n227 0.228786
R31939 C9_N_btm.n280 C9_N_btm.n227 0.228786
R31940 C9_N_btm.n389 C9_N_btm.n388 0.228786
R31941 C9_N_btm.n390 C9_N_btm.n389 0.228786
R31942 C9_N_btm.n391 C9_N_btm.n226 0.228786
R31943 C9_N_btm.n230 C9_N_btm.n226 0.228786
R31944 C9_N_btm.n372 C9_N_btm.n225 0.228786
R31945 C9_N_btm.n392 C9_N_btm.n225 0.228786
R31946 C9_N_btm.n393 C9_N_btm.n224 0.228786
R31947 C9_N_btm.n371 C9_N_btm.n224 0.228786
R31948 C9_N_btm.n208 C9_N_btm.n207 0.228786
R31949 C9_N_btm.n394 C9_N_btm.n208 0.228786
R31950 C9_N_btm.n396 C9_N_btm.n395 0.228786
R31951 C9_N_btm.n397 C9_N_btm.n396 0.228786
R31952 C9_N_btm.n209 C9_N_btm.n205 0.228786
R31953 C9_N_btm.n223 C9_N_btm.n209 0.228786
R31954 C9_N_btm.n222 C9_N_btm.n221 0.228786
R31955 C9_N_btm.n221 C9_N_btm.n220 0.228786
R31956 C9_N_btm.n219 C9_N_btm.n211 0.228786
R31957 C9_N_btm.n211 C9_N_btm.n210 0.228786
R31958 C9_N_btm.n214 C9_N_btm.n213 0.228786
R31959 C9_N_btm.n216 C9_N_btm.n215 0.228786
R31960 C9_N_btm.n215 C9_N_btm.n214 0.228786
R31961 C9_N_btm.n191 C9_N_btm.n190 0.228786
R31962 C9_N_btm.n192 C9_N_btm.n191 0.228786
R31963 C9_N_btm.n431 C9_N_btm.n430 0.228786
R31964 C9_N_btm.n432 C9_N_btm.n431 0.228786
R31965 C9_N_btm.n433 C9_N_btm.n189 0.228786
R31966 C9_N_btm.n193 C9_N_btm.n189 0.228786
R31967 C9_N_btm.n416 C9_N_btm.n187 0.228786
R31968 C9_N_btm.n435 C9_N_btm.n187 0.228786
R31969 C9_N_btm.n436 C9_N_btm.n186 0.228786
R31970 C9_N_btm.n415 C9_N_btm.n186 0.228786
R31971 C9_N_btm.n173 C9_N_btm.n172 0.228786
R31972 C9_N_btm.n437 C9_N_btm.n173 0.228786
R31973 C9_N_btm.n439 C9_N_btm.n438 0.228786
R31974 C9_N_btm.n440 C9_N_btm.n439 0.228786
R31975 C9_N_btm.n174 C9_N_btm.n170 0.228786
R31976 C9_N_btm.n175 C9_N_btm.n174 0.228786
R31977 C9_N_btm.n183 C9_N_btm.n182 0.228786
R31978 C9_N_btm.n182 C9_N_btm.n181 0.228786
R31979 C9_N_btm.n180 C9_N_btm.n179 0.228786
R31980 C9_N_btm.n179 C9_N_btm.n178 0.228786
R31981 C9_N_btm.n157 C9_N_btm.n156 0.228786
R31982 C9_N_btm.n158 C9_N_btm.n157 0.228786
R31983 C9_N_btm.n459 C9_N_btm.n458 0.228786
R31984 C9_N_btm.n460 C9_N_btm.n459 0.228786
R31985 C9_N_btm.n461 C9_N_btm.n155 0.228786
R31986 C9_N_btm.n159 C9_N_btm.n155 0.228786
R31987 C9_N_btm.n154 C9_N_btm.n146 0.228786
R31988 C9_N_btm.n146 C9_N_btm.n144 0.228786
R31989 C9_N_btm.n160 C9_N_btm.n159 0.228786
R31990 C9_N_btm.n448 C9_N_btm.n160 0.228786
R31991 C9_N_btm.n457 C9_N_btm.n161 0.228786
R31992 C9_N_btm.n458 C9_N_btm.n457 0.228786
R31993 C9_N_btm.n456 C9_N_btm.n158 0.228786
R31994 C9_N_btm.n456 C9_N_btm.n455 0.228786
R31995 C9_N_btm.n454 C9_N_btm.n162 0.228786
R31996 C9_N_btm.n180 C9_N_btm.n162 0.228786
R31997 C9_N_btm.n181 C9_N_btm.n169 0.228786
R31998 C9_N_btm.n169 C9_N_btm.n164 0.228786
R31999 C9_N_btm.n443 C9_N_btm.n442 0.228786
R32000 C9_N_btm.n442 C9_N_btm.n170 0.228786
R32001 C9_N_btm.n441 C9_N_btm.n440 0.228786
R32002 C9_N_btm.n441 C9_N_btm.n168 0.228786
R32003 C9_N_btm.n412 C9_N_btm.n171 0.228786
R32004 C9_N_btm.n172 C9_N_btm.n171 0.228786
R32005 C9_N_btm.n415 C9_N_btm.n414 0.228786
R32006 C9_N_btm.n414 C9_N_btm.n413 0.228786
R32007 C9_N_btm.n418 C9_N_btm.n417 0.228786
R32008 C9_N_btm.n417 C9_N_btm.n416 0.228786
R32009 C9_N_btm.n194 C9_N_btm.n193 0.228786
R32010 C9_N_btm.n407 C9_N_btm.n194 0.228786
R32011 C9_N_btm.n429 C9_N_btm.n195 0.228786
R32012 C9_N_btm.n430 C9_N_btm.n429 0.228786
R32013 C9_N_btm.n428 C9_N_btm.n192 0.228786
R32014 C9_N_btm.n428 C9_N_btm.n427 0.228786
R32015 C9_N_btm.n217 C9_N_btm.n198 0.228786
R32016 C9_N_btm.n426 C9_N_btm.n196 0.228786
R32017 C9_N_btm.n216 C9_N_btm.n196 0.228786
R32018 C9_N_btm.n218 C9_N_btm.n217 0.228786
R32019 C9_N_btm.n219 C9_N_btm.n218 0.228786
R32020 C9_N_btm.n220 C9_N_btm.n204 0.228786
R32021 C9_N_btm.n402 C9_N_btm.n201 0.228786
R32022 C9_N_btm.n204 C9_N_btm.n201 0.228786
R32023 C9_N_btm.n400 C9_N_btm.n399 0.228786
R32024 C9_N_btm.n399 C9_N_btm.n205 0.228786
R32025 C9_N_btm.n398 C9_N_btm.n397 0.228786
R32026 C9_N_btm.n398 C9_N_btm.n203 0.228786
R32027 C9_N_btm.n376 C9_N_btm.n206 0.228786
R32028 C9_N_btm.n207 C9_N_btm.n206 0.228786
R32029 C9_N_btm.n371 C9_N_btm.n369 0.228786
R32030 C9_N_btm.n375 C9_N_btm.n369 0.228786
R32031 C9_N_btm.n374 C9_N_btm.n373 0.228786
R32032 C9_N_btm.n373 C9_N_btm.n372 0.228786
R32033 C9_N_btm.n231 C9_N_btm.n230 0.228786
R32034 C9_N_btm.n370 C9_N_btm.n231 0.228786
R32035 C9_N_btm.n386 C9_N_btm.n385 0.228786
R32036 C9_N_btm.n387 C9_N_btm.n232 0.228786
R32037 C9_N_btm.n388 C9_N_btm.n387 0.228786
R32038 C9_N_btm.n386 C9_N_btm.n229 0.228786
R32039 C9_N_btm.n229 C9_N_btm.n228 0.228786
R32040 C9_N_btm.n246 C9_N_btm.n245 0.228786
R32041 C9_N_btm.n245 C9_N_btm.n233 0.228786
R32042 C9_N_btm.n234 C9_N_btm.n233 0.228786
R32043 C9_N_btm.n360 C9_N_btm.n238 0.228786
R32044 C9_N_btm.n359 C9_N_btm.n358 0.228786
R32045 C9_N_btm.n358 C9_N_btm.n357 0.228786
R32046 C9_N_btm.n242 C9_N_btm.n238 0.228786
R32047 C9_N_btm.n355 C9_N_btm.n242 0.228786
R32048 C9_N_btm.n357 C9_N_btm.n356 0.228786
R32049 C9_N_btm.n356 C9_N_btm.n244 0.228786
R32050 C9_N_btm.n355 C9_N_btm.n354 0.228786
R32051 C9_N_btm.n354 C9_N_btm.n353 0.228786
R32052 C9_N_btm.n248 C9_N_btm.n244 0.228786
R32053 C9_N_btm.n351 C9_N_btm.n248 0.228786
R32054 C9_N_btm.n353 C9_N_btm.n352 0.228786
R32055 C9_N_btm.n352 C9_N_btm.n251 0.228786
R32056 C9_N_btm.n351 C9_N_btm.n350 0.228786
R32057 C9_N_btm.n350 C9_N_btm.n349 0.228786
R32058 C9_N_btm.n255 C9_N_btm.n251 0.228786
R32059 C9_N_btm.n347 C9_N_btm.n255 0.228786
R32060 C9_N_btm.n349 C9_N_btm.n348 0.228786
R32061 C9_N_btm.n348 C9_N_btm.n257 0.228786
R32062 C9_N_btm.n347 C9_N_btm.n346 0.228786
R32063 C9_N_btm.n346 C9_N_btm.n345 0.228786
R32064 C9_N_btm.n260 C9_N_btm.n257 0.228786
R32065 C9_N_btm.n343 C9_N_btm.n260 0.228786
R32066 C9_N_btm.n345 C9_N_btm.n344 0.228786
R32067 C9_N_btm.n344 C9_N_btm.n263 0.228786
R32068 C9_N_btm.n343 C9_N_btm.n342 0.228786
R32069 C9_N_btm.n342 C9_N_btm.n341 0.228786
R32070 C9_N_btm.n267 C9_N_btm.n263 0.228786
R32071 C9_N_btm.n339 C9_N_btm.n267 0.228786
R32072 C9_N_btm.n341 C9_N_btm.n340 0.228786
R32073 C9_N_btm.n340 C9_N_btm.n269 0.228786
R32074 C9_N_btm.n339 C9_N_btm.n338 0.228786
R32075 C9_N_btm.n338 C9_N_btm.n337 0.228786
R32076 C9_N_btm.n272 C9_N_btm.n269 0.228786
R32077 C9_N_btm.n335 C9_N_btm.n272 0.228786
R32078 C9_N_btm.n337 C9_N_btm.n336 0.228786
R32079 C9_N_btm.n336 C9_N_btm.n275 0.228786
R32080 C9_N_btm.n335 C9_N_btm.n334 0.228786
R32081 C9_N_btm.n334 C9_N_btm.n333 0.228786
R32082 C9_N_btm.n279 C9_N_btm.n275 0.228786
R32083 C9_N_btm.n302 C9_N_btm.n279 0.228786
R32084 C9_N_btm.n333 C9_N_btm.n332 0.228786
R32085 C9_N_btm.n278 C9_N_btm.n277 0.228786
R32086 C9_N_btm.n277 C9_N_btm.n276 0.228786
R32087 C9_N_btm.n330 C9_N_btm.n329 0.228786
R32088 C9_N_btm.n329 C9_N_btm.n328 0.228786
R32089 C9_N_btm.n327 C9_N_btm.n276 0.228786
R32090 C9_N_btm.n327 C9_N_btm.n326 0.228786
R32091 C9_N_btm.n328 C9_N_btm.n325 0.228786
R32092 C9_N_btm.n325 C9_N_btm.n324 0.228786
R32093 C9_N_btm.n326 C9_N_btm.n268 0.228786
R32094 C9_N_btm.n268 C9_N_btm.n266 0.228786
R32095 C9_N_btm.n324 C9_N_btm.n323 0.228786
R32096 C9_N_btm.n323 C9_N_btm.n322 0.228786
R32097 C9_N_btm.n266 C9_N_btm.n265 0.228786
R32098 C9_N_btm.n265 C9_N_btm.n264 0.228786
R32099 C9_N_btm.n322 C9_N_btm.n321 0.228786
R32100 C9_N_btm.n321 C9_N_btm.n320 0.228786
R32101 C9_N_btm.n319 C9_N_btm.n264 0.228786
R32102 C9_N_btm.n319 C9_N_btm.n318 0.228786
R32103 C9_N_btm.n320 C9_N_btm.n317 0.228786
R32104 C9_N_btm.n317 C9_N_btm.n316 0.228786
R32105 C9_N_btm.n318 C9_N_btm.n256 0.228786
R32106 C9_N_btm.n256 C9_N_btm.n254 0.228786
R32107 C9_N_btm.n316 C9_N_btm.n315 0.228786
R32108 C9_N_btm.n315 C9_N_btm.n314 0.228786
R32109 C9_N_btm.n254 C9_N_btm.n253 0.228786
R32110 C9_N_btm.n253 C9_N_btm.n252 0.228786
R32111 C9_N_btm.n314 C9_N_btm.n313 0.228786
R32112 C9_N_btm.n313 C9_N_btm.n312 0.228786
R32113 C9_N_btm.n311 C9_N_btm.n252 0.228786
R32114 C9_N_btm.n311 C9_N_btm.n310 0.228786
R32115 C9_N_btm.n312 C9_N_btm.n309 0.228786
R32116 C9_N_btm.n309 C9_N_btm.n308 0.228786
R32117 C9_N_btm.n310 C9_N_btm.n243 0.228786
R32118 C9_N_btm.n243 C9_N_btm.n241 0.228786
R32119 C9_N_btm.n308 C9_N_btm.n307 0.228786
R32120 C9_N_btm.n307 C9_N_btm.n306 0.228786
R32121 C9_N_btm.n241 C9_N_btm.n240 0.228786
R32122 C9_N_btm.n240 C9_N_btm.n239 0.228786
R32123 C9_N_btm.n306 C9_N_btm.n305 0.228786
R32124 C9_N_btm.n303 C9_N_btm.n239 0.228786
R32125 C9_N_btm.n359 C9_N_btm.n237 0.228786
R32126 C9_N_btm.n361 C9_N_btm.n360 0.228786
R32127 C9_N_btm.n235 C9_N_btm.n234 0.228786
R32128 C9_N_btm.n385 C9_N_btm.n384 0.228786
R32129 C9_N_btm.n383 C9_N_btm.n232 0.228786
R32130 C9_N_btm.n370 C9_N_btm.n365 0.228786
R32131 C9_N_btm.n374 C9_N_btm.n366 0.228786
R32132 C9_N_btm.n378 C9_N_btm.n375 0.228786
R32133 C9_N_btm.n377 C9_N_btm.n376 0.228786
R32134 C9_N_btm.n203 C9_N_btm.n202 0.228786
R32135 C9_N_btm.n401 C9_N_btm.n400 0.228786
R32136 C9_N_btm.n403 C9_N_btm.n402 0.228786
R32137 C9_N_btm.n199 C9_N_btm.n198 0.228786
R32138 C9_N_btm.n426 C9_N_btm.n425 0.228786
R32139 C9_N_btm.n427 C9_N_btm.n197 0.228786
R32140 C9_N_btm.n405 C9_N_btm.n195 0.228786
R32141 C9_N_btm.n420 C9_N_btm.n407 0.228786
R32142 C9_N_btm.n419 C9_N_btm.n418 0.228786
R32143 C9_N_btm.n413 C9_N_btm.n408 0.228786
R32144 C9_N_btm.n412 C9_N_btm.n411 0.228786
R32145 C9_N_btm.n168 C9_N_btm.n167 0.228786
R32146 C9_N_btm.n444 C9_N_btm.n443 0.228786
R32147 C9_N_btm.n165 C9_N_btm.n164 0.228786
R32148 C9_N_btm.n454 C9_N_btm.n453 0.228786
R32149 C9_N_btm.n455 C9_N_btm.n163 0.228786
R32150 C9_N_btm.n447 C9_N_btm.n161 0.228786
R32151 C9_N_btm.n144 C9_N_btm.n143 0.228786
R32152 C9_N_btm.n477 C9_N_btm.n476 0.228786
R32153 C9_N_btm.n145 C9_N_btm.n141 0.228786
R32154 C9_N_btm.n481 C9_N_btm.n49 0.228786
R32155 C9_N_btm.n148 C9_N_btm.n49 0.228786
R32156 C9_N_btm.n483 C9_N_btm.n47 0.228786
R32157 C9_N_btm.n467 C9_N_btm.n47 0.228786
R32158 C9_N_btm.n485 C9_N_btm.n45 0.228786
R32159 C9_N_btm.n466 C9_N_btm.n45 0.228786
R32160 C9_N_btm.n487 C9_N_btm.n41 0.228786
R32161 C9_N_btm.n41 C9_N_btm.n40 0.228786
R32162 C9_N_btm.n490 C9_N_btm.n489 0.228786
R32163 C9_N_btm.n491 C9_N_btm.n490 0.228786
R32164 C9_N_btm.n492 C9_N_btm.n39 0.228786
R32165 C9_N_btm.n493 C9_N_btm.n492 0.228786
R32166 C9_N_btm.n491 C9_N_btm.n36 0.228786
R32167 C9_N_btm.n36 C9_N_btm.n33 0.228786
R32168 C9_N_btm.n494 C9_N_btm.n493 0.228786
R32169 C9_N_btm.n495 C9_N_btm.n494 0.228786
R32170 C9_N_btm.n496 C9_N_btm.n33 0.228786
R32171 C9_N_btm.n497 C9_N_btm.n496 0.228786
R32172 C9_N_btm.n495 C9_N_btm.n32 0.228786
R32173 C9_N_btm.n32 C9_N_btm.n31 0.228786
R32174 C9_N_btm.n498 C9_N_btm.n497 0.228786
R32175 C9_N_btm.n499 C9_N_btm.n498 0.228786
R32176 C9_N_btm.n500 C9_N_btm.n31 0.228786
R32177 C9_N_btm.n501 C9_N_btm.n500 0.228786
R32178 C9_N_btm.n499 C9_N_btm.n28 0.228786
R32179 C9_N_btm.n28 C9_N_btm.n25 0.228786
R32180 C9_N_btm.n502 C9_N_btm.n501 0.228786
R32181 C9_N_btm.n503 C9_N_btm.n502 0.228786
R32182 C9_N_btm.n504 C9_N_btm.n25 0.228786
R32183 C9_N_btm.n505 C9_N_btm.n504 0.228786
R32184 C9_N_btm.n503 C9_N_btm.n24 0.228786
R32185 C9_N_btm.n24 C9_N_btm.n23 0.228786
R32186 C9_N_btm.n506 C9_N_btm.n505 0.228786
R32187 C9_N_btm.n507 C9_N_btm.n506 0.228786
R32188 C9_N_btm.n508 C9_N_btm.n23 0.228786
R32189 C9_N_btm.n509 C9_N_btm.n508 0.228786
R32190 C9_N_btm.n507 C9_N_btm.n20 0.228786
R32191 C9_N_btm.n20 C9_N_btm.n17 0.228786
R32192 C9_N_btm.n510 C9_N_btm.n509 0.228786
R32193 C9_N_btm.n511 C9_N_btm.n510 0.228786
R32194 C9_N_btm.n512 C9_N_btm.n17 0.228786
R32195 C9_N_btm.n513 C9_N_btm.n512 0.228786
R32196 C9_N_btm.n511 C9_N_btm.n16 0.228786
R32197 C9_N_btm.n104 C9_N_btm.n103 0.208893
R32198 C9_N_btm.n67 C9_N_btm.n66 0.208893
R32199 C9_N_btm.n302 C9_N_btm.n301 0.208893
R32200 C9_N_btm.n304 C9_N_btm.n236 0.208893
R32201 C9_N_btm.n424 C9_N_btm.n404 0.208893
R32202 C9_N_btm.n451 C9_N_btm.n450 0.208893
R32203 C9_N_btm.n185 C9_N_btm.n184 0.208893
R32204 C9_N_btm.n434 C9_N_btm.n188 0.208893
R32205 C9_N_btm.n332 C9_N_btm.n331 0.208893
R32206 C9_N_btm.n102 C9_N_btm.n16 0.09425
R32207 C9_N_btm.n103 C9_N_btm.n102 0.09425
R32208 C9_N_btm.n101 C9_N_btm.n18 0.09425
R32209 C9_N_btm.n105 C9_N_btm.n101 0.09425
R32210 C9_N_btm.n107 C9_N_btm.n98 0.09425
R32211 C9_N_btm.n106 C9_N_btm.n99 0.09425
R32212 C9_N_btm.n106 C9_N_btm.n100 0.09425
R32213 C9_N_btm.n94 C9_N_btm.n21 0.09425
R32214 C9_N_btm.n107 C9_N_btm.n94 0.09425
R32215 C9_N_btm.n510 C9_N_btm.n19 0.09425
R32216 C9_N_btm.n99 C9_N_btm.n19 0.09425
R32217 C9_N_btm.n508 C9_N_btm.n22 0.09425
R32218 C9_N_btm.n109 C9_N_btm.n22 0.09425
R32219 C9_N_btm.n111 C9_N_btm.n110 0.09425
R32220 C9_N_btm.n110 C9_N_btm.n93 0.09425
R32221 C9_N_btm.n109 C9_N_btm.n108 0.09425
R32222 C9_N_btm.n108 C9_N_btm.n97 0.09425
R32223 C9_N_btm.n96 C9_N_btm.n93 0.09425
R32224 C9_N_btm.n115 C9_N_btm.n91 0.09425
R32225 C9_N_btm.n113 C9_N_btm.n92 0.09425
R32226 C9_N_btm.n95 C9_N_btm.n92 0.09425
R32227 C9_N_btm.n114 C9_N_btm.n26 0.09425
R32228 C9_N_btm.n115 C9_N_btm.n114 0.09425
R32229 C9_N_btm.n112 C9_N_btm.n24 0.09425
R32230 C9_N_btm.n113 C9_N_btm.n112 0.09425
R32231 C9_N_btm.n502 C9_N_btm.n27 0.09425
R32232 C9_N_btm.n89 C9_N_btm.n27 0.09425
R32233 C9_N_btm.n88 C9_N_btm.n29 0.09425
R32234 C9_N_btm.n117 C9_N_btm.n88 0.09425
R32235 C9_N_btm.n116 C9_N_btm.n89 0.09425
R32236 C9_N_btm.n116 C9_N_btm.n90 0.09425
R32237 C9_N_btm.n117 C9_N_btm.n82 0.09425
R32238 C9_N_btm.n120 C9_N_btm.n81 0.09425
R32239 C9_N_btm.n118 C9_N_btm.n87 0.09425
R32240 C9_N_btm.n119 C9_N_btm.n118 0.09425
R32241 C9_N_btm.n86 C9_N_btm.n83 0.09425
R32242 C9_N_btm.n86 C9_N_btm.n81 0.09425
R32243 C9_N_btm.n500 C9_N_btm.n30 0.09425
R32244 C9_N_btm.n87 C9_N_btm.n30 0.09425
R32245 C9_N_btm.n84 C9_N_btm.n32 0.09425
R32246 C9_N_btm.n85 C9_N_btm.n84 0.09425
R32247 C9_N_btm.n79 C9_N_btm.n34 0.09425
R32248 C9_N_btm.n123 C9_N_btm.n79 0.09425
R32249 C9_N_btm.n85 C9_N_btm.n80 0.09425
R32250 C9_N_btm.n121 C9_N_btm.n80 0.09425
R32251 C9_N_btm.n123 C9_N_btm.n122 0.09425
R32252 C9_N_btm.n125 C9_N_btm.n76 0.09425
R32253 C9_N_btm.n124 C9_N_btm.n77 0.09425
R32254 C9_N_btm.n124 C9_N_btm.n78 0.09425
R32255 C9_N_btm.n57 C9_N_btm.n37 0.09425
R32256 C9_N_btm.n125 C9_N_btm.n57 0.09425
R32257 C9_N_btm.n494 C9_N_btm.n35 0.09425
R32258 C9_N_btm.n77 C9_N_btm.n35 0.09425
R32259 C9_N_btm.n492 C9_N_btm.n38 0.09425
R32260 C9_N_btm.n127 C9_N_btm.n38 0.09425
R32261 C9_N_btm.n129 C9_N_btm.n128 0.09425
R32262 C9_N_btm.n128 C9_N_btm.n56 0.09425
R32263 C9_N_btm.n127 C9_N_btm.n126 0.09425
R32264 C9_N_btm.n126 C9_N_btm.n75 0.09425
R32265 C9_N_btm.n74 C9_N_btm.n56 0.09425
R32266 C9_N_btm.n71 C9_N_btm.n58 0.09425
R32267 C9_N_btm.n72 C9_N_btm.n55 0.09425
R32268 C9_N_btm.n73 C9_N_btm.n72 0.09425
R32269 C9_N_btm.n131 C9_N_btm.n54 0.09425
R32270 C9_N_btm.n71 C9_N_btm.n54 0.09425
R32271 C9_N_btm.n130 C9_N_btm.n42 0.09425
R32272 C9_N_btm.n130 C9_N_btm.n55 0.09425
R32273 C9_N_btm.n488 C9_N_btm.n43 0.09425
R32274 C9_N_btm.n131 C9_N_btm.n43 0.09425
R32275 C9_N_btm.n484 C9_N_btm.n46 0.09425
R32276 C9_N_btm.n135 C9_N_btm.n46 0.09425
R32277 C9_N_btm.n486 C9_N_btm.n44 0.09425
R32278 C9_N_btm.n133 C9_N_btm.n44 0.09425
R32279 C9_N_btm.n135 C9_N_btm.n134 0.09425
R32280 C9_N_btm.n134 C9_N_btm.n52 0.09425
R32281 C9_N_btm.n133 C9_N_btm.n132 0.09425
R32282 C9_N_btm.n132 C9_N_btm.n53 0.09425
R32283 C9_N_btm.n60 C9_N_btm.n52 0.09425
R32284 C9_N_btm.n69 C9_N_btm.n60 0.09425
R32285 C9_N_btm.n70 C9_N_btm.n53 0.09425
R32286 C9_N_btm.n70 C9_N_btm.n59 0.09425
R32287 C9_N_btm.n69 C9_N_btm.n68 0.09425
R32288 C9_N_btm.n65 C9_N_btm.n61 0.09425
R32289 C9_N_btm.n66 C9_N_btm.n63 0.09425
R32290 C9_N_btm.n64 C9_N_btm.n51 0.09425
R32291 C9_N_btm.n65 C9_N_btm.n64 0.09425
R32292 C9_N_btm.n62 C9_N_btm.n50 0.09425
R32293 C9_N_btm.n63 C9_N_btm.n62 0.09425
R32294 C9_N_btm.n137 C9_N_btm.n136 0.09425
R32295 C9_N_btm.n136 C9_N_btm.n51 0.09425
R32296 C9_N_btm.n139 C9_N_btm.n138 0.09425
R32297 C9_N_btm.n138 C9_N_btm.n50 0.09425
R32298 C9_N_btm.n482 C9_N_btm.n48 0.09425
R32299 C9_N_btm.n137 C9_N_btm.n48 0.09425
R32300 C9_N_btm.n140 C9_N_btm.n139 0.09425
R32301 C9_N_btm.n480 C9_N_btm.n140 0.09425
R32302 C9_N_btm.n448 C9_N_btm.n143 0.09425
R32303 C9_N_btm.n148 C9_N_btm.n47 0.09425
R32304 C9_N_btm.n467 C9_N_btm.n45 0.09425
R32305 C9_N_btm.n466 C9_N_btm.n41 0.09425
R32306 C9_N_btm.n490 C9_N_btm.n40 0.09425
R32307 C9_N_btm.n465 C9_N_btm.n40 0.09425
R32308 C9_N_btm.n469 C9_N_btm.n465 0.09425
R32309 C9_N_btm.n464 C9_N_btm.n463 0.09425
R32310 C9_N_btm.n471 C9_N_btm.n464 0.09425
R32311 C9_N_btm.n472 C9_N_btm.n150 0.09425
R32312 C9_N_btm.n472 C9_N_btm.n151 0.09425
R32313 C9_N_btm.n471 C9_N_btm.n470 0.09425
R32314 C9_N_btm.n470 C9_N_btm.n469 0.09425
R32315 C9_N_btm.n468 C9_N_btm.n151 0.09425
R32316 C9_N_btm.n468 C9_N_btm.n466 0.09425
R32317 C9_N_btm.n473 C9_N_btm.n149 0.09425
R32318 C9_N_btm.n467 C9_N_btm.n149 0.09425
R32319 C9_N_btm.n145 C9_N_btm.n49 0.09425
R32320 C9_N_btm.n476 C9_N_btm.n144 0.09425
R32321 C9_N_btm.n476 C9_N_btm.n145 0.09425
R32322 C9_N_btm.n475 C9_N_btm.n474 0.09425
R32323 C9_N_btm.n474 C9_N_btm.n148 0.09425
R32324 C9_N_btm.n154 C9_N_btm.n147 0.09425
R32325 C9_N_btm.n473 C9_N_btm.n147 0.09425
R32326 C9_N_btm.n461 C9_N_btm.n152 0.09425
R32327 C9_N_btm.n152 C9_N_btm.n150 0.09425
R32328 C9_N_btm.n462 C9_N_btm.n153 0.09425
R32329 C9_N_btm.n463 C9_N_btm.n462 0.09425
R32330 C9_N_btm.n460 C9_N_btm.n156 0.09425
R32331 C9_N_btm.n461 C9_N_btm.n460 0.09425
R32332 C9_N_btm.n177 C9_N_btm.n176 0.09425
R32333 C9_N_btm.n176 C9_N_btm.n153 0.09425
R32334 C9_N_btm.n183 C9_N_btm.n178 0.09425
R32335 C9_N_btm.n178 C9_N_btm.n156 0.09425
R32336 C9_N_btm.n184 C9_N_btm.n177 0.09425
R32337 C9_N_btm.n183 C9_N_btm.n175 0.09425
R32338 C9_N_btm.n438 C9_N_btm.n437 0.09425
R32339 C9_N_btm.n437 C9_N_btm.n436 0.09425
R32340 C9_N_btm.n436 C9_N_btm.n435 0.09425
R32341 C9_N_btm.n432 C9_N_btm.n190 0.09425
R32342 C9_N_btm.n433 C9_N_btm.n432 0.09425
R32343 C9_N_btm.n212 C9_N_btm.n188 0.09425
R32344 C9_N_btm.n213 C9_N_btm.n212 0.09425
R32345 C9_N_btm.n213 C9_N_btm.n210 0.09425
R32346 C9_N_btm.n222 C9_N_btm.n210 0.09425
R32347 C9_N_btm.n223 C9_N_btm.n222 0.09425
R32348 C9_N_btm.n395 C9_N_btm.n223 0.09425
R32349 C9_N_btm.n395 C9_N_btm.n394 0.09425
R32350 C9_N_btm.n394 C9_N_btm.n393 0.09425
R32351 C9_N_btm.n393 C9_N_btm.n392 0.09425
R32352 C9_N_btm.n392 C9_N_btm.n391 0.09425
R32353 C9_N_btm.n332 C9_N_btm.n302 0.09425
R32354 C9_N_btm.n300 C9_N_btm.n279 0.09425
R32355 C9_N_btm.n299 C9_N_btm.n298 0.09425
R32356 C9_N_btm.n336 C9_N_btm.n274 0.09425
R32357 C9_N_btm.n297 C9_N_btm.n274 0.09425
R32358 C9_N_btm.n296 C9_N_btm.n273 0.09425
R32359 C9_N_btm.n338 C9_N_btm.n271 0.09425
R32360 C9_N_btm.n295 C9_N_btm.n271 0.09425
R32361 C9_N_btm.n294 C9_N_btm.n270 0.09425
R32362 C9_N_btm.n292 C9_N_btm.n267 0.09425
R32363 C9_N_btm.n293 C9_N_btm.n292 0.09425
R32364 C9_N_btm.n291 C9_N_btm.n290 0.09425
R32365 C9_N_btm.n344 C9_N_btm.n262 0.09425
R32366 C9_N_btm.n289 C9_N_btm.n262 0.09425
R32367 C9_N_btm.n288 C9_N_btm.n261 0.09425
R32368 C9_N_btm.n346 C9_N_btm.n259 0.09425
R32369 C9_N_btm.n287 C9_N_btm.n259 0.09425
R32370 C9_N_btm.n286 C9_N_btm.n258 0.09425
R32371 C9_N_btm.n284 C9_N_btm.n255 0.09425
R32372 C9_N_btm.n285 C9_N_btm.n284 0.09425
R32373 C9_N_btm.n283 C9_N_btm.n282 0.09425
R32374 C9_N_btm.n280 C9_N_btm.n249 0.09425
R32375 C9_N_btm.n352 C9_N_btm.n250 0.09425
R32376 C9_N_btm.n281 C9_N_btm.n250 0.09425
R32377 C9_N_btm.n354 C9_N_btm.n247 0.09425
R32378 C9_N_btm.n247 C9_N_btm.n227 0.09425
R32379 C9_N_btm.n246 C9_N_btm.n228 0.09425
R32380 C9_N_btm.n389 C9_N_btm.n228 0.09425
R32381 C9_N_btm.n390 C9_N_btm.n227 0.09425
R32382 C9_N_btm.n391 C9_N_btm.n390 0.09425
R32383 C9_N_btm.n388 C9_N_btm.n229 0.09425
R32384 C9_N_btm.n388 C9_N_btm.n230 0.09425
R32385 C9_N_btm.n389 C9_N_btm.n226 0.09425
R32386 C9_N_btm.n226 C9_N_btm.n225 0.09425
R32387 C9_N_btm.n372 C9_N_btm.n230 0.09425
R32388 C9_N_btm.n372 C9_N_btm.n371 0.09425
R32389 C9_N_btm.n225 C9_N_btm.n224 0.09425
R32390 C9_N_btm.n224 C9_N_btm.n208 0.09425
R32391 C9_N_btm.n371 C9_N_btm.n207 0.09425
R32392 C9_N_btm.n397 C9_N_btm.n207 0.09425
R32393 C9_N_btm.n396 C9_N_btm.n208 0.09425
R32394 C9_N_btm.n396 C9_N_btm.n209 0.09425
R32395 C9_N_btm.n397 C9_N_btm.n205 0.09425
R32396 C9_N_btm.n220 C9_N_btm.n205 0.09425
R32397 C9_N_btm.n221 C9_N_btm.n209 0.09425
R32398 C9_N_btm.n221 C9_N_btm.n211 0.09425
R32399 C9_N_btm.n220 C9_N_btm.n219 0.09425
R32400 C9_N_btm.n219 C9_N_btm.n215 0.09425
R32401 C9_N_btm.n214 C9_N_btm.n211 0.09425
R32402 C9_N_btm.n214 C9_N_btm.n190 0.09425
R32403 C9_N_btm.n218 C9_N_btm.n216 0.09425
R32404 C9_N_btm.n216 C9_N_btm.n192 0.09425
R32405 C9_N_btm.n215 C9_N_btm.n191 0.09425
R32406 C9_N_btm.n431 C9_N_btm.n191 0.09425
R32407 C9_N_btm.n430 C9_N_btm.n192 0.09425
R32408 C9_N_btm.n430 C9_N_btm.n193 0.09425
R32409 C9_N_btm.n431 C9_N_btm.n189 0.09425
R32410 C9_N_btm.n189 C9_N_btm.n187 0.09425
R32411 C9_N_btm.n416 C9_N_btm.n193 0.09425
R32412 C9_N_btm.n416 C9_N_btm.n415 0.09425
R32413 C9_N_btm.n187 C9_N_btm.n186 0.09425
R32414 C9_N_btm.n186 C9_N_btm.n173 0.09425
R32415 C9_N_btm.n415 C9_N_btm.n172 0.09425
R32416 C9_N_btm.n440 C9_N_btm.n172 0.09425
R32417 C9_N_btm.n439 C9_N_btm.n173 0.09425
R32418 C9_N_btm.n439 C9_N_btm.n174 0.09425
R32419 C9_N_btm.n440 C9_N_btm.n170 0.09425
R32420 C9_N_btm.n181 C9_N_btm.n170 0.09425
R32421 C9_N_btm.n182 C9_N_btm.n174 0.09425
R32422 C9_N_btm.n182 C9_N_btm.n179 0.09425
R32423 C9_N_btm.n181 C9_N_btm.n180 0.09425
R32424 C9_N_btm.n180 C9_N_btm.n158 0.09425
R32425 C9_N_btm.n179 C9_N_btm.n157 0.09425
R32426 C9_N_btm.n459 C9_N_btm.n157 0.09425
R32427 C9_N_btm.n458 C9_N_btm.n158 0.09425
R32428 C9_N_btm.n458 C9_N_btm.n159 0.09425
R32429 C9_N_btm.n459 C9_N_btm.n155 0.09425
R32430 C9_N_btm.n155 C9_N_btm.n154 0.09425
R32431 C9_N_btm.n159 C9_N_btm.n146 0.09425
R32432 C9_N_btm.n475 C9_N_btm.n146 0.09425
R32433 C9_N_btm.n457 C9_N_btm.n160 0.09425
R32434 C9_N_btm.n160 C9_N_btm.n144 0.09425
R32435 C9_N_btm.n455 C9_N_btm.n161 0.09425
R32436 C9_N_btm.n448 C9_N_btm.n161 0.09425
R32437 C9_N_btm.n456 C9_N_btm.n162 0.09425
R32438 C9_N_btm.n457 C9_N_btm.n456 0.09425
R32439 C9_N_btm.n454 C9_N_btm.n164 0.09425
R32440 C9_N_btm.n455 C9_N_btm.n454 0.09425
R32441 C9_N_btm.n442 C9_N_btm.n169 0.09425
R32442 C9_N_btm.n169 C9_N_btm.n162 0.09425
R32443 C9_N_btm.n443 C9_N_btm.n168 0.09425
R32444 C9_N_btm.n443 C9_N_btm.n164 0.09425
R32445 C9_N_btm.n441 C9_N_btm.n171 0.09425
R32446 C9_N_btm.n442 C9_N_btm.n441 0.09425
R32447 C9_N_btm.n413 C9_N_btm.n412 0.09425
R32448 C9_N_btm.n412 C9_N_btm.n168 0.09425
R32449 C9_N_btm.n417 C9_N_btm.n414 0.09425
R32450 C9_N_btm.n414 C9_N_btm.n171 0.09425
R32451 C9_N_btm.n418 C9_N_btm.n407 0.09425
R32452 C9_N_btm.n418 C9_N_btm.n413 0.09425
R32453 C9_N_btm.n429 C9_N_btm.n194 0.09425
R32454 C9_N_btm.n417 C9_N_btm.n194 0.09425
R32455 C9_N_btm.n427 C9_N_btm.n195 0.09425
R32456 C9_N_btm.n407 C9_N_btm.n195 0.09425
R32457 C9_N_btm.n428 C9_N_btm.n196 0.09425
R32458 C9_N_btm.n429 C9_N_btm.n428 0.09425
R32459 C9_N_btm.n402 C9_N_btm.n198 0.09425
R32460 C9_N_btm.n426 C9_N_btm.n198 0.09425
R32461 C9_N_btm.n427 C9_N_btm.n426 0.09425
R32462 C9_N_btm.n217 C9_N_btm.n201 0.09425
R32463 C9_N_btm.n217 C9_N_btm.n196 0.09425
R32464 C9_N_btm.n399 C9_N_btm.n204 0.09425
R32465 C9_N_btm.n218 C9_N_btm.n204 0.09425
R32466 C9_N_btm.n400 C9_N_btm.n203 0.09425
R32467 C9_N_btm.n400 C9_N_btm.n201 0.09425
R32468 C9_N_btm.n398 C9_N_btm.n206 0.09425
R32469 C9_N_btm.n399 C9_N_btm.n398 0.09425
R32470 C9_N_btm.n376 C9_N_btm.n375 0.09425
R32471 C9_N_btm.n376 C9_N_btm.n203 0.09425
R32472 C9_N_btm.n373 C9_N_btm.n369 0.09425
R32473 C9_N_btm.n369 C9_N_btm.n206 0.09425
R32474 C9_N_btm.n374 C9_N_btm.n370 0.09425
R32475 C9_N_btm.n375 C9_N_btm.n374 0.09425
R32476 C9_N_btm.n387 C9_N_btm.n231 0.09425
R32477 C9_N_btm.n373 C9_N_btm.n231 0.09425
R32478 C9_N_btm.n385 C9_N_btm.n234 0.09425
R32479 C9_N_btm.n385 C9_N_btm.n232 0.09425
R32480 C9_N_btm.n370 C9_N_btm.n232 0.09425
R32481 C9_N_btm.n386 C9_N_btm.n233 0.09425
R32482 C9_N_btm.n387 C9_N_btm.n386 0.09425
R32483 C9_N_btm.n245 C9_N_btm.n242 0.09425
R32484 C9_N_btm.n245 C9_N_btm.n229 0.09425
R32485 C9_N_btm.n360 C9_N_btm.n234 0.09425
R32486 C9_N_btm.n359 C9_N_btm.n239 0.09425
R32487 C9_N_btm.n360 C9_N_btm.n359 0.09425
R32488 C9_N_btm.n358 C9_N_btm.n238 0.09425
R32489 C9_N_btm.n238 C9_N_btm.n233 0.09425
R32490 C9_N_btm.n357 C9_N_btm.n241 0.09425
R32491 C9_N_btm.n357 C9_N_btm.n242 0.09425
R32492 C9_N_btm.n356 C9_N_btm.n355 0.09425
R32493 C9_N_btm.n355 C9_N_btm.n246 0.09425
R32494 C9_N_btm.n310 C9_N_btm.n244 0.09425
R32495 C9_N_btm.n354 C9_N_btm.n244 0.09425
R32496 C9_N_btm.n353 C9_N_btm.n248 0.09425
R32497 C9_N_btm.n353 C9_N_btm.n249 0.09425
R32498 C9_N_btm.n351 C9_N_btm.n252 0.09425
R32499 C9_N_btm.n352 C9_N_btm.n351 0.09425
R32500 C9_N_btm.n350 C9_N_btm.n251 0.09425
R32501 C9_N_btm.n283 C9_N_btm.n251 0.09425
R32502 C9_N_btm.n349 C9_N_btm.n254 0.09425
R32503 C9_N_btm.n349 C9_N_btm.n255 0.09425
R32504 C9_N_btm.n348 C9_N_btm.n347 0.09425
R32505 C9_N_btm.n347 C9_N_btm.n258 0.09425
R32506 C9_N_btm.n318 C9_N_btm.n257 0.09425
R32507 C9_N_btm.n346 C9_N_btm.n257 0.09425
R32508 C9_N_btm.n345 C9_N_btm.n260 0.09425
R32509 C9_N_btm.n345 C9_N_btm.n261 0.09425
R32510 C9_N_btm.n343 C9_N_btm.n264 0.09425
R32511 C9_N_btm.n344 C9_N_btm.n343 0.09425
R32512 C9_N_btm.n342 C9_N_btm.n263 0.09425
R32513 C9_N_btm.n291 C9_N_btm.n263 0.09425
R32514 C9_N_btm.n341 C9_N_btm.n266 0.09425
R32515 C9_N_btm.n341 C9_N_btm.n267 0.09425
R32516 C9_N_btm.n340 C9_N_btm.n339 0.09425
R32517 C9_N_btm.n339 C9_N_btm.n270 0.09425
R32518 C9_N_btm.n326 C9_N_btm.n269 0.09425
R32519 C9_N_btm.n338 C9_N_btm.n269 0.09425
R32520 C9_N_btm.n337 C9_N_btm.n272 0.09425
R32521 C9_N_btm.n337 C9_N_btm.n273 0.09425
R32522 C9_N_btm.n335 C9_N_btm.n276 0.09425
R32523 C9_N_btm.n336 C9_N_btm.n335 0.09425
R32524 C9_N_btm.n334 C9_N_btm.n275 0.09425
R32525 C9_N_btm.n299 C9_N_btm.n275 0.09425
R32526 C9_N_btm.n333 C9_N_btm.n278 0.09425
R32527 C9_N_btm.n333 C9_N_btm.n279 0.09425
R32528 C9_N_btm.n330 C9_N_btm.n277 0.09425
R32529 C9_N_btm.n334 C9_N_btm.n277 0.09425
R32530 C9_N_btm.n329 C9_N_btm.n276 0.09425
R32531 C9_N_btm.n328 C9_N_btm.n327 0.09425
R32532 C9_N_btm.n327 C9_N_btm.n272 0.09425
R32533 C9_N_btm.n326 C9_N_btm.n325 0.09425
R32534 C9_N_btm.n324 C9_N_btm.n268 0.09425
R32535 C9_N_btm.n340 C9_N_btm.n268 0.09425
R32536 C9_N_btm.n323 C9_N_btm.n266 0.09425
R32537 C9_N_btm.n322 C9_N_btm.n265 0.09425
R32538 C9_N_btm.n342 C9_N_btm.n265 0.09425
R32539 C9_N_btm.n321 C9_N_btm.n264 0.09425
R32540 C9_N_btm.n320 C9_N_btm.n319 0.09425
R32541 C9_N_btm.n319 C9_N_btm.n260 0.09425
R32542 C9_N_btm.n318 C9_N_btm.n317 0.09425
R32543 C9_N_btm.n316 C9_N_btm.n256 0.09425
R32544 C9_N_btm.n348 C9_N_btm.n256 0.09425
R32545 C9_N_btm.n315 C9_N_btm.n254 0.09425
R32546 C9_N_btm.n314 C9_N_btm.n253 0.09425
R32547 C9_N_btm.n350 C9_N_btm.n253 0.09425
R32548 C9_N_btm.n313 C9_N_btm.n252 0.09425
R32549 C9_N_btm.n312 C9_N_btm.n311 0.09425
R32550 C9_N_btm.n311 C9_N_btm.n248 0.09425
R32551 C9_N_btm.n310 C9_N_btm.n309 0.09425
R32552 C9_N_btm.n308 C9_N_btm.n243 0.09425
R32553 C9_N_btm.n356 C9_N_btm.n243 0.09425
R32554 C9_N_btm.n307 C9_N_btm.n241 0.09425
R32555 C9_N_btm.n306 C9_N_btm.n240 0.09425
R32556 C9_N_btm.n358 C9_N_btm.n240 0.09425
R32557 C9_N_btm.n305 C9_N_btm.n239 0.09425
R32558 C9_N_btm.n303 C9_N_btm.n237 0.09425
R32559 C9_N_btm.n361 C9_N_btm.n237 0.09425
R32560 C9_N_btm.n362 C9_N_btm.n236 0.09425
R32561 C9_N_btm.n363 C9_N_btm.n362 0.09425
R32562 C9_N_btm.n361 C9_N_btm.n235 0.09425
R32563 C9_N_btm.n384 C9_N_btm.n235 0.09425
R32564 C9_N_btm.n364 C9_N_btm.n363 0.09425
R32565 C9_N_btm.n382 C9_N_btm.n364 0.09425
R32566 C9_N_btm.n384 C9_N_btm.n383 0.09425
R32567 C9_N_btm.n383 C9_N_btm.n365 0.09425
R32568 C9_N_btm.n382 C9_N_btm.n381 0.09425
R32569 C9_N_btm.n381 C9_N_btm.n380 0.09425
R32570 C9_N_btm.n366 C9_N_btm.n365 0.09425
R32571 C9_N_btm.n378 C9_N_btm.n366 0.09425
R32572 C9_N_btm.n380 C9_N_btm.n379 0.09425
R32573 C9_N_btm.n379 C9_N_btm.n368 0.09425
R32574 C9_N_btm.n378 C9_N_btm.n377 0.09425
R32575 C9_N_btm.n377 C9_N_btm.n202 0.09425
R32576 C9_N_btm.n368 C9_N_btm.n367 0.09425
R32577 C9_N_btm.n367 C9_N_btm.n200 0.09425
R32578 C9_N_btm.n401 C9_N_btm.n202 0.09425
R32579 C9_N_btm.n402 C9_N_btm.n401 0.09425
R32580 C9_N_btm.n403 C9_N_btm.n200 0.09425
R32581 C9_N_btm.n425 C9_N_btm.n199 0.09425
R32582 C9_N_btm.n425 C9_N_btm.n197 0.09425
R32583 C9_N_btm.n424 C9_N_btm.n423 0.09425
R32584 C9_N_btm.n423 C9_N_btm.n422 0.09425
R32585 C9_N_btm.n405 C9_N_btm.n197 0.09425
R32586 C9_N_btm.n420 C9_N_btm.n405 0.09425
R32587 C9_N_btm.n422 C9_N_btm.n421 0.09425
R32588 C9_N_btm.n421 C9_N_btm.n406 0.09425
R32589 C9_N_btm.n420 C9_N_btm.n419 0.09425
R32590 C9_N_btm.n419 C9_N_btm.n408 0.09425
R32591 C9_N_btm.n409 C9_N_btm.n406 0.09425
R32592 C9_N_btm.n410 C9_N_btm.n409 0.09425
R32593 C9_N_btm.n411 C9_N_btm.n408 0.09425
R32594 C9_N_btm.n411 C9_N_btm.n167 0.09425
R32595 C9_N_btm.n410 C9_N_btm.n166 0.09425
R32596 C9_N_btm.n445 C9_N_btm.n166 0.09425
R32597 C9_N_btm.n444 C9_N_btm.n167 0.09425
R32598 C9_N_btm.n444 C9_N_btm.n165 0.09425
R32599 C9_N_btm.n446 C9_N_btm.n445 0.09425
R32600 C9_N_btm.n452 C9_N_btm.n446 0.09425
R32601 C9_N_btm.n453 C9_N_btm.n165 0.09425
R32602 C9_N_btm.n453 C9_N_btm.n163 0.09425
R32603 C9_N_btm.n452 C9_N_btm.n451 0.09425
R32604 C9_N_btm.n447 C9_N_btm.n163 0.09425
R32605 C9_N_btm.n449 C9_N_btm.n142 0.09425
R32606 C9_N_btm.n478 C9_N_btm.n142 0.09425
R32607 C9_N_btm.n477 C9_N_btm.n143 0.09425
R32608 C9_N_btm.n477 C9_N_btm.n141 0.09425
R32609 C9_N_btm.n479 C9_N_btm.n478 0.09425
R32610 C9_N_btm.n480 C9_N_btm.n479 0.09425
R32611 C9_N_btm.n481 C9_N_btm.n141 0.09425
R32612 C9_N_btm.n482 C9_N_btm.n481 0.09425
R32613 C9_N_btm.n483 C9_N_btm.n49 0.09425
R32614 C9_N_btm.n484 C9_N_btm.n483 0.09425
R32615 C9_N_btm.n485 C9_N_btm.n47 0.09425
R32616 C9_N_btm.n486 C9_N_btm.n485 0.09425
R32617 C9_N_btm.n487 C9_N_btm.n45 0.09425
R32618 C9_N_btm.n488 C9_N_btm.n487 0.09425
R32619 C9_N_btm.n489 C9_N_btm.n41 0.09425
R32620 C9_N_btm.n489 C9_N_btm.n42 0.09425
R32621 C9_N_btm.n490 C9_N_btm.n39 0.09425
R32622 C9_N_btm.n129 C9_N_btm.n39 0.09425
R32623 C9_N_btm.n492 C9_N_btm.n491 0.09425
R32624 C9_N_btm.n493 C9_N_btm.n36 0.09425
R32625 C9_N_btm.n493 C9_N_btm.n37 0.09425
R32626 C9_N_btm.n494 C9_N_btm.n33 0.09425
R32627 C9_N_btm.n496 C9_N_btm.n495 0.09425
R32628 C9_N_btm.n495 C9_N_btm.n34 0.09425
R32629 C9_N_btm.n497 C9_N_btm.n32 0.09425
R32630 C9_N_btm.n498 C9_N_btm.n31 0.09425
R32631 C9_N_btm.n83 C9_N_btm.n31 0.09425
R32632 C9_N_btm.n500 C9_N_btm.n499 0.09425
R32633 C9_N_btm.n501 C9_N_btm.n28 0.09425
R32634 C9_N_btm.n501 C9_N_btm.n29 0.09425
R32635 C9_N_btm.n502 C9_N_btm.n25 0.09425
R32636 C9_N_btm.n504 C9_N_btm.n503 0.09425
R32637 C9_N_btm.n503 C9_N_btm.n26 0.09425
R32638 C9_N_btm.n505 C9_N_btm.n24 0.09425
R32639 C9_N_btm.n506 C9_N_btm.n23 0.09425
R32640 C9_N_btm.n111 C9_N_btm.n23 0.09425
R32641 C9_N_btm.n508 C9_N_btm.n507 0.09425
R32642 C9_N_btm.n509 C9_N_btm.n20 0.09425
R32643 C9_N_btm.n509 C9_N_btm.n21 0.09425
R32644 C9_N_btm.n510 C9_N_btm.n17 0.09425
R32645 C9_N_btm.n512 C9_N_btm.n511 0.09425
R32646 C9_N_btm.n511 C9_N_btm.n18 0.09425
R32647 C9_N_btm.n513 C9_N_btm.n16 0.09425
R32648 C9_N_btm.n438 C9_N_btm.n185 0.047875
R32649 C9_N_btm.n435 C9_N_btm.n434 0.047875
R32650 C9_N_btm.n404 C9_N_btm.n403 0.047875
R32651 C9_N_btm.n450 C9_N_btm.n449 0.047875
R32652 C9_N_btm.n105 C9_N_btm.n104 0.0342289
R32653 C9_N_btm.n67 C9_N_btm.n61 0.0342289
R32654 C9_N_btm.n185 C9_N_btm.n175 0.0342289
R32655 C9_N_btm.n434 C9_N_btm.n433 0.0342289
R32656 C9_N_btm.n301 C9_N_btm.n300 0.0342289
R32657 C9_N_btm.n331 C9_N_btm.n278 0.0342289
R32658 C9_N_btm.n304 C9_N_btm.n303 0.0342289
R32659 C9_N_btm.n404 C9_N_btm.n199 0.0342289
R32660 C9_N_btm.n450 C9_N_btm.n447 0.0342289
R32661 a_17538_32519.n1 a_17538_32519.t4 1415.15
R32662 a_17538_32519.n1 a_17538_32519.t5 1320.68
R32663 a_17538_32519.n3 a_17538_32519.n2 296.139
R32664 a_17538_32519.n2 a_17538_32519.n1 280.685
R32665 a_17538_32519.n2 a_17538_32519.n0 269.182
R32666 a_17538_32519.t1 a_17538_32519.n3 26.5955
R32667 a_17538_32519.n3 a_17538_32519.t0 26.5955
R32668 a_17538_32519.n0 a_17538_32519.t2 24.9236
R32669 a_17538_32519.n0 a_17538_32519.t3 24.9236
R32670 a_20205_31679.n1 a_20205_31679.t4 601.154
R32671 a_20205_31679.n2 a_20205_31679.n1 287.752
R32672 a_20205_31679.n1 a_20205_31679.n0 277.568
R32673 a_20205_31679.t1 a_20205_31679.n2 26.5955
R32674 a_20205_31679.n2 a_20205_31679.t0 26.5955
R32675 a_20205_31679.n0 a_20205_31679.t2 24.9236
R32676 a_20205_31679.n0 a_20205_31679.t3 24.9236
R32677 a_n3420_39616.n4 a_n3420_39616.t11 1415.15
R32678 a_n3420_39616.n4 a_n3420_39616.t10 1320.68
R32679 a_n3420_39616.n8 a_n3420_39616.n7 360.399
R32680 a_n3420_39616.n5 a_n3420_39616.n4 245.97
R32681 a_n3420_39616.n3 a_n3420_39616.t9 241.536
R32682 a_n3420_39616.n2 a_n3420_39616.n1 232.862
R32683 a_n3420_39616.n9 a_n3420_39616.n8 203.161
R32684 a_n3420_39616.n3 a_n3420_39616.t8 169.237
R32685 a_n3420_39616.n5 a_n3420_39616.n3 166.983
R32686 a_n3420_39616.n2 a_n3420_39616.n0 95.6721
R32687 a_n3420_39616.n6 a_n3420_39616.n2 60.5918
R32688 a_n3420_39616.n7 a_n3420_39616.t2 27.5805
R32689 a_n3420_39616.n7 a_n3420_39616.t1 27.5805
R32690 a_n3420_39616.n9 a_n3420_39616.t0 27.5805
R32691 a_n3420_39616.t3 a_n3420_39616.n9 27.5805
R32692 a_n3420_39616.n1 a_n3420_39616.t7 25.8467
R32693 a_n3420_39616.n1 a_n3420_39616.t4 25.8467
R32694 a_n3420_39616.n0 a_n3420_39616.t6 25.8467
R32695 a_n3420_39616.n0 a_n3420_39616.t5 25.8467
R32696 a_n3420_39616.n8 a_n3420_39616.n6 22.6489
R32697 a_n3420_39616.n6 a_n3420_39616.n5 9.3005
R32698 a_n1925_46634.n0 a_n1925_46634.t4 276.464
R32699 a_n1925_46634.n1 a_n1925_46634.t2 209.291
R32700 a_n1925_46634.n2 a_n1925_46634.n0 205.827
R32701 a_n1925_46634.n0 a_n1925_46634.t5 196.131
R32702 a_n1925_46634.n3 a_n1925_46634.n2 194.331
R32703 a_n1925_46634.n1 a_n1925_46634.t3 174.583
R32704 a_n1925_46634.n2 a_n1925_46634.n1 50.3011
R32705 a_n1925_46634.t0 a_n1925_46634.n3 39.4005
R32706 a_n1925_46634.n3 a_n1925_46634.t1 37.4305
R32707 a_n3674_39304.n3 a_n3674_39304.n2 296.139
R32708 a_n3674_39304.n2 a_n3674_39304.n0 269.182
R32709 a_n3674_39304.n1 a_n3674_39304.t5 235.821
R32710 a_n3674_39304.n2 a_n3674_39304.n1 231.439
R32711 a_n3674_39304.n1 a_n3674_39304.t4 163.52
R32712 a_n3674_39304.n3 a_n3674_39304.t0 26.5955
R32713 a_n3674_39304.t1 a_n3674_39304.n3 26.5955
R32714 a_n3674_39304.n0 a_n3674_39304.t3 24.9236
R32715 a_n3674_39304.n0 a_n3674_39304.t2 24.9236
R32716 a_n4315_30879.n4 a_n4315_30879.t12 756.547
R32717 a_n4315_30879.n18 a_n4315_30879.t8 756.226
R32718 a_n4315_30879.n17 a_n4315_30879.t20 756.226
R32719 a_n4315_30879.n16 a_n4315_30879.t22 756.226
R32720 a_n4315_30879.n15 a_n4315_30879.t16 756.226
R32721 a_n4315_30879.n14 a_n4315_30879.t10 756.226
R32722 a_n4315_30879.n13 a_n4315_30879.t17 756.226
R32723 a_n4315_30879.n12 a_n4315_30879.t23 756.226
R32724 a_n4315_30879.n11 a_n4315_30879.t15 756.226
R32725 a_n4315_30879.n10 a_n4315_30879.t21 756.226
R32726 a_n4315_30879.n9 a_n4315_30879.t25 756.226
R32727 a_n4315_30879.n8 a_n4315_30879.t11 756.226
R32728 a_n4315_30879.n7 a_n4315_30879.t24 756.226
R32729 a_n4315_30879.n6 a_n4315_30879.t9 756.226
R32730 a_n4315_30879.n5 a_n4315_30879.t14 756.226
R32731 a_n4315_30879.n4 a_n4315_30879.t13 756.226
R32732 a_n4315_30879.n23 a_n4315_30879.n22 340.637
R32733 a_n4315_30879.n3 a_n4315_30879.t19 241.536
R32734 a_n4315_30879.n22 a_n4315_30879.n21 195.577
R32735 a_n4315_30879.n19 a_n4315_30879.n3 174.202
R32736 a_n4315_30879.n3 a_n4315_30879.t18 169.237
R32737 a_n4315_30879.n2 a_n4315_30879.n0 137.189
R32738 a_n4315_30879.n2 a_n4315_30879.n1 98.787
R32739 a_n4315_30879.n19 a_n4315_30879.n18 66.0013
R32740 a_n4315_30879.n20 a_n4315_30879.n2 38.9679
R32741 a_n4315_30879.n21 a_n4315_30879.t2 26.5955
R32742 a_n4315_30879.n21 a_n4315_30879.t1 26.5955
R32743 a_n4315_30879.t3 a_n4315_30879.n23 26.5955
R32744 a_n4315_30879.n23 a_n4315_30879.t0 26.5955
R32745 a_n4315_30879.n22 a_n4315_30879.n20 26.0391
R32746 a_n4315_30879.n0 a_n4315_30879.t6 24.9236
R32747 a_n4315_30879.n0 a_n4315_30879.t4 24.9236
R32748 a_n4315_30879.n1 a_n4315_30879.t7 24.9236
R32749 a_n4315_30879.n1 a_n4315_30879.t5 24.9236
R32750 a_n4315_30879.n20 a_n4315_30879.n19 9.30997
R32751 a_n4315_30879.n5 a_n4315_30879.n4 0.3205
R32752 a_n4315_30879.n6 a_n4315_30879.n5 0.3205
R32753 a_n4315_30879.n7 a_n4315_30879.n6 0.3205
R32754 a_n4315_30879.n8 a_n4315_30879.n7 0.3205
R32755 a_n4315_30879.n9 a_n4315_30879.n8 0.3205
R32756 a_n4315_30879.n10 a_n4315_30879.n9 0.3205
R32757 a_n4315_30879.n11 a_n4315_30879.n10 0.3205
R32758 a_n4315_30879.n12 a_n4315_30879.n11 0.3205
R32759 a_n4315_30879.n13 a_n4315_30879.n12 0.3205
R32760 a_n4315_30879.n14 a_n4315_30879.n13 0.3205
R32761 a_n4315_30879.n15 a_n4315_30879.n14 0.3205
R32762 a_n4315_30879.n16 a_n4315_30879.n15 0.3205
R32763 a_n4315_30879.n17 a_n4315_30879.n16 0.3205
R32764 a_n4315_30879.n18 a_n4315_30879.n17 0.303833
R32765 a_n3420_37984.n4 a_n3420_37984.t9 639.304
R32766 a_n3420_37984.n7 a_n3420_37984.n6 360.399
R32767 a_n3420_37984.n3 a_n3420_37984.t10 241.536
R32768 a_n3420_37984.n2 a_n3420_37984.n1 232.862
R32769 a_n3420_37984.n8 a_n3420_37984.n7 203.161
R32770 a_n3420_37984.n3 a_n3420_37984.t8 169.237
R32771 a_n3420_37984.n4 a_n3420_37984.n3 167.149
R32772 a_n3420_37984.n2 a_n3420_37984.n0 95.6721
R32773 a_n3420_37984.n5 a_n3420_37984.n2 60.5918
R32774 a_n3420_37984.n6 a_n3420_37984.t2 27.5805
R32775 a_n3420_37984.n6 a_n3420_37984.t0 27.5805
R32776 a_n3420_37984.n8 a_n3420_37984.t1 27.5805
R32777 a_n3420_37984.t3 a_n3420_37984.n8 27.5805
R32778 a_n3420_37984.n1 a_n3420_37984.t7 25.8467
R32779 a_n3420_37984.n1 a_n3420_37984.t4 25.8467
R32780 a_n3420_37984.n0 a_n3420_37984.t6 25.8467
R32781 a_n3420_37984.n0 a_n3420_37984.t5 25.8467
R32782 a_n3420_37984.n7 a_n3420_37984.n5 22.6489
R32783 a_n3420_37984.n5 a_n3420_37984.n4 9.3012
R32784 a_13507_46334.t0 a_13507_46334.n11 340.885
R32785 a_13507_46334.n0 a_13507_46334.t4 323.55
R32786 a_13507_46334.n3 a_13507_46334.t13 293.969
R32787 a_13507_46334.n5 a_13507_46334.t2 276.464
R32788 a_13507_46334.n1 a_13507_46334.t1 233.881
R32789 a_13507_46334.n2 a_13507_46334.t3 231.835
R32790 a_13507_46334.n8 a_13507_46334.t5 224.984
R32791 a_13507_46334.n7 a_13507_46334.t6 224.984
R32792 a_13507_46334.n4 a_13507_46334.n3 218.953
R32793 a_13507_46334.n5 a_13507_46334.t12 196.131
R32794 a_13507_46334.n0 a_13507_46334.t7 195.017
R32795 a_13507_46334.n8 a_13507_46334.t10 187.714
R32796 a_13507_46334.n7 a_13507_46334.t9 187.714
R32797 a_13507_46334.n9 a_13507_46334.n7 182.264
R32798 a_13507_46334.n9 a_13507_46334.n8 181.147
R32799 a_13507_46334.n6 a_13507_46334.n5 168.401
R32800 a_13507_46334.n4 a_13507_46334.n2 163.881
R32801 a_13507_46334.n1 a_13507_46334.n0 159.168
R32802 a_13507_46334.n2 a_13507_46334.t11 157.07
R32803 a_13507_46334.n3 a_13507_46334.t8 138.338
R32804 a_13507_46334.n6 a_13507_46334.n4 23.0348
R32805 a_13507_46334.n11 a_13507_46334.n10 20.8566
R32806 a_13507_46334.n11 a_13507_46334.n1 8.88939
R32807 a_13507_46334.n10 a_13507_46334.n9 4.46393
R32808 a_13507_46334.n10 a_13507_46334.n6 4.0544
R32809 a_5934_30871.n0 a_5934_30871.t4 645.846
R32810 a_5934_30871.n0 a_5934_30871.t6 641.817
R32811 a_5934_30871.n5 a_5934_30871.n4 380.32
R32812 a_5934_30871.n1 a_5934_30871.t7 260.322
R32813 a_5934_30871.n4 a_5934_30871.n3 185
R32814 a_5934_30871.n2 a_5934_30871.n1 177.923
R32815 a_5934_30871.n1 a_5934_30871.t5 175.169
R32816 a_5934_30871.n2 a_5934_30871.n0 125.263
R32817 a_5934_30871.n5 a_5934_30871.t0 26.5955
R32818 a_5934_30871.t1 a_5934_30871.n5 26.5955
R32819 a_5934_30871.n3 a_5934_30871.t3 24.9236
R32820 a_5934_30871.n3 a_5934_30871.t2 24.9236
R32821 a_5934_30871.n4 a_5934_30871.n2 16.3764
R32822 a_n2956_39304.n3 a_n2956_39304.n2 380.32
R32823 a_n2956_39304.n2 a_n2956_39304.n0 252.547
R32824 a_n2956_39304.n0 a_n2956_39304.t5 228.649
R32825 a_n2956_39304.n2 a_n2956_39304.n1 185
R32826 a_n2956_39304.n0 a_n2956_39304.t4 156.35
R32827 a_n2956_39304.t1 a_n2956_39304.n3 26.5955
R32828 a_n2956_39304.n3 a_n2956_39304.t0 26.5955
R32829 a_n2956_39304.n1 a_n2956_39304.t3 24.9236
R32830 a_n2956_39304.n1 a_n2956_39304.t2 24.9236
R32831 a_n4318_39304.n3 a_n4318_39304.n2 287.752
R32832 a_n4318_39304.n2 a_n4318_39304.n0 277.568
R32833 a_n4318_39304.n1 a_n4318_39304.t5 235.821
R32834 a_n4318_39304.n2 a_n4318_39304.n1 235.444
R32835 a_n4318_39304.n1 a_n4318_39304.t4 163.52
R32836 a_n4318_39304.t1 a_n4318_39304.n3 26.5955
R32837 a_n4318_39304.n3 a_n4318_39304.t0 26.5955
R32838 a_n4318_39304.n0 a_n4318_39304.t3 24.9236
R32839 a_n4318_39304.n0 a_n4318_39304.t2 24.9236
R32840 a_19692_46634.n3 a_19692_46634.n2 433.394
R32841 a_19692_46634.n1 a_19692_46634.t4 329.902
R32842 a_19692_46634.n2 a_19692_46634.t7 272.062
R32843 a_19692_46634.n0 a_19692_46634.t11 231.017
R32844 a_19692_46634.n9 a_19692_46634.t2 223.441
R32845 a_19692_46634.n5 a_19692_46634.t8 212.081
R32846 a_19692_46634.n6 a_19692_46634.t6 212.081
R32847 a_19692_46634.n8 a_19692_46634.n7 211.43
R32848 a_19692_46634.n2 a_19692_46634.t12 206.19
R32849 a_19692_46634.n4 a_19692_46634.n0 180.732
R32850 a_19692_46634.n3 a_19692_46634.n1 178.274
R32851 a_19692_46634.n10 a_19692_46634.n9 175.648
R32852 a_19692_46634.n0 a_19692_46634.t10 158.716
R32853 a_19692_46634.n1 a_19692_46634.t3 148.35
R32854 a_19692_46634.n5 a_19692_46634.t9 139.78
R32855 a_19692_46634.n6 a_19692_46634.t5 139.78
R32856 a_19692_46634.n7 a_19692_46634.n5 31.4035
R32857 a_19692_46634.n7 a_19692_46634.n6 31.4035
R32858 a_19692_46634.t0 a_19692_46634.n10 24.9236
R32859 a_19692_46634.n10 a_19692_46634.t1 24.9236
R32860 a_19692_46634.n8 a_19692_46634.n4 18.2368
R32861 a_19692_46634.n9 a_19692_46634.n8 17.2467
R32862 a_19692_46634.n4 a_19692_46634.n3 9.3005
R32863 a_15227_44166.n19 a_15227_44166.t13 471.289
R32864 a_15227_44166.n23 a_15227_44166.n22 380.32
R32865 a_15227_44166.n6 a_15227_44166.t9 327.99
R32866 a_15227_44166.n1 a_15227_44166.t11 267.065
R32867 a_15227_44166.n10 a_15227_44166.t25 256.728
R32868 a_15227_44166.n3 a_15227_44166.t15 256.716
R32869 a_15227_44166.n5 a_15227_44166.t12 241.536
R32870 a_15227_44166.n2 a_15227_44166.t7 241.536
R32871 a_15227_44166.n0 a_15227_44166.t14 236.18
R32872 a_15227_44166.n7 a_15227_44166.t16 212.081
R32873 a_15227_44166.n8 a_15227_44166.t5 212.081
R32874 a_15227_44166.n6 a_15227_44166.t17 199.457
R32875 a_15227_44166.n15 a_15227_44166.t18 196.549
R32876 a_15227_44166.n4 a_15227_44166.n2 192.591
R32877 a_15227_44166.n12 a_15227_44166.n6 189.279
R32878 a_15227_44166.n11 a_15227_44166.n10 185.749
R32879 a_15227_44166.n22 a_15227_44166.n21 185
R32880 a_15227_44166.n13 a_15227_44166.n5 179.663
R32881 a_15227_44166.n4 a_15227_44166.n3 179.017
R32882 a_15227_44166.n11 a_15227_44166.n9 174.653
R32883 a_15227_44166.n18 a_15227_44166.n0 173.488
R32884 a_15227_44166.n5 a_15227_44166.t4 169.237
R32885 a_15227_44166.n2 a_15227_44166.t10 169.237
R32886 a_15227_44166.n17 a_15227_44166.n1 167.506
R32887 a_15227_44166.n16 a_15227_44166.n15 167.506
R32888 a_15227_44166.n0 a_15227_44166.t22 163.881
R32889 a_15227_44166.n20 a_15227_44166.n19 162.514
R32890 a_15227_44166.n10 a_15227_44166.t20 161.275
R32891 a_15227_44166.n3 a_15227_44166.t21 161.275
R32892 a_15227_44166.n19 a_15227_44166.t6 148.35
R32893 a_15227_44166.n1 a_15227_44166.t23 148.35
R32894 a_15227_44166.n15 a_15227_44166.t19 148.35
R32895 a_15227_44166.n7 a_15227_44166.t8 139.78
R32896 a_15227_44166.n8 a_15227_44166.t24 139.78
R32897 a_15227_44166.n9 a_15227_44166.n8 37.246
R32898 a_15227_44166.n23 a_15227_44166.t0 26.5955
R32899 a_15227_44166.t1 a_15227_44166.n23 26.5955
R32900 a_15227_44166.n21 a_15227_44166.t2 24.9236
R32901 a_15227_44166.n21 a_15227_44166.t3 24.9236
R32902 a_15227_44166.n22 a_15227_44166.n20 24.7881
R32903 a_15227_44166.n9 a_15227_44166.n7 24.1005
R32904 a_15227_44166.n20 a_15227_44166.n18 20.9466
R32905 a_15227_44166.n18 a_15227_44166.n17 18.5527
R32906 a_15227_44166.n14 a_15227_44166.n13 8.95242
R32907 a_15227_44166.n16 a_15227_44166.n14 8.41275
R32908 a_15227_44166.n12 a_15227_44166.n11 6.7972
R32909 a_15227_44166.n14 a_15227_44166.n4 5.58292
R32910 a_15227_44166.n13 a_15227_44166.n12 2.39885
R32911 a_15227_44166.n17 a_15227_44166.n16 1.93748
R32912 a_19479_31679.n1 a_19479_31679.t4 595
R32913 a_19479_31679.n2 a_19479_31679.n1 380.32
R32914 a_19479_31679.n1 a_19479_31679.n0 185
R32915 a_19479_31679.n2 a_19479_31679.t0 26.5955
R32916 a_19479_31679.t1 a_19479_31679.n2 26.5955
R32917 a_19479_31679.n0 a_19479_31679.t2 24.9236
R32918 a_19479_31679.n0 a_19479_31679.t3 24.9236
R32919 a_1273_38525.t9 a_1273_38525.n5 542.547
R32920 a_1273_38525.n8 a_1273_38525.t9 542.081
R32921 a_1273_38525.n11 a_1273_38525.n0 344.094
R32922 a_1273_38525.n12 a_1273_38525.n11 313.916
R32923 a_1273_38525.n7 a_1273_38525.t12 270.545
R32924 a_1273_38525.n3 a_1273_38525.n1 230.554
R32925 a_1273_38525.n3 a_1273_38525.n2 200.375
R32926 a_1273_38525.n4 a_1273_38525.t11 199.597
R32927 a_1273_38525.n6 a_1273_38525.t13 199.572
R32928 a_1273_38525.n4 a_1273_38525.t8 197.951
R32929 a_1273_38525.n6 a_1273_38525.t10 197.947
R32930 a_1273_38525.n0 a_1273_38525.t2 26.5955
R32931 a_1273_38525.n0 a_1273_38525.t0 26.5955
R32932 a_1273_38525.t3 a_1273_38525.n12 26.5955
R32933 a_1273_38525.n12 a_1273_38525.t1 26.5955
R32934 a_1273_38525.n1 a_1273_38525.t7 24.9236
R32935 a_1273_38525.n1 a_1273_38525.t5 24.9236
R32936 a_1273_38525.n2 a_1273_38525.t4 24.9236
R32937 a_1273_38525.n2 a_1273_38525.t6 24.9236
R32938 a_1273_38525.n10 a_1273_38525.n9 21.1224
R32939 a_1273_38525.n11 a_1273_38525.n10 9.56818
R32940 a_1273_38525.n10 a_1273_38525.n3 8.79242
R32941 a_1273_38525.n8 a_1273_38525.n7 4.16605
R32942 a_1273_38525.n7 a_1273_38525.n6 2.52511
R32943 a_1273_38525.n9 a_1273_38525.n5 1.76521
R32944 a_1273_38525.n5 a_1273_38525.n4 1.27548
R32945 a_1273_38525.n9 a_1273_38525.n8 0.473054
R32946 a_13717_47436.t0 a_13717_47436.n1 461.301
R32947 a_13717_47436.n1 a_13717_47436.n0 270.363
R32948 a_13717_47436.n0 a_13717_47436.t2 241.536
R32949 a_13717_47436.n1 a_13717_47436.t1 216.155
R32950 a_13717_47436.n0 a_13717_47436.t3 169.237
R32951 a_3754_38470.n3 a_3754_38470.t9 542.561
R32952 a_3754_38470.n1 a_3754_38470.t8 542.561
R32953 a_3754_38470.n0 a_3754_38470.t10 542.561
R32954 a_3754_38470.n6 a_3754_38470.t7 542.545
R32955 a_3754_38470.n3 a_3754_38470.t4 542.081
R32956 a_3754_38470.n5 a_3754_38470.t5 542.081
R32957 a_3754_38470.n1 a_3754_38470.t3 542.081
R32958 a_3754_38470.n0 a_3754_38470.t6 542.081
R32959 a_3754_38470.n8 a_3754_38470.t1 100.382
R32960 a_3754_38470.t0 a_3754_38470.n8 44.988
R32961 a_3754_38470.n7 a_3754_38470.t2 44.0791
R32962 a_3754_38470.n8 a_3754_38470.n7 18.1307
R32963 a_3754_38470.n7 a_3754_38470.n6 2.16717
R32964 a_3754_38470.n4 a_3754_38470.n2 1.438
R32965 a_3754_38470.n4 a_3754_38470.n3 0.703
R32966 a_3754_38470.n2 a_3754_38470.n0 0.588
R32967 a_3754_38470.n2 a_3754_38470.n1 0.463
R32968 a_3754_38470.n5 a_3754_38470.n4 0.348
R32969 a_3754_38470.n6 a_3754_38470.n5 0.0155
R32970 VIN_P.n2 VIN_P.t12 92.1604
R32971 VIN_P.n4 VIN_P.t2 91.0227
R32972 VIN_P.n8 VIN_P.t1 90.7102
R32973 VIN_P.n7 VIN_P.t8 90.7102
R32974 VIN_P.n6 VIN_P.t6 90.7102
R32975 VIN_P.n5 VIN_P.t15 90.7102
R32976 VIN_P.n2 VIN_P.t11 90.6265
R32977 VIN_P.n3 VIN_P.t7 90.6219
R32978 VIN_P.n11 VIN_P.t13 47.4586
R32979 VIN_P.n10 VIN_P.n9 37.5586
R32980 VIN_P.n14 VIN_P.n13 29.098
R32981 VIN_P.n0 VIN_P.t9 25.3459
R32982 VIN_P.n0 VIN_P.t10 25.1217
R32983 VIN_P.n14 VIN_P.n0 20.9238
R32984 VIN_P VIN_P.n14 20.705
R32985 VIN_P.n13 VIN_P.t4 16.5266
R32986 VIN_P.n12 VIN_P.n1 14.0516
R32987 VIN_P.n12 VIN_P.n11 11.2899
R32988 VIN_P.n9 VIN_P.t3 9.9005
R32989 VIN_P.n9 VIN_P.t14 9.9005
R32990 VIN_P.n1 VIN_P.t0 2.4755
R32991 VIN_P.n1 VIN_P.t5 2.4755
R32992 VIN_P.n3 VIN_P.n2 1.6255
R32993 VIN_P.n4 VIN_P.n3 1.2505
R32994 VIN_P.n10 VIN_P.n8 0.8755
R32995 VIN_P.n6 VIN_P.n5 0.563
R32996 VIN_P.n7 VIN_P.n6 0.563
R32997 VIN_P.n8 VIN_P.n7 0.563
R32998 VIN_P.n11 VIN_P.n10 0.453625
R32999 VIN_P.n13 VIN_P.n12 0.438
R33000 VIN_P.n5 VIN_P.n4 0.2505
R33001 a_2711_45572.n6 a_2711_45572.t8 276.464
R33002 a_2711_45572.n1 a_2711_45572.t4 276.464
R33003 a_2711_45572.n4 a_2711_45572.t11 241.536
R33004 a_2711_45572.n2 a_2711_45572.t7 241.536
R33005 a_2711_45572.n9 a_2711_45572.n8 241.043
R33006 a_2711_45572.n6 a_2711_45572.t5 196.131
R33007 a_2711_45572.n1 a_2711_45572.t10 196.131
R33008 a_2711_45572.n3 a_2711_45572.n1 193.419
R33009 a_2711_45572.n5 a_2711_45572.n4 191.45
R33010 a_2711_45572.n4 a_2711_45572.t9 169.237
R33011 a_2711_45572.n2 a_2711_45572.t6 169.237
R33012 a_2711_45572.n7 a_2711_45572.n6 162.685
R33013 a_2711_45572.n3 a_2711_45572.n2 162.56
R33014 a_2711_45572.n8 a_2711_45572.n0 100.132
R33015 a_2711_45572.n9 a_2711_45572.t0 26.5955
R33016 a_2711_45572.t1 a_2711_45572.n9 26.5955
R33017 a_2711_45572.n0 a_2711_45572.t2 24.9236
R33018 a_2711_45572.n0 a_2711_45572.t3 24.9236
R33019 a_2711_45572.n7 a_2711_45572.n5 16.1995
R33020 a_2711_45572.n8 a_2711_45572.n7 15.5863
R33021 a_2711_45572.n5 a_2711_45572.n3 14.6088
R33022 a_n1057_35014.n17 a_n1057_35014.n16 21.0497
R33023 a_n1057_35014.n16 a_n1057_35014.n15 20.1816
R33024 a_n1057_35014.t4 a_n1057_35014.n1 9.23464
R33025 a_n1057_35014.n12 a_n1057_35014.t4 9.23464
R33026 a_n1057_35014.t6 a_n1057_35014.n5 9.23464
R33027 a_n1057_35014.n6 a_n1057_35014.t6 9.23464
R33028 a_n1057_35014.n5 a_n1057_35014.t5 9.23464
R33029 a_n1057_35014.t5 a_n1057_35014.n3 9.23464
R33030 a_n1057_35014.n12 a_n1057_35014.t7 9.23464
R33031 a_n1057_35014.t7 a_n1057_35014.n0 9.23464
R33032 a_n1057_35014.n16 a_n1057_35014.n14 8.608
R33033 a_n1057_35014.n13 a_n1057_35014.n1 7.21068
R33034 a_n1057_35014.n7 a_n1057_35014.n6 6.97092
R33035 a_n1057_35014.n14 a_n1057_35014.n0 6.82709
R33036 a_n1057_35014.n10 a_n1057_35014.n1 5.37709
R33037 a_n1057_35014.n15 a_n1057_35014.t2 4.9505
R33038 a_n1057_35014.n15 a_n1057_35014.t3 4.9505
R33039 a_n1057_35014.n17 a_n1057_35014.t0 4.9505
R33040 a_n1057_35014.t1 a_n1057_35014.n17 4.9505
R33041 a_n1057_35014.n6 a_n1057_35014.n4 4.2698
R33042 a_n1057_35014.n4 a_n1057_35014.n3 4.2697
R33043 a_n1057_35014.n8 a_n1057_35014.n3 3.69104
R33044 a_n1057_35014.n13 a_n1057_35014.n12 3.36698
R33045 a_n1057_35014.n8 a_n1057_35014.n7 3.27414
R33046 a_n1057_35014.n10 a_n1057_35014.n9 3.26815
R33047 a_n1057_35014.n9 a_n1057_35014.n8 3.08441
R33048 a_n1057_35014.n5 a_n1057_35014.n4 2.53338
R33049 a_n1057_35014.n7 a_n1057_35014.n2 2.24497
R33050 a_n1057_35014.n11 a_n1057_35014.n10 2.23901
R33051 a_n1057_35014.n9 a_n1057_35014.n0 2.15966
R33052 a_n1057_35014.n5 a_n1057_35014.n2 1.07382
R33053 a_n1057_35014.n11 a_n1057_35014.n2 0.911512
R33054 a_n1057_35014.n12 a_n1057_35014.n11 0.623492
R33055 a_n1057_35014.n14 a_n1057_35014.n13 0.34925
R33056 a_8696_44636.t0 a_8696_44636.n7 427.791
R33057 a_8696_44636.n1 a_8696_44636.t5 267.065
R33058 a_8696_44636.n6 a_8696_44636.n0 232.155
R33059 a_8696_44636.n0 a_8696_44636.t4 212.081
R33060 a_8696_44636.n7 a_8696_44636.t1 209.923
R33061 a_8696_44636.n2 a_8696_44636.t9 185.376
R33062 a_8696_44636.n4 a_8696_44636.t2 185.168
R33063 a_8696_44636.n3 a_8696_44636.n2 182.799
R33064 a_8696_44636.n3 a_8696_44636.n1 172.006
R33065 a_8696_44636.n5 a_8696_44636.n4 167.286
R33066 a_8696_44636.n1 a_8696_44636.t6 148.35
R33067 a_8696_44636.n0 a_8696_44636.t3 139.78
R33068 a_8696_44636.n2 a_8696_44636.t7 137.177
R33069 a_8696_44636.n4 a_8696_44636.t8 136.969
R33070 a_8696_44636.n7 a_8696_44636.n6 19.824
R33071 a_8696_44636.n5 a_8696_44636.n3 1.84871
R33072 a_8696_44636.n6 a_8696_44636.n5 1.28189
R33073 a_n443_42852.t12 a_n443_42852.t14 378.255
R33074 a_n443_42852.n6 a_n443_42852.t21 334.723
R33075 a_n443_42852.n4 a_n443_42852.t12 331.243
R33076 a_n443_42852.n21 a_n443_42852.n20 248.087
R33077 a_n443_42852.n16 a_n443_42852.t15 241.536
R33078 a_n443_42852.n8 a_n443_42852.t19 231.835
R33079 a_n443_42852.n7 a_n443_42852.n5 229.064
R33080 a_n443_42852.n10 a_n443_42852.t10 212.081
R33081 a_n443_42852.n11 a_n443_42852.t25 212.081
R33082 a_n443_42852.n20 a_n443_42852.n19 208.508
R33083 a_n443_42852.n6 a_n443_42852.t11 206.19
R33084 a_n443_42852.n5 a_n443_42852.t22 196.549
R33085 a_n443_42852.n12 a_n443_42852.n11 194.022
R33086 a_n443_42852.n7 a_n443_42852.n6 193.534
R33087 a_n443_42852.n4 a_n443_42852.n3 188.665
R33088 a_n443_42852.n9 a_n443_42852.n8 174.601
R33089 a_n443_42852.n17 a_n443_42852.n16 172.821
R33090 a_n443_42852.n16 a_n443_42852.t23 169.237
R33091 a_n443_42852.n15 a_n443_42852.n14 162.837
R33092 a_n443_42852.n8 a_n443_42852.t24 157.07
R33093 a_n443_42852.n5 a_n443_42852.t20 148.35
R33094 a_n443_42852.n3 a_n443_42852.t17 142.994
R33095 a_n443_42852.n10 a_n443_42852.t9 139.78
R33096 a_n443_42852.n11 a_n443_42852.t8 139.78
R33097 a_n443_42852.n2 a_n443_42852.n0 137.575
R33098 a_n443_42852.n14 a_n443_42852.t18 137.177
R33099 a_n443_42852.n3 a_n443_42852.t13 126.927
R33100 a_n443_42852.n14 a_n443_42852.t16 121.109
R33101 a_n443_42852.n2 a_n443_42852.n1 99.1749
R33102 a_n443_42852.n11 a_n443_42852.n10 61.346
R33103 a_n443_42852.n18 a_n443_42852.n2 36.0958
R33104 a_n443_42852.n19 a_n443_42852.t2 26.5955
R33105 a_n443_42852.n19 a_n443_42852.t0 26.5955
R33106 a_n443_42852.t3 a_n443_42852.n21 26.5955
R33107 a_n443_42852.n21 a_n443_42852.t1 26.5955
R33108 a_n443_42852.n0 a_n443_42852.t4 24.9236
R33109 a_n443_42852.n0 a_n443_42852.t6 24.9236
R33110 a_n443_42852.n1 a_n443_42852.t7 24.9236
R33111 a_n443_42852.n1 a_n443_42852.t5 24.9236
R33112 a_n443_42852.n13 a_n443_42852.n4 18.1682
R33113 a_n443_42852.n20 a_n443_42852.n18 17.2539
R33114 a_n443_42852.n12 a_n443_42852.n9 13.5127
R33115 a_n443_42852.n18 a_n443_42852.n17 12.2632
R33116 a_n443_42852.n15 a_n443_42852.n13 6.72933
R33117 a_n443_42852.n13 a_n443_42852.n12 5.55076
R33118 a_n443_42852.n9 a_n443_42852.n7 5.45754
R33119 a_n443_42852.n17 a_n443_42852.n15 0.309894
R33120 a_n1741_47186.n7 a_n1741_47186.n6 386.012
R33121 a_n1741_47186.n6 a_n1741_47186.n5 314.791
R33122 a_n1741_47186.n4 a_n1741_47186.n3 307.005
R33123 a_n1741_47186.n1 a_n1741_47186.t9 276.464
R33124 a_n1741_47186.n2 a_n1741_47186.n1 204.091
R33125 a_n1741_47186.n1 a_n1741_47186.t8 196.131
R33126 a_n1741_47186.n2 a_n1741_47186.n0 188.492
R33127 a_n1741_47186.n6 a_n1741_47186.n4 45.177
R33128 a_n1741_47186.n4 a_n1741_47186.n2 30.0611
R33129 a_n1741_47186.n3 a_n1741_47186.t3 27.5805
R33130 a_n1741_47186.n3 a_n1741_47186.t2 27.5805
R33131 a_n1741_47186.n5 a_n1741_47186.t7 27.5805
R33132 a_n1741_47186.n5 a_n1741_47186.t6 27.5805
R33133 a_n1741_47186.t1 a_n1741_47186.n7 27.5805
R33134 a_n1741_47186.n7 a_n1741_47186.t0 27.5805
R33135 a_n1741_47186.n0 a_n1741_47186.t4 25.8467
R33136 a_n1741_47186.n0 a_n1741_47186.t5 25.8467
R33137 COMP_P.n9 COMP_P.n8 321.861
R33138 COMP_P.n2 COMP_P.n1 244.067
R33139 COMP_P.n5 COMP_P.n3 236.589
R33140 COMP_P.n8 COMP_P.t11 230.155
R33141 COMP_P.n7 COMP_P.t10 224.984
R33142 COMP_P.n2 COMP_P.n0 204.893
R33143 COMP_P.n9 COMP_P.n7 203.353
R33144 COMP_P.n5 COMP_P.n4 200.321
R33145 COMP_P.n7 COMP_P.t9 187.714
R33146 COMP_P.n8 COMP_P.t8 157.856
R33147 COMP_P.n6 COMP_P.n2 30.0599
R33148 COMP_P.n6 COMP_P.n5 27.5565
R33149 COMP_P.n0 COMP_P.t1 26.5955
R33150 COMP_P.n0 COMP_P.t0 26.5955
R33151 COMP_P.n1 COMP_P.t3 26.5955
R33152 COMP_P.n1 COMP_P.t2 26.5955
R33153 COMP_P.n3 COMP_P.t4 24.9236
R33154 COMP_P.n3 COMP_P.t7 24.9236
R33155 COMP_P.n4 COMP_P.t6 24.9236
R33156 COMP_P.n4 COMP_P.t5 24.9236
R33157 COMP_P COMP_P.n6 14.4099
R33158 COMP_P COMP_P.n9 0.96925
R33159 DATA[2].n3 DATA[2].n2 647.148
R33160 DATA[2].n5 DATA[2].n4 200.262
R33161 DATA[2].n3 DATA[2].n1 194.441
R33162 DATA[2].n6 DATA[2].n0 185
R33163 DATA[2].n6 DATA[2].n5 58.6278
R33164 DATA[2].n5 DATA[2].n3 50.5705
R33165 DATA[2].n0 DATA[2].t7 40.0005
R33166 DATA[2].n0 DATA[2].t4 40.0005
R33167 DATA[2].n4 DATA[2].t6 40.0005
R33168 DATA[2].n4 DATA[2].t5 40.0005
R33169 DATA[2].n1 DATA[2].t3 27.5805
R33170 DATA[2].n1 DATA[2].t1 27.5805
R33171 DATA[2].n2 DATA[2].t0 27.5805
R33172 DATA[2].n2 DATA[2].t2 27.5805
R33173 DATA[2] DATA[2].n6 15.0895
R33174 SMPL_ON_P.n0 SMPL_ON_P.t8 260.322
R33175 SMPL_ON_P.n6 SMPL_ON_P.n4 244.069
R33176 SMPL_ON_P.n3 SMPL_ON_P.n1 236.589
R33177 SMPL_ON_P.n6 SMPL_ON_P.n5 204.893
R33178 SMPL_ON_P.n3 SMPL_ON_P.n2 200.321
R33179 SMPL_ON_P SMPL_ON_P.n0 192.925
R33180 SMPL_ON_P.n0 SMPL_ON_P.t9 175.169
R33181 SMPL_ON_P SMPL_ON_P.n7 96.1034
R33182 SMPL_ON_P.n7 SMPL_ON_P.n6 27.3804
R33183 SMPL_ON_P.n4 SMPL_ON_P.t0 26.5955
R33184 SMPL_ON_P.n4 SMPL_ON_P.t2 26.5955
R33185 SMPL_ON_P.n5 SMPL_ON_P.t3 26.5955
R33186 SMPL_ON_P.n5 SMPL_ON_P.t1 26.5955
R33187 SMPL_ON_P.n1 SMPL_ON_P.t5 24.9236
R33188 SMPL_ON_P.n1 SMPL_ON_P.t7 24.9236
R33189 SMPL_ON_P.n2 SMPL_ON_P.t4 24.9236
R33190 SMPL_ON_P.n2 SMPL_ON_P.t6 24.9236
R33191 SMPL_ON_P.n7 SMPL_ON_P.n3 24.8775
R33192 a_5742_30871.n1 a_5742_30871.t6 444.502
R33193 a_5742_30871.n0 a_5742_30871.t8 444.502
R33194 a_5742_30871.n7 a_5742_30871.n6 380.32
R33195 a_5742_30871.n1 a_5742_30871.t4 356.68
R33196 a_5742_30871.n0 a_5742_30871.t5 356.68
R33197 a_5742_30871.n3 a_5742_30871.t9 260.322
R33198 a_5742_30871.n2 a_5742_30871.n0 201.839
R33199 a_5742_30871.n2 a_5742_30871.n1 197.06
R33200 a_5742_30871.n6 a_5742_30871.n5 185
R33201 a_5742_30871.n3 a_5742_30871.t7 175.169
R33202 a_5742_30871.n4 a_5742_30871.n3 173.249
R33203 a_5742_30871.n4 a_5742_30871.n2 133.296
R33204 a_5742_30871.n7 a_5742_30871.t0 26.5955
R33205 a_5742_30871.t1 a_5742_30871.n7 26.5955
R33206 a_5742_30871.n5 a_5742_30871.t3 24.9236
R33207 a_5742_30871.n5 a_5742_30871.t2 24.9236
R33208 a_5742_30871.n6 a_5742_30871.n4 16.921
R33209 a_n2661_44458.n1 a_n2661_44458.t1 308.543
R33210 a_n2661_44458.n2 a_n2661_44458.n1 300.805
R33211 a_n2661_44458.n0 a_n2661_44458.t3 276.464
R33212 a_n2661_44458.n1 a_n2661_44458.n0 199.28
R33213 a_n2661_44458.n0 a_n2661_44458.t4 196.131
R33214 a_n2661_44458.n4 a_n2661_44458.n3 118.201
R33215 a_n2661_44458.n2 a_n2661_44458.t2 46.4362
R33216 a_n2661_44458.n3 a_n2661_44458.t0 28.7596
R33217 a_n2661_44458.n3 a_n2661_44458.n2 28.1434
R33218 w_10694_33990.n64 w_10694_33990.n7 15667.1
R33219 w_10694_33990.n61 w_10694_33990.n7 15667.1
R33220 w_10694_33990.n61 w_10694_33990.n9 15667.1
R33221 w_10694_33990.n33 w_10694_33990.n9 12324.7
R33222 w_10694_33990.n42 w_10694_33990.n22 3017.65
R33223 w_10694_33990.n44 w_10694_33990.n22 3017.65
R33224 w_10694_33990.n44 w_10694_33990.n23 3017.65
R33225 w_10694_33990.n34 w_10694_33990.n24 1757.65
R33226 w_10694_33990.n33 w_10694_33990.n6 1757.65
R33227 w_10694_33990.n60 w_10694_33990.n59 1671.15
R33228 w_10694_33990.n58 w_10694_33990.n10 1494.32
R33229 w_10694_33990.n64 w_10694_33990.n6 1464.71
R33230 w_10694_33990.n42 w_10694_33990.n24 1080
R33231 w_10694_33990.n65 w_10694_33990.n5 965.874
R33232 w_10694_33990.n37 w_10694_33990.t0 905.04
R33233 w_10694_33990.t2 w_10694_33990.n61 849.226
R33234 w_10694_33990.n63 w_10694_33990.t7 842.11
R33235 w_10694_33990.t0 w_10694_33990.n36 812.54
R33236 w_10694_33990.t7 w_10694_33990.n62 788.865
R33237 w_10694_33990.n62 w_10694_33990.t2 788.865
R33238 w_10694_33990.n15 w_10694_33990.n10 692.707
R33239 w_10694_33990.n59 w_10694_33990.n5 673.366
R33240 w_10694_33990.n15 w_10694_33990.n3 621.929
R33241 w_10694_33990.n37 w_10694_33990.n24 557.648
R33242 w_10694_33990.n37 w_10694_33990.n33 557.648
R33243 w_10694_33990.n35 w_10694_33990.n34 557.648
R33244 w_10694_33990.n35 w_10694_33990.n6 557.648
R33245 w_10694_33990.n45 w_10694_33990.n21 298.877
R33246 w_10694_33990.n32 w_10694_33990.n25 280.202
R33247 w_10694_33990.n46 w_10694_33990.n20 277.776
R33248 w_10694_33990.t1 w_10694_33990.n69 228.215
R33249 w_10694_33990.n66 w_10694_33990.n3 187.482
R33250 w_10694_33990.n40 w_10694_33990.n39 187.482
R33251 w_10694_33990.n60 w_10694_33990.n58 169.53
R33252 w_10694_33990.n66 w_10694_33990.n65 156.236
R33253 w_10694_33990.t12 w_10694_33990.n22 137.529
R33254 w_10694_33990.n41 w_10694_33990.n40 115.201
R33255 w_10694_33990.n36 w_10694_33990.n8 103.859
R33256 w_10694_33990.n38 w_10694_33990.n37 92.5005
R33257 w_10694_33990.n35 w_10694_33990.n4 92.5005
R33258 w_10694_33990.n36 w_10694_33990.n35 92.5005
R33259 w_10694_33990.t16 w_10694_33990.n8 75.2024
R33260 w_10694_33990.t10 w_10694_33990.t12 73.6677
R33261 w_10694_33990.t14 w_10694_33990.t16 73.6677
R33262 w_10694_33990.n14 w_10694_33990.t6 67.9353
R33263 w_10694_33990.t8 w_10694_33990.n11 67.9353
R33264 w_10694_33990.n54 w_10694_33990.t4 67.9353
R33265 w_10694_33990.t9 w_10694_33990.n51 67.9353
R33266 w_10694_33990.n27 w_10694_33990.t13 65.4041
R33267 w_10694_33990.n18 w_10694_33990.t17 62.5643
R33268 w_10694_33990.n34 w_10694_33990.n23 60.0005
R33269 w_10694_33990.n13 w_10694_33990.n12 59.5338
R33270 w_10694_33990.n53 w_10694_33990.n52 59.5338
R33271 w_10694_33990.n40 w_10694_33990.n38 59.4829
R33272 w_10694_33990.n38 w_10694_33990.n3 59.4829
R33273 w_10694_33990.n39 w_10694_33990.n4 59.4829
R33274 w_10694_33990.n66 w_10694_33990.n4 59.4829
R33275 w_10694_33990.n27 w_10694_33990.n26 56.8163
R33276 w_10694_33990.n43 w_10694_33990.t10 36.8341
R33277 w_10694_33990.n43 w_10694_33990.t14 36.8341
R33278 w_10694_33990.n63 w_10694_33990.n8 35.2823
R33279 w_10694_33990.n45 w_10694_33990.n44 26.4291
R33280 w_10694_33990.n44 w_10694_33990.n43 26.4291
R33281 w_10694_33990.n42 w_10694_33990.n41 26.4291
R33282 w_10694_33990.n43 w_10694_33990.n42 26.4291
R33283 w_10694_33990.n25 w_10694_33990.n20 20.4805
R33284 w_10694_33990.n41 w_10694_33990.n32 16.9417
R33285 w_10694_33990.n68 w_10694_33990.n1 15.2505
R33286 w_10694_33990.n22 w_10694_33990.n20 13.2148
R33287 w_10694_33990.n23 w_10694_33990.n21 13.2148
R33288 w_10694_33990.n23 w_10694_33990.n8 13.2148
R33289 w_10694_33990.n12 w_10694_33990.t8 8.40197
R33290 w_10694_33990.n12 w_10694_33990.t5 8.40197
R33291 w_10694_33990.n52 w_10694_33990.t9 8.40197
R33292 w_10694_33990.n52 w_10694_33990.t3 8.40197
R33293 w_10694_33990.n46 w_10694_33990.n45 8.2968
R33294 w_10694_33990.n26 w_10694_33990.t11 8.12675
R33295 w_10694_33990.n26 w_10694_33990.t15 8.12675
R33296 w_10694_33990.n56 w_10694_33990.n16 7.19895
R33297 w_10694_33990.n61 w_10694_33990.n60 7.11588
R33298 w_10694_33990.n65 w_10694_33990.n64 7.11588
R33299 w_10694_33990.n64 w_10694_33990.n63 7.11588
R33300 w_10694_33990.n55 w_10694_33990.n17 7.06493
R33301 w_10694_33990.n39 w_10694_33990.n21 6.4005
R33302 w_10694_33990.n28 w_10694_33990.n27 2.72081
R33303 w_10694_33990.n50 w_10694_33990.n17 2.33711
R33304 w_10694_33990.n29 w_10694_33990.n16 2.12421
R33305 w_10694_33990.n59 w_10694_33990.n7 1.8505
R33306 w_10694_33990.n62 w_10694_33990.n7 1.8505
R33307 w_10694_33990.n10 w_10694_33990.n9 1.8505
R33308 w_10694_33990.n62 w_10694_33990.n9 1.8505
R33309 w_10694_33990.n47 w_10694_33990.n46 1.5505
R33310 w_10694_33990.n32 w_10694_33990.n31 1.5505
R33311 w_10694_33990.n47 w_10694_33990.n19 1.26012
R33312 w_10694_33990.n25 w_10694_33990.n19 1.03383
R33313 w_10694_33990.n67 w_10694_33990.n66 1.03383
R33314 w_10694_33990.n58 w_10694_33990.n57 1.03383
R33315 w_10694_33990.n48 w_10694_33990.n18 1.00774
R33316 w_10694_33990.n53 w_10694_33990.n51 0.984766
R33317 w_10694_33990.n54 w_10694_33990.n53 0.984766
R33318 w_10694_33990.n13 w_10694_33990.n11 0.984766
R33319 w_10694_33990.n14 w_10694_33990.n13 0.984766
R33320 w_10694_33990.n31 w_10694_33990.n19 0.937356
R33321 w_10694_33990.n56 w_10694_33990.n55 0.741479
R33322 w_10694_33990.n48 w_10694_33990.n47 0.543562
R33323 w_10694_33990.n30 w_10694_33990.n29 0.494823
R33324 w_10694_33990.n31 w_10694_33990.n30 0.44251
R33325 w_10694_33990.n30 w_10694_33990.n28 0.428803
R33326 w_10694_33990.n49 w_10694_33990.n1 0.286876
R33327 w_10694_33990.n50 w_10694_33990.n49 0.260002
R33328 w_10694_33990.n29 w_10694_33990.n0 0.253077
R33329 w_10694_33990.n17 w_10694_33990.n5 0.227329
R33330 w_10694_33990.n16 w_10694_33990.n15 0.227329
R33331 w_10694_33990.n49 w_10694_33990.n48 0.192353
R33332 w_10694_33990.n2 w_10694_33990.n1 0.178335
R33333 w_10694_33990.n69 w_10694_33990.n68 0.0711522
R33334 w_10694_33990.n2 w_10694_33990.n0 0.0700876
R33335 w_10694_33990.n28 w_10694_33990.n18 0.057539
R33336 w_10694_33990.n55 w_10694_33990.n54 0.0348823
R33337 w_10694_33990.n57 w_10694_33990.n14 0.0334254
R33338 w_10694_33990.n51 w_10694_33990.n50 0.0330539
R33339 w_10694_33990.n11 w_10694_33990.n2 0.0325513
R33340 w_10694_33990.n69 w_10694_33990.n0 0.0303913
R33341 w_10694_33990.n68 w_10694_33990.n67 0.0136119
R33342 w_10694_33990.n57 w_10694_33990.n56 0.00195688
R33343 w_10694_33990.n67 w_10694_33990.n2 0.0016655
R33344 a_17364_32525.n1 a_17364_32525.t4 1687.01
R33345 a_17364_32525.n2 a_17364_32525.n1 287.752
R33346 a_17364_32525.n1 a_17364_32525.n0 277.568
R33347 a_17364_32525.t1 a_17364_32525.n2 26.5955
R33348 a_17364_32525.n2 a_17364_32525.t0 26.5955
R33349 a_17364_32525.n0 a_17364_32525.t2 24.9236
R33350 a_17364_32525.n0 a_17364_32525.t3 24.9236
R33351 VDAC_N.n0 VDAC_N.t20 946.489
R33352 VDAC_N.n10 VDAC_N.t23 946.489
R33353 VDAC_N.n3 VDAC_N.t9 946.489
R33354 VDAC_N.n2 VDAC_N.t15 945.755
R33355 VDAC_N.n1 VDAC_N.t12 945.755
R33356 VDAC_N.n0 VDAC_N.t16 945.755
R33357 VDAC_N.n12 VDAC_N.t22 945.755
R33358 VDAC_N.n11 VDAC_N.t17 945.755
R33359 VDAC_N.n10 VDAC_N.t21 945.755
R33360 VDAC_N.n9 VDAC_N.t19 945.755
R33361 VDAC_N.n8 VDAC_N.t13 945.755
R33362 VDAC_N.n7 VDAC_N.t11 945.755
R33363 VDAC_N.n6 VDAC_N.t10 945.755
R33364 VDAC_N.n5 VDAC_N.t8 945.755
R33365 VDAC_N.n4 VDAC_N.t18 945.755
R33366 VDAC_N.n3 VDAC_N.t14 945.755
R33367 VDAC_N.n22 VDAC_N.n14 20.1582
R33368 VDAC_N.n17 VDAC_N.n15 14.894
R33369 VDAC_N.n20 VDAC_N.n18 14.894
R33370 VDAC_N.n20 VDAC_N.n19 14.394
R33371 VDAC_N.n17 VDAC_N.n16 14.394
R33372 VDAC_N.n22 VDAC_N.n21 12.9266
R33373 VDAC_N.n6 VDAC_N.n5 6.84978
R33374 VDAC_N.n14 VDAC_N.n13 3.02654
R33375 VDAC_N.n14 VDAC_N.n2 2.75535
R33376 VDAC_N.n19 VDAC_N.t4 2.4755
R33377 VDAC_N.n19 VDAC_N.t6 2.4755
R33378 VDAC_N.n16 VDAC_N.t2 2.4755
R33379 VDAC_N.n16 VDAC_N.t5 2.4755
R33380 VDAC_N.n15 VDAC_N.t0 2.4755
R33381 VDAC_N.n15 VDAC_N.t3 2.4755
R33382 VDAC_N.n18 VDAC_N.t1 2.4755
R33383 VDAC_N.n18 VDAC_N.t7 2.4755
R33384 VDAC_N VDAC_N.n22 1.81269
R33385 VDAC_N.n13 VDAC_N.n9 1.04597
R33386 VDAC_N.n13 VDAC_N.n12 0.929304
R33387 VDAC_N.n1 VDAC_N.n0 0.733109
R33388 VDAC_N.n2 VDAC_N.n1 0.733109
R33389 VDAC_N.n11 VDAC_N.n10 0.733109
R33390 VDAC_N.n12 VDAC_N.n11 0.733109
R33391 VDAC_N.n4 VDAC_N.n3 0.733109
R33392 VDAC_N.n5 VDAC_N.n4 0.733109
R33393 VDAC_N.n7 VDAC_N.n6 0.733109
R33394 VDAC_N.n8 VDAC_N.n7 0.733109
R33395 VDAC_N.n9 VDAC_N.n8 0.733109
R33396 VDAC_N.n21 VDAC_N.n17 0.21925
R33397 VDAC_N.n21 VDAC_N.n20 0.188
R33398 a_5700_37509.n16 a_5700_37509.t1 120.882
R33399 a_5700_37509.n15 a_5700_37509.t3 120.57
R33400 a_5700_37509.n17 a_5700_37509.n16 104.317
R33401 a_5700_37509.n9 a_5700_37509.n7 39.965
R33402 a_5700_37509.n2 a_5700_37509.n0 39.792
R33403 a_5700_37509.n13 a_5700_37509.n12 39.6681
R33404 a_5700_37509.n11 a_5700_37509.n10 39.6681
R33405 a_5700_37509.n9 a_5700_37509.n8 39.6681
R33406 a_5700_37509.n6 a_5700_37509.n5 39.4951
R33407 a_5700_37509.n4 a_5700_37509.n3 39.4951
R33408 a_5700_37509.n2 a_5700_37509.n1 39.4951
R33409 a_5700_37509.t0 a_5700_37509.n17 16.253
R33410 a_5700_37509.n17 a_5700_37509.t2 16.253
R33411 a_5700_37509.n14 a_5700_37509.n13 14.9015
R33412 a_5700_37509.n15 a_5700_37509.n14 14.0786
R33413 a_5700_37509.n12 a_5700_37509.t15 4.76133
R33414 a_5700_37509.n12 a_5700_37509.t11 4.76133
R33415 a_5700_37509.n10 a_5700_37509.t16 4.76133
R33416 a_5700_37509.n10 a_5700_37509.t17 4.76133
R33417 a_5700_37509.n8 a_5700_37509.t8 4.76133
R33418 a_5700_37509.n8 a_5700_37509.t4 4.76133
R33419 a_5700_37509.n7 a_5700_37509.t5 4.76133
R33420 a_5700_37509.n7 a_5700_37509.t19 4.76133
R33421 a_5700_37509.n5 a_5700_37509.t18 4.76133
R33422 a_5700_37509.n5 a_5700_37509.t10 4.76133
R33423 a_5700_37509.n3 a_5700_37509.t7 4.76133
R33424 a_5700_37509.n3 a_5700_37509.t14 4.76133
R33425 a_5700_37509.n1 a_5700_37509.t6 4.76133
R33426 a_5700_37509.n1 a_5700_37509.t13 4.76133
R33427 a_5700_37509.n0 a_5700_37509.t9 4.76133
R33428 a_5700_37509.n0 a_5700_37509.t12 4.76133
R33429 a_5700_37509.n14 a_5700_37509.n6 1.96925
R33430 a_5700_37509.n11 a_5700_37509.n9 0.313
R33431 a_5700_37509.n13 a_5700_37509.n11 0.313
R33432 a_5700_37509.n4 a_5700_37509.n2 0.313
R33433 a_5700_37509.n6 a_5700_37509.n4 0.313
R33434 a_5700_37509.n16 a_5700_37509.n15 0.297375
R33435 C1_N_btm.n2 C1_N_btm.t0 102.406
R33436 C1_N_btm.n1 C1_N_btm.t2 101.787
R33437 C1_N_btm.n0 C1_N_btm.t1 54.9098
R33438 C1_N_btm.n0 C1_N_btm.t3 47.3635
R33439 C1_N_btm C1_N_btm.n2 46.0109
R33440 C1_N_btm.n2 C1_N_btm.n1 8.33383
R33441 C1_N_btm.n1 C1_N_btm.n0 7.99529
R33442 a_n4318_38216.n3 a_n4318_38216.n2 287.752
R33443 a_n4318_38216.n2 a_n4318_38216.n0 277.568
R33444 a_n4318_38216.n2 a_n4318_38216.n1 237.011
R33445 a_n4318_38216.n1 a_n4318_38216.t4 235.821
R33446 a_n4318_38216.n1 a_n4318_38216.t5 163.52
R33447 a_n4318_38216.n3 a_n4318_38216.t0 26.5955
R33448 a_n4318_38216.t1 a_n4318_38216.n3 26.5955
R33449 a_n4318_38216.n0 a_n4318_38216.t2 24.9236
R33450 a_n4318_38216.n0 a_n4318_38216.t3 24.9236
R33451 a_n1435_47204.t0 a_n1435_47204.n1 457.955
R33452 a_n1435_47204.n1 a_n1435_47204.n0 303.106
R33453 a_n1435_47204.n0 a_n1435_47204.t3 241.536
R33454 a_n1435_47204.n1 a_n1435_47204.t1 216.155
R33455 a_n1435_47204.n0 a_n1435_47204.t2 169.237
R33456 C1_P_btm.n2 C1_P_btm.t0 102.406
R33457 C1_P_btm.n1 C1_P_btm.t2 101.787
R33458 C1_P_btm.n0 C1_P_btm.t3 54.9098
R33459 C1_P_btm.n0 C1_P_btm.t1 47.3635
R33460 C1_P_btm C1_P_btm.n2 46.0422
R33461 C1_P_btm.n2 C1_P_btm.n1 8.33383
R33462 C1_P_btm.n1 C1_P_btm.n0 7.99529
R33463 a_5932_42308.n1 a_5932_42308.t4 580.756
R33464 a_5932_42308.n1 a_5932_42308.t6 578.977
R33465 a_5932_42308.n5 a_5932_42308.n4 380.32
R33466 a_5932_42308.n0 a_5932_42308.t5 260.322
R33467 a_5932_42308.n4 a_5932_42308.n3 185
R33468 a_5932_42308.n2 a_5932_42308.n0 175.847
R33469 a_5932_42308.n0 a_5932_42308.t7 175.169
R33470 a_5932_42308.n2 a_5932_42308.n1 106.338
R33471 a_5932_42308.t1 a_5932_42308.n5 26.5955
R33472 a_5932_42308.n5 a_5932_42308.t0 26.5955
R33473 a_5932_42308.n3 a_5932_42308.t3 24.9236
R33474 a_5932_42308.n3 a_5932_42308.t2 24.9236
R33475 a_5932_42308.n4 a_5932_42308.n2 21.4679
R33476 C3_N_btm.n1 C3_N_btm.t2 101.516
R33477 C3_N_btm.n2 C3_N_btm.t0 100.142
R33478 C3_N_btm.n0 C3_N_btm.t1 54.9311
R33479 C3_N_btm.n0 C3_N_btm.t3 47.3635
R33480 C3_N_btm C3_N_btm.n2 46.1255
R33481 C3_N_btm.n2 C3_N_btm.n1 9.7505
R33482 C3_N_btm.n1 C3_N_btm.n0 7.43279
R33483 a_11453_44696.t0 a_11453_44696.n4 728.274
R33484 a_11453_44696.t0 a_11453_44696.n0 685.292
R33485 a_11453_44696.n0 a_11453_44696.t1 289.469
R33486 a_11453_44696.n1 a_11453_44696.t4 276.464
R33487 a_11453_44696.n2 a_11453_44696.t2 254.256
R33488 a_11453_44696.n3 a_11453_44696.n1 207.054
R33489 a_11453_44696.n1 a_11453_44696.t3 196.131
R33490 a_11453_44696.n3 a_11453_44696.n2 182.899
R33491 a_11453_44696.n2 a_11453_44696.t5 181.956
R33492 a_11453_44696.n4 a_11453_44696.n0 15.826
R33493 a_11453_44696.n4 a_11453_44696.n3 15.2583
R33494 DATA[1].n4 DATA[1].n3 647.148
R33495 DATA[1].n5 DATA[1].n1 243.627
R33496 DATA[1].n4 DATA[1].n2 194.441
R33497 DATA[1].n6 DATA[1].n0 185
R33498 DATA[1].n5 DATA[1].n4 50.5705
R33499 DATA[1].n0 DATA[1].t6 40.0005
R33500 DATA[1].n0 DATA[1].t4 40.0005
R33501 DATA[1].n1 DATA[1].t5 40.0005
R33502 DATA[1].n1 DATA[1].t7 40.0005
R33503 DATA[1].n2 DATA[1].t0 27.5805
R33504 DATA[1].n2 DATA[1].t2 27.5805
R33505 DATA[1].n3 DATA[1].t3 27.5805
R33506 DATA[1].n3 DATA[1].t1 27.5805
R33507 DATA[1].n6 DATA[1].n5 15.262
R33508 DATA[1] DATA[1].n6 15.0895
R33509 a_4361_42308.t0 a_4361_42308.n1 463.529
R33510 a_4361_42308.n0 a_4361_42308.t3 276.464
R33511 a_4361_42308.n1 a_4361_42308.t1 254.047
R33512 a_4361_42308.n1 a_4361_42308.n0 207.708
R33513 a_4361_42308.n0 a_4361_42308.t2 196.131
R33514 a_n4318_40392.n3 a_n4318_40392.n2 296.139
R33515 a_n4318_40392.n2 a_n4318_40392.n0 269.182
R33516 a_n4318_40392.n1 a_n4318_40392.t4 235.821
R33517 a_n4318_40392.n2 a_n4318_40392.n1 224.416
R33518 a_n4318_40392.n1 a_n4318_40392.t5 163.52
R33519 a_n4318_40392.t1 a_n4318_40392.n3 26.5955
R33520 a_n4318_40392.n3 a_n4318_40392.t0 26.5955
R33521 a_n4318_40392.n0 a_n4318_40392.t2 24.9236
R33522 a_n4318_40392.n0 a_n4318_40392.t3 24.9236
R33523 a_n2661_46634.n0 a_n2661_46634.t3 276.464
R33524 a_n2661_46634.n1 a_n2661_46634.n0 218.47
R33525 a_n2661_46634.n2 a_n2661_46634.n1 196.846
R33526 a_n2661_46634.n0 a_n2661_46634.t4 196.131
R33527 a_n2661_46634.n1 a_n2661_46634.t1 193.519
R33528 a_n2661_46634.n2 a_n2661_46634.t2 26.5955
R33529 a_n2661_46634.t0 a_n2661_46634.n2 26.5955
R33530 a_413_45260.t0 a_413_45260.n3 386.269
R33531 a_413_45260.n2 a_413_45260.n0 292.861
R33532 a_413_45260.n0 a_413_45260.t3 276.464
R33533 a_413_45260.n1 a_413_45260.t2 230.155
R33534 a_413_45260.n0 a_413_45260.t4 196.131
R33535 a_413_45260.n2 a_413_45260.n1 178.494
R33536 a_413_45260.n1 a_413_45260.t5 157.856
R33537 a_413_45260.n3 a_413_45260.t1 131.219
R33538 a_413_45260.n3 a_413_45260.n2 20.6467
R33539 VDAC_Pi VDAC_Pi.t9 388.01
R33540 VDAC_Pi.n3 VDAC_Pi.t10 234.685
R33541 VDAC_Pi.n2 VDAC_Pi.n0 104.316
R33542 VDAC_Pi.n2 VDAC_Pi.n1 104.019
R33543 VDAC_Pi.n3 VDAC_Pi.t8 50.2666
R33544 VDAC_Pi.n8 VDAC_Pi.n7 37.3277
R33545 VDAC_Pi.n6 VDAC_Pi.n5 37.3277
R33546 VDAC_Pi.n1 VDAC_Pi.t2 16.253
R33547 VDAC_Pi.n1 VDAC_Pi.t1 16.253
R33548 VDAC_Pi.n0 VDAC_Pi.t3 16.253
R33549 VDAC_Pi.n0 VDAC_Pi.t0 16.253
R33550 VDAC_Pi VDAC_Pi.n8 14.5151
R33551 VDAC_Pi.n7 VDAC_Pi.t6 9.9005
R33552 VDAC_Pi.n7 VDAC_Pi.t7 9.9005
R33553 VDAC_Pi.n5 VDAC_Pi.t4 9.9005
R33554 VDAC_Pi.n5 VDAC_Pi.t5 9.9005
R33555 VDAC_Pi.n4 VDAC_Pi.n3 6.15675
R33556 VDAC_Pi.n4 VDAC_Pi.n2 1.46925
R33557 VDAC_Pi.n6 VDAC_Pi.n4 0.359875
R33558 VDAC_Pi.n8 VDAC_Pi.n6 0.297375
R33559 a_7174_31319.n0 a_7174_31319.t4 569.808
R33560 a_7174_31319.n0 a_7174_31319.t5 567.279
R33561 a_7174_31319.n3 a_7174_31319.n2 380.32
R33562 a_7174_31319.n2 a_7174_31319.n0 196.883
R33563 a_7174_31319.n2 a_7174_31319.n1 185
R33564 a_7174_31319.n3 a_7174_31319.t0 26.5955
R33565 a_7174_31319.t1 a_7174_31319.n3 26.5955
R33566 a_7174_31319.n1 a_7174_31319.t3 24.9236
R33567 a_7174_31319.n1 a_7174_31319.t2 24.9236
R33568 a_20447_31679.n1 a_20447_31679.t4 601.816
R33569 a_20447_31679.n2 a_20447_31679.n1 287.752
R33570 a_20447_31679.n1 a_20447_31679.n0 277.568
R33571 a_20447_31679.n2 a_20447_31679.t0 26.5955
R33572 a_20447_31679.t1 a_20447_31679.n2 26.5955
R33573 a_20447_31679.n0 a_20447_31679.t3 24.9236
R33574 a_20447_31679.n0 a_20447_31679.t2 24.9236
R33575 a_n357_42282.n10 a_n357_42282.t15 722.096
R33576 a_n357_42282.n8 a_n357_42282.t11 722.096
R33577 a_n357_42282.n6 a_n357_42282.t13 722.096
R33578 a_n357_42282.n4 a_n357_42282.t17 722.096
R33579 a_n357_42282.n2 a_n357_42282.t14 722.096
R33580 a_n357_42282.n15 a_n357_42282.n14 380.32
R33581 a_n357_42282.n0 a_n357_42282.t8 276.464
R33582 a_n357_42282.n1 a_n357_42282.t9 241.536
R33583 a_n357_42282.n0 a_n357_42282.t7 196.131
R33584 a_n357_42282.n3 a_n357_42282.n1 194.608
R33585 a_n357_42282.n14 a_n357_42282.n13 185
R33586 a_n357_42282.n5 a_n357_42282.n4 182.524
R33587 a_n357_42282.n11 a_n357_42282.n10 176.232
R33588 a_n357_42282.n9 a_n357_42282.n8 176.232
R33589 a_n357_42282.n7 a_n357_42282.n6 176.232
R33590 a_n357_42282.n3 a_n357_42282.n2 173.22
R33591 a_n357_42282.n12 a_n357_42282.n0 169.312
R33592 a_n357_42282.n1 a_n357_42282.t4 169.237
R33593 a_n357_42282.n10 a_n357_42282.t6 162.963
R33594 a_n357_42282.n8 a_n357_42282.t12 162.963
R33595 a_n357_42282.n6 a_n357_42282.t5 162.963
R33596 a_n357_42282.n4 a_n357_42282.t16 162.963
R33597 a_n357_42282.n2 a_n357_42282.t10 162.963
R33598 a_n357_42282.n15 a_n357_42282.t0 26.5955
R33599 a_n357_42282.t1 a_n357_42282.n15 26.5955
R33600 a_n357_42282.n13 a_n357_42282.t3 24.9236
R33601 a_n357_42282.n13 a_n357_42282.t2 24.9236
R33602 a_n357_42282.n14 a_n357_42282.n12 17.6554
R33603 a_n357_42282.n11 a_n357_42282.n9 7.49073
R33604 a_n357_42282.n12 a_n357_42282.n11 6.36053
R33605 a_n357_42282.n7 a_n357_42282.n5 4.3198
R33606 a_n357_42282.n5 a_n357_42282.n3 4.2171
R33607 a_n357_42282.n9 a_n357_42282.n7 1.14887
R33608 a_n4318_37592.n3 a_n4318_37592.n2 296.139
R33609 a_n4318_37592.n2 a_n4318_37592.n0 269.182
R33610 a_n4318_37592.n2 a_n4318_37592.n1 244.493
R33611 a_n4318_37592.n1 a_n4318_37592.t4 235.821
R33612 a_n4318_37592.n1 a_n4318_37592.t5 163.52
R33613 a_n4318_37592.t1 a_n4318_37592.n3 26.5955
R33614 a_n4318_37592.n3 a_n4318_37592.t0 26.5955
R33615 a_n4318_37592.n0 a_n4318_37592.t3 24.9236
R33616 a_n4318_37592.n0 a_n4318_37592.t2 24.9236
R33617 a_19721_31679.n1 a_19721_31679.t4 593.259
R33618 a_19721_31679.n2 a_19721_31679.n1 380.32
R33619 a_19721_31679.n1 a_19721_31679.n0 185
R33620 a_19721_31679.t1 a_19721_31679.n2 26.5955
R33621 a_19721_31679.n2 a_19721_31679.t0 26.5955
R33622 a_19721_31679.n0 a_19721_31679.t2 24.9236
R33623 a_19721_31679.n0 a_19721_31679.t3 24.9236
R33624 C2_N_btm.n1 C2_N_btm.t3 101.621
R33625 C2_N_btm.n2 C2_N_btm.t1 98.936
R33626 C2_N_btm.n0 C2_N_btm.t2 54.9311
R33627 C2_N_btm C2_N_btm.n2 50.6047
R33628 C2_N_btm.n0 C2_N_btm.t0 47.3635
R33629 C2_N_btm.n1 C2_N_btm.n0 7.71404
R33630 C2_N_btm.n2 C2_N_btm.n1 7.20883
R33631 a_n4064_38528.n4 a_n4064_38528.t8 698.881
R33632 a_n4064_38528.n7 a_n4064_38528.n6 360.399
R33633 a_n4064_38528.n3 a_n4064_38528.t10 241.536
R33634 a_n4064_38528.n2 a_n4064_38528.n1 232.862
R33635 a_n4064_38528.n8 a_n4064_38528.n7 203.161
R33636 a_n4064_38528.n4 a_n4064_38528.n3 172.543
R33637 a_n4064_38528.n3 a_n4064_38528.t9 169.237
R33638 a_n4064_38528.n2 a_n4064_38528.n0 95.6721
R33639 a_n4064_38528.n5 a_n4064_38528.n2 61.9632
R33640 a_n4064_38528.n6 a_n4064_38528.t1 27.5805
R33641 a_n4064_38528.n6 a_n4064_38528.t2 27.5805
R33642 a_n4064_38528.t3 a_n4064_38528.n8 27.5805
R33643 a_n4064_38528.n8 a_n4064_38528.t0 27.5805
R33644 a_n4064_38528.n1 a_n4064_38528.t4 25.8467
R33645 a_n4064_38528.n1 a_n4064_38528.t5 25.8467
R33646 a_n4064_38528.n0 a_n4064_38528.t6 25.8467
R33647 a_n4064_38528.n0 a_n4064_38528.t7 25.8467
R33648 a_n4064_38528.n7 a_n4064_38528.n5 21.2775
R33649 a_n4064_38528.n5 a_n4064_38528.n4 9.3005
R33650 C5_P_btm.n1 C5_P_btm.t2 101.204
R33651 C5_P_btm.n2 C5_P_btm.t0 98.0923
R33652 C5_P_btm C5_P_btm.n2 55.9172
R33653 C5_P_btm.n0 C5_P_btm.t3 54.9311
R33654 C5_P_btm.n0 C5_P_btm.t1 47.3635
R33655 C5_P_btm.n2 C5_P_btm.n1 8.08383
R33656 C5_P_btm.n1 C5_P_btm.n0 6.87029
R33657 a_3357_43084.n2 a_3357_43084.n0 281.579
R33658 a_3357_43084.n0 a_3357_43084.t3 276.464
R33659 a_3357_43084.n4 a_3357_43084.n3 259.058
R33660 a_3357_43084.n1 a_3357_43084.t6 230.155
R33661 a_3357_43084.n0 a_3357_43084.t4 196.131
R33662 a_3357_43084.n2 a_3357_43084.n1 178.806
R33663 a_3357_43084.n1 a_3357_43084.t5 157.856
R33664 a_3357_43084.n3 a_3357_43084.t1 131.308
R33665 a_3357_43084.t0 a_3357_43084.n4 26.5955
R33666 a_3357_43084.n4 a_3357_43084.t2 26.5955
R33667 a_3357_43084.n3 a_3357_43084.n2 20.6941
R33668 a_1666_39587.n0 a_1666_39587.t6 440.495
R33669 a_1666_39587.n4 a_1666_39587.t2 239.103
R33670 a_1666_39587.n1 a_1666_39587.t4 230.576
R33671 a_1666_39587.n0 a_1666_39587.t5 191.952
R33672 a_1666_39587.n2 a_1666_39587.n1 174.456
R33673 a_1666_39587.n1 a_1666_39587.t3 158.275
R33674 a_1666_39587.n3 a_1666_39587.t1 85.1701
R33675 a_1666_39587.t0 a_1666_39587.n4 61.169
R33676 a_1666_39587.n2 a_1666_39587.n0 5.84425
R33677 a_1666_39587.n3 a_1666_39587.n2 4.5005
R33678 a_1666_39587.n4 a_1666_39587.n3 2.04495
R33679 DATA[0].n6 DATA[0].n5 585
R33680 DATA[0].n2 DATA[0].n0 243.627
R33681 DATA[0].n2 DATA[0].n1 200.262
R33682 DATA[0].n4 DATA[0].n3 194.441
R33683 DATA[0].n6 DATA[0].n4 62.148
R33684 DATA[0].n4 DATA[0].n2 50.5705
R33685 DATA[0].n0 DATA[0].t7 40.0005
R33686 DATA[0].n0 DATA[0].t5 40.0005
R33687 DATA[0].n1 DATA[0].t6 40.0005
R33688 DATA[0].n1 DATA[0].t4 40.0005
R33689 DATA[0].n5 DATA[0].t0 27.5805
R33690 DATA[0].n5 DATA[0].t1 27.5805
R33691 DATA[0].n3 DATA[0].t2 27.5805
R33692 DATA[0].n3 DATA[0].t3 27.5805
R33693 DATA[0] DATA[0].n6 23.6347
R33694 C3_P_btm.n1 C3_P_btm.t0 101.516
R33695 C3_P_btm.n2 C3_P_btm.t2 100.142
R33696 C3_P_btm.n0 C3_P_btm.t1 54.9311
R33697 C3_P_btm.n0 C3_P_btm.t3 47.3635
R33698 C3_P_btm C3_P_btm.n2 46.1567
R33699 C3_P_btm.n2 C3_P_btm.n1 9.7505
R33700 C3_P_btm.n1 C3_P_btm.n0 7.43279
R33701 a_2982_43646.n4 a_2982_43646.n3 677.66
R33702 a_2982_43646.n5 a_2982_43646.n4 291.856
R33703 a_2982_43646.n1 a_2982_43646.t7 276.464
R33704 a_2982_43646.n2 a_2982_43646.n1 217.475
R33705 a_2982_43646.n1 a_2982_43646.t6 196.131
R33706 a_2982_43646.n2 a_2982_43646.n0 190.487
R33707 a_2982_43646.n4 a_2982_43646.n2 54.5624
R33708 a_2982_43646.n3 a_2982_43646.t5 27.5805
R33709 a_2982_43646.n3 a_2982_43646.t4 27.5805
R33710 a_2982_43646.n5 a_2982_43646.t0 27.5805
R33711 a_2982_43646.t1 a_2982_43646.n5 27.5805
R33712 a_2982_43646.n0 a_2982_43646.t2 25.8467
R33713 a_2982_43646.n0 a_2982_43646.t3 25.8467
R33714 a_5649_42852.n1 a_5649_42852.t1 362.774
R33715 a_5649_42852.t0 a_5649_42852.n1 317.154
R33716 a_5649_42852.n1 a_5649_42852.n0 282.308
R33717 a_5649_42852.n0 a_5649_42852.t3 276.464
R33718 a_5649_42852.n0 a_5649_42852.t2 196.131
R33719 a_6945_45028.n0 a_6945_45028.t4 276.464
R33720 a_6945_45028.n2 a_6945_45028.n1 254.679
R33721 a_6945_45028.n1 a_6945_45028.n0 217.331
R33722 a_6945_45028.n0 a_6945_45028.t3 196.131
R33723 a_6945_45028.n1 a_6945_45028.t1 135.579
R33724 a_6945_45028.t0 a_6945_45028.n2 26.5955
R33725 a_6945_45028.n2 a_6945_45028.t2 26.5955
R33726 a_n4064_37440.n4 a_n4064_37440.t9 636.116
R33727 a_n4064_37440.n7 a_n4064_37440.n6 360.399
R33728 a_n4064_37440.n3 a_n4064_37440.t10 241.536
R33729 a_n4064_37440.n2 a_n4064_37440.n1 232.862
R33730 a_n4064_37440.n8 a_n4064_37440.n7 203.161
R33731 a_n4064_37440.n4 a_n4064_37440.n3 172.543
R33732 a_n4064_37440.n3 a_n4064_37440.t8 169.237
R33733 a_n4064_37440.n2 a_n4064_37440.n0 95.6721
R33734 a_n4064_37440.n5 a_n4064_37440.n2 61.9632
R33735 a_n4064_37440.n6 a_n4064_37440.t1 27.5805
R33736 a_n4064_37440.n6 a_n4064_37440.t0 27.5805
R33737 a_n4064_37440.t3 a_n4064_37440.n8 27.5805
R33738 a_n4064_37440.n8 a_n4064_37440.t2 27.5805
R33739 a_n4064_37440.n1 a_n4064_37440.t7 25.8467
R33740 a_n4064_37440.n1 a_n4064_37440.t6 25.8467
R33741 a_n4064_37440.n0 a_n4064_37440.t5 25.8467
R33742 a_n4064_37440.n0 a_n4064_37440.t4 25.8467
R33743 a_n4064_37440.n7 a_n4064_37440.n5 21.2775
R33744 a_n4064_37440.n5 a_n4064_37440.n4 9.3005
R33745 a_n2956_37592.n3 a_n2956_37592.n2 287.752
R33746 a_n2956_37592.n2 a_n2956_37592.n0 277.568
R33747 a_n2956_37592.n2 a_n2956_37592.n1 262.291
R33748 a_n2956_37592.n1 a_n2956_37592.t4 228.649
R33749 a_n2956_37592.n1 a_n2956_37592.t5 156.35
R33750 a_n2956_37592.n3 a_n2956_37592.t0 26.5955
R33751 a_n2956_37592.t1 a_n2956_37592.n3 26.5955
R33752 a_n2956_37592.n0 a_n2956_37592.t2 24.9236
R33753 a_n2956_37592.n0 a_n2956_37592.t3 24.9236
R33754 C7_N_btm C7_N_btm.n3 60.4693
R33755 C7_N_btm.n3 C7_N_btm.t0 53.6613
R33756 C7_N_btm.n1 C7_N_btm.n0 52.9499
R33757 C7_N_btm.n1 C7_N_btm.t4 23.6451
R33758 C7_N_btm.n2 C7_N_btm.t1 23.6328
R33759 C7_N_btm.n2 C7_N_btm.n1 11.2505
R33760 C7_N_btm.n3 C7_N_btm.n2 8.41717
R33761 C7_N_btm.n0 C7_N_btm.t2 3.57113
R33762 C7_N_btm.n0 C7_N_btm.t3 3.57113
R33763 DATA[4].n3 DATA[4].n2 647.148
R33764 DATA[4].n5 DATA[4].n4 200.262
R33765 DATA[4].n3 DATA[4].n1 194.441
R33766 DATA[4].n6 DATA[4].n0 185
R33767 DATA[4].n6 DATA[4].n5 58.6278
R33768 DATA[4].n5 DATA[4].n3 50.5705
R33769 DATA[4].n0 DATA[4].t6 40.0005
R33770 DATA[4].n0 DATA[4].t7 40.0005
R33771 DATA[4].n4 DATA[4].t5 40.0005
R33772 DATA[4].n4 DATA[4].t4 40.0005
R33773 DATA[4].n1 DATA[4].t1 27.5805
R33774 DATA[4].n1 DATA[4].t3 27.5805
R33775 DATA[4].n2 DATA[4].t2 27.5805
R33776 DATA[4].n2 DATA[4].t0 27.5805
R33777 DATA[4] DATA[4].n6 16.205
R33778 a_n2661_45546.n0 a_n2661_45546.t3 276.464
R33779 a_n2661_45546.n2 a_n2661_45546.n1 259.058
R33780 a_n2661_45546.n1 a_n2661_45546.n0 207.364
R33781 a_n2661_45546.n0 a_n2661_45546.t4 196.131
R33782 a_n2661_45546.n1 a_n2661_45546.t1 131.308
R33783 a_n2661_45546.n2 a_n2661_45546.t2 26.5955
R33784 a_n2661_45546.t0 a_n2661_45546.n2 26.5955
R33785 a_n3674_38216.n3 a_n3674_38216.n2 380.32
R33786 a_n3674_38216.n0 a_n3674_38216.t4 235.821
R33787 a_n3674_38216.n2 a_n3674_38216.n0 234.791
R33788 a_n3674_38216.n2 a_n3674_38216.n1 185
R33789 a_n3674_38216.n0 a_n3674_38216.t5 163.52
R33790 a_n3674_38216.n3 a_n3674_38216.t0 26.5955
R33791 a_n3674_38216.t1 a_n3674_38216.n3 26.5955
R33792 a_n3674_38216.n1 a_n3674_38216.t2 24.9236
R33793 a_n3674_38216.n1 a_n3674_38216.t3 24.9236
R33794 a_14401_32519.n1 a_14401_32519.t5 444.502
R33795 a_14401_32519.n1 a_14401_32519.t4 356.68
R33796 a_14401_32519.n2 a_14401_32519.n1 302.296
R33797 a_14401_32519.n3 a_14401_32519.n2 287.752
R33798 a_14401_32519.n2 a_14401_32519.n0 277.568
R33799 a_14401_32519.n3 a_14401_32519.t0 26.5955
R33800 a_14401_32519.t1 a_14401_32519.n3 26.5955
R33801 a_14401_32519.n0 a_14401_32519.t2 24.9236
R33802 a_14401_32519.n0 a_14401_32519.t3 24.9236
R33803 a_n3420_38528.n4 a_n3420_38528.t8 639.018
R33804 a_n3420_38528.n7 a_n3420_38528.n6 360.399
R33805 a_n3420_38528.n3 a_n3420_38528.t9 241.536
R33806 a_n3420_38528.n2 a_n3420_38528.n1 232.862
R33807 a_n3420_38528.n8 a_n3420_38528.n7 203.161
R33808 a_n3420_38528.n3 a_n3420_38528.t10 169.237
R33809 a_n3420_38528.n4 a_n3420_38528.n3 166.983
R33810 a_n3420_38528.n2 a_n3420_38528.n0 95.6721
R33811 a_n3420_38528.n5 a_n3420_38528.n2 60.5918
R33812 a_n3420_38528.n6 a_n3420_38528.t1 27.5805
R33813 a_n3420_38528.n6 a_n3420_38528.t2 27.5805
R33814 a_n3420_38528.n8 a_n3420_38528.t0 27.5805
R33815 a_n3420_38528.t3 a_n3420_38528.n8 27.5805
R33816 a_n3420_38528.n1 a_n3420_38528.t7 25.8467
R33817 a_n3420_38528.n1 a_n3420_38528.t4 25.8467
R33818 a_n3420_38528.n0 a_n3420_38528.t6 25.8467
R33819 a_n3420_38528.n0 a_n3420_38528.t5 25.8467
R33820 a_n3420_38528.n7 a_n3420_38528.n5 22.6489
R33821 a_n3420_38528.n5 a_n3420_38528.n4 9.3005
R33822 a_n2956_38216.n3 a_n2956_38216.n2 380.32
R33823 a_n2956_38216.n2 a_n2956_38216.n0 251.31
R33824 a_n2956_38216.n0 a_n2956_38216.t5 228.649
R33825 a_n2956_38216.n2 a_n2956_38216.n1 185
R33826 a_n2956_38216.n0 a_n2956_38216.t4 156.35
R33827 a_n2956_38216.n3 a_n2956_38216.t0 26.5955
R33828 a_n2956_38216.t1 a_n2956_38216.n3 26.5955
R33829 a_n2956_38216.n1 a_n2956_38216.t2 24.9236
R33830 a_n2956_38216.n1 a_n2956_38216.t3 24.9236
R33831 a_n2293_45546.n0 a_n2293_45546.t4 276.464
R33832 a_n2293_45546.n3 a_n2293_45546.n2 244.631
R33833 a_n2293_45546.n2 a_n2293_45546.t1 209.291
R33834 a_n2293_45546.n1 a_n2293_45546.n0 202.655
R33835 a_n2293_45546.n0 a_n2293_45546.t5 196.131
R33836 a_n2293_45546.n1 a_n2293_45546.t2 169.752
R33837 a_n2293_45546.t0 a_n2293_45546.n3 39.4005
R33838 a_n2293_45546.n3 a_n2293_45546.t3 37.4305
R33839 a_n2293_45546.n2 a_n2293_45546.n1 4.33281
R33840 a_14209_32519.n1 a_14209_32519.t4 736.798
R33841 a_14209_32519.n2 a_14209_32519.n1 380.32
R33842 a_14209_32519.n1 a_14209_32519.n0 185
R33843 a_14209_32519.t1 a_14209_32519.n2 26.5955
R33844 a_14209_32519.n2 a_14209_32519.t0 26.5955
R33845 a_14209_32519.n0 a_14209_32519.t3 24.9236
R33846 a_14209_32519.n0 a_14209_32519.t2 24.9236
R33847 CLK CLK.n3 242.577
R33848 CLK.n3 CLK.t1 184.768
R33849 CLK.n2 CLK.t7 184.768
R33850 CLK.n1 CLK.t5 184.768
R33851 CLK.n0 CLK.t2 184.768
R33852 CLK.n3 CLK.t0 146.208
R33853 CLK.n2 CLK.t6 146.208
R33854 CLK.n1 CLK.t3 146.208
R33855 CLK.n0 CLK.t4 146.208
R33856 CLK.n3 CLK.n2 40.6397
R33857 CLK.n2 CLK.n1 40.6397
R33858 CLK.n1 CLK.n0 40.6397
R33859 a_9313_44734.n2 a_9313_44734.n1 398.971
R33860 a_9313_44734.n0 a_9313_44734.t3 276.464
R33861 a_9313_44734.n1 a_9313_44734.n0 211.371
R33862 a_9313_44734.n1 a_9313_44734.t1 209.923
R33863 a_9313_44734.n0 a_9313_44734.t4 196.131
R33864 a_9313_44734.n2 a_9313_44734.t2 56.9025
R33865 a_9313_44734.t0 a_9313_44734.n2 46.4362
R33866 a_9145_43396.n0 a_9145_43396.t2 334.723
R33867 a_9145_43396.t0 a_9145_43396.n1 325.793
R33868 a_9145_43396.n1 a_9145_43396.t1 303.44
R33869 a_9145_43396.n1 a_9145_43396.n0 217.119
R33870 a_9145_43396.n0 a_9145_43396.t3 206.19
R33871 C4_P_btm.n1 C4_P_btm.t0 101.361
R33872 C4_P_btm.n2 C4_P_btm.t2 98.3735
R33873 C4_P_btm.n0 C4_P_btm.t3 54.9311
R33874 C4_P_btm C4_P_btm.n2 52.9172
R33875 C4_P_btm.n0 C4_P_btm.t1 47.3635
R33876 C4_P_btm.n2 C4_P_btm.n1 8.08383
R33877 C4_P_btm.n1 C4_P_btm.n0 7.15154
R33878 a_n3420_37440.n4 a_n3420_37440.t9 640.486
R33879 a_n3420_37440.n7 a_n3420_37440.n6 360.399
R33880 a_n3420_37440.n3 a_n3420_37440.t8 241.536
R33881 a_n3420_37440.n2 a_n3420_37440.n1 232.862
R33882 a_n3420_37440.n8 a_n3420_37440.n7 203.161
R33883 a_n3420_37440.n3 a_n3420_37440.t10 169.237
R33884 a_n3420_37440.n4 a_n3420_37440.n3 166.983
R33885 a_n3420_37440.n2 a_n3420_37440.n0 95.6721
R33886 a_n3420_37440.n5 a_n3420_37440.n2 60.5918
R33887 a_n3420_37440.n6 a_n3420_37440.t1 27.5805
R33888 a_n3420_37440.n6 a_n3420_37440.t2 27.5805
R33889 a_n3420_37440.n8 a_n3420_37440.t0 27.5805
R33890 a_n3420_37440.t3 a_n3420_37440.n8 27.5805
R33891 a_n3420_37440.n1 a_n3420_37440.t7 25.8467
R33892 a_n3420_37440.n1 a_n3420_37440.t4 25.8467
R33893 a_n3420_37440.n0 a_n3420_37440.t6 25.8467
R33894 a_n3420_37440.n0 a_n3420_37440.t5 25.8467
R33895 a_n3420_37440.n7 a_n3420_37440.n5 22.6489
R33896 a_n3420_37440.n5 a_n3420_37440.n4 9.3005
R33897 a_n2810_45572.n3 a_n2810_45572.n2 296.139
R33898 a_n2810_45572.n2 a_n2810_45572.n0 269.182
R33899 a_n2810_45572.n2 a_n2810_45572.n1 261.625
R33900 a_n2810_45572.n1 a_n2810_45572.t5 228.649
R33901 a_n2810_45572.n1 a_n2810_45572.t4 156.35
R33902 a_n2810_45572.t1 a_n2810_45572.n3 26.5955
R33903 a_n2810_45572.n3 a_n2810_45572.t0 26.5955
R33904 a_n2810_45572.n0 a_n2810_45572.t3 24.9236
R33905 a_n2810_45572.n0 a_n2810_45572.t2 24.9236
R33906 a_n2661_43922.n0 a_n2661_43922.t3 276.464
R33907 a_n2661_43922.n2 a_n2661_43922.n1 259.06
R33908 a_n2661_43922.n1 a_n2661_43922.n0 204.612
R33909 a_n2661_43922.n0 a_n2661_43922.t4 196.131
R33910 a_n2661_43922.n1 a_n2661_43922.t1 131.308
R33911 a_n2661_43922.n2 a_n2661_43922.t2 26.5955
R33912 a_n2661_43922.t0 a_n2661_43922.n2 26.5955
R33913 a_4338_37500.t0 a_4338_37500.n4 258.05
R33914 a_4338_37500.n4 a_4338_37500.n3 53.4434
R33915 a_4338_37500.n1 a_4338_37500.t5 47.8126
R33916 a_4338_37500.n2 a_4338_37500.t2 47.5157
R33917 a_4338_37500.n1 a_4338_37500.n0 37.6157
R33918 a_4338_37500.n3 a_4338_37500.t6 10.4216
R33919 a_4338_37500.n3 a_4338_37500.t1 10.4216
R33920 a_4338_37500.n0 a_4338_37500.t3 9.9005
R33921 a_4338_37500.n0 a_4338_37500.t4 9.9005
R33922 a_4338_37500.n4 a_4338_37500.n2 2.8755
R33923 a_4338_37500.n2 a_4338_37500.n1 0.313
R33924 RST_Z.n0 RST_Z.t3 751.299
R33925 RST_Z.n0 RST_Z.t5 403.308
R33926 RST_Z.n3 RST_Z.t1 260.322
R33927 RST_Z.n1 RST_Z.t0 230.576
R33928 RST_Z.n3 RST_Z.t2 175.169
R33929 RST_Z RST_Z.n3 171.161
R33930 RST_Z.n2 RST_Z.n1 167.165
R33931 RST_Z.n1 RST_Z.t4 158.275
R33932 RST_Z RST_Z.n2 147.383
R33933 RST_Z.n2 RST_Z.n0 36.9629
R33934 CAL_P.n5 CAL_P.n4 601.129
R33935 CAL_P.n5 CAL_P.t1 251.643
R33936 CAL_P CAL_P.t5 137
R33937 CAL_P.n4 CAL_P.t2 77.3934
R33938 CAL_P.n4 CAL_P.t0 77.3934
R33939 CAL_P.n1 CAL_P.t4 36.3712
R33940 CAL_P.t6 CAL_P.n0 36.2721
R33941 CAL_P.n2 CAL_P.t4 35.5162
R33942 CAL_P.n3 CAL_P.t6 35.4454
R33943 CAL_P.n2 CAL_P.t3 31.2287
R33944 CAL_P.t3 CAL_P.n1 31.2287
R33945 CAL_P CAL_P.n6 23.5275
R33946 CAL_P.n6 CAL_P.n5 8.34425
R33947 CAL_P.n6 CAL_P.n3 7.5005
R33948 CAL_P.n6 CAL_P.n0 5.95883
R33949 CAL_P.n1 CAL_P.n0 0.0713333
R33950 CAL_P.n3 CAL_P.n2 0.0713333
R33951 C5_N_btm.n1 C5_N_btm.t2 101.204
R33952 C5_N_btm.n2 C5_N_btm.t0 98.0923
R33953 C5_N_btm C5_N_btm.n2 55.9797
R33954 C5_N_btm.n0 C5_N_btm.t3 54.9311
R33955 C5_N_btm.n0 C5_N_btm.t1 47.3635
R33956 C5_N_btm.n2 C5_N_btm.n1 8.08383
R33957 C5_N_btm.n1 C5_N_btm.n0 6.87029
R33958 a_19963_31679.n1 a_19963_31679.t4 592.938
R33959 a_19963_31679.n2 a_19963_31679.n1 296.139
R33960 a_19963_31679.n1 a_19963_31679.n0 269.182
R33961 a_19963_31679.t1 a_19963_31679.n2 26.5955
R33962 a_19963_31679.n2 a_19963_31679.t0 26.5955
R33963 a_19963_31679.n0 a_19963_31679.t3 24.9236
R33964 a_19963_31679.n0 a_19963_31679.t2 24.9236
R33965 a_n2293_46634.n0 a_n2293_46634.t3 276.464
R33966 a_n2293_46634.n1 a_n2293_46634.n0 233.769
R33967 a_n2293_46634.n1 a_n2293_46634.t1 199.456
R33968 a_n2293_46634.n0 a_n2293_46634.t4 196.131
R33969 a_n2293_46634.n2 a_n2293_46634.n1 190.911
R33970 a_n2293_46634.n2 a_n2293_46634.t2 26.5955
R33971 a_n2293_46634.t0 a_n2293_46634.n2 26.5955
R33972 a_n2293_46098.n1 a_n2293_46098.t1 377.127
R33973 a_n2293_46098.t0 a_n2293_46098.n1 327.82
R33974 a_n2293_46098.n0 a_n2293_46098.t3 276.464
R33975 a_n2293_46098.n1 a_n2293_46098.n0 220.982
R33976 a_n2293_46098.n0 a_n2293_46098.t2 196.131
R33977 a_11341_43940.n2 a_11341_43940.n1 285.519
R33978 a_11341_43940.n0 a_11341_43940.t4 276.464
R33979 a_11341_43940.n1 a_11341_43940.n0 213.929
R33980 a_11341_43940.n1 a_11341_43940.t1 196.238
R33981 a_11341_43940.n0 a_11341_43940.t3 196.131
R33982 a_11341_43940.n2 a_11341_43940.t2 127.066
R33983 a_11341_43940.t0 a_11341_43940.n2 27.5805
R33984 a_13678_32519.n1 a_13678_32519.t4 678.686
R33985 a_13678_32519.n2 a_13678_32519.n1 380.32
R33986 a_13678_32519.n1 a_13678_32519.n0 185
R33987 a_13678_32519.t1 a_13678_32519.n2 26.5955
R33988 a_13678_32519.n2 a_13678_32519.t0 26.5955
R33989 a_13678_32519.n0 a_13678_32519.t3 24.9236
R33990 a_13678_32519.n0 a_13678_32519.t2 24.9236
R33991 C0_dummy_N_btm.n0 C0_dummy_N_btm.t0 104.561
R33992 C0_dummy_N_btm.n0 C0_dummy_N_btm.t1 62.8375
R33993 C0_dummy_N_btm C0_dummy_N_btm.n0 46.6776
R33994 a_8685_43396.n0 a_8685_43396.t3 330.12
R33995 a_8685_43396.t0 a_8685_43396.n1 279.577
R33996 a_8685_43396.n1 a_8685_43396.n0 225.47
R33997 a_8685_43396.n0 a_8685_43396.t2 201.587
R33998 a_8685_43396.n1 a_8685_43396.t1 130.916
R33999 a_n356_44636.n2 a_n356_44636.n0 459.668
R34000 a_n356_44636.n1 a_n356_44636.t5 329.902
R34001 a_n356_44636.t0 a_n356_44636.n3 295.594
R34002 a_n356_44636.n0 a_n356_44636.t2 272.062
R34003 a_n356_44636.n0 a_n356_44636.t4 206.19
R34004 a_n356_44636.n2 a_n356_44636.n1 152
R34005 a_n356_44636.n1 a_n356_44636.t3 148.35
R34006 a_n356_44636.n3 a_n356_44636.n2 147.788
R34007 a_n356_44636.n3 a_n356_44636.t1 129.046
R34008 a_n2312_38680.n3 a_n2312_38680.n2 380.32
R34009 a_n2312_38680.n2 a_n2312_38680.n0 267.74
R34010 a_n2312_38680.n0 a_n2312_38680.t5 228.649
R34011 a_n2312_38680.n2 a_n2312_38680.n1 185
R34012 a_n2312_38680.n0 a_n2312_38680.t4 156.35
R34013 a_n2312_38680.n3 a_n2312_38680.t0 26.5955
R34014 a_n2312_38680.t1 a_n2312_38680.n3 26.5955
R34015 a_n2312_38680.n1 a_n2312_38680.t2 24.9236
R34016 a_n2312_38680.n1 a_n2312_38680.t3 24.9236
R34017 a_n2109_47186.t0 a_n2109_47186.n1 463.529
R34018 a_n2109_47186.n0 a_n2109_47186.t3 276.464
R34019 a_n2109_47186.n1 a_n2109_47186.t1 254.047
R34020 a_n2109_47186.n1 a_n2109_47186.n0 225.118
R34021 a_n2109_47186.n0 a_n2109_47186.t2 196.131
R34022 C2_P_btm.n1 C2_P_btm.t3 101.621
R34023 C2_P_btm.n2 C2_P_btm.t1 98.936
R34024 C2_P_btm.n0 C2_P_btm.t2 54.9311
R34025 C2_P_btm C2_P_btm.n2 50.3859
R34026 C2_P_btm.n0 C2_P_btm.t0 47.3635
R34027 C2_P_btm.n1 C2_P_btm.n0 7.71404
R34028 C2_P_btm.n2 C2_P_btm.n1 7.20883
R34029 a_n4318_38680.n3 a_n4318_38680.n2 380.32
R34030 a_n4318_38680.n2 a_n4318_38680.n0 238.207
R34031 a_n4318_38680.n0 a_n4318_38680.t4 235.821
R34032 a_n4318_38680.n2 a_n4318_38680.n1 185
R34033 a_n4318_38680.n0 a_n4318_38680.t5 163.52
R34034 a_n4318_38680.n3 a_n4318_38680.t0 26.5955
R34035 a_n4318_38680.t1 a_n4318_38680.n3 26.5955
R34036 a_n4318_38680.n1 a_n4318_38680.t2 24.9236
R34037 a_n4318_38680.n1 a_n4318_38680.t3 24.9236
R34038 a_n2661_42282.t0 a_n2661_42282.n1 392.938
R34039 a_n2661_42282.n0 a_n2661_42282.t3 276.464
R34040 a_n2661_42282.n1 a_n2661_42282.t1 257.678
R34041 a_n2661_42282.n1 a_n2661_42282.n0 241.732
R34042 a_n2661_42282.n0 a_n2661_42282.t2 196.131
R34043 SINGLE_ENDED.n0 SINGLE_ENDED.t0 260.322
R34044 SINGLE_ENDED.n0 SINGLE_ENDED.t1 175.169
R34045 SINGLE_ENDED SINGLE_ENDED.n0 173.482
R34046 C0_dummy_P_btm.n0 C0_dummy_P_btm.t0 104.561
R34047 C0_dummy_P_btm.n0 C0_dummy_P_btm.t1 62.8375
R34048 C0_dummy_P_btm C0_dummy_P_btm.n0 46.6776
R34049 C8_P_btm C8_P_btm.n8 64.7297
R34050 C8_P_btm.n8 C8_P_btm.n7 43.4801
R34051 C8_P_btm.n2 C8_P_btm.n1 33.0333
R34052 C8_P_btm.n2 C8_P_btm.n0 32.3614
R34053 C8_P_btm.n4 C8_P_btm.n2 21.6828
R34054 C8_P_btm.n4 C8_P_btm.n3 20.8888
R34055 C8_P_btm.n6 C8_P_btm.n5 20.8766
R34056 C8_P_btm.n6 C8_P_btm.n4 11.2088
R34057 C8_P_btm.n7 C8_P_btm.t5 9.9005
R34058 C8_P_btm.n7 C8_P_btm.t4 9.9005
R34059 C8_P_btm.n8 C8_P_btm.n6 8.45883
R34060 C8_P_btm C8_P_btm.n250 5.72472
R34061 C8_P_btm.n0 C8_P_btm.t0 3.57113
R34062 C8_P_btm.n0 C8_P_btm.t1 3.57113
R34063 C8_P_btm.n1 C8_P_btm.t2 3.57113
R34064 C8_P_btm.n1 C8_P_btm.t3 3.57113
R34065 C8_P_btm.n3 C8_P_btm.t6 2.4755
R34066 C8_P_btm.n3 C8_P_btm.t7 2.4755
R34067 C8_P_btm.n5 C8_P_btm.t9 2.4755
R34068 C8_P_btm.n5 C8_P_btm.t8 2.4755
R34069 C8_P_btm.n160 C8_P_btm.n130 0.276161
R34070 C8_P_btm.n41 C8_P_btm.n40 0.276161
R34071 C8_P_btm.n53 C8_P_btm.n51 0.276161
R34072 C8_P_btm.n177 C8_P_btm.n176 0.276161
R34073 C8_P_btm.n155 C8_P_btm.n154 0.276161
R34074 C8_P_btm.n39 C8_P_btm.n34 0.228786
R34075 C8_P_btm.n38 C8_P_btm.n35 0.228786
R34076 C8_P_btm.n52 C8_P_btm.n11 0.228786
R34077 C8_P_btm.n55 C8_P_btm.n54 0.228786
R34078 C8_P_btm.n12 C8_P_btm.n11 0.228786
R34079 C8_P_btm.n14 C8_P_btm.n12 0.228786
R34080 C8_P_btm.n56 C8_P_btm.n55 0.228786
R34081 C8_P_btm.n57 C8_P_btm.n56 0.228786
R34082 C8_P_btm.n15 C8_P_btm.n14 0.228786
R34083 C8_P_btm.n59 C8_P_btm.n15 0.228786
R34084 C8_P_btm.n58 C8_P_btm.n57 0.228786
R34085 C8_P_btm.n61 C8_P_btm.n58 0.228786
R34086 C8_P_btm.n60 C8_P_btm.n59 0.228786
R34087 C8_P_btm.n60 C8_P_btm.n19 0.228786
R34088 C8_P_btm.n62 C8_P_btm.n61 0.228786
R34089 C8_P_btm.n63 C8_P_btm.n62 0.228786
R34090 C8_P_btm.n20 C8_P_btm.n19 0.228786
R34091 C8_P_btm.n22 C8_P_btm.n20 0.228786
R34092 C8_P_btm.n64 C8_P_btm.n63 0.228786
R34093 C8_P_btm.n64 C8_P_btm.n44 0.228786
R34094 C8_P_btm.n23 C8_P_btm.n22 0.228786
R34095 C8_P_btm.n37 C8_P_btm.n23 0.228786
R34096 C8_P_btm.n70 C8_P_btm.n37 0.228786
R34097 C8_P_btm.n69 C8_P_btm.n68 0.228786
R34098 C8_P_btm.n69 C8_P_btm.n36 0.228786
R34099 C8_P_btm.n27 C8_P_btm.n26 0.228786
R34100 C8_P_btm.n71 C8_P_btm.n70 0.228786
R34101 C8_P_btm.n72 C8_P_btm.n71 0.228786
R34102 C8_P_btm.n233 C8_P_btm.n28 0.228786
R34103 C8_P_btm.n73 C8_P_btm.n27 0.228786
R34104 C8_P_btm.n74 C8_P_btm.n73 0.228786
R34105 C8_P_btm.n75 C8_P_btm.n28 0.228786
R34106 C8_P_btm.n76 C8_P_btm.n75 0.228786
R34107 C8_P_btm.n77 C8_P_btm.n29 0.228786
R34108 C8_P_btm.n231 C8_P_btm.n29 0.228786
R34109 C8_P_btm.n229 C8_P_btm.n228 0.228786
R34110 C8_P_btm.n227 C8_P_btm.n32 0.228786
R34111 C8_P_btm.n226 C8_P_btm.n78 0.228786
R34112 C8_P_btm.n225 C8_P_btm.n224 0.228786
R34113 C8_P_btm.n223 C8_P_btm.n79 0.228786
R34114 C8_P_btm.n86 C8_P_btm.n81 0.228786
R34115 C8_P_btm.n213 C8_P_btm.n212 0.228786
R34116 C8_P_btm.n211 C8_P_btm.n85 0.228786
R34117 C8_P_btm.n210 C8_P_btm.n87 0.228786
R34118 C8_P_btm.n209 C8_P_btm.n208 0.228786
R34119 C8_P_btm.n207 C8_P_btm.n88 0.228786
R34120 C8_P_btm.n95 C8_P_btm.n90 0.228786
R34121 C8_P_btm.n198 C8_P_btm.n197 0.228786
R34122 C8_P_btm.n196 C8_P_btm.n94 0.228786
R34123 C8_P_btm.n195 C8_P_btm.n96 0.228786
R34124 C8_P_btm.n194 C8_P_btm.n193 0.228786
R34125 C8_P_btm.n192 C8_P_btm.n97 0.228786
R34126 C8_P_btm.n108 C8_P_btm.n99 0.228786
R34127 C8_P_btm.n114 C8_P_btm.n106 0.228786
R34128 C8_P_btm.n113 C8_P_btm.n112 0.228786
R34129 C8_P_btm.n111 C8_P_btm.n110 0.228786
R34130 C8_P_btm.n183 C8_P_btm.n104 0.228786
R34131 C8_P_btm.n119 C8_P_btm.n117 0.228786
R34132 C8_P_btm.n117 C8_P_btm.n105 0.228786
R34133 C8_P_btm.n182 C8_P_btm.n102 0.228786
R34134 C8_P_btm.n182 C8_P_btm.n181 0.228786
R34135 C8_P_btm.n180 C8_P_btm.n105 0.228786
R34136 C8_P_btm.n180 C8_P_btm.n179 0.228786
R34137 C8_P_btm.n179 C8_P_btm.n115 0.228786
R34138 C8_P_btm.n178 C8_P_btm.n107 0.228786
R34139 C8_P_btm.n176 C8_P_btm.n175 0.228786
R34140 C8_P_btm.n174 C8_P_btm.n173 0.228786
R34141 C8_P_btm.n118 C8_P_btm.n116 0.228786
R34142 C8_P_btm.n172 C8_P_btm.n171 0.228786
R34143 C8_P_btm.n170 C8_P_btm.n169 0.228786
R34144 C8_P_btm.n169 C8_P_btm.n168 0.228786
R34145 C8_P_btm.n141 C8_P_btm.n139 0.228786
R34146 C8_P_btm.n124 C8_P_btm.n123 0.228786
R34147 C8_P_btm.n126 C8_P_btm.n124 0.228786
R34148 C8_P_btm.n149 C8_P_btm.n138 0.228786
R34149 C8_P_btm.n151 C8_P_btm.n150 0.228786
R34150 C8_P_btm.n136 C8_P_btm.n127 0.228786
R34151 C8_P_btm.n136 C8_P_btm.n135 0.228786
R34152 C8_P_btm.n135 C8_P_btm.n131 0.228786
R34153 C8_P_btm.n152 C8_P_btm.n133 0.228786
R34154 C8_P_btm.n157 C8_P_btm.n156 0.228786
R34155 C8_P_btm.n159 C8_P_btm.n158 0.228786
R34156 C8_P_btm.n159 C8_P_btm.n129 0.228786
R34157 C8_P_btm.n161 C8_P_btm.n160 0.228786
R34158 C8_P_btm.n162 C8_P_btm.n161 0.228786
R34159 C8_P_btm.n129 C8_P_btm.n128 0.228786
R34160 C8_P_btm.n164 C8_P_btm.n128 0.228786
R34161 C8_P_btm.n163 C8_P_btm.n162 0.228786
R34162 C8_P_btm.n163 C8_P_btm.n125 0.228786
R34163 C8_P_btm.n165 C8_P_btm.n164 0.228786
R34164 C8_P_btm.n166 C8_P_btm.n165 0.228786
R34165 C8_P_btm.n125 C8_P_btm.n122 0.228786
R34166 C8_P_btm.n168 C8_P_btm.n122 0.228786
R34167 C8_P_btm.n167 C8_P_btm.n166 0.228786
R34168 C8_P_btm.n167 C8_P_btm.n121 0.228786
R34169 C8_P_btm.n140 C8_P_btm.n123 0.228786
R34170 C8_P_btm.n140 C8_P_btm.n120 0.228786
R34171 C8_P_btm.n143 C8_P_btm.n141 0.228786
R34172 C8_P_btm.n143 C8_P_btm.n142 0.228786
R34173 C8_P_btm.n186 C8_P_btm.n100 0.228786
R34174 C8_P_btm.n191 C8_P_btm.n190 0.228786
R34175 C8_P_btm.n189 C8_P_btm.n98 0.228786
R34176 C8_P_btm.n188 C8_P_btm.n187 0.228786
R34177 C8_P_btm.n93 C8_P_btm.n92 0.228786
R34178 C8_P_btm.n200 C8_P_btm.n199 0.228786
R34179 C8_P_btm.n201 C8_P_btm.n91 0.228786
R34180 C8_P_btm.n206 C8_P_btm.n205 0.228786
R34181 C8_P_btm.n204 C8_P_btm.n89 0.228786
R34182 C8_P_btm.n203 C8_P_btm.n202 0.228786
R34183 C8_P_btm.n84 C8_P_btm.n83 0.228786
R34184 C8_P_btm.n215 C8_P_btm.n214 0.228786
R34185 C8_P_btm.n216 C8_P_btm.n82 0.228786
R34186 C8_P_btm.n222 C8_P_btm.n221 0.228786
R34187 C8_P_btm.n220 C8_P_btm.n80 0.228786
R34188 C8_P_btm.n219 C8_P_btm.n217 0.228786
R34189 C8_P_btm.n218 C8_P_btm.n30 0.228786
R34190 C8_P_btm.n230 C8_P_btm.n31 0.228786
R34191 C8_P_btm.n235 C8_P_btm.n234 0.228786
R34192 C8_P_btm.n237 C8_P_btm.n24 0.228786
R34193 C8_P_btm.n236 C8_P_btm.n21 0.228786
R34194 C8_P_btm.n239 C8_P_btm.n238 0.228786
R34195 C8_P_btm.n241 C8_P_btm.n18 0.228786
R34196 C8_P_btm.n240 C8_P_btm.n17 0.228786
R34197 C8_P_btm.n243 C8_P_btm.n242 0.228786
R34198 C8_P_btm.n245 C8_P_btm.n16 0.228786
R34199 C8_P_btm.n244 C8_P_btm.n13 0.228786
R34200 C8_P_btm.n247 C8_P_btm.n246 0.228786
R34201 C8_P_btm.n249 C8_P_btm.n10 0.228786
R34202 C8_P_btm.n248 C8_P_btm.n9 0.228786
R34203 C8_P_btm.n74 C8_P_btm.n33 0.228786
R34204 C8_P_btm.n72 C8_P_btm.n34 0.228786
R34205 C8_P_btm.n36 C8_P_btm.n35 0.228786
R34206 C8_P_btm.n42 C8_P_btm.n41 0.228786
R34207 C8_P_btm.n43 C8_P_btm.n42 0.228786
R34208 C8_P_btm.n67 C8_P_btm.n43 0.228786
R34209 C8_P_btm.n68 C8_P_btm.n44 0.228786
R34210 C8_P_btm.n67 C8_P_btm.n66 0.228786
R34211 C8_P_btm.n66 C8_P_btm.n65 0.228786
R34212 C8_P_btm.n65 C8_P_btm.n45 0.228786
R34213 C8_P_btm.n46 C8_P_btm.n45 0.228786
R34214 C8_P_btm.n47 C8_P_btm.n46 0.228786
R34215 C8_P_btm.n48 C8_P_btm.n47 0.228786
R34216 C8_P_btm.n49 C8_P_btm.n48 0.228786
R34217 C8_P_btm.n50 C8_P_btm.n49 0.228786
R34218 C8_P_btm.n51 C8_P_btm.n50 0.228786
R34219 C8_P_btm.n26 C8_P_btm.n24 0.228786
R34220 C8_P_btm.n234 C8_P_btm.n233 0.228786
R34221 C8_P_btm.n232 C8_P_btm.n231 0.228786
R34222 C8_P_btm.n230 C8_P_btm.n229 0.228786
R34223 C8_P_btm.n32 C8_P_btm.n30 0.228786
R34224 C8_P_btm.n217 C8_P_btm.n78 0.228786
R34225 C8_P_btm.n224 C8_P_btm.n80 0.228786
R34226 C8_P_btm.n223 C8_P_btm.n222 0.228786
R34227 C8_P_btm.n82 C8_P_btm.n81 0.228786
R34228 C8_P_btm.n214 C8_P_btm.n213 0.228786
R34229 C8_P_btm.n85 C8_P_btm.n84 0.228786
R34230 C8_P_btm.n202 C8_P_btm.n87 0.228786
R34231 C8_P_btm.n208 C8_P_btm.n89 0.228786
R34232 C8_P_btm.n207 C8_P_btm.n206 0.228786
R34233 C8_P_btm.n91 C8_P_btm.n90 0.228786
R34234 C8_P_btm.n199 C8_P_btm.n198 0.228786
R34235 C8_P_btm.n94 C8_P_btm.n93 0.228786
R34236 C8_P_btm.n187 C8_P_btm.n96 0.228786
R34237 C8_P_btm.n193 C8_P_btm.n98 0.228786
R34238 C8_P_btm.n192 C8_P_btm.n191 0.228786
R34239 C8_P_btm.n100 C8_P_btm.n99 0.228786
R34240 C8_P_btm.n111 C8_P_btm.n109 0.228786
R34241 C8_P_btm.n181 C8_P_btm.n106 0.228786
R34242 C8_P_btm.n112 C8_P_btm.n104 0.228786
R34243 C8_P_btm.n110 C8_P_btm.n101 0.228786
R34244 C8_P_btm.n184 C8_P_btm.n183 0.228786
R34245 C8_P_btm.n120 C8_P_btm.n119 0.228786
R34246 C8_P_btm.n142 C8_P_btm.n102 0.228786
R34247 C8_P_btm.n174 C8_P_btm.n107 0.228786
R34248 C8_P_btm.n175 C8_P_btm.n116 0.228786
R34249 C8_P_btm.n173 C8_P_btm.n172 0.228786
R34250 C8_P_btm.n170 C8_P_btm.n118 0.228786
R34251 C8_P_btm.n171 C8_P_btm.n121 0.228786
R34252 C8_P_btm.n144 C8_P_btm.n103 0.228786
R34253 C8_P_btm.n145 C8_P_btm.n144 0.228786
R34254 C8_P_btm.n146 C8_P_btm.n145 0.228786
R34255 C8_P_btm.n139 C8_P_btm.n138 0.228786
R34256 C8_P_btm.n147 C8_P_btm.n146 0.228786
R34257 C8_P_btm.n148 C8_P_btm.n147 0.228786
R34258 C8_P_btm.n127 C8_P_btm.n126 0.228786
R34259 C8_P_btm.n150 C8_P_btm.n149 0.228786
R34260 C8_P_btm.n148 C8_P_btm.n137 0.228786
R34261 C8_P_btm.n137 C8_P_btm.n134 0.228786
R34262 C8_P_btm.n154 C8_P_btm.n153 0.228786
R34263 C8_P_btm.n153 C8_P_btm.n134 0.228786
R34264 C8_P_btm.n152 C8_P_btm.n151 0.228786
R34265 C8_P_btm.n157 C8_P_btm.n131 0.228786
R34266 C8_P_btm.n133 C8_P_btm.n132 0.228786
R34267 C8_P_btm.n184 C8_P_btm.n103 0.228786
R34268 C8_P_btm.n236 C8_P_btm.n235 0.228786
R34269 C8_P_btm.n238 C8_P_btm.n237 0.228786
R34270 C8_P_btm.n21 C8_P_btm.n18 0.228786
R34271 C8_P_btm.n240 C8_P_btm.n239 0.228786
R34272 C8_P_btm.n242 C8_P_btm.n241 0.228786
R34273 C8_P_btm.n17 C8_P_btm.n16 0.228786
R34274 C8_P_btm.n244 C8_P_btm.n243 0.228786
R34275 C8_P_btm.n246 C8_P_btm.n245 0.228786
R34276 C8_P_btm.n13 C8_P_btm.n10 0.228786
R34277 C8_P_btm.n248 C8_P_btm.n247 0.228786
R34278 C8_P_btm.n250 C8_P_btm.n249 0.228786
R34279 C8_P_btm.n177 C8_P_btm.n115 0.208893
R34280 C8_P_btm.n156 C8_P_btm.n130 0.208893
R34281 C8_P_btm.n234 C8_P_btm.n25 0.208893
R34282 C8_P_btm.n40 C8_P_btm.n39 0.208893
R34283 C8_P_btm.n53 C8_P_btm.n52 0.208893
R34284 C8_P_btm.n156 C8_P_btm.n155 0.208893
R34285 C8_P_btm.n185 C8_P_btm.n184 0.208893
R34286 C8_P_btm.n171 C8_P_btm.n120 0.09425
R34287 C8_P_btm.n142 C8_P_btm.n119 0.09425
R34288 C8_P_btm.n183 C8_P_btm.n101 0.09425
R34289 C8_P_btm.n110 C8_P_btm.n100 0.09425
R34290 C8_P_btm.n70 C8_P_btm.n26 0.09425
R34291 C8_P_btm.n72 C8_P_btm.n35 0.09425
R34292 C8_P_btm.n74 C8_P_btm.n34 0.09425
R34293 C8_P_btm.n76 C8_P_btm.n33 0.09425
R34294 C8_P_btm.n39 C8_P_btm.n33 0.09425
R34295 C8_P_btm.n38 C8_P_btm.n34 0.09425
R34296 C8_P_btm.n41 C8_P_btm.n35 0.09425
R34297 C8_P_btm.n42 C8_P_btm.n36 0.09425
R34298 C8_P_btm.n68 C8_P_btm.n37 0.09425
R34299 C8_P_btm.n68 C8_P_btm.n67 0.09425
R34300 C8_P_btm.n66 C8_P_btm.n44 0.09425
R34301 C8_P_btm.n63 C8_P_btm.n45 0.09425
R34302 C8_P_btm.n61 C8_P_btm.n47 0.09425
R34303 C8_P_btm.n57 C8_P_btm.n49 0.09425
R34304 C8_P_btm.n55 C8_P_btm.n51 0.09425
R34305 C8_P_btm.n52 C8_P_btm.n9 0.09425
R34306 C8_P_btm.n54 C8_P_btm.n11 0.09425
R34307 C8_P_btm.n247 C8_P_btm.n12 0.09425
R34308 C8_P_btm.n55 C8_P_btm.n12 0.09425
R34309 C8_P_btm.n56 C8_P_btm.n14 0.09425
R34310 C8_P_btm.n56 C8_P_btm.n50 0.09425
R34311 C8_P_btm.n245 C8_P_btm.n15 0.09425
R34312 C8_P_btm.n57 C8_P_btm.n15 0.09425
R34313 C8_P_btm.n59 C8_P_btm.n58 0.09425
R34314 C8_P_btm.n58 C8_P_btm.n48 0.09425
R34315 C8_P_btm.n60 C8_P_btm.n17 0.09425
R34316 C8_P_btm.n61 C8_P_btm.n60 0.09425
R34317 C8_P_btm.n62 C8_P_btm.n19 0.09425
R34318 C8_P_btm.n62 C8_P_btm.n46 0.09425
R34319 C8_P_btm.n239 C8_P_btm.n20 0.09425
R34320 C8_P_btm.n63 C8_P_btm.n20 0.09425
R34321 C8_P_btm.n64 C8_P_btm.n22 0.09425
R34322 C8_P_btm.n65 C8_P_btm.n64 0.09425
R34323 C8_P_btm.n237 C8_P_btm.n23 0.09425
R34324 C8_P_btm.n44 C8_P_btm.n23 0.09425
R34325 C8_P_btm.n70 C8_P_btm.n69 0.09425
R34326 C8_P_btm.n69 C8_P_btm.n43 0.09425
R34327 C8_P_btm.n233 C8_P_btm.n27 0.09425
R34328 C8_P_btm.n71 C8_P_btm.n27 0.09425
R34329 C8_P_btm.n71 C8_P_btm.n36 0.09425
R34330 C8_P_btm.n231 C8_P_btm.n28 0.09425
R34331 C8_P_btm.n73 C8_P_btm.n28 0.09425
R34332 C8_P_btm.n73 C8_P_btm.n72 0.09425
R34333 C8_P_btm.n75 C8_P_btm.n29 0.09425
R34334 C8_P_btm.n75 C8_P_btm.n74 0.09425
R34335 C8_P_btm.n228 C8_P_btm.n77 0.09425
R34336 C8_P_btm.n77 C8_P_btm.n76 0.09425
R34337 C8_P_btm.n229 C8_P_btm.n32 0.09425
R34338 C8_P_btm.n229 C8_P_btm.n29 0.09425
R34339 C8_P_btm.n227 C8_P_btm.n226 0.09425
R34340 C8_P_btm.n228 C8_P_btm.n227 0.09425
R34341 C8_P_btm.n224 C8_P_btm.n78 0.09425
R34342 C8_P_btm.n78 C8_P_btm.n32 0.09425
R34343 C8_P_btm.n225 C8_P_btm.n79 0.09425
R34344 C8_P_btm.n226 C8_P_btm.n225 0.09425
R34345 C8_P_btm.n223 C8_P_btm.n81 0.09425
R34346 C8_P_btm.n224 C8_P_btm.n223 0.09425
R34347 C8_P_btm.n212 C8_P_btm.n86 0.09425
R34348 C8_P_btm.n86 C8_P_btm.n79 0.09425
R34349 C8_P_btm.n213 C8_P_btm.n85 0.09425
R34350 C8_P_btm.n213 C8_P_btm.n81 0.09425
R34351 C8_P_btm.n211 C8_P_btm.n210 0.09425
R34352 C8_P_btm.n212 C8_P_btm.n211 0.09425
R34353 C8_P_btm.n208 C8_P_btm.n87 0.09425
R34354 C8_P_btm.n87 C8_P_btm.n85 0.09425
R34355 C8_P_btm.n209 C8_P_btm.n88 0.09425
R34356 C8_P_btm.n207 C8_P_btm.n90 0.09425
R34357 C8_P_btm.n208 C8_P_btm.n207 0.09425
R34358 C8_P_btm.n197 C8_P_btm.n95 0.09425
R34359 C8_P_btm.n95 C8_P_btm.n88 0.09425
R34360 C8_P_btm.n198 C8_P_btm.n94 0.09425
R34361 C8_P_btm.n198 C8_P_btm.n90 0.09425
R34362 C8_P_btm.n196 C8_P_btm.n195 0.09425
R34363 C8_P_btm.n197 C8_P_btm.n196 0.09425
R34364 C8_P_btm.n193 C8_P_btm.n96 0.09425
R34365 C8_P_btm.n96 C8_P_btm.n94 0.09425
R34366 C8_P_btm.n194 C8_P_btm.n97 0.09425
R34367 C8_P_btm.n195 C8_P_btm.n194 0.09425
R34368 C8_P_btm.n192 C8_P_btm.n99 0.09425
R34369 C8_P_btm.n193 C8_P_btm.n192 0.09425
R34370 C8_P_btm.n108 C8_P_btm.n97 0.09425
R34371 C8_P_btm.n109 C8_P_btm.n108 0.09425
R34372 C8_P_btm.n115 C8_P_btm.n114 0.09425
R34373 C8_P_btm.n179 C8_P_btm.n106 0.09425
R34374 C8_P_btm.n112 C8_P_btm.n106 0.09425
R34375 C8_P_btm.n114 C8_P_btm.n113 0.09425
R34376 C8_P_btm.n113 C8_P_btm.n109 0.09425
R34377 C8_P_btm.n112 C8_P_btm.n111 0.09425
R34378 C8_P_btm.n111 C8_P_btm.n99 0.09425
R34379 C8_P_btm.n181 C8_P_btm.n104 0.09425
R34380 C8_P_btm.n110 C8_P_btm.n104 0.09425
R34381 C8_P_btm.n184 C8_P_btm.n102 0.09425
R34382 C8_P_btm.n173 C8_P_btm.n117 0.09425
R34383 C8_P_btm.n117 C8_P_btm.n102 0.09425
R34384 C8_P_btm.n182 C8_P_btm.n105 0.09425
R34385 C8_P_btm.n183 C8_P_btm.n182 0.09425
R34386 C8_P_btm.n180 C8_P_btm.n107 0.09425
R34387 C8_P_btm.n181 C8_P_btm.n180 0.09425
R34388 C8_P_btm.n179 C8_P_btm.n178 0.09425
R34389 C8_P_btm.n176 C8_P_btm.n107 0.09425
R34390 C8_P_btm.n175 C8_P_btm.n174 0.09425
R34391 C8_P_btm.n174 C8_P_btm.n105 0.09425
R34392 C8_P_btm.n173 C8_P_btm.n116 0.09425
R34393 C8_P_btm.n172 C8_P_btm.n118 0.09425
R34394 C8_P_btm.n172 C8_P_btm.n119 0.09425
R34395 C8_P_btm.n171 C8_P_btm.n170 0.09425
R34396 C8_P_btm.n169 C8_P_btm.n121 0.09425
R34397 C8_P_btm.n133 C8_P_btm.n131 0.09425
R34398 C8_P_btm.n135 C8_P_btm.n129 0.09425
R34399 C8_P_btm.n149 C8_P_btm.n126 0.09425
R34400 C8_P_btm.n145 C8_P_btm.n141 0.09425
R34401 C8_P_btm.n139 C8_P_btm.n123 0.09425
R34402 C8_P_btm.n146 C8_P_btm.n139 0.09425
R34403 C8_P_btm.n166 C8_P_btm.n124 0.09425
R34404 C8_P_btm.n138 C8_P_btm.n124 0.09425
R34405 C8_P_btm.n147 C8_P_btm.n138 0.09425
R34406 C8_P_btm.n149 C8_P_btm.n148 0.09425
R34407 C8_P_btm.n150 C8_P_btm.n137 0.09425
R34408 C8_P_btm.n151 C8_P_btm.n136 0.09425
R34409 C8_P_btm.n151 C8_P_btm.n134 0.09425
R34410 C8_P_btm.n164 C8_P_btm.n127 0.09425
R34411 C8_P_btm.n150 C8_P_btm.n127 0.09425
R34412 C8_P_btm.n152 C8_P_btm.n135 0.09425
R34413 C8_P_btm.n153 C8_P_btm.n152 0.09425
R34414 C8_P_btm.n154 C8_P_btm.n133 0.09425
R34415 C8_P_btm.n158 C8_P_btm.n157 0.09425
R34416 C8_P_btm.n157 C8_P_btm.n132 0.09425
R34417 C8_P_btm.n160 C8_P_btm.n159 0.09425
R34418 C8_P_btm.n159 C8_P_btm.n131 0.09425
R34419 C8_P_btm.n161 C8_P_btm.n129 0.09425
R34420 C8_P_btm.n162 C8_P_btm.n128 0.09425
R34421 C8_P_btm.n136 C8_P_btm.n128 0.09425
R34422 C8_P_btm.n164 C8_P_btm.n163 0.09425
R34423 C8_P_btm.n165 C8_P_btm.n125 0.09425
R34424 C8_P_btm.n165 C8_P_btm.n126 0.09425
R34425 C8_P_btm.n166 C8_P_btm.n122 0.09425
R34426 C8_P_btm.n168 C8_P_btm.n167 0.09425
R34427 C8_P_btm.n167 C8_P_btm.n123 0.09425
R34428 C8_P_btm.n140 C8_P_btm.n121 0.09425
R34429 C8_P_btm.n141 C8_P_btm.n140 0.09425
R34430 C8_P_btm.n143 C8_P_btm.n120 0.09425
R34431 C8_P_btm.n144 C8_P_btm.n143 0.09425
R34432 C8_P_btm.n142 C8_P_btm.n103 0.09425
R34433 C8_P_btm.n190 C8_P_btm.n186 0.09425
R34434 C8_P_btm.n191 C8_P_btm.n100 0.09425
R34435 C8_P_btm.n191 C8_P_btm.n98 0.09425
R34436 C8_P_btm.n190 C8_P_btm.n189 0.09425
R34437 C8_P_btm.n189 C8_P_btm.n188 0.09425
R34438 C8_P_btm.n187 C8_P_btm.n98 0.09425
R34439 C8_P_btm.n187 C8_P_btm.n93 0.09425
R34440 C8_P_btm.n188 C8_P_btm.n92 0.09425
R34441 C8_P_btm.n200 C8_P_btm.n92 0.09425
R34442 C8_P_btm.n199 C8_P_btm.n93 0.09425
R34443 C8_P_btm.n199 C8_P_btm.n91 0.09425
R34444 C8_P_btm.n201 C8_P_btm.n200 0.09425
R34445 C8_P_btm.n205 C8_P_btm.n201 0.09425
R34446 C8_P_btm.n206 C8_P_btm.n91 0.09425
R34447 C8_P_btm.n206 C8_P_btm.n89 0.09425
R34448 C8_P_btm.n205 C8_P_btm.n204 0.09425
R34449 C8_P_btm.n204 C8_P_btm.n203 0.09425
R34450 C8_P_btm.n202 C8_P_btm.n89 0.09425
R34451 C8_P_btm.n202 C8_P_btm.n84 0.09425
R34452 C8_P_btm.n203 C8_P_btm.n83 0.09425
R34453 C8_P_btm.n215 C8_P_btm.n83 0.09425
R34454 C8_P_btm.n214 C8_P_btm.n84 0.09425
R34455 C8_P_btm.n214 C8_P_btm.n82 0.09425
R34456 C8_P_btm.n216 C8_P_btm.n215 0.09425
R34457 C8_P_btm.n221 C8_P_btm.n216 0.09425
R34458 C8_P_btm.n222 C8_P_btm.n82 0.09425
R34459 C8_P_btm.n222 C8_P_btm.n80 0.09425
R34460 C8_P_btm.n221 C8_P_btm.n220 0.09425
R34461 C8_P_btm.n220 C8_P_btm.n219 0.09425
R34462 C8_P_btm.n217 C8_P_btm.n80 0.09425
R34463 C8_P_btm.n217 C8_P_btm.n30 0.09425
R34464 C8_P_btm.n219 C8_P_btm.n218 0.09425
R34465 C8_P_btm.n218 C8_P_btm.n31 0.09425
R34466 C8_P_btm.n230 C8_P_btm.n30 0.09425
R34467 C8_P_btm.n231 C8_P_btm.n230 0.09425
R34468 C8_P_btm.n233 C8_P_btm.n232 0.09425
R34469 C8_P_btm.n234 C8_P_btm.n26 0.09425
R34470 C8_P_btm.n235 C8_P_btm.n24 0.09425
R34471 C8_P_btm.n37 C8_P_btm.n24 0.09425
R34472 C8_P_btm.n237 C8_P_btm.n236 0.09425
R34473 C8_P_btm.n238 C8_P_btm.n21 0.09425
R34474 C8_P_btm.n238 C8_P_btm.n22 0.09425
R34475 C8_P_btm.n239 C8_P_btm.n18 0.09425
R34476 C8_P_btm.n241 C8_P_btm.n240 0.09425
R34477 C8_P_btm.n240 C8_P_btm.n19 0.09425
R34478 C8_P_btm.n242 C8_P_btm.n17 0.09425
R34479 C8_P_btm.n243 C8_P_btm.n16 0.09425
R34480 C8_P_btm.n59 C8_P_btm.n16 0.09425
R34481 C8_P_btm.n245 C8_P_btm.n244 0.09425
R34482 C8_P_btm.n246 C8_P_btm.n13 0.09425
R34483 C8_P_btm.n246 C8_P_btm.n14 0.09425
R34484 C8_P_btm.n247 C8_P_btm.n10 0.09425
R34485 C8_P_btm.n249 C8_P_btm.n248 0.09425
R34486 C8_P_btm.n248 C8_P_btm.n11 0.09425
R34487 C8_P_btm.n250 C8_P_btm.n9 0.09425
R34488 C8_P_btm.n210 C8_P_btm.n209 0.0816039
R34489 C8_P_btm.n186 C8_P_btm.n185 0.047875
R34490 C8_P_btm.n31 C8_P_btm.n25 0.047875
R34491 C8_P_btm.n54 C8_P_btm.n53 0.0342289
R34492 C8_P_btm.n155 C8_P_btm.n132 0.0342289
R34493 C8_P_btm.n185 C8_P_btm.n101 0.0342289
R34494 C8_P_btm.n40 C8_P_btm.n38 0.0342289
R34495 C8_P_btm.n178 C8_P_btm.n177 0.0342289
R34496 C8_P_btm.n158 C8_P_btm.n130 0.0342289
R34497 C8_P_btm.n232 C8_P_btm.n25 0.0342289
R34498 a_5342_30871.n2 a_5342_30871.t6 1421.83
R34499 a_5342_30871.n1 a_5342_30871.t5 1421.83
R34500 a_5342_30871.n2 a_5342_30871.t9 1320.68
R34501 a_5342_30871.n1 a_5342_30871.t4 1320.68
R34502 a_5342_30871.n7 a_5342_30871.n6 380.32
R34503 a_5342_30871.n0 a_5342_30871.t8 260.322
R34504 a_5342_30871.n3 a_5342_30871.n2 194.02
R34505 a_5342_30871.n3 a_5342_30871.n1 192.049
R34506 a_5342_30871.n6 a_5342_30871.n5 185
R34507 a_5342_30871.n0 a_5342_30871.t7 175.169
R34508 a_5342_30871.n4 a_5342_30871.n0 172.587
R34509 a_5342_30871.n4 a_5342_30871.n3 68.7679
R34510 a_5342_30871.t1 a_5342_30871.n7 26.5955
R34511 a_5342_30871.n7 a_5342_30871.t0 26.5955
R34512 a_5342_30871.n5 a_5342_30871.t3 24.9236
R34513 a_5342_30871.n5 a_5342_30871.t2 24.9236
R34514 a_5342_30871.n6 a_5342_30871.n4 20.9746
R34515 START.n0 START.t0 260.322
R34516 START.n0 START.t1 175.169
R34517 START START.n0 175.018
R34518 EN_OFFSET_CAL.n0 EN_OFFSET_CAL.t0 260.322
R34519 EN_OFFSET_CAL EN_OFFSET_CAL.n0 175.327
R34520 EN_OFFSET_CAL.n0 EN_OFFSET_CAL.t1 175.169
C0 a_2479_44172# a_2905_42968# 0.163227f
C1 a_n863_45724# a_n452_44636# 0.01836f
C2 C3_N_btm VDD 0.26836f
C3 a_18597_46090# a_19123_46287# 0.188676f
C4 a_18479_47436# a_20107_46660# 0.019527f
C5 C7_P_btm VIN_P 1.52449f
C6 C7_N_btm C8_N_btm 31.072699f
C7 C6_N_btm C9_N_btm 0.165353f
C8 C5_N_btm C10_N_btm 0.51798f
C9 C9_P_btm VREF 7.369471f
C10 C10_P_btm VREF_GND 10.3207f
C11 a_20301_43646# a_20556_43646# 0.114664f
C12 a_n2661_45010# a_n23_44458# 0.049334f
C13 a_2479_44172# VDD 0.431428f
C14 a_13720_44458# a_13857_44734# 0.126609f
C15 a_4007_47204# VDD 0.41212f
C16 a_14537_43396# a_15682_43940# 0.01288f
C17 a_12465_44636# a_14180_45002# 0.015526f
C18 a_2998_44172# a_3600_43914# 0.012242f
C19 a_15368_46634# VDD 0.324877f
C20 a_2382_45260# a_3681_42891# 0.067836f
C21 a_3316_45546# a_3175_45822# 0.05019f
C22 a_n2104_42282# VDD 0.280329f
C23 a_5343_44458# a_8292_43218# 0.01105f
C24 a_17715_44484# a_17767_44458# 0.07408f
C25 a_7754_38470# VDD 0.302129f
C26 VDAC_P C6_P_btm 55.214397f
C27 a_15681_43442# a_15781_43660# 0.167615f
C28 a_2680_45002# VDD 0.145087f
C29 a_22959_45572# a_22959_45036# 0.026152f
C30 a_n863_45724# a_n809_44244# 0.016179f
C31 a_5807_45002# a_14275_46494# 0.013842f
C32 a_15743_43084# a_22400_42852# 0.010325f
C33 a_5257_43370# a_6194_45824# 0.029055f
C34 a_n2497_47436# a_375_42282# 0.018989f
C35 COMP_P a_n1329_42308# 0.232443f
C36 a_n229_43646# VDD 0.278436f
C37 a_2864_46660# VDD 0.076834f
C38 a_10057_43914# a_10555_44260# 0.041594f
C39 a_1467_44172# a_1427_43646# 0.104539f
C40 a_20708_46348# VDD 0.093079f
C41 a_1138_42852# a_949_44458# 0.013552f
C42 a_11415_45002# a_14539_43914# 0.010769f
C43 a_21496_47436# a_20916_46384# 0.113102f
C44 a_4574_45260# a_4558_45348# 0.19344f
C45 a_7499_43078# a_5883_43914# 0.100372f
C46 a_9049_44484# a_8701_44490# 0.100038f
C47 a_20916_46384# a_21363_46634# 0.017401f
C48 a_15743_43084# a_22223_42860# 0.021215f
C49 a_5518_44484# VDD 0.40715f
C50 a_13059_46348# a_13351_46090# 0.074689f
C51 a_5807_45002# a_6194_45824# 0.02442f
C52 a_n2157_46122# a_n1991_46122# 0.614266f
C53 a_n863_45724# a_n2293_42282# 0.028166f
C54 a_16922_45042# a_20269_44172# 0.010825f
C55 a_14815_43914# a_14673_44172# 0.173231f
C56 a_n2497_47436# a_4181_44734# 0.01129f
C57 a_18597_46090# a_20193_45348# 0.021804f
C58 a_3877_44458# a_3065_45002# 0.287919f
C59 a_18579_44172# a_19319_43548# 0.031277f
C60 a_8162_45546# a_7499_43078# 0.021916f
C61 a_11415_45002# a_14309_45028# 0.040538f
C62 a_18479_47436# a_19386_47436# 0.219411f
C63 a_18780_47178# a_18597_46090# 0.175179f
C64 a_13070_42354# VDD 0.18656f
C65 a_22485_38105# a_22527_39145# 0.984424f
C66 a_1568_43370# a_1756_43548# 0.094732f
C67 a_2479_44172# a_2075_43172# 0.034186f
C68 a_8746_45002# a_8560_45348# 0.044092f
C69 C2_N_btm VDD 0.268945f
C70 a_18597_46090# a_18285_46348# 0.012666f
C71 C8_P_btm VIN_P 0.907642f
C72 C6_N_btm C8_N_btm 0.163943f
C73 C4_N_btm C10_N_btm 0.703336f
C74 C5_N_btm C9_N_btm 0.150576f
C75 C10_P_btm VREF 14.773f
C76 a_21259_43561# a_21487_43396# 0.08444f
C77 a_17339_46660# a_19095_43396# 0.049229f
C78 a_2127_44172# VDD 0.138239f
C79 a_3815_47204# VDD 0.260661f
C80 a_14537_43396# a_14955_43940# 0.104291f
C81 a_22223_45036# a_22315_44484# 0.011923f
C82 a_n1549_44318# a_n1453_44318# 0.013793f
C83 a_14976_45028# VDD 0.484864f
C84 a_n699_43396# a_n1557_42282# 0.02911f
C85 a_10586_45546# a_10907_45822# 0.05477f
C86 a_3218_45724# a_3175_45822# 0.132424f
C87 a_18051_46116# VDD 0.189782f
C88 a_22629_37990# a_22725_37990# 0.087835f
C89 VDAC_P C7_P_btm 0.11042p
C90 a_2382_45260# VDD 1.6285f
C91 a_7499_43078# a_11541_44484# 0.048175f
C92 a_12251_46660# a_12347_46660# 0.013793f
C93 a_n2661_46098# a_1138_42852# 0.020229f
C94 a_15433_44458# VDD 0.201121f
C95 a_5257_43370# a_5907_45546# 0.064039f
C96 a_20835_44721# a_21145_44484# 0.013793f
C97 a_3524_46660# VDD 0.278519f
C98 a_18989_43940# a_18451_43940# 0.114286f
C99 a_11189_46129# a_10907_45822# 0.021145f
C100 a_19511_42282# a_20712_42282# 0.05034f
C101 a_19900_46494# VDD 0.279179f
C102 a_1138_42852# a_742_44458# 0.040731f
C103 a_10907_45822# a_11136_45572# 0.080042f
C104 a_1169_39587# VDD 0.531695f
C105 a_8953_45546# a_9028_43914# 0.01093f
C106 a_7499_43078# a_8701_44490# 0.011795f
C107 a_10249_46116# a_6755_46942# 0.068878f
C108 a_5343_44458# VDD 0.49245f
C109 a_5807_45002# a_5907_45546# 0.013402f
C110 a_13059_46348# a_12594_46348# 0.03479f
C111 a_n2157_46122# a_n1853_46287# 0.617317f
C112 a_16922_45042# a_19862_44208# 0.038132f
C113 a_13059_46348# a_15037_45618# 0.064109f
C114 a_8162_45546# a_8568_45546# 0.078784f
C115 a_18479_47436# a_18597_46090# 0.473843f
C116 a_12563_42308# VDD 0.254292f
C117 a_22485_38105# a_22589_40055# 0.212168f
C118 a_19862_44208# a_15743_43084# 0.022478f
C119 a_2479_44172# a_1847_42826# 0.141223f
C120 C1_N_btm VDD 0.264503f
C121 a_12465_44636# a_13059_46348# 0.163448f
C122 C9_P_btm VIN_P 1.82823f
C123 C4_N_btm C9_N_btm 0.154834f
C124 C3_N_btm C10_N_btm 0.321945f
C125 C5_N_btm C8_N_btm 0.145019f
C126 C6_N_btm C7_N_btm 26.0771f
C127 a_453_43940# VDD 0.225569f
C128 a_13076_44458# a_13468_44734# 0.016359f
C129 a_3785_47178# VDD 0.387755f
C130 SMPL_ON_N a_22537_40625# 0.028814f
C131 a_11827_44484# a_22315_44484# 0.013f
C132 a_18494_42460# a_20512_43084# 0.115057f
C133 a_12465_44636# a_13556_45296# 0.248126f
C134 a_2889_44172# a_2998_44172# 0.179664f
C135 a_n1549_44318# a_n1644_44306# 0.049827f
C136 a_2957_45546# a_3175_45822# 0.08213f
C137 a_10586_45546# a_10210_45822# 0.042978f
C138 a_n2472_42282# VDD 0.278905f
C139 a_22629_38406# a_22737_37285# 0.08753f
C140 VDAC_P C8_P_btm 0.220914p
C141 a_2274_45254# VDD 0.256655f
C142 a_375_42282# a_626_44172# 0.017957f
C143 a_n2661_46098# a_1176_45822# 0.144277f
C144 a_5807_45002# a_13925_46122# 0.027158f
C145 a_14815_43914# VDD 0.307386f
C146 a_3065_45002# a_3905_42865# 0.034773f
C147 a_1823_45246# a_n2293_42282# 0.03994f
C148 a_5257_43370# a_5263_45724# 0.088982f
C149 a_8199_44636# a_9625_46129# 0.011574f
C150 a_8016_46348# a_9823_46155# 0.048283f
C151 a_n1736_42282# a_n1329_42308# 0.050456f
C152 a_3699_46634# VDD 0.347281f
C153 a_8199_44636# a_9159_45572# 0.049711f
C154 a_17303_42282# a_22397_42558# 0.012536f
C155 a_19511_42282# a_20107_42308# 0.043647f
C156 a_20075_46420# VDD 0.347847f
C157 a_8199_44636# a_9672_43914# 0.043804f
C158 a_4743_44484# VDD 0.266843f
C159 a_18597_46090# a_19511_42282# 0.156698f
C160 a_18479_47436# a_20193_45348# 0.021013f
C161 a_3877_44458# a_2382_45260# 0.395451f
C162 a_1823_45246# a_3775_45552# 0.070347f
C163 a_11415_45002# a_11652_45724# 0.128811f
C164 a_n1736_43218# VDD 0.082445f
C165 a_14456_42282# a_14113_42308# 0.038993f
C166 a_18479_47436# a_18780_47178# 0.056304f
C167 a_11633_42558# VDD 0.193501f
C168 C0_N_btm VDD 1.02806f
C169 a_12891_46348# a_12816_46660# 0.024711f
C170 a_5807_45002# a_8270_45546# 0.029164f
C171 C10_P_btm VIN_P 3.66034f
C172 C4_N_btm C8_N_btm 0.145646f
C173 C3_N_btm C9_N_btm 0.137552f
C174 C2_N_btm C10_N_btm 0.327137f
C175 C5_N_btm C7_N_btm 0.151416f
C176 a_21753_35474# VIN_N 0.029412f
C177 a_5111_44636# a_5518_44484# 0.124556f
C178 a_1414_42308# VDD 0.657887f
C179 a_13076_44458# a_13213_44734# 0.126609f
C180 a_3381_47502# VDD 0.197761f
C181 a_12465_44636# a_9482_43914# 0.069673f
C182 a_12281_43396# VDD 0.341026f
C183 a_4921_42308# a_5755_42308# 0.175841f
C184 a_2675_43914# a_2998_44172# 0.173844f
C185 a_15009_46634# VDD 0.205396f
C186 a_12891_46348# a_13213_44734# 0.052195f
C187 a_n2302_39866# a_n2302_39072# 0.052227f
C188 a_11459_47204# a_11735_46660# 0.010464f
C189 VDAC_P C9_P_btm 0.441881p
C190 a_1667_45002# VDD 0.315476f
C191 a_n2661_46098# a_1208_46090# 0.023477f
C192 a_5807_45002# a_13759_46122# 0.022269f
C193 a_3065_45002# a_3600_43914# 0.011102f
C194 a_8016_46348# a_9569_46155# 0.044705f
C195 a_8199_44636# a_8953_45546# 0.71291f
C196 a_2959_46660# VDD 0.19762f
C197 a_18287_44626# a_19328_44172# 0.011011f
C198 a_10405_44172# a_10867_43940# 0.022925f
C199 a_19335_46494# VDD 0.198512f
C200 a_6547_43396# a_6643_43396# 0.013793f
C201 a_8016_46348# a_10405_44172# 0.098226f
C202 a_7927_46660# a_8035_47026# 0.057222f
C203 a_10554_47026# a_10249_46116# 0.023301f
C204 a_16823_43084# a_16795_42852# 0.065873f
C205 a_n699_43396# VDD 0.922998f
C206 a_7499_43078# a_10555_44260# 0.03816f
C207 a_22959_43948# VDD 0.297936f
C208 SMPL_ON_N VIN_N 0.525208f
C209 a_13575_42558# a_14113_42308# 0.11418f
C210 a_19279_43940# a_19319_43548# 0.023499f
C211 a_22959_46660# VDD 0.299681f
C212 a_11551_42558# VDD 0.192086f
C213 a_n2833_47464# a_n2840_46634# 0.019713f
C214 a_22485_38105# a_22537_40625# 0.0722f
C215 a_18597_46090# a_17339_46660# 0.018491f
C216 a_12891_46348# a_12991_46634# 0.018656f
C217 a_3699_46634# a_3877_44458# 0.087244f
C218 a_19998_34978# VIN_N 0.37444f
C219 C3_N_btm C8_N_btm 0.134581f
C220 C2_N_btm C9_N_btm 0.141891f
C221 C1_N_btm C10_N_btm 0.31753f
C222 C5_N_btm C6_N_btm 22.305399f
C223 C4_N_btm C7_N_btm 0.145303f
C224 EN_VIN_BSTR_N VCM 0.927954f
C225 a_5147_45002# a_5518_44484# 0.064422f
C226 a_5111_44636# a_5343_44458# 0.477401f
C227 a_1467_44172# VDD 0.391994f
C228 a_13556_45296# a_14955_43940# 0.059957f
C229 a_2675_43914# a_2889_44172# 0.083573f
C230 a_n1899_43946# a_n1644_44306# 0.06121f
C231 a_14084_46812# VDD 0.087769f
C232 a_n2840_42282# VDD 0.294987f
C233 a_19240_46482# VDD 0.077608f
C234 a_7227_45028# a_6709_45028# 0.115677f
C235 VDAC_Ni VDD 0.288547f
C236 a_22629_38406# a_22629_37990# 0.32625f
C237 VDAC_P C10_P_btm 0.883474p
C238 a_327_44734# VDD 0.667364f
C239 a_n2661_46098# a_805_46414# 0.044109f
C240 a_13857_44734# VDD 0.18416f
C241 a_3065_45002# a_2998_44172# 0.024536f
C242 a_2382_45260# a_3905_42865# 0.291572f
C243 a_8016_46348# a_9625_46129# 0.128435f
C244 a_n1809_43762# VDD 0.142403f
C245 a_3177_46902# VDD 0.200982f
C246 a_133_42852# VDD 0.184203f
C247 a_19511_42282# a_19647_42308# 0.038787f
C248 a_10405_44172# a_10651_43940# 0.014272f
C249 a_19553_46090# VDD 0.204238f
C250 a_n2302_39866# VDD 0.361509f
C251 a_8016_46348# a_9672_43914# 0.074243f
C252 a_7927_46660# a_7832_46660# 0.049827f
C253 a_8145_46902# a_8035_47026# 0.097745f
C254 a_10623_46897# a_10249_46116# 0.032312f
C255 a_10467_46802# a_6755_46942# 0.256039f
C256 a_12891_46348# a_11415_45002# 0.059955f
C257 a_16823_43084# a_16414_43172# 0.024882f
C258 a_n2472_46090# a_n2157_46122# 0.080495f
C259 a_15493_43940# VDD 1.4617f
C260 a_11415_45002# a_11322_45546# 0.527707f
C261 a_13575_42558# a_13657_42558# 0.171361f
C262 a_16922_45042# a_20749_43396# 0.106779f
C263 a_1823_45246# a_2809_45028# 0.076288f
C264 a_18143_47464# a_18479_47436# 0.238309f
C265 a_22485_38105# a_22589_40599# 0.132855f
C266 a_1209_43370# a_1049_43396# 0.194938f
C267 a_15493_43940# a_16137_43396# 0.043956f
C268 a_13059_46348# a_13483_43940# 0.124566f
C269 C2_N_btm C8_N_btm 0.138777f
C270 C1_N_btm C9_N_btm 0.132506f
C271 C0_N_btm C10_N_btm 0.365593f
C272 C4_N_btm C6_N_btm 0.143514f
C273 C3_N_btm C7_N_btm 0.134911f
C274 EN_VIN_BSTR_N VREF_GND 0.857366f
C275 a_5147_45002# a_5343_44458# 0.063193f
C276 a_5111_44636# a_4743_44484# 0.02485f
C277 a_16019_45002# a_16237_45028# 0.053167f
C278 a_17339_46660# a_18285_46348# 0.184197f
C279 a_1115_44172# VDD 0.165092f
C280 a_14543_43071# a_14635_42282# 0.075815f
C281 a_3160_47472# VDD 0.256092f
C282 a_13607_46688# VDD 0.209568f
C283 a_n1761_44111# a_n1644_44306# 0.170098f
C284 a_3877_44458# a_n699_43396# 0.061672f
C285 a_16375_45002# VDD 1.14948f
C286 a_7227_45028# a_7229_43940# 0.019397f
C287 a_7754_38636# VDD 0.036155f
C288 CAL_P a_22629_37990# 0.205295f
C289 a_22629_38406# a_22725_38406# 0.090011f
C290 a_n2661_46098# a_472_46348# 0.065456f
C291 a_12251_46660# a_12359_47026# 0.057222f
C292 a_2382_45260# a_3600_43914# 0.158274f
C293 a_18479_45785# a_15493_43940# 0.016583f
C294 a_14035_46660# a_14180_46482# 0.157972f
C295 a_8016_46348# a_8953_45546# 0.060003f
C296 a_n2012_43396# VDD 0.08228f
C297 a_19279_43940# a_21398_44850# 0.183186f
C298 a_2609_46660# VDD 0.312974f
C299 a_19778_44110# a_19741_43940# 0.054731f
C300 a_8199_44636# a_8192_45572# 0.04905f
C301 a_18985_46122# VDD 0.253642f
C302 a_10405_44172# a_10555_43940# 0.018661f
C303 a_15143_45578# a_15037_45618# 0.13675f
C304 a_12465_44636# a_5807_45002# 0.59474f
C305 a_7499_43078# a_5343_44458# 0.050528f
C306 a_7577_46660# a_8035_47026# 0.027606f
C307 a_10467_46802# a_10249_46116# 0.12624f
C308 a_10428_46928# a_6755_46942# 0.155315f
C309 a_10623_46897# a_10554_47026# 0.209641f
C310 a_2779_44458# VDD 0.38604f
C311 a_14035_46660# a_13925_46122# 0.207108f
C312 a_19466_46812# a_19335_46494# 0.017838f
C313 a_22223_43948# VDD 0.254313f
C314 a_13291_42460# a_14635_42282# 0.111986f
C315 a_18597_46090# a_11827_44484# 0.039373f
C316 a_n13_43084# VDD 0.260551f
C317 a_11323_42473# VDD 0.205172f
C318 a_22485_38105# CAL_N 0.072058f
C319 a_2684_37794# a_2113_38308# 0.468006f
C320 en_comp comp_n 0.026386f
C321 a_458_43396# a_1049_43396# 0.052073f
C322 C0_P_btm VDD 1.02806f
C323 C1_N_btm C8_N_btm 0.129306f
C324 C0_N_btm C9_N_btm 0.146135f
C325 C0_dummy_N_btm C10_N_btm 0.749362f
C326 C4_N_btm C5_N_btm 18.6196f
C327 C3_N_btm C6_N_btm 0.133742f
C328 C2_N_btm C7_N_btm 0.138288f
C329 a_1568_43370# a_1793_42852# 0.011559f
C330 a_8953_45546# a_8791_43396# 0.012124f
C331 a_5111_44636# a_n699_43396# 0.016349f
C332 a_644_44056# VDD 0.147321f
C333 a_14543_43071# a_13291_42460# 0.107887f
C334 a_2905_45572# VDD 1.22598f
C335 a_1431_47204# DATA[1] 0.334099f
C336 a_12816_46660# VDD 0.293798f
C337 a_895_43940# a_2675_43914# 0.099822f
C338 a_n2065_43946# a_n1644_44306# 0.090164f
C339 a_6755_46942# a_11827_44484# 0.529579f
C340 a_20753_42852# VDD 0.193909f
C341 a_7227_45028# a_7276_45260# 0.098279f
C342 a_11415_45002# a_14673_44172# 0.229077f
C343 a_n37_45144# VDD 0.138f
C344 a_22223_45572# a_22223_45036# 0.026152f
C345 a_n746_45260# a_310_45028# 0.378188f
C346 a_n2661_46098# a_376_46348# 0.060405f
C347 a_12469_46902# a_12359_47026# 0.097745f
C348 a_12251_46660# a_12156_46660# 0.049827f
C349 a_13213_44734# VDD 0.184239f
C350 a_2382_45260# a_2998_44172# 0.045272f
C351 a_8349_46414# a_8199_44636# 0.032352f
C352 a_104_43370# VDD 0.252393f
C353 a_17701_42308# a_17531_42308# 0.109201f
C354 a_2443_46660# VDD 0.413663f
C355 a_6755_46942# a_15595_45028# 0.012879f
C356 a_18819_46122# VDD 0.453432f
C357 a_20894_47436# a_20843_47204# 0.134298f
C358 a_n2946_39866# VDD 0.393552f
C359 a_16223_45938# VDD 0.132317f
C360 a_10807_43548# a_10341_42308# 0.099222f
C361 a_3065_45002# a_3429_45260# 0.037292f
C362 a_10467_46802# a_10554_47026# 0.07009f
C363 a_10428_46928# a_10249_46116# 0.704177f
C364 a_7577_46660# a_7832_46660# 0.056391f
C365 a_949_44458# VDD 1.2275f
C366 a_19700_43370# a_19339_43156# 0.012115f
C367 a_11827_44484# a_20193_45348# 0.051742f
C368 a_12465_44636# a_14495_45572# 0.019417f
C369 a_14035_46660# a_13759_46122# 0.162408f
C370 SMPL_ON_N EN_OFFSET_CAL 0.066251f
C371 a_n1076_43230# VDD 0.292942f
C372 COMP_P a_1169_39587# 0.388738f
C373 a_13070_42354# a_13333_42558# 0.011552f
C374 a_22591_46660# VDD 0.251892f
C375 a_10723_42308# VDD 0.223902f
C376 a_458_43396# a_1209_43370# 0.0172f
C377 a_12465_44636# a_14513_46634# 0.01549f
C378 C1_P_btm VDD 0.264503f
C379 a_12891_46348# a_11901_46660# 0.028795f
C380 a_2959_46660# a_3055_46660# 0.013793f
C381 EN_VIN_BSTR_N VIN_N 1.41696f
C382 C3_N_btm C5_N_btm 0.135528f
C383 C0_N_btm C8_N_btm 0.146541f
C384 C0_dummy_N_btm C9_N_btm 0.111645f
C385 C2_N_btm C6_N_btm 0.137206f
C386 C1_N_btm C7_N_btm 0.128479f
C387 EN_VIN_BSTR_P VCM 0.929382f
C388 a_1568_43370# a_1709_42852# 0.015873f
C389 a_175_44278# VDD 0.20887f
C390 a_2952_47436# VDD 0.089131f
C391 a_9482_43914# a_12429_44172# 0.0636f
C392 a_1239_47204# DATA[1] 0.01925f
C393 a_8199_44636# a_8034_45724# 0.127067f
C394 a_4933_42558# a_4921_42308# 0.012385f
C395 a_5379_42460# a_6171_42473# 0.110293f
C396 a_12991_46634# VDD 0.357655f
C397 a_1414_42308# a_3600_43914# 0.012293f
C398 a_2479_44172# a_2675_43914# 0.061502f
C399 a_18597_46090# a_19279_43940# 0.021978f
C400 a_997_45618# a_1260_45572# 0.010598f
C401 a_n2946_39866# a_n2946_39072# 0.052227f
C402 a_n143_45144# VDD 0.092f
C403 a_n746_45260# a_n1099_45572# 0.015931f
C404 a_n2661_46098# a_n1076_46494# 0.037593f
C405 a_11901_46660# a_12359_47026# 0.034619f
C406 a_13635_43156# a_14543_43071# 0.013803f
C407 a_6298_44484# a_8103_44636# 0.016067f
C408 a_5343_44458# a_5883_43914# 0.042199f
C409 a_8016_46348# a_8199_44636# 0.33718f
C410 a_17701_42308# a_17303_42282# 0.049097f
C411 a_20835_44721# a_21398_44850# 0.049827f
C412 a_20766_44850# a_20980_44850# 0.097745f
C413 a_n2661_46098# VDD 0.979859f
C414 a_18494_42460# a_19319_43548# 0.016978f
C415 a_17303_42282# a_21613_42308# 0.061584f
C416 a_17957_46116# VDD 0.138777f
C417 a_742_44458# a_2905_42968# 0.15065f
C418 a_9672_43914# a_9801_43940# 0.062574f
C419 a_16020_45572# VDD 0.077625f
C420 a_10807_43548# a_10922_42852# 0.010566f
C421 a_10150_46912# a_10249_46116# 0.066949f
C422 a_10467_46802# a_10623_46897# 0.107482f
C423 a_7715_46873# a_7832_46660# 0.157972f
C424 a_9863_46634# a_6755_46942# 0.014818f
C425 a_10428_46928# a_10554_47026# 0.181217f
C426 a_742_44458# VDD 1.3845f
C427 a_15743_43084# a_19164_43230# 0.0353f
C428 a_12465_44636# a_13249_42308# 0.541909f
C429 a_19466_46812# a_18985_46122# 0.033782f
C430 a_21115_43940# VDD 0.145936f
C431 a_18479_47436# a_11827_44484# 0.035345f
C432 a_18597_46090# a_21101_45002# 0.033595f
C433 a_n901_43156# VDD 0.475947f
C434 a_9803_42558# a_10149_42308# 0.013377f
C435 a_13070_42354# a_13249_42558# 0.010303f
C436 a_11415_45002# VDD 1.84504f
C437 a_16375_45002# a_16147_45260# 1.01554f
C438 a_10533_42308# VDD 0.216201f
C439 a_12465_44636# a_14180_46812# 0.026945f
C440 C2_P_btm VDD 0.268945f
C441 C2_N_btm C5_N_btm 0.13795f
C442 C3_N_btm C4_N_btm 9.61674f
C443 C1_N_btm C6_N_btm 0.127656f
C444 C0_dummy_N_btm C8_N_btm 0.234177f
C445 C0_N_btm C7_N_btm 0.140846f
C446 EN_VIN_BSTR_P VREF_GND 0.857366f
C447 a_n984_44318# VDD 0.281427f
C448 a_2553_47502# VDD 0.150286f
C449 a_20193_45348# a_19279_43940# 0.021458f
C450 a_9482_43914# a_11750_44172# 0.020902f
C451 a_1209_47178# DATA[1] 0.076054f
C452 a_8349_46414# a_8034_45724# 0.05863f
C453 a_9885_43646# VDD 0.190473f
C454 a_12251_46660# VDD 0.195617f
C455 a_2479_44172# a_895_43940# 0.318312f
C456 a_1414_42308# a_2998_44172# 0.447595f
C457 a_2127_44172# a_2675_43914# 0.090298f
C458 a_4007_47204# a_4700_47436# 0.010942f
C459 a_8333_44056# a_8147_43396# 0.011009f
C460 a_17339_46660# a_18579_44172# 0.016577f
C461 a_1823_45246# a_3363_44484# 0.046566f
C462 a_22537_39537# a_22629_37990# 0.490939f
C463 a_n467_45028# VDD 0.385804f
C464 a_n2661_46098# a_n901_46420# 0.054328f
C465 a_11901_46660# a_12156_46660# 0.06121f
C466 a_15368_46634# a_15559_46634# 0.022471f
C467 a_3681_42891# a_n2293_42282# 0.012859f
C468 a_13635_43156# a_13460_43230# 0.234322f
C469 a_22959_46660# a_22959_46124# 0.026152f
C470 a_8016_46348# a_8349_46414# 0.232167f
C471 a_n447_43370# VDD 0.204801f
C472 a_20835_44721# a_20980_44850# 0.057222f
C473 a_20679_44626# a_21398_44850# 0.086708f
C474 a_1799_45572# VDD 0.381212f
C475 a_12594_46348# a_13904_45546# 0.077346f
C476 a_11415_45002# a_18479_45785# 0.047896f
C477 a_18189_46348# VDD 0.211855f
C478 a_1414_42308# a_1568_43370# 0.01352f
C479 a_1467_44172# a_1756_43548# 0.100052f
C480 a_19787_47423# a_19594_46812# 0.108653f
C481 a_n3690_39616# VDD 0.358567f
C482 a_7754_38470# a_8530_39574# 0.143675f
C483 a_17478_45572# VDD 0.411207f
C484 a_10807_43548# a_10991_42826# 0.01427f
C485 a_2680_45002# a_3065_45002# 0.13328f
C486 a_2382_45260# a_3429_45260# 0.011518f
C487 a_10150_46912# a_10554_47026# 0.051162f
C488 a_7411_46660# a_7832_46660# 0.086708f
C489 a_8492_46660# a_6755_46942# 0.024647f
C490 a_9863_46634# a_10249_46116# 0.027588f
C491 a_10428_46928# a_10623_46897# 0.21686f
C492 a_15743_43084# a_19339_43156# 0.128224f
C493 a_n452_44636# VDD 0.112149f
C494 a_19466_46812# a_18819_46122# 0.02948f
C495 a_20935_43940# VDD 0.184334f
C496 a_12465_44636# CLK 0.795478f
C497 a_2747_46873# VDD 0.626468f
C498 a_22223_47212# EN_OFFSET_CAL 0.011048f
C499 a_n699_43396# a_2998_44172# 0.127437f
C500 a_n967_45348# a_n1557_42282# 0.092498f
C501 a_18597_46090# a_21005_45260# 0.034207f
C502 a_n1641_43230# VDD 0.203991f
C503 a_20202_43084# VDD 0.987622f
C504 a_15493_43940# a_15781_43660# 0.049304f
C505 C3_P_btm VDD 0.26836f
C506 a_12891_46348# a_11735_46660# 0.034334f
C507 C2_N_btm C4_N_btm 7.72909f
C508 C1_N_btm C5_N_btm 0.127408f
C509 C0_N_btm C6_N_btm 0.139059f
C510 C0_dummy_N_btm C7_N_btm 0.119061f
C511 a_5837_45028# VDD 0.191549f
C512 a_15743_43084# a_22591_43396# 0.016556f
C513 a_n2661_46098# a_n1736_46482# 0.024986f
C514 a_n809_44244# VDD 0.47719f
C515 a_8016_46348# a_8034_45724# 0.254614f
C516 a_14955_43396# VDD 0.401358f
C517 a_5267_42460# a_5755_42308# 0.055455f
C518 a_2127_44172# a_895_43940# 0.132679f
C519 a_1414_42308# a_2889_44172# 0.128883f
C520 a_12469_46902# VDD 0.203316f
C521 a_18479_47436# a_19279_43940# 0.017993f
C522 a_18597_46090# a_20835_44721# 0.012854f
C523 a_14383_46116# VDD 0.132317f
C524 a_7754_38968# VDD 0.041093f
C525 a_5691_45260# a_5837_45028# 0.171361f
C526 a_21513_45002# a_11827_44484# 0.010541f
C527 a_n2661_46098# a_n1641_46494# 0.035694f
C528 a_11813_46116# a_12156_46660# 0.157972f
C529 a_16795_42852# a_17303_42282# 0.010298f
C530 a_n1352_43396# VDD 0.288329f
C531 a_20640_44752# a_21398_44850# 0.056391f
C532 a_16922_45042# a_20974_43370# 0.077191f
C533 a_12594_46348# a_13527_45546# 0.100424f
C534 a_8199_44636# a_10907_45822# 0.081841f
C535 a_6755_46942# a_14537_43396# 0.120241f
C536 a_n2293_42282# VDD 0.464485f
C537 a_19332_42282# a_19647_42308# 0.084365f
C538 a_1467_44172# a_1568_43370# 0.055004f
C539 a_9028_43914# a_9420_43940# 0.016359f
C540 a_17715_44484# VDD 0.526119f
C541 a_742_44458# a_1847_42826# 0.372436f
C542 a_13904_45546# a_14033_45822# 0.062574f
C543 a_18479_47436# a_20916_46384# 0.014237f
C544 a_19386_47436# a_19594_46812# 0.069651f
C545 a_19787_47423# a_19321_45002# 0.029499f
C546 a_15861_45028# VDD 0.690795f
C547 a_8791_43396# a_9396_43370# 0.011032f
C548 a_10807_43548# a_10796_42968# 0.030352f
C549 a_2382_45260# a_3065_45002# 0.632538f
C550 a_10428_46928# a_10467_46802# 0.820079f
C551 a_8667_46634# a_6755_46942# 0.011524f
C552 a_19594_46812# a_19551_46910# 0.07027f
C553 a_n1352_44484# VDD 0.276725f
C554 a_20623_43914# VDD 0.258478f
C555 a_14537_43396# a_15037_43940# 0.018234f
C556 a_19335_46494# a_19443_46116# 0.057222f
C557 a_n1423_42826# VDD 0.211036f
C558 a_22365_46825# VDD 0.193587f
C559 a_17339_46660# a_11827_44484# 0.031147f
C560 a_9885_42558# VDD 0.18767f
C561 a_2112_39137# VDAC_Pi 0.01062f
C562 a_15493_43940# a_15681_43442# 0.03571f
C563 a_3775_45552# VDD 0.089667f
C564 C4_P_btm VDD 0.265463f
C565 a_n746_45260# a_167_45260# 0.234425f
C566 C0_dummy_N_btm C6_N_btm 0.1194f
C567 C2_N_btm C3_N_btm 5.99608f
C568 C0_N_btm C5_N_btm 0.138093f
C569 C1_N_btm C4_N_btm 0.128167f
C570 a_5093_45028# VDD 0.168437f
C571 a_19466_46812# a_11415_45002# 0.037852f
C572 a_12891_46348# a_12839_46116# 0.038804f
C573 a_12895_43230# a_13003_42852# 0.057222f
C574 a_n1549_44318# VDD 0.200608f
C575 a_11827_44484# a_18579_44172# 0.045146f
C576 a_9482_43914# a_10949_43914# 0.025292f
C577 a_327_47204# DATA[0] 0.353891f
C578 a_7920_46348# a_8034_45724# 0.032141f
C579 a_15095_43370# VDD 0.169652f
C580 a_5267_42460# a_5421_42558# 0.010303f
C581 a_2127_44172# a_2479_44172# 0.168988f
C582 a_453_43940# a_895_43940# 0.420851f
C583 a_1414_42308# a_2675_43914# 0.305556f
C584 a_11901_46660# VDD 0.57548f
C585 a_7640_43914# a_7499_43940# 0.049504f
C586 a_18597_46090# a_20679_44626# 0.025074f
C587 a_18189_46348# a_18175_45572# 0.018402f
C588 a_22400_42852# RST_Z 0.059672f
C589 a_3785_47178# a_4700_47436# 0.090466f
C590 a_3815_47204# a_4007_47204# 0.224415f
C591 a_9313_45822# a_8270_45546# 0.0271f
C592 a_22527_39145# a_22737_36887# 0.011525f
C593 a_22537_39537# a_22629_38406# 0.198762f
C594 a_8199_44636# a_9801_43940# 0.048015f
C595 a_21513_45002# a_21359_45002# 0.289039f
C596 a_n746_45260# a_n863_45724# 0.664707f
C597 a_n2661_46098# a_n1423_46090# 0.021984f
C598 a_14976_45028# a_15368_46634# 0.097092f
C599 a_11735_46660# a_12156_46660# 0.086708f
C600 a_13113_42826# a_13460_43230# 0.051162f
C601 a_5343_44458# a_6298_44484# 0.128602f
C602 a_18597_46090# a_20528_45572# 0.03478f
C603 a_7920_46348# a_8016_46348# 0.318386f
C604 a_n1177_43370# VDD 0.354704f
C605 a_20640_44752# a_20980_44850# 0.027606f
C606 a_5111_44636# a_9885_43646# 0.010527f
C607 a_17767_44458# a_17973_43940# 0.012863f
C608 a_12594_46348# a_13163_45724# 0.053634f
C609 a_11415_45002# a_16147_45260# 0.058206f
C610 a_8199_44636# a_10210_45822# 0.012124f
C611 a_22959_42860# VDD 0.30747f
C612 a_19332_42282# a_19511_42282# 0.174683f
C613 a_n1761_44111# a_n1557_42282# 0.018977f
C614 a_9028_43914# a_9165_43940# 0.126609f
C615 a_17583_46090# VDD 0.23578f
C616 VDAC_Pi a_6886_37412# 0.259481f
C617 a_19386_47436# a_19321_45002# 0.086877f
C618 a_n4334_39616# VDD 0.385881f
C619 a_10807_43548# a_10835_43094# 0.02952f
C620 a_18494_42460# a_20107_42308# 0.035023f
C621 a_2382_45260# a_2680_45002# 0.023953f
C622 a_7927_46660# a_6755_46942# 0.036549f
C623 a_10150_46912# a_10467_46802# 0.102355f
C624 a_n1177_44458# VDD 0.347966f
C625 a_13249_42308# a_13483_43940# 0.193724f
C626 a_20567_45036# a_20193_45348# 0.037561f
C627 a_11827_44484# a_22223_45036# 0.179208f
C628 a_20365_43914# VDD 0.261299f
C629 a_n699_43396# a_2675_43914# 0.015641f
C630 a_18479_47436# a_21005_45260# 0.015257f
C631 a_19553_46090# a_19443_46116# 0.097745f
C632 a_n1991_42858# VDD 0.575656f
C633 a_7499_43078# a_10723_42308# 0.029878f
C634 a_7227_45028# VDD 0.501104f
C635 EN_VIN_BSTR_P VIN_P 1.41696f
C636 C5_P_btm VDD 0.267489f
C637 a_18597_46090# a_16388_46812# 0.011997f
C638 C1_N_btm C3_N_btm 8.06688f
C639 C0_dummy_N_btm C5_N_btm 0.11375f
C640 C0_N_btm C4_N_btm 0.138331f
C641 a_5009_45028# VDD 0.151712f
C642 a_13113_42826# a_13003_42852# 0.097745f
C643 a_n1331_43914# VDD 0.203823f
C644 a_2124_47436# VDD 0.086403f
C645 SMPL_ON_P VIN_P 0.525401f
C646 a_20193_45348# a_20679_44626# 0.017743f
C647 a_16922_45042# a_20512_43084# 0.055985f
C648 a_9482_43914# a_10729_43914# 0.047853f
C649 a_n785_47204# DATA[0] 0.598846f
C650 a_14205_43396# VDD 0.311811f
C651 a_5267_42460# a_5337_42558# 0.011552f
C652 a_5379_42460# a_4921_42308# 0.033756f
C653 a_1414_42308# a_895_43940# 0.208524f
C654 a_11813_46116# VDD 0.434656f
C655 a_18597_46090# a_20640_44752# 0.027095f
C656 a_18189_46348# a_16147_45260# 0.129202f
C657 a_5066_45546# a_9159_45572# 0.040307f
C658 a_n3690_39616# a_n3690_39392# 0.052468f
C659 a_22400_42852# VDD 0.888056f
C660 a_3785_47178# a_4007_47204# 0.106797f
C661 a_20512_43084# a_15743_43084# 0.761578f
C662 a_17478_45572# a_16147_45260# 0.050291f
C663 a_22527_39145# a_22737_37285# 0.012249f
C664 a_22581_37893# a_22629_37990# 0.333805f
C665 a_22537_39537# CAL_P 0.024815f
C666 VDAC_N EN_VIN_BSTR_N 0.341739f
C667 a_n967_45348# VDD 0.556063f
C668 en_comp RST_Z 4.35406f
C669 a_8746_45002# a_10617_44484# 0.01623f
C670 a_4927_45028# a_5093_45028# 0.143754f
C671 a_5111_44636# a_5837_45028# 0.019542f
C672 a_15595_45028# a_16019_45002# 0.017418f
C673 a_n2661_46098# a_n1991_46122# 0.025798f
C674 a_12545_42858# a_13460_43230# 0.118423f
C675 a_5343_44458# a_5518_44484# 0.054464f
C676 a_n1917_43396# VDD 0.204644f
C677 a_19279_43940# a_18579_44172# 0.372064f
C678 a_12594_46348# a_12791_45546# 0.026771f
C679 a_22223_42860# VDD 0.250812f
C680 a_15682_46116# VDD 1.25004f
C681 a_n863_45724# a_n2293_45010# 0.090522f
C682 a_7754_39964# a_6886_37412# 0.035115f
C683 a_18597_46090# a_19321_45002# 0.024487f
C684 a_18479_47436# a_20843_47204# 0.021416f
C685 a_16680_45572# VDD 0.275078f
C686 a_6547_43396# a_6655_43762# 0.057222f
C687 a_21381_43940# a_15743_43084# 0.02274f
C688 a_2274_45254# a_2680_45002# 0.076507f
C689 a_8145_46902# a_6755_46942# 0.02566f
C690 a_9863_46634# a_10467_46802# 0.043587f
C691 a_10150_46912# a_10428_46928# 0.118759f
C692 a_18783_43370# a_18817_42826# 0.012757f
C693 a_n13_43084# a_133_43172# 0.013377f
C694 a_n1917_44484# VDD 0.186988f
C695 a_18494_42460# a_20193_45348# 0.116597f
C696 a_20269_44172# VDD 0.169009f
C697 a_18985_46122# a_19443_46116# 0.027606f
C698 a_1823_45246# a_4099_45572# 0.047087f
C699 a_n1853_43023# VDD 0.370563f
C700 a_7499_43078# a_10533_42308# 0.225871f
C701 a_16763_47508# a_17591_47464# 0.010417f
C702 a_6598_45938# VDD 0.204705f
C703 C6_P_btm VDD 0.210613f
C704 C0_dummy_N_btm C4_N_btm 0.113156f
C705 C1_N_btm C2_N_btm 5.24136f
C706 C0_N_btm C3_N_btm 0.409238f
C707 a_2959_46660# a_3067_47026# 0.057222f
C708 a_2809_45028# VDD 0.189682f
C709 a_3065_45002# a_n699_43396# 0.020711f
C710 a_16388_46812# a_18285_46348# 0.028532f
C711 a_12545_42858# a_13003_42852# 0.027606f
C712 a_n1899_43946# VDD 0.475205f
C713 a_1431_47204# VDD 0.423871f
C714 a_20193_45348# a_20640_44752# 0.017592f
C715 a_9482_43914# a_10405_44172# 0.01085f
C716 a_8975_43940# a_10617_44484# 0.025058f
C717 a_n23_47502# DATA[0] 0.022435f
C718 a_8953_45546# a_5066_45546# 0.191859f
C719 a_20075_46420# a_20708_46348# 0.017547f
C720 a_14358_43442# VDD 0.170277f
C721 a_5267_42460# a_4921_42308# 0.04229f
C722 a_1467_44172# a_895_43940# 0.017277f
C723 a_1414_42308# a_2479_44172# 0.110442f
C724 a_11735_46660# VDD 0.407307f
C725 a_n699_43396# a_458_43396# 0.064001f
C726 a_742_44458# a_1756_43548# 0.152145f
C727 a_18479_47436# a_20679_44626# 0.018117f
C728 a_17715_44484# a_16147_45260# 0.020415f
C729 a_3785_47178# a_3815_47204# 0.270823f
C730 a_15861_45028# a_16147_45260# 0.146279f
C731 a_17478_45572# a_17786_45822# 0.017351f
C732 VDAC_P EN_VIN_BSTR_P 0.340512f
C733 en_comp VDD 4.30454f
C734 a_4927_45028# a_5009_45028# 0.096132f
C735 a_5111_44636# a_5093_45028# 0.021262f
C736 a_14537_43396# a_16751_45260# 0.011362f
C737 a_n2661_46098# a_n1853_46287# 0.019613f
C738 a_6755_46942# a_13059_46348# 0.239671f
C739 a_10617_44484# VDD 0.141193f
C740 a_12545_42858# a_13635_43156# 0.041762f
C741 a_13113_42826# a_12895_43230# 0.209641f
C742 a_n1699_43638# VDD 0.210236f
C743 a_8199_44636# a_8697_45822# 0.067739f
C744 a_6755_46942# a_13556_45296# 0.103107f
C745 a_19321_45002# a_20193_45348# 0.489018f
C746 a_22165_42308# VDD 0.336187f
C747 a_18479_47436# a_19594_46812# 0.108004f
C748 a_16855_45546# VDD 0.339227f
C749 a_6547_43396# a_6452_43396# 0.049827f
C750 a_6765_43638# a_6655_43762# 0.097745f
C751 a_18494_42460# a_19647_42308# 0.030348f
C752 a_2274_45254# a_2382_45260# 0.130215f
C753 a_9863_46634# a_10428_46928# 0.042509f
C754 a_7577_46660# a_6755_46942# 0.035922f
C755 a_n1699_44726# VDD 0.198612f
C756 a_19862_44208# VDD 0.588967f
C757 a_n699_43396# a_2479_44172# 0.063139f
C758 a_n2157_42858# VDD 0.424058f
C759 a_16763_47508# a_16588_47582# 0.233657f
C760 a_9803_42558# VDD 0.253745f
C761 a_n2302_38778# a_n2302_37984# 0.052227f
C762 a_6667_45809# VDD 0.195842f
C763 a_3177_46902# a_3067_47026# 0.097745f
C764 a_3699_46634# a_3524_46660# 0.233657f
C765 a_2959_46660# a_2864_46660# 0.049827f
C766 C7_P_btm VDD 0.121904f
C767 C0_dummy_N_btm C3_N_btm 0.087354f
C768 C0_N_btm C2_N_btm 0.827449f
C769 a_n1761_44111# VDD 0.620042f
C770 a_1239_47204# VDD 0.278979f
C771 a_11827_44484# a_19279_43940# 0.078733f
C772 a_20193_45348# a_20362_44736# 0.013057f
C773 a_9482_43914# a_9672_43914# 0.122568f
C774 a_10057_43914# a_10617_44484# 0.033364f
C775 a_20075_46420# a_19900_46494# 0.233657f
C776 a_14579_43548# VDD 0.278225f
C777 a_n699_43396# a_n229_43646# 0.043893f
C778 a_742_44458# a_1568_43370# 0.525694f
C779 a_1115_44172# a_895_43940# 0.029554f
C780 a_1414_42308# a_2127_44172# 0.091064f
C781 a_11186_47026# VDD 0.077608f
C782 a_18479_47436# a_20640_44752# 0.018112f
C783 a_3381_47502# a_3815_47204# 0.021997f
C784 a_12839_46116# VDD 0.347766f
C785 a_10586_45546# CLK 0.125859f
C786 a_7754_39300# VDD 0.048307f
C787 a_22527_39145# a_22629_37990# 0.172129f
C788 a_22537_40625# a_22737_36887# 0.011861f
C789 a_22589_40055# a_22725_37990# 0.016815f
C790 a_22581_37893# a_22629_38406# 0.236891f
C791 a_15415_45028# a_15595_45028# 0.185422f
C792 a_15009_46634# a_14976_45028# 0.071873f
C793 a_n2661_46098# a_n2157_46122# 0.227082f
C794 a_15743_43084# a_15597_42852# 0.055955f
C795 a_12379_42858# a_13460_43230# 0.102325f
C796 a_12545_42858# a_12895_43230# 0.215953f
C797 a_18597_46090# a_20623_45572# 0.046479f
C798 a_n2267_43396# VDD 0.570924f
C799 a_491_47026# VDD 0.132552f
C800 a_12465_44636# a_14539_43914# 0.054102f
C801 a_12594_46348# a_12427_45724# 0.040872f
C802 a_6755_46942# a_9482_43914# 0.01168f
C803 a_21671_42860# VDD 0.229963f
C804 a_14840_46494# VDD 0.275785f
C805 a_n863_45724# a_n2661_45010# 0.345234f
C806 a_18479_47436# a_19321_45002# 0.262984f
C807 a_16115_45572# VDD 0.194492f
C808 a_6197_43396# a_6655_43762# 0.027317f
C809 a_20193_45348# a_17303_42282# 0.013391f
C810 a_18494_42460# a_19511_42282# 0.047119f
C811 a_13059_46348# a_13565_43940# 0.011241f
C812 a_9863_46634# a_10150_46912# 0.233657f
C813 a_7715_46873# a_6755_46942# 0.089466f
C814 a_7411_46660# a_6969_46634# 0.033891f
C815 a_n2267_44484# VDD 0.289888f
C816 a_19778_44110# a_20193_45348# 0.020562f
C817 a_19478_44306# VDD 0.127794f
C818 a_n2472_42826# VDD 0.229608f
C819 a_7499_43078# a_9885_42558# 0.020607f
C820 a_9223_42460# VDD 0.205797f
C821 a_17973_43940# a_17499_43370# 0.018568f
C822 a_6511_45714# VDD 0.405279f
C823 a_2609_46660# a_3067_47026# 0.027317f
C824 a_n1550_35448# VIN_P 0.37444f
C825 C8_P_btm VDD 0.19922f
C826 C0_dummy_N_btm C2_N_btm 7.14548f
C827 C0_N_btm C1_N_btm 11.2332f
C828 a_2382_45260# a_n699_43396# 0.075387f
C829 a_7927_46660# a_8349_46414# 0.01072f
C830 a_12281_43396# a_12563_42308# 0.173003f
C831 a_n2065_43946# VDD 0.4213f
C832 a_1209_47178# VDD 0.38145f
C833 a_9482_43914# a_9028_43914# 0.092045f
C834 a_10440_44484# a_10617_44484# 0.134298f
C835 a_n746_45260# DATA[0] 0.03466f
C836 a_8199_44636# a_5066_45546# 0.178583f
C837 a_13667_43396# VDD 0.402378f
C838 a_1414_42308# a_453_43940# 0.248504f
C839 a_644_44056# a_895_43940# 0.106452f
C840 a_10768_47026# VDD 0.132317f
C841 a_380_45546# a_603_45572# 0.011458f
C842 a_22589_40055# a_22629_37990# 0.234448f
C843 a_22581_37893# CAL_P 0.026818f
C844 a_9049_44484# a_9159_44484# 0.031707f
C845 a_12379_42858# a_13635_43156# 0.043475f
C846 a_12545_42858# a_13113_42826# 0.178024f
C847 a_18597_46090# a_20841_45814# 0.024341f
C848 a_11415_45002# a_22223_46124# 0.011454f
C849 a_n2129_43609# VDD 0.400674f
C850 a_288_46660# VDD 0.079457f
C851 a_14539_43914# a_15682_43940# 0.161926f
C852 a_12594_46348# a_11962_45724# 0.177228f
C853 a_12005_46116# a_12427_45724# 0.01091f
C854 a_19321_45002# a_19113_45348# 0.147788f
C855 a_21195_42852# VDD 0.285496f
C856 a_n967_45348# a_n961_42308# 0.174237f
C857 a_15015_46420# VDD 0.337162f
C858 a_10210_45822# a_10907_45822# 0.013775f
C859 a_7754_38636# a_7754_38470# 0.296258f
C860 VDAC_Pi a_3726_37500# 1.17174f
C861 a_n2302_40160# VDD 0.428934f
C862 a_16333_45814# VDD 0.201203f
C863 a_6197_43396# a_6452_43396# 0.06121f
C864 a_7411_46660# a_6755_46942# 0.265786f
C865 a_n2129_44697# VDD 1.4165f
C866 a_21101_45002# a_21359_45002# 0.22264f
C867 a_n2293_42282# COMP_P 0.026882f
C868 a_18479_47436# a_19778_44110# 0.038618f
C869 a_n2840_42826# VDD 0.302305f
C870 a_8791_42308# VDD 0.226318f
C871 a_17737_43940# a_17499_43370# 0.013048f
C872 a_104_43370# a_458_43396# 0.07022f
C873 a_6472_45840# VDD 0.257073f
C874 a_2609_46660# a_2864_46660# 0.055869f
C875 a_3177_46902# a_3524_46660# 0.051162f
C876 a_n2002_35448# VIN_P 0.029412f
C877 C9_P_btm VDD 0.345685f
C878 C0_dummy_N_btm C1_N_btm 1.24905f
C879 a_14537_43396# a_11827_44484# 0.076354f
C880 a_16388_46812# a_17339_46660# 0.24887f
C881 a_12891_46348# a_12638_46436# 0.13727f
C882 a_12895_43230# a_12991_43230# 0.013793f
C883 a_n2472_43914# VDD 0.236691f
C884 a_327_47204# VDD 0.367528f
C885 a_19553_46090# a_19900_46494# 0.051162f
C886 a_10695_43548# VDD 0.201247f
C887 a_3823_42558# a_3905_42558# 0.171361f
C888 a_1467_44172# a_453_43940# 0.05905f
C889 a_380_45546# a_509_45572# 0.010132f
C890 a_1848_45724# a_1609_45822# 0.042695f
C891 a_n4334_39616# a_n4334_39392# 0.052468f
C892 a_18707_42852# VDD 0.132317f
C893 a_22581_37893# a_22944_39857# 0.011943f
C894 a_22589_40599# a_22737_37285# 0.010048f
C895 a_22527_39145# a_22629_38406# 0.123152f
C896 a_22537_40625# a_22725_37990# 0.010408f
C897 a_22589_40055# a_22725_38406# 0.010302f
C898 a_22889_38993# a_22537_39537# 0.033924f
C899 a_n1761_44111# a_n473_42460# 0.110251f
C900 a_n745_45366# VDD 0.20887f
C901 a_4558_45348# a_5009_45028# 0.013349f
C902 a_n2661_46098# a_n2472_46090# 0.094589f
C903 a_12379_42858# a_12895_43230# 0.109156f
C904 a_n699_43396# a_4743_44484# 0.235328f
C905 a_18597_46090# a_20273_45572# 0.048762f
C906 a_n2433_43396# VDD 0.416276f
C907 a_20766_44850# a_19279_43940# 0.021466f
C908 a_1983_46706# VDD 0.119964f
C909 a_14539_43914# a_14955_43940# 0.064683f
C910 a_626_44172# a_648_43396# 0.04847f
C911 a_16375_45002# a_18051_46116# 0.038793f
C912 a_21356_42826# VDD 0.225688f
C913 a_18057_42282# a_18310_42308# 0.011913f
C914 a_n967_45348# a_n1329_42308# 0.033651f
C915 a_14275_46494# VDD 0.196859f
C916 a_7754_39964# a_3726_37500# 0.030605f
C917 a_15765_45572# VDD 0.249471f
C918 a_19319_43548# a_19268_43646# 0.17076f
C919 a_6293_42852# a_6452_43396# 0.157972f
C920 a_7287_43370# a_7112_43396# 0.234322f
C921 a_18525_43370# a_18083_42858# 0.016073f
C922 a_n1641_43230# a_n1533_42852# 0.057222f
C923 a_n2433_44484# VDD 0.40658f
C924 a_19328_44172# VDD 0.263964f
C925 a_n699_43396# a_1414_42308# 0.104607f
C926 a_742_44458# a_895_43940# 0.025021f
C927 a_22959_47212# VDD 0.245964f
C928 a_19335_46494# a_19431_46494# 0.013793f
C929 a_5066_45546# a_8034_45724# 0.242476f
C930 a_11551_42558# a_11633_42558# 0.171361f
C931 a_10057_43914# a_10695_43548# 0.148476f
C932 a_8199_44636# a_9482_43914# 0.276776f
C933 a_16241_47178# a_16588_47582# 0.051162f
C934 a_8685_42308# VDD 0.286875f
C935 a_6194_45824# VDD 0.274689f
C936 a_21363_45546# a_21513_45002# 0.06363f
C937 a_5807_45002# a_6755_46942# 1.47519f
C938 a_2609_46660# a_3524_46660# 0.118759f
C939 a_2443_46660# a_2864_46660# 0.090164f
C940 C10_P_btm VDD 2.40001f
C941 C0_dummy_N_btm C0_N_btm 7.97415f
C942 a_19268_43646# a_19095_43396# 0.032587f
C943 a_12895_43230# a_12800_43218# 0.049827f
C944 a_n2840_43914# VDD 0.304745f
C945 a_n785_47204# VDD 0.452945f
C946 a_11827_44484# a_20679_44626# 0.030022f
C947 a_21101_45002# a_20766_44850# 0.01337f
C948 a_n452_47436# DATA[0] 0.039965f
C949 a_18985_46122# a_19900_46494# 0.118759f
C950 a_8016_46348# a_5066_45546# 0.054471f
C951 a_9803_43646# VDD 0.261557f
C952 a_1755_42282# a_6481_42558# 0.012532f
C953 a_1467_44172# a_1414_42308# 0.335735f
C954 a_1115_44172# a_453_43940# 0.150214f
C955 a_1138_42852# a_n2661_45010# 0.017849f
C956 a_n2302_39866# a_n2216_39866# 0.011479f
C957 a_14539_43914# a_17333_42852# 0.072085f
C958 a_7754_39632# RST_Z 0.030938f
C959 a_22581_37893# a_22848_39857# 0.01318f
C960 a_22537_40625# a_22629_37990# 0.130478f
C961 a_22589_40055# a_22629_38406# 0.1922f
C962 a_22613_38993# a_22537_39537# 0.049665f
C963 a_12293_43646# a_12281_43396# 0.01129f
C964 a_12891_46348# a_13351_46090# 0.019821f
C965 a_n2661_46098# a_n2840_46090# 0.170439f
C966 a_383_46660# a_805_46414# 0.01072f
C967 a_12379_42858# a_13113_42826# 0.06628f
C968 a_12089_42308# a_12545_42858# 0.261463f
C969 a_18479_47436# a_20841_45814# 0.011134f
C970 a_18597_46090# a_20107_45572# 0.069963f
C971 a_22365_46825# a_22223_46124# 0.011912f
C972 a_22400_42852# COMP_P 0.595635f
C973 a_20835_44721# a_19279_43940# 0.036128f
C974 a_12465_44636# a_13720_44458# 0.019702f
C975 a_20922_43172# VDD 0.192467f
C976 a_18727_42674# a_18214_42558# 0.035505f
C977 a_18057_42282# a_18220_42308# 0.01135f
C978 a_18907_42674# a_19332_42282# 0.017308f
C979 a_14493_46090# VDD 0.203567f
C980 a_n2472_45546# a_n2472_45002# 0.026152f
C981 a_n4334_40480# VDD 0.390668f
C982 a_2905_45572# a_3524_46660# 0.011982f
C983 a_15903_45785# VDD 0.291109f
C984 a_19319_43548# a_15743_43084# 0.035611f
C985 a_6031_43396# a_6452_43396# 0.086708f
C986 a_n1423_42826# a_n1533_42852# 0.097745f
C987 a_5147_45002# a_5708_44484# 0.055267f
C988 a_18494_42460# a_11827_44484# 0.031498f
C989 a_18911_45144# a_19113_45348# 0.054737f
C990 a_21005_45260# a_21101_45002# 0.419086f
C991 a_18451_43940# VDD 0.172318f
C992 a_n699_43396# a_1467_44172# 0.030347f
C993 a_742_44458# a_2479_44172# 0.019563f
C994 SMPL_ON_N RST_Z 2.43362f
C995 a_19335_46494# a_19240_46482# 0.049827f
C996 a_7499_43078# a_9803_42558# 0.158876f
C997 a_8325_42308# VDD 0.313956f
C998 a_15673_47210# a_16588_47582# 0.125324f
C999 a_n2946_38778# a_n2946_37984# 0.052227f
C1000 a_15682_43940# a_16759_43396# 0.013707f
C1001 a_5907_45546# VDD 0.390381f
C1002 a_5807_45002# a_10249_46116# 0.041839f
C1003 a_3177_46902# a_2959_46660# 0.209641f
C1004 a_2609_46660# a_3699_46634# 0.042415f
C1005 a_2443_46660# a_3524_46660# 0.102325f
C1006 a_21753_35474# VDD 0.525301f
C1007 a_15743_43084# a_19095_43396# 0.012939f
C1008 a_n23_47502# VDD 0.152616f
C1009 a_11827_44484# a_20640_44752# 0.016882f
C1010 a_19778_44110# a_18579_44172# 0.268475f
C1011 a_5883_43914# a_9159_44484# 0.049132f
C1012 a_n815_47178# DATA[0] 0.068508f
C1013 a_18985_46122# a_20075_46420# 0.042415f
C1014 a_18819_46122# a_19900_46494# 0.102355f
C1015 a_19553_46090# a_19335_46494# 0.209641f
C1016 a_7920_46348# a_5066_45546# 0.04093f
C1017 a_8270_45546# a_8746_45002# 0.017581f
C1018 a_3318_42354# a_3581_42558# 0.011552f
C1019 a_5267_42460# a_5379_42460# 0.156424f
C1020 a_644_44056# a_453_43940# 0.077973f
C1021 a_1115_44172# a_1414_42308# 0.134389f
C1022 a_n356_45724# a_n23_45546# 0.360492f
C1023 a_3160_47472# a_3381_47502# 0.099936f
C1024 a_2905_45572# a_3785_47178# 0.013619f
C1025 a_14180_46482# VDD 0.077608f
C1026 a_742_44458# a_1793_42852# 0.010622f
C1027 a_7754_39632# VDD 0.205733f
C1028 a_22589_40599# a_22629_37990# 0.021352f
C1029 a_22581_37893# a_22537_39537# 1.00904f
C1030 a_22613_38993# a_22889_38993# 0.237336f
C1031 a_14537_43396# a_14797_45144# 0.082443f
C1032 a_12891_46348# a_12594_46348# 0.088156f
C1033 a_6755_46942# a_14513_46634# 0.036712f
C1034 a_12379_42858# a_12545_42858# 0.810394f
C1035 a_18479_47436# a_20273_45572# 0.028755f
C1036 a_n2840_43370# VDD 0.246858f
C1037 a_20679_44626# a_19279_43940# 0.279785f
C1038 a_20835_44721# a_20766_44850# 0.209641f
C1039 a_948_46660# VDD 0.278482f
C1040 a_9482_43914# a_9396_43370# 0.011522f
C1041 a_19321_45002# a_11827_44484# 0.037739f
C1042 a_12465_44636# a_13076_44458# 0.01224f
C1043 a_19987_42826# VDD 0.588466f
C1044 a_18057_42282# a_18214_42558# 0.18824f
C1045 en_comp COMP_P 1.91962f
C1046 a_15493_43940# a_22959_43948# 0.182001f
C1047 a_13925_46122# VDD 0.251868f
C1048 a_12465_44636# a_12891_46348# 0.033919f
C1049 a_15599_45572# VDD 0.390565f
C1050 a_6765_43638# a_7112_43396# 0.051162f
C1051 a_18494_42460# a_18214_42558# 0.012583f
C1052 a_8667_46634# a_8492_46660# 0.233657f
C1053 a_n1991_42858# a_n1533_42852# 0.034619f
C1054 a_18326_43940# VDD 0.129408f
C1055 a_12465_44636# SINGLE_ENDED 0.067716f
C1056 SMPL_ON_N VDD 0.497737f
C1057 a_17957_46116# a_18051_46116# 0.062574f
C1058 a_22959_43396# VDD 0.303237f
C1059 a_7499_43078# a_9223_42460# 0.013802f
C1060 a_8016_46348# a_9482_43914# 0.293982f
C1061 a_13059_46348# a_11827_44484# 0.495367f
C1062 a_7227_45028# a_7230_45938# 0.170618f
C1063 a_8270_45546# a_8975_43940# 0.207334f
C1064 a_16241_47178# a_16023_47582# 0.209641f
C1065 a_15673_47210# a_16763_47508# 0.042509f
C1066 a_2112_39137# a_2113_38308# 0.478223f
C1067 a_n447_43370# a_n229_43646# 0.08213f
C1068 a_5263_45724# VDD 0.202719f
C1069 C7_P_btm C7_N_btm 0.028901f
C1070 C6_P_btm C6_N_btm 0.019861f
C1071 C5_P_btm C5_N_btm 0.03705f
C1072 C4_P_btm C4_N_btm 0.02642f
C1073 C3_P_btm C3_N_btm 2.90911f
C1074 C2_P_btm C2_N_btm 0.026726f
C1075 C1_P_btm C1_N_btm 0.065833f
C1076 C0_P_btm C0_N_btm 0.044249f
C1077 C0_dummy_P_btm C0_dummy_N_btm 0.033338f
C1078 a_19998_34978# VDD 0.319197f
C1079 a_2443_46660# a_3699_46634# 0.043475f
C1080 a_2609_46660# a_2959_46660# 0.216095f
C1081 a_n746_45260# a_376_46348# 0.010981f
C1082 a_18783_43370# a_19095_43396# 0.038241f
C1083 a_13556_45296# a_11827_44484# 0.05613f
C1084 a_14976_45028# a_11415_45002# 0.039578f
C1085 a_n1991_42858# a_n1736_42282# 0.0101f
C1086 a_12545_42858# a_12800_43218# 0.05936f
C1087 a_22959_44484# VDD 0.303517f
C1088 a_21359_45002# a_20640_44752# 0.013689f
C1089 a_18494_42460# a_19279_43940# 0.137363f
C1090 a_6419_46155# a_5066_45546# 0.038923f
C1091 a_18819_46122# a_20075_46420# 0.043567f
C1092 a_18985_46122# a_19335_46494# 0.210876f
C1093 a_3318_42354# a_3497_42558# 0.010303f
C1094 a_1755_42282# a_6171_42473# 0.065035f
C1095 a_175_44278# a_453_43940# 0.112594f
C1096 a_1115_44172# a_1467_44172# 0.115277f
C1097 a_8270_45546# VDD 1.26092f
C1098 a_2905_45572# a_3381_47502# 0.208262f
C1099 a_14539_43914# a_17701_42308# 0.039977f
C1100 a_n863_45724# a_2304_45348# 0.091195f
C1101 a_2747_46873# a_2864_46660# 0.174836f
C1102 a_22537_40625# a_22629_38406# 0.066321f
C1103 a_22581_37893# a_22889_38993# 0.112329f
C1104 a_14358_43442# a_14621_43646# 0.011552f
C1105 a_5691_45260# a_5837_45348# 0.013377f
C1106 a_14180_45002# a_14797_45144# 0.070624f
C1107 a_6755_46942# a_14180_46812# 0.063843f
C1108 a_13607_46688# a_14084_46812# 0.014875f
C1109 a_12379_42858# a_12089_42308# 0.16885f
C1110 a_2779_44458# a_n699_43396# 0.025176f
C1111 a_8953_45546# a_8952_43230# 0.01883f
C1112 a_18479_47436# a_20107_45572# 0.025968f
C1113 a_5204_45822# a_5497_46414# 0.099282f
C1114 a_19615_44636# a_18579_44172# 0.158449f
C1115 a_20679_44626# a_20766_44850# 0.052825f
C1116 a_20640_44752# a_19279_43940# 0.22152f
C1117 a_1123_46634# VDD 0.469393f
C1118 a_5111_44636# a_9803_43646# 0.118936f
C1119 a_12465_44636# a_12883_44458# 0.017889f
C1120 a_19164_43230# VDD 0.278643f
C1121 a_18727_42674# a_18907_42674# 0.185422f
C1122 a_13759_46122# VDD 0.399995f
C1123 a_22485_38105# RST_Z 0.036748f
C1124 a_6197_43396# a_7112_43396# 0.118423f
C1125 a_2479_44172# a_n2293_42282# 0.059476f
C1126 a_18494_42460# a_19332_42282# 0.040916f
C1127 a_15743_43084# a_15567_42826# 0.215954f
C1128 a_n2840_44458# VDD 0.247948f
C1129 a_19778_44110# a_11827_44484# 0.029054f
C1130 a_20567_45036# a_21005_45260# 0.015494f
C1131 a_18079_43940# VDD 0.162408f
C1132 a_n2293_42282# a_n2104_42282# 0.058363f
C1133 a_21811_47423# SINGLE_ENDED 0.215228f
C1134 a_22731_47423# VDD 0.196667f
C1135 a_12465_44636# START 0.065727f
C1136 a_18189_46348# a_18051_46116# 0.045453f
C1137 a_18985_46122# a_19240_46482# 0.05936f
C1138 a_11323_42473# a_11551_42558# 0.062483f
C1139 a_19321_45002# a_19279_43940# 0.019898f
C1140 a_15673_47210# a_16023_47582# 0.228897f
C1141 a_15507_47210# a_16588_47582# 0.102325f
C1142 a_4099_45572# VDD 0.296272f
C1143 a_20623_45572# a_20719_45572# 0.013793f
C1144 a_2609_46660# a_3177_46902# 0.17072f
C1145 a_2443_46660# a_2959_46660# 0.110816f
C1146 a_19250_34978# VDD 0.323729f
C1147 a_9482_43914# a_11827_44484# 0.031913f
C1148 a_7715_46873# a_7920_46348# 0.080253f
C1149 a_10922_42852# a_11136_42852# 0.097745f
C1150 a_12089_42308# a_12800_43218# 0.15794f
C1151 a_n746_45260# VDD 1.41433f
C1152 a_11827_44484# a_20159_44458# 0.012941f
C1153 a_7499_43078# a_10695_43548# 0.124597f
C1154 a_18819_46122# a_19335_46494# 0.108964f
C1155 a_6165_46155# a_5066_45546# 0.041118f
C1156 a_18985_46122# a_19553_46090# 0.16939f
C1157 a_n699_43396# a_104_43370# 0.21575f
C1158 a_6755_46942# CLK 0.031541f
C1159 a_10586_45546# a_11962_45724# 0.137051f
C1160 a_12465_44636# a_14673_44172# 0.101564f
C1161 a_n2946_39866# a_n2860_39866# 0.011479f
C1162 a_14539_43914# a_17595_43084# 0.141972f
C1163 a_5907_45546# a_5111_44636# 0.01337f
C1164 a_16115_45572# a_16211_45572# 0.013793f
C1165 a_11415_45002# a_14815_43914# 0.070306f
C1166 a_7754_39964# RST_Z 0.843939f
C1167 VDAC_Pi VDD 0.591846f
C1168 a_22589_40599# a_22629_38406# 0.032572f
C1169 a_22527_39145# a_22537_39537# 0.351623f
C1170 a_22581_37893# a_22613_38993# 0.275268f
C1171 a_14358_43442# a_14537_43646# 0.010303f
C1172 a_n2109_45247# VDD 0.266396f
C1173 a_21363_45546# a_21359_45002# 0.01738f
C1174 a_14180_45002# a_14537_43396# 0.143922f
C1175 a_6755_46942# a_14035_46660# 0.040006f
C1176 a_n13_43084# a_133_42852# 0.171361f
C1177 a_13249_42308# a_13565_43940# 0.048533f
C1178 a_5164_46348# a_5497_46414# 0.203417f
C1179 a_383_46660# VDD 0.198466f
C1180 a_20679_44626# a_20835_44721# 0.105995f
C1181 a_20362_44736# a_19279_43940# 0.039759f
C1182 a_20640_44752# a_20766_44850# 0.17072f
C1183 a_12465_44636# a_12607_44458# 0.186652f
C1184 a_19339_43156# VDD 0.338297f
C1185 a_13351_46090# VDD 0.238036f
C1186 a_14955_43940# a_15301_44260# 0.013377f
C1187 a_22223_43948# a_15493_43940# 0.051823f
C1188 a_11525_45546# a_11778_45572# 0.011913f
C1189 a_22485_38105# VDD 1.31335f
C1190 a_2905_45572# a_3177_46902# 0.014554f
C1191 a_3160_47472# a_2609_46660# 0.018687f
C1192 a_6765_43638# a_6547_43396# 0.209641f
C1193 a_6197_43396# a_7287_43370# 0.041762f
C1194 a_18494_42460# a_18907_42674# 0.11494f
C1195 a_8145_46902# a_8492_46660# 0.051162f
C1196 a_5807_45002# a_17339_46660# 0.02927f
C1197 a_n1641_43230# a_n1545_43230# 0.013793f
C1198 a_17973_43940# VDD 0.265874f
C1199 a_742_44458# a_1414_42308# 0.052151f
C1200 a_22223_47212# VDD 0.236555f
C1201 a_18443_44721# a_18753_44484# 0.013793f
C1202 a_18989_43940# a_18579_44172# 0.035827f
C1203 a_18597_46090# a_16922_45042# 0.028931f
C1204 a_18819_46122# a_19240_46482# 0.089677f
C1205 a_22591_43396# VDD 0.280354f
C1206 a_20731_47026# VDD 0.132317f
C1207 a_2382_45260# a_n2293_42282# 0.080755f
C1208 a_6598_45938# a_6812_45938# 0.097745f
C1209 a_6667_45809# a_7230_45938# 0.049827f
C1210 a_15507_47210# a_16763_47508# 0.043475f
C1211 a_3175_45822# VDD 0.193907f
C1212 a_18597_46090# a_15743_43084# 0.023066f
C1213 C0_P_btm C0_dummy_P_btm 7.97415f
C1214 a_2443_46660# a_3177_46902# 0.053479f
C1215 a_22591_44484# VDD 0.223346f
C1216 a_10991_42826# a_11136_42852# 0.057222f
C1217 a_12379_42858# a_12800_43218# 0.089677f
C1218 a_19778_44110# a_19279_43940# 0.020911f
C1219 SMPL_ON_P CLK_DATA 0.200962f
C1220 a_18819_46122# a_19553_46090# 0.052547f
C1221 a_5497_46414# a_5066_45546# 0.05403f
C1222 a_10249_46116# CLK 0.063525f
C1223 a_644_44056# a_1115_44172# 0.013441f
C1224 a_13059_46348# a_14797_45144# 0.066603f
C1225 a_10586_45546# a_11652_45724# 0.046802f
C1226 a_2905_45572# a_3160_47472# 0.54473f
C1227 a_14539_43914# a_16795_42852# 0.037061f
C1228 a_310_45028# a_375_42282# 0.078376f
C1229 a_7754_39964# VDD 0.848281f
C1230 CAL_N a_22629_38406# 0.204616f
C1231 a_22589_40055# a_22537_39537# 0.035975f
C1232 a_22527_39145# a_22889_38993# 0.010853f
C1233 a_n2293_45010# VDD 1.885f
C1234 a_4927_45028# a_5365_45348# 0.013015f
C1235 a_6755_46942# a_13885_46660# 0.078788f
C1236 a_n2497_47436# a_n863_45724# 0.337007f
C1237 a_742_44458# a_n699_43396# 0.047576f
C1238 a_3877_44458# a_4099_45572# 0.01632f
C1239 a_5164_46348# a_5204_45822# 0.132894f
C1240 a_20974_43370# VDD 0.550101f
C1241 a_20159_44458# a_19279_43940# 0.06519f
C1242 a_20640_44752# a_20835_44721# 0.20669f
C1243 a_20362_44736# a_20766_44850# 0.051162f
C1244 a_601_46902# VDD 0.204253f
C1245 a_8270_45546# a_5111_44636# 0.035253f
C1246 a_18599_43230# VDD 0.197104f
C1247 a_12594_46348# VDD 1.03351f
C1248 a_12891_46348# a_13483_43940# 0.062818f
C1249 a_11525_45546# a_11688_45572# 0.011381f
C1250 a_2905_45572# a_2609_46660# 0.027251f
C1251 a_3160_47472# a_2443_46660# 0.019074f
C1252 a_15037_45618# VDD 0.08759f
C1253 a_6197_43396# a_6547_43396# 0.216095f
C1254 a_6031_43396# a_7112_43396# 0.101963f
C1255 a_18494_42460# a_18727_42674# 0.031761f
C1256 a_7577_46660# a_8492_46660# 0.118423f
C1257 a_n1641_43230# a_n1736_43218# 0.049827f
C1258 a_16922_45042# a_20193_45348# 0.328274f
C1259 a_17737_43940# VDD 0.285511f
C1260 a_n2293_42282# a_n2472_42282# 0.163758f
C1261 a_949_44458# a_1115_44172# 0.016355f
C1262 a_742_44458# a_1467_44172# 0.018499f
C1263 a_21496_47436# SINGLE_ENDED 0.055146f
C1264 a_12465_44636# VDD 0.773277f
C1265 a_20528_46660# VDD 0.077608f
C1266 a_20193_45348# a_15743_43084# 0.060559f
C1267 a_6511_45714# a_7230_45938# 0.088127f
C1268 a_6667_45809# a_6812_45938# 0.057222f
C1269 a_15673_47210# a_16241_47178# 0.183195f
C1270 a_15507_47210# a_16023_47582# 0.109156f
C1271 a_8515_42308# VDD 0.194691f
C1272 a_n3690_38528# a_n3690_38304# 0.052468f
C1273 a_15682_43940# a_16243_43396# 0.013782f
C1274 C1_P_btm C0_dummy_P_btm 1.24905f
C1275 a_2443_46660# a_2609_46660# 0.579196f
C1276 EN_VIN_BSTR_N VDD 1.19259f
C1277 a_16388_46812# a_16721_46634# 0.222024f
C1278 a_22485_44484# VDD 0.258874f
C1279 a_10796_42968# a_11136_42852# 0.027606f
C1280 a_n452_47436# VDD 0.092189f
C1281 a_5204_45822# a_5066_45546# 0.402457f
C1282 a_18819_46122# a_18985_46122# 0.749955f
C1283 a_n699_43396# a_n447_43370# 0.040315f
C1284 a_10554_47026# CLK 0.014924f
C1285 a_13249_42308# a_13291_42460# 0.068754f
C1286 a_5066_45546# a_8697_45822# 0.033513f
C1287 a_3316_45546# a_3503_45724# 0.024901f
C1288 a_310_45028# a_509_45822# 0.039722f
C1289 a_10586_45546# a_11525_45546# 0.115475f
C1290 a_13059_46348# a_14537_43396# 0.30244f
C1291 a_2952_47436# a_3160_47472# 0.192116f
C1292 a_16877_42852# VDD 0.192454f
C1293 a_2747_46873# a_2959_46660# 0.010672f
C1294 a_22527_39145# a_22613_38993# 0.12129f
C1295 a_22589_40055# a_22889_38993# 0.19183f
C1296 CAL_N CAL_P 5.92093f
C1297 a_n2472_45002# VDD 0.217954f
C1298 a_2680_45002# a_2809_45028# 0.062574f
C1299 a_13556_45296# a_14537_43396# 0.590856f
C1300 a_171_46873# a_376_46348# 0.080253f
C1301 a_11309_47204# a_11387_46155# 0.061891f
C1302 a_16137_43396# a_16877_42852# 0.010276f
C1303 a_11827_44484# a_18989_43940# 0.054716f
C1304 a_8199_44636# a_9127_43156# 0.01079f
C1305 a_5068_46348# a_5204_45822# 0.20685f
C1306 a_20640_44752# a_20679_44626# 0.582607f
C1307 a_33_46660# VDD 0.272723f
C1308 a_13249_42308# a_13460_43230# 0.014543f
C1309 a_11189_46129# a_11525_45546# 0.085926f
C1310 a_19321_45002# a_20567_45036# 0.205038f
C1311 a_5807_45002# a_11827_44484# 0.022597f
C1312 a_18817_42826# VDD 0.204624f
C1313 a_8199_44636# CLK 0.231904f
C1314 a_12005_46116# VDD 0.518463f
C1315 a_21115_43940# a_15493_43940# 0.0516f
C1316 a_n2840_45546# a_n2840_45002# 0.026152f
C1317 a_2905_45572# a_2443_46660# 0.026052f
C1318 a_16588_47582# a_5807_45002# 0.040789f
C1319 a_3754_38802# VDAC_Ni 0.301032f
C1320 a_14033_45822# VDD 0.195067f
C1321 a_6031_43396# a_7287_43370# 0.042271f
C1322 a_6197_43396# a_6765_43638# 0.17072f
C1323 a_18494_42460# a_18057_42282# 0.085802f
C1324 a_9313_45822# a_9569_46155# 0.019679f
C1325 a_7577_46660# a_8667_46634# 0.041879f
C1326 a_8145_46902# a_7927_46660# 0.209641f
C1327 a_19778_44110# a_21005_45260# 0.135527f
C1328 a_15682_43940# VDD 1.22657f
C1329 a_21811_47423# VDD 0.201359f
C1330 a_167_45260# a_2277_45546# 0.214157f
C1331 a_17957_46116# a_16375_45002# 0.017118f
C1332 a_22223_43396# VDD 0.279195f
C1333 a_22000_46634# VDD 0.257047f
C1334 a_167_45260# a_626_44172# 0.04273f
C1335 a_8199_44636# a_10951_45334# 0.237774f
C1336 a_6472_45840# a_7230_45938# 0.05936f
C1337 a_8953_45546# a_8953_45002# 0.023516f
C1338 a_19321_45002# a_20679_44626# 0.023087f
C1339 C2_P_btm C0_dummy_P_btm 7.14548f
C1340 C1_P_btm C0_P_btm 11.2332f
C1341 a_n2497_47436# a_1823_45246# 0.025359f
C1342 a_16751_45260# a_17023_45118# 0.13675f
C1343 a_17609_46634# a_18280_46660# 0.094543f
C1344 a_5257_43370# a_6419_46155# 0.186651f
C1345 a_20512_43084# VDD 0.317257f
C1346 a_n2157_42858# a_n2104_42282# 0.011248f
C1347 a_n815_47178# VDD 0.380339f
C1348 a_5164_46348# a_5066_45546# 0.096188f
C1349 a_11415_45002# a_16375_45002# 0.080382f
C1350 a_8270_45546# a_7499_43078# 0.063428f
C1351 a_10623_46897# CLK 0.016177f
C1352 a_13059_46348# a_14180_45002# 0.073427f
C1353 a_n1099_45572# a_509_45822# 0.026885f
C1354 a_3218_45724# a_3503_45724# 0.099872f
C1355 a_10586_45546# a_11322_45546# 0.220166f
C1356 a_2952_47436# a_2905_45572# 0.318161f
C1357 a_16245_42852# VDD 0.205729f
C1358 a_18579_44172# a_19700_43370# 0.175511f
C1359 a_n863_45724# a_626_44172# 0.097275f
C1360 a_22537_40625# a_22537_39537# 0.604835f
C1361 a_22527_39145# a_22581_37893# 0.076507f
C1362 a_19321_45002# a_19594_46812# 0.267862f
C1363 a_n2661_45010# VDD 0.842431f
C1364 a_2382_45260# a_2809_45028# 0.034331f
C1365 a_9482_43914# a_14537_43396# 0.040878f
C1366 a_5807_45002# a_6419_46155# 0.072498f
C1367 a_11309_47204# a_11133_46155# 0.040357f
C1368 a_12991_46634# a_12816_46660# 0.233657f
C1369 a_16137_43396# a_16245_42852# 0.016079f
C1370 a_10922_42852# a_10341_42308# 0.053077f
C1371 a_8953_45546# a_8037_42858# 0.017317f
C1372 a_5068_46348# a_5164_46348# 0.31819f
C1373 a_21381_43940# VDD 0.344882f
C1374 a_20362_44736# a_20679_44626# 0.102355f
C1375 a_171_46873# VDD 0.539781f
C1376 a_11189_46129# a_11322_45546# 0.05577f
C1377 a_19321_45002# a_18494_42460# 0.084551f
C1378 a_18249_42858# VDD 0.250132f
C1379 a_20935_43940# a_15493_43940# 0.037795f
C1380 a_17339_46660# a_18287_44626# 0.018815f
C1381 a_11322_45546# a_11136_45572# 0.044092f
C1382 a_16763_47508# a_5807_45002# 0.127783f
C1383 a_6031_43396# a_6547_43396# 0.105995f
C1384 a_n143_45144# a_n37_45144# 0.13675f
C1385 a_20202_43084# a_15493_43940# 0.02138f
C1386 a_9313_45822# a_9625_46129# 0.018694f
C1387 a_7411_46660# a_8492_46660# 0.102325f
C1388 a_7577_46660# a_7927_46660# 0.206455f
C1389 a_16137_43396# a_18249_42858# 0.021561f
C1390 a_n1991_42858# a_n1736_43218# 0.064178f
C1391 a_n901_43156# a_n13_43084# 0.014329f
C1392 a_7229_43940# a_7640_43914# 0.177622f
C1393 a_19778_44110# a_20567_45036# 0.044967f
C1394 a_9313_45822# a_9159_45572# 0.051702f
C1395 a_14955_43940# VDD 0.253201f
C1396 a_18989_43940# a_19279_43940# 0.053948f
C1397 a_18287_44626# a_18579_44172# 0.107662f
C1398 a_21177_47436# SINGLE_ENDED 0.057266f
C1399 a_17957_46116# a_18243_46436# 0.010132f
C1400 a_18189_46348# a_16375_45002# 0.165328f
C1401 a_167_45260# a_1609_45822# 0.141505f
C1402 a_21188_46660# VDD 0.284105f
C1403 a_16922_45042# a_21259_43561# 0.108631f
C1404 a_8199_44636# a_10775_45002# 0.064568f
C1405 a_6472_45840# a_6812_45938# 0.027606f
C1406 a_19321_45002# a_20640_44752# 0.034599f
C1407 a_15811_47375# a_15673_47210# 0.281607f
C1408 a_15507_47210# a_16241_47178# 0.06628f
C1409 a_7963_42308# VDD 0.266057f
C1410 a_n1917_43396# a_n1821_43396# 0.013793f
C1411 a_15493_43940# a_14955_43396# 0.013181f
C1412 a_20623_45572# a_20731_45938# 0.057222f
C1413 C3_P_btm C0_dummy_P_btm 0.087354f
C1414 EN_VIN_BSTR_N C10_N_btm 0.320569f
C1415 C2_P_btm C0_P_btm 0.827449f
C1416 a_n2661_46098# a_2443_46660# 0.063999f
C1417 a_n217_35014# VDD 0.296751f
C1418 a_n2497_47436# a_1138_42852# 0.144386f
C1419 a_15811_47375# a_16388_46812# 0.010369f
C1420 a_16751_45260# a_16922_45042# 0.12103f
C1421 SMPL_ON_N COMP_P 2.13156f
C1422 a_17609_46634# a_17639_46660# 0.094289f
C1423 a_5257_43370# a_6165_46155# 0.11382f
C1424 a_10341_42308# a_11554_42852# 0.170124f
C1425 a_n1605_47204# VDD 0.20224f
C1426 a_5518_44484# a_5708_44484# 0.045837f
C1427 a_5068_46348# a_5066_45546# 0.04842f
C1428 a_8270_45546# a_8568_45546# 0.015327f
C1429 a_n699_43396# a_n1177_43370# 0.060973f
C1430 a_10467_46802# CLK 0.028547f
C1431 a_380_45546# a_509_45822# 0.062574f
C1432 a_n863_45724# a_1609_45822# 0.117311f
C1433 a_3218_45724# a_3316_45546# 0.162813f
C1434 a_10586_45546# a_10490_45724# 0.235237f
C1435 a_22589_40055# a_22581_37893# 0.461959f
C1436 a_22589_40599# a_22537_39537# 0.380009f
C1437 a_2747_46873# a_2609_46660# 0.347674f
C1438 a_9313_45822# a_6755_46942# 0.031706f
C1439 a_n2840_45002# VDD 0.289706f
C1440 a_20273_45572# a_21101_45002# 0.014321f
C1441 a_13556_45296# a_13777_45326# 0.101558f
C1442 a_9482_43914# a_14180_45002# 0.022677f
C1443 a_5807_45002# a_6165_46155# 0.039202f
C1444 a_11309_47204# a_11189_46129# 0.03753f
C1445 a_10991_42826# a_10341_42308# 0.035667f
C1446 a_742_44458# a_949_44458# 0.185221f
C1447 a_19741_43940# VDD 0.153579f
C1448 a_20159_44458# a_20679_44626# 0.043567f
C1449 a_20362_44736# a_20640_44752# 0.118759f
C1450 a_n133_46660# VDD 0.483405f
C1451 a_7640_43914# a_7845_44172# 0.021949f
C1452 a_11189_46129# a_10490_45724# 0.03271f
C1453 a_17333_42852# VDD 0.525529f
C1454 a_11387_46155# VDD 0.099732f
C1455 a_20623_43914# a_15493_43940# 0.040969f
C1456 en_comp a_n2472_42282# 0.018838f
C1457 a_10490_45724# a_11136_45572# 0.048799f
C1458 a_17339_46660# a_18248_44752# 0.019889f
C1459 a_7754_38968# a_7754_38636# 0.296258f
C1460 a_6031_43396# a_6765_43638# 0.053479f
C1461 a_6293_42852# a_6197_43396# 0.213423f
C1462 a_13249_42308# a_11827_44484# 0.029876f
C1463 a_9313_45822# a_8953_45546# 0.038855f
C1464 a_6540_46812# a_6755_46942# 0.057503f
C1465 a_7577_46660# a_8145_46902# 0.170059f
C1466 a_7411_46660# a_8667_46634# 0.043475f
C1467 a_16137_43396# a_17333_42852# 0.01487f
C1468 a_n1853_43023# a_n1736_43218# 0.183149f
C1469 a_n901_43156# a_n1076_43230# 0.234322f
C1470 a_19778_44110# a_18494_42460# 0.04586f
C1471 a_11415_45002# a_22591_46660# 0.172844f
C1472 a_15368_46634# a_15015_46420# 0.012546f
C1473 a_14976_45028# a_14840_46494# 0.010576f
C1474 a_13483_43940# VDD 0.219591f
C1475 a_21496_47436# VDD 0.198362f
C1476 a_20990_47178# SINGLE_ENDED 0.067698f
C1477 a_17957_46116# a_18147_46436# 0.011458f
C1478 a_17715_44484# a_16375_45002# 0.026655f
C1479 a_10533_42308# a_10723_42308# 0.23663f
C1480 a_21363_46634# VDD 0.357368f
C1481 a_167_45260# a_375_42282# 0.017297f
C1482 a_17339_46660# a_16922_45042# 0.02918f
C1483 a_16375_45002# a_15861_45028# 0.029833f
C1484 a_8199_44636# a_8953_45002# 0.12099f
C1485 a_8270_45546# a_5883_43914# 0.20967f
C1486 a_6755_46942# a_14539_43914# 0.094724f
C1487 a_2905_45572# a_2747_46873# 0.010677f
C1488 a_15507_47210# a_15673_47210# 0.81159f
C1489 a_20623_45572# a_20528_45572# 0.049827f
C1490 a_20841_45814# a_20731_45938# 0.097745f
C1491 a_21363_45546# a_21188_45572# 0.233657f
C1492 C4_P_btm C0_dummy_P_btm 0.113156f
C1493 EN_VIN_BSTR_N C9_N_btm 0.226529f
C1494 C2_P_btm C1_P_btm 5.24136f
C1495 C3_P_btm C0_P_btm 0.409238f
C1496 EN_VIN_BSTR_P VDD 0.917665f
C1497 a_17339_46660# a_15743_43084# 0.450316f
C1498 SMPL_ON_P VDD 0.613427f
C1499 a_18494_42460# a_20159_44458# 0.024732f
C1500 a_5343_44458# a_5708_44484# 0.048542f
C1501 a_8270_45546# a_8162_45546# 0.170838f
C1502 a_8035_47026# VDD 0.132317f
C1503 a_10428_46928# CLK 0.032943f
C1504 a_14539_43914# a_15037_43940# 0.054182f
C1505 a_13059_46348# a_13556_45296# 0.274813f
C1506 a_15597_42852# VDD 0.239357f
C1507 a_n863_45724# a_375_42282# 0.451905f
C1508 CAL_N a_22537_39537# 0.02334f
C1509 a_22589_40055# a_22848_40081# 0.010269f
C1510 a_2747_46873# a_2443_46660# 0.129886f
C1511 a_3754_39964# VDD 0.033808f
C1512 a_9803_43646# a_10149_43396# 0.013377f
C1513 a_9482_43914# a_13777_45326# 0.206086f
C1514 a_12469_46902# a_12816_46660# 0.051162f
C1515 a_10796_42968# a_10341_42308# 0.65943f
C1516 a_10991_42826# a_10922_42852# 0.209641f
C1517 a_11827_44484# a_18287_44626# 0.024541f
C1518 a_8953_45546# a_7871_42858# 0.017048f
C1519 a_20159_44458# a_20640_44752# 0.042415f
C1520 a_7640_43914# a_7542_44172# 0.20977f
C1521 a_19321_45002# a_19778_44110# 0.568668f
C1522 a_17303_42282# a_17531_42308# 0.04615f
C1523 a_18083_42858# VDD 0.408512f
C1524 a_11133_46155# VDD 0.176249f
C1525 a_20365_43914# a_15493_43940# 0.048673f
C1526 a_22775_42308# VDD 0.426061f
C1527 a_16023_47582# a_16131_47204# 0.057222f
C1528 a_6031_43396# a_6197_43396# 0.581047f
C1529 a_7411_46660# a_7927_46660# 0.105839f
C1530 a_n2157_42858# a_n1736_43218# 0.089677f
C1531 a_16409_43396# a_16795_42852# 0.010927f
C1532 a_7715_46873# a_5066_45546# 0.020181f
C1533 a_14976_45028# a_15015_46420# 0.012921f
C1534 a_12429_44172# VDD 0.169047f
C1535 a_20894_47436# SINGLE_ENDED 0.044283f
C1536 a_1823_45246# a_1609_45822# 0.35471f
C1537 a_21855_43396# VDD 0.289066f
C1538 COMP_P a_22485_38105# 0.062482f
C1539 a_20623_46660# VDD 0.194217f
C1540 a_1138_42852# a_626_44172# 0.010739f
C1541 a_8199_44636# a_8191_45002# 0.234072f
C1542 a_8270_45546# a_8701_44490# 0.015888f
C1543 a_6755_46942# a_16112_44458# 0.023983f
C1544 a_19466_46812# a_19929_45028# 0.012303f
C1545 a_19321_45002# a_20159_44458# 0.065041f
C1546 a_2952_47436# a_2747_46873# 0.078913f
C1547 a_15507_47210# a_15811_47375# 0.170975f
C1548 a_n4334_38528# a_n4334_38304# 0.052468f
C1549 a_n2302_38778# a_n2216_38778# 0.011479f
C1550 a_7227_42308# VDD 0.296912f
C1551 a_n1917_43396# a_n1809_43762# 0.057222f
C1552 a_20273_45572# a_20731_45938# 0.034619f
C1553 C5_P_btm C0_dummy_P_btm 0.11375f
C1554 EN_VIN_BSTR_N C8_N_btm 0.090252f
C1555 C3_P_btm C1_P_btm 8.06688f
C1556 C4_P_btm C0_P_btm 0.138331f
C1557 a_17339_46660# a_18783_43370# 0.02025f
C1558 a_15227_46910# a_13059_46348# 0.043664f
C1559 a_10991_42826# a_11554_42852# 0.049827f
C1560 a_n2472_42826# a_n2472_42282# 0.025171f
C1561 a_n2497_47436# CLK_DATA 0.026654f
C1562 a_18189_46348# a_17957_46116# 0.038851f
C1563 a_2713_42308# a_2903_42308# 0.23738f
C1564 a_7832_46660# VDD 0.077608f
C1565 a_2957_45546# a_3218_45724# 0.063846f
C1566 a_13059_46348# a_9482_43914# 0.448068f
C1567 a_10586_45546# VDD 0.582083f
C1568 a_22589_40055# a_22527_39145# 0.130029f
C1569 a_22537_40625# a_22581_37893# 0.656829f
C1570 a_9482_43914# a_13556_45296# 0.726155f
C1571 a_11901_46660# a_12816_46660# 0.125324f
C1572 a_10796_42968# a_10922_42852# 0.170059f
C1573 a_10835_43094# a_10341_42308# 0.541777f
C1574 a_3539_42460# a_3905_42558# 0.015463f
C1575 a_11415_45002# a_18189_46348# 0.028334f
C1576 a_20159_44458# a_20362_44736# 0.233657f
C1577 a_13249_42308# a_12545_42858# 0.030353f
C1578 a_19321_45002# a_18911_45144# 0.050257f
C1579 a_10355_46116# a_10490_45724# 0.01084f
C1580 a_17701_42308# VDD 0.243354f
C1581 a_11189_46129# VDD 0.944289f
C1582 a_13483_43940# a_13829_44260# 0.013377f
C1583 a_20935_43940# a_21115_43940# 0.185422f
C1584 a_20269_44172# a_15493_43940# 0.051355f
C1585 a_21613_42308# VDD 0.27399f
C1586 a_6031_43396# a_6293_42852# 0.163953f
C1587 a_10907_45822# CLK 0.035046f
C1588 a_9313_45822# a_8199_44636# 0.015956f
C1589 a_7411_46660# a_8145_46902# 0.053385f
C1590 a_7715_46873# a_7577_46660# 0.205227f
C1591 a_5807_45002# a_16721_46634# 0.112018f
C1592 a_16547_43609# a_16795_42852# 0.081093f
C1593 a_n1423_42826# a_n1076_43230# 0.051162f
C1594 a_16137_43396# a_17701_42308# 0.025497f
C1595 a_5205_44484# a_6109_44484# 0.029986f
C1596 a_16922_45042# a_11827_44484# 0.032223f
C1597 a_22365_46825# a_22591_46660# 0.08571f
C1598 a_20202_43084# a_11415_45002# 0.041726f
C1599 a_11750_44172# VDD 0.131662f
C1600 a_21177_47436# VDD 0.179587f
C1601 a_n699_43396# a_n1761_44111# 0.018554f
C1602 a_10545_42558# a_10533_42308# 0.011812f
C1603 a_20841_46902# VDD 0.20446f
C1604 a_19321_45002# a_19615_44636# 0.035767f
C1605 a_8016_46348# a_8953_45002# 0.016464f
C1606 a_2553_47502# a_2747_46873# 0.14563f
C1607 a_6761_42308# VDD 0.259312f
C1608 a_n1917_43396# a_n2012_43396# 0.049827f
C1609 a_n1699_43638# a_n1809_43762# 0.097745f
C1610 a_20841_45814# a_21188_45572# 0.051162f
C1611 a_20273_45572# a_20528_45572# 0.064178f
C1612 C6_P_btm C0_dummy_P_btm 0.1194f
C1613 C4_P_btm C1_P_btm 0.128167f
C1614 C5_P_btm C0_P_btm 0.138093f
C1615 C3_P_btm C2_P_btm 5.99608f
C1616 EN_VIN_BSTR_N C7_N_btm 0.115875f
C1617 a_n467_45028# a_n452_44636# 0.092885f
C1618 a_17339_46660# a_18525_43370# 0.060382f
C1619 a_5257_43370# a_5164_46348# 0.02844f
C1620 a_10991_42826# a_11301_43218# 0.013793f
C1621 a_10796_42968# a_11554_42852# 0.056391f
C1622 a_n1920_47178# VDD 0.229556f
C1623 a_n2833_47464# CLK_DATA 0.331592f
C1624 a_n809_44244# a_n984_44318# 0.234322f
C1625 a_310_45028# a_n23_45546# 0.022295f
C1626 a_13059_46348# a_13348_45260# 0.010157f
C1627 a_18579_44172# a_18525_43370# 0.012789f
C1628 a_22589_40599# a_22581_37893# 0.365664f
C1629 CAL_N a_22613_38993# 0.010642f
C1630 a_13017_45260# a_14180_45002# 0.079928f
C1631 a_13348_45260# a_13556_45296# 0.189446f
C1632 a_11901_46660# a_12991_46634# 0.042415f
C1633 a_12469_46902# a_12251_46660# 0.209641f
C1634 a_10796_42968# a_10991_42826# 0.206455f
C1635 a_10835_43094# a_10922_42852# 0.053385f
C1636 a_11827_44484# a_17970_44736# 0.012326f
C1637 a_n467_45028# a_n809_44244# 0.010788f
C1638 a_4419_46090# a_4704_46090# 0.016592f
C1639 a_11415_45002# a_17715_44484# 0.032854f
C1640 a_18533_43940# VDD 0.182147f
C1641 a_n1021_46688# VDD 0.226043f
C1642 a_11415_45002# a_15861_45028# 0.041647f
C1643 a_17595_43084# VDD 0.168112f
C1644 a_19862_44208# a_15493_43940# 0.534481f
C1645 a_21887_42336# VDD 0.210392f
C1646 a_15673_47210# a_5807_45002# 0.011029f
C1647 a_16241_47178# a_16131_47204# 0.097745f
C1648 a_7411_46660# a_7577_46660# 0.634781f
C1649 a_5807_45002# a_16388_46812# 0.235518f
C1650 a_n1853_43023# a_n13_43084# 0.109925f
C1651 a_n1991_42858# a_n1076_43230# 0.123255f
C1652 a_16547_43609# a_16414_43172# 0.143695f
C1653 a_15009_46634# a_15015_46420# 0.012232f
C1654 a_5257_43370# a_5066_45546# 0.053231f
C1655 a_10807_43548# VDD 0.68049f
C1656 a_20990_47178# VDD 0.210484f
C1657 a_19787_47423# START 0.220891f
C1658 a_15368_46634# a_15599_45572# 0.100853f
C1659 a_1176_45822# a_1609_45822# 0.010535f
C1660 a_20273_46660# VDD 0.247553f
C1661 a_n2267_43396# a_n1809_43762# 0.034619f
C1662 a_20273_45572# a_21188_45572# 0.125324f
C1663 a_20107_45572# a_20528_45572# 0.086377f
C1664 a_13249_42308# a_14537_43396# 0.020089f
C1665 C7_P_btm C0_dummy_P_btm 0.119061f
C1666 a_n1550_35448# VDD 0.366274f
C1667 C4_P_btm C2_P_btm 7.72909f
C1668 C5_P_btm C1_P_btm 0.127408f
C1669 C6_P_btm C0_P_btm 0.139059f
C1670 EN_VIN_BSTR_N C6_N_btm 0.118916f
C1671 a_15743_43084# a_16823_43084# 0.031733f
C1672 a_17339_46660# a_18429_43548# 0.033468f
C1673 a_5807_45002# a_5066_45546# 0.027744f
C1674 a_22315_44484# VDD 0.213791f
C1675 a_10835_43094# a_11554_42852# 0.086334f
C1676 a_19778_44110# a_19615_44636# 0.012379f
C1677 a_16922_45042# a_19279_43940# 0.018289f
C1678 a_5883_43914# a_9241_44734# 0.010354f
C1679 a_17715_44484# a_18189_46348# 0.014348f
C1680 a_17583_46090# a_17957_46116# 0.092344f
C1681 a_1755_42282# a_5379_42460# 0.045501f
C1682 a_2725_42558# a_2713_42308# 0.01129f
C1683 a_n967_45348# a_n1076_43230# 0.019022f
C1684 a_n699_43396# a_n2129_43609# 0.062898f
C1685 a_10586_45546# a_10053_45546# 0.024917f
C1686 a_17715_44484# a_17478_45572# 0.017416f
C1687 a_310_45028# a_n356_45724# 0.12349f
C1688 a_n1099_45572# a_n23_45546# 0.042611f
C1689 a_15861_45028# a_17478_45572# 0.080824f
C1690 a_5807_45002# a_19321_45002# 0.376188f
C1691 CAL_N a_22581_37893# 0.023534f
C1692 a_22537_40625# a_22527_39145# 0.245895f
C1693 a_22959_45572# VDD 0.304443f
C1694 a_20107_45572# a_18494_42460# 0.010062f
C1695 a_13017_45260# a_13777_45326# 0.195607f
C1696 a_13348_45260# a_9482_43914# 0.352976f
C1697 a_11735_46660# a_12816_46660# 0.102325f
C1698 a_11901_46660# a_12251_46660# 0.219633f
C1699 a_10835_43094# a_10991_42826# 0.105839f
C1700 a_10518_42984# a_10922_42852# 0.051162f
C1701 a_8375_44464# VDD 0.086619f
C1702 a_11827_44484# a_17767_44458# 0.014019f
C1703 a_18597_46090# a_19431_45546# 0.062716f
C1704 a_19319_43548# VDD 0.561461f
C1705 a_10057_43914# a_10807_43548# 0.039192f
C1706 a_6109_44484# a_6453_43914# 0.165572f
C1707 a_13249_42308# a_12379_42858# 0.029761f
C1708 a_16795_42852# VDD 0.179044f
C1709 a_10355_46116# VDD 0.222751f
C1710 a_20623_43914# a_20935_43940# 0.040559f
C1711 a_19478_44306# a_15493_43940# 0.025498f
C1712 a_21335_42336# VDD 0.199586f
C1713 a_15673_47210# a_16131_47204# 0.034619f
C1714 a_5343_44458# a_8325_42308# 0.014133f
C1715 a_9313_45822# a_8016_46348# 0.02464f
C1716 a_5807_45002# a_13059_46348# 0.1145f
C1717 a_7411_46660# a_7715_46873# 0.162909f
C1718 a_16137_43396# a_16795_42852# 0.010001f
C1719 a_n1853_43023# a_n1076_43230# 0.040291f
C1720 a_n1991_42858# a_n901_43156# 0.041762f
C1721 a_n1423_42826# a_n1641_43230# 0.209641f
C1722 a_5205_44484# a_5289_44734# 0.011388f
C1723 a_22365_46825# a_20202_43084# 0.115624f
C1724 a_10949_43914# VDD 0.797824f
C1725 a_20894_47436# VDD 0.188358f
C1726 a_19386_47436# START 0.042951f
C1727 a_13059_46348# a_15143_45578# 0.262261f
C1728 a_5807_45002# a_13556_45296# 0.017285f
C1729 a_7845_44172# a_8333_44056# 0.065494f
C1730 a_20411_46873# VDD 0.348821f
C1731 a_n2946_38778# a_n2860_38778# 0.011479f
C1732 a_n2267_43396# a_n2012_43396# 0.064178f
C1733 a_n1177_43370# a_n447_43370# 0.010921f
C1734 a_20841_45814# a_20623_45572# 0.209641f
C1735 a_20273_45572# a_21363_45546# 0.042415f
C1736 a_20107_45572# a_21188_45572# 0.102355f
C1737 a_13249_42308# a_14180_45002# 0.014749f
C1738 a_n2002_35448# VDD 0.522945f
C1739 a_12891_46348# a_6755_46942# 0.025465f
C1740 C5_P_btm C2_P_btm 0.13795f
C1741 C4_P_btm C3_P_btm 9.61674f
C1742 C7_P_btm C0_P_btm 0.140846f
C1743 C6_P_btm C1_P_btm 0.127656f
C1744 EN_VIN_BSTR_N C5_N_btm 0.115337f
C1745 C8_P_btm C0_dummy_P_btm 0.234177f
C1746 a_n2840_42826# a_n2840_42282# 0.025171f
C1747 a_n2288_47178# VDD 0.29372f
C1748 a_18479_45785# a_19319_43548# 0.102555f
C1749 a_n699_43396# a_3363_44484# 0.07346f
C1750 a_n1331_43914# a_n984_44318# 0.051162f
C1751 a_n1079_45724# a_n1013_45572# 0.010598f
C1752 a_13059_46348# a_13017_45260# 0.022433f
C1753 a_17715_44484# a_15861_45028# 0.184272f
C1754 a_n1099_45572# a_n356_45724# 0.070228f
C1755 a_18504_43218# VDD 0.077608f
C1756 a_n2302_40160# a_n2302_39866# 0.050477f
C1757 a_22589_40599# a_22527_39145# 1.41544f
C1758 a_22537_40625# a_22589_40055# 0.076642f
C1759 a_15095_43370# a_14955_43396# 0.130374f
C1760 a_13017_45260# a_13556_45296# 0.049621f
C1761 a_13159_45002# a_9482_43914# 0.020865f
C1762 a_11901_46660# a_12469_46902# 0.175891f
C1763 a_11735_46660# a_12991_46634# 0.043475f
C1764 a_10835_43094# a_10796_42968# 0.671797f
C1765 a_7640_43914# VDD 0.196713f
C1766 a_n2293_45010# a_895_43940# 0.283316f
C1767 a_11827_44484# a_16979_44734# 0.012885f
C1768 a_n1177_44458# a_n452_44636# 0.011059f
C1769 a_5807_45002# a_19778_44110# 0.032504f
C1770 a_16414_43172# VDD 0.201389f
C1771 a_9823_46155# VDD 0.102474f
C1772 VREF_GND VCM 2.79113f
C1773 a_22959_47212# a_22959_46660# 0.025171f
C1774 a_16137_43396# a_16414_43172# 0.179708f
C1775 a_n1853_43023# a_n901_43156# 0.081949f
C1776 a_n2157_42858# a_n1076_43230# 0.102325f
C1777 a_n1991_42858# a_n1641_43230# 0.229804f
C1778 a_5205_44484# a_5205_44734# 0.015405f
C1779 a_18587_45118# a_18911_45144# 0.010993f
C1780 a_10729_43914# VDD 0.681371f
C1781 a_19787_47423# VDD 0.256911f
C1782 a_18597_46090# START 0.020125f
C1783 a_1823_45246# a_3905_42558# 0.010516f
C1784 a_3147_46376# a_3316_45546# 0.012262f
C1785 a_5807_45002# a_9482_43914# 0.018229f
C1786 a_21487_43396# VDD 0.222231f
C1787 a_20107_46660# VDD 0.442554f
C1788 a_n2129_43609# a_n2012_43396# 0.183186f
C1789 a_n1177_43370# a_n1352_43396# 0.233657f
C1790 a_20273_45572# a_20623_45572# 0.219856f
C1791 a_20107_45572# a_21363_45546# 0.043567f
C1792 a_11309_47204# a_6755_46942# 0.09972f
C1793 a_5807_45002# a_7715_46873# 0.029268f
C1794 C5_P_btm C3_P_btm 0.135528f
C1795 C8_P_btm C0_P_btm 0.146541f
C1796 C7_P_btm C1_P_btm 0.128479f
C1797 C6_P_btm C2_P_btm 0.137206f
C1798 EN_VIN_BSTR_N C4_N_btm 0.116925f
C1799 C9_P_btm C0_dummy_P_btm 0.111645f
C1800 a_21398_44850# VDD 0.077608f
C1801 a_n2497_47436# VDD 1.33346f
C1802 a_17583_46090# a_17715_44484# 0.22771f
C1803 a_n1899_43946# a_n984_44318# 0.118759f
C1804 a_380_45546# a_n356_45724# 0.088749f
C1805 a_16115_45572# a_16223_45938# 0.057222f
C1806 CAL_N a_22527_39145# 0.010004f
C1807 a_22589_40599# a_22589_40055# 0.086408f
C1808 a_22591_45572# VDD 0.314172f
C1809 a_10695_43548# a_10849_43646# 0.010303f
C1810 a_14205_43396# a_14955_43396# 0.157423f
C1811 SMPL_ON_P COMP_P 0.03194f
C1812 a_13017_45260# a_9482_43914# 0.048717f
C1813 a_13159_45002# a_13348_45260# 0.105274f
C1814 a_10623_46897# a_10933_46660# 0.013793f
C1815 a_11735_46660# a_12251_46660# 0.105995f
C1816 a_6755_46942# a_12156_46660# 0.013732f
C1817 a_9804_47204# a_9823_46155# 0.063581f
C1818 a_10518_42984# a_10796_42968# 0.118759f
C1819 a_6109_44484# VDD 0.243629f
C1820 a_11827_44484# a_14539_43914# 0.044058f
C1821 a_n1177_44458# a_n1352_44484# 0.233657f
C1822 a_18911_45144# a_18989_43940# 0.016276f
C1823 a_n2104_46634# VDD 0.286113f
C1824 a_10057_43914# a_10729_43914# 0.063518f
C1825 a_15567_42826# VDD 0.163583f
C1826 a_9569_46155# VDD 0.19288f
C1827 a_12429_44172# a_12603_44260# 0.011572f
C1828 a_19862_44208# a_21115_43940# 0.064973f
C1829 a_19328_44172# a_15493_43940# 0.062184f
C1830 a_20365_43914# a_20623_43914# 0.22264f
C1831 a_11962_45724# a_11682_45822# 0.014813f
C1832 a_6755_46942# a_14673_44172# 0.050772f
C1833 a_20712_42282# VDD 0.282526f
C1834 a_7754_39964# a_7754_38470# 0.241119f
C1835 a_3754_39134# a_3754_38802# 0.296258f
C1836 a_n967_45348# a_n955_45028# 0.014419f
C1837 VREF VCM 44.262398f
C1838 a_n1853_43023# a_n1641_43230# 0.036072f
C1839 a_n2157_42858# a_n901_43156# 0.043475f
C1840 a_n1991_42858# a_n1423_42826# 0.186387f
C1841 a_327_44734# a_556_44484# 0.033015f
C1842 a_7499_43078# a_11750_44172# 0.195997f
C1843 a_10405_44172# VDD 0.408512f
C1844 a_19386_47436# VDD 0.121241f
C1845 a_18780_47178# START 0.01578f
C1846 a_18479_47436# SINGLE_ENDED 0.040779f
C1847 a_n967_45348# a_n1352_43396# 0.010028f
C1848 a_3147_46376# a_3218_45724# 0.0111f
C1849 a_13059_46348# a_13249_42308# 0.306398f
C1850 a_20556_43646# VDD 0.34939f
C1851 a_19551_46910# VDD 0.226848f
C1852 a_7845_44172# a_7911_44260# 0.010598f
C1853 a_6171_42473# VDD 0.184622f
C1854 a_n1761_44111# a_n901_43156# 0.013702f
C1855 a_n2433_43396# a_n2012_43396# 0.089677f
C1856 a_13249_42308# a_13556_45296# 0.059719f
C1857 a_20107_45572# a_20623_45572# 0.103168f
C1858 a_20273_45572# a_20841_45814# 0.175891f
C1859 a_11309_47204# a_10249_46116# 0.033926f
C1860 C8_P_btm C1_P_btm 0.129306f
C1861 C9_P_btm C0_P_btm 0.146135f
C1862 C5_P_btm C4_P_btm 18.6196f
C1863 C7_P_btm C2_P_btm 0.138288f
C1864 C6_P_btm C3_P_btm 0.133742f
C1865 EN_VIN_BSTR_N C3_N_btm 0.100325f
C1866 C10_P_btm C0_dummy_P_btm 0.749362f
C1867 a_18429_43548# a_16823_43084# 0.130506f
C1868 a_5009_45028# a_5093_45028# 0.092725f
C1869 a_14180_46812# a_13059_46348# 0.074456f
C1870 a_20980_44850# VDD 0.132317f
C1871 a_2779_44458# a_3363_44484# 0.020864f
C1872 a_n2833_47464# VDD 0.461379f
C1873 a_6969_46634# VDD 0.154507f
C1874 a_n1761_44111# a_n984_44318# 0.056404f
C1875 a_n1899_43946# a_n809_44244# 0.042737f
C1876 a_n1331_43914# a_n1549_44318# 0.209641f
C1877 a_n967_45348# a_n1423_42826# 0.010397f
C1878 a_n452_45724# a_n356_45724# 0.318161f
C1879 a_375_42282# a_564_42282# 0.022891f
C1880 a_5745_43940# a_5829_43940# 0.092725f
C1881 a_16115_45572# a_16020_45572# 0.049827f
C1882 a_16333_45814# a_16223_45938# 0.097745f
C1883 a_n2302_37984# VDD 0.350854f
C1884 a_3726_37500# CAL_P 0.102027f
C1885 a_10695_43548# a_10765_43646# 0.011552f
C1886 a_14205_43396# a_15095_43370# 0.086245f
C1887 a_13017_45260# a_13348_45260# 0.044101f
C1888 a_11735_46660# a_12469_46902# 0.053479f
C1889 a_11813_46116# a_11901_46660# 0.211542f
C1890 a_9804_47204# a_9569_46155# 0.040648f
C1891 a_10083_42826# a_10796_42968# 0.042737f
C1892 a_10518_42984# a_10835_43094# 0.102355f
C1893 a_3539_42460# a_3823_42558# 0.07742f
C1894 a_n2661_45010# a_895_43940# 0.020382f
C1895 a_18597_46090# a_18341_45572# 0.010006f
C1896 a_10057_43914# a_10405_44172# 0.028414f
C1897 a_375_42282# a_n1557_42282# 0.450989f
C1898 a_8953_45546# a_8746_45002# 0.020026f
C1899 a_9625_46129# VDD 0.996485f
C1900 a_12429_44172# a_12495_44260# 0.012714f
C1901 a_19862_44208# a_20935_43940# 0.03846f
C1902 a_18451_43940# a_15493_43940# 0.051906f
C1903 a_14539_43914# a_16823_43084# 0.058282f
C1904 a_10053_45546# a_10306_45572# 0.011897f
C1905 a_20107_42308# VDD 0.284252f
C1906 a_n2497_47436# a_3877_44458# 0.024435f
C1907 a_n2302_37984# a_n2302_37690# 0.050477f
C1908 a_22959_43948# a_22959_43396# 0.025171f
C1909 a_20202_43084# a_19862_44208# 0.058613f
C1910 a_n863_45724# a_n23_44458# 0.056041f
C1911 VIN_N VCM 1.7189f
C1912 VREF VREF_GND 44.051197f
C1913 a_16237_45028# VDD 0.248452f
C1914 a_n1853_43023# a_n1423_42826# 0.022091f
C1915 a_n2157_42858# a_n1641_43230# 0.110532f
C1916 a_18315_45260# a_18587_45118# 0.13675f
C1917 a_16922_45042# a_18494_42460# 0.242236f
C1918 a_7499_43078# a_10807_43548# 0.119721f
C1919 a_9672_43914# VDD 0.150499f
C1920 a_18597_46090# VDD 0.930122f
C1921 a_18479_47436# START 0.313639f
C1922 a_n967_45348# a_n1177_43370# 0.013627f
C1923 a_19123_46287# VDD 0.336379f
C1924 a_18494_42460# a_15743_43084# 0.027791f
C1925 en_comp a_n2293_42282# 0.026f
C1926 a_22959_44484# a_22959_43948# 0.026152f
C1927 a_5755_42308# VDD 0.229304f
C1928 a_2112_39137# a_2684_37794# 0.091415f
C1929 a_2277_45546# VDD 0.209584f
C1930 a_n1699_43638# a_n1352_43396# 0.051162f
C1931 a_13249_42308# a_9482_43914# 0.061734f
C1932 a_20107_45572# a_20841_45814# 0.053479f
C1933 a_22725_37990# VDD 0.085163f
C1934 a_n2497_47436# a_n1641_46494# 0.020605f
C1935 a_5807_45002# a_5257_43370# 0.683815f
C1936 C8_P_btm C2_P_btm 0.138777f
C1937 C9_P_btm C1_P_btm 0.132506f
C1938 C10_P_btm C0_P_btm 0.365593f
C1939 C7_P_btm C3_P_btm 0.134911f
C1940 C6_P_btm C4_P_btm 0.143514f
C1941 EN_VIN_BSTR_N C2_N_btm 0.118072f
C1942 a_626_44172# VDD 0.621601f
C1943 a_17324_43396# a_16823_43084# 0.038999f
C1944 a_n967_45348# a_n1177_44458# 0.012502f
C1945 a_14035_46660# a_13059_46348# 0.072321f
C1946 a_15682_46116# a_17583_46090# 0.013015f
C1947 a_6755_46942# VDD 1.05713f
C1948 a_n1761_44111# a_n809_44244# 0.038277f
C1949 a_n2065_43946# a_n984_44318# 0.102325f
C1950 a_n1899_43946# a_n1549_44318# 0.218775f
C1951 a_n967_45348# a_n1991_42858# 0.034664f
C1952 a_15765_45572# a_16223_45938# 0.027606f
C1953 a_8953_45546# a_8975_43940# 0.02155f
C1954 a_22589_40599# a_22537_40625# 1.96968f
C1955 a_13017_45260# a_13159_45002# 0.160415f
C1956 a_3429_45260# a_3495_45348# 0.010598f
C1957 a_11735_46660# a_11901_46660# 0.579036f
C1958 a_9804_47204# a_9625_46129# 0.037672f
C1959 a_10083_42826# a_10835_43094# 0.043619f
C1960 a_3539_42460# a_3318_42354# 0.161793f
C1961 a_n2293_45010# a_453_43940# 0.181603f
C1962 a_n1699_44726# a_n1352_44484# 0.051162f
C1963 a_15037_43940# VDD 0.190221f
C1964 a_8975_43940# a_9028_43914# 0.184602f
C1965 a_10057_43914# a_9672_43914# 0.143523f
C1966 a_19321_45002# a_16922_45042# 0.493823f
C1967 a_8199_44636# a_10490_45724# 0.019372f
C1968 a_15279_43071# VDD 0.189193f
C1969 a_17124_42282# a_17303_42282# 0.172579f
C1970 a_8953_45546# VDD 1.32809f
C1971 a_19862_44208# a_20623_43914# 0.023134f
C1972 a_18326_43940# a_15493_43940# 0.075033f
C1973 a_20269_44172# a_20365_43914# 0.419086f
C1974 a_11525_45546# a_11682_45822# 0.18824f
C1975 a_10053_45546# a_10216_45572# 0.011381f
C1976 a_16023_47582# a_16119_47582# 0.013793f
C1977 a_7754_39300# a_7754_38968# 0.296258f
C1978 a_3877_44458# a_6969_46634# 0.101189f
C1979 VIN_P VCM 1.7189f
C1980 VIN_N VREF_GND 16.4969f
C1981 a_20193_45348# VDD 0.793111f
C1982 a_n2157_42858# a_n1423_42826# 0.07009f
C1983 a_n1853_43023# a_n1991_42858# 0.237526f
C1984 a_7499_43078# a_10949_43914# 0.152939f
C1985 a_9028_43914# VDD 0.17194f
C1986 a_22223_42860# a_22400_42852# 0.154104f
C1987 a_20922_43172# a_20753_42852# 0.08213f
C1988 a_18989_43940# a_19006_44850# 0.168452f
C1989 a_18780_47178# VDD 0.245515f
C1990 a_13059_46348# a_13527_45546# 0.017655f
C1991 a_20301_43646# VDD 0.296691f
C1992 a_9803_42558# a_9885_42558# 0.171361f
C1993 a_18285_46348# VDD 0.259614f
C1994 a_22959_46124# a_22959_45572# 0.025171f
C1995 a_1609_45822# VDD 0.270106f
C1996 a_n2129_43609# a_n447_43370# 0.119518f
C1997 a_n2267_43396# a_n1352_43396# 0.124988f
C1998 a_20107_45572# a_20273_45572# 0.667378f
C1999 a_22629_37990# VDD 0.079474f
C2000 a_9804_47204# a_6755_46942# 0.028571f
C2001 a_1983_46706# a_n2661_46098# 0.147223f
C2002 C8_P_btm C3_P_btm 0.134581f
C2003 C9_P_btm C2_P_btm 0.141891f
C2004 C10_P_btm C1_P_btm 0.31753f
C2005 C7_P_btm C4_P_btm 0.145303f
C2006 C6_P_btm C5_P_btm 22.305399f
C2007 EN_VIN_BSTR_N C1_N_btm 0.110046f
C2008 a_17499_43370# a_16823_43084# 0.064861f
C2009 a_10249_46116# VDD 1.03004f
C2010 a_n1761_44111# a_n1549_44318# 0.033724f
C2011 a_n2065_43946# a_n809_44244# 0.043475f
C2012 a_n1899_43946# a_n1331_43914# 0.171939f
C2013 a_n967_45348# a_n1853_43023# 0.021497f
C2014 a_1431_47204# a_2124_47436# 0.010942f
C2015 a_15765_45572# a_16020_45572# 0.056391f
C2016 a_6545_47178# a_6755_46942# 0.022995f
C2017 a_n2946_37984# VDD 0.38275f
C2018 a_22223_45572# VDD 0.287831f
C2019 a_14579_43548# a_15095_43370# 0.109081f
C2020 a_14358_43442# a_14205_43396# 0.163543f
C2021 a_7499_43078# a_7640_43914# 0.021219f
C2022 a_11735_46660# a_11813_46116# 0.162547f
C2023 a_10083_42826# a_10518_42984# 0.234322f
C2024 a_20202_43084# a_21195_42852# 0.018373f
C2025 a_n2661_45010# a_2127_44172# 0.096614f
C2026 a_n967_45348# a_n1899_43946# 0.025102f
C2027 a_n2129_44697# a_n452_44636# 0.079904f
C2028 a_n2267_44484# a_n1352_44484# 0.118759f
C2029 a_n746_45260# a_327_44734# 0.256943f
C2030 a_5807_45002# a_14495_45572# 0.012666f
C2031 a_13565_43940# VDD 0.175245f
C2032 a_n2472_46634# VDD 0.287589f
C2033 a_8199_44636# a_8746_45002# 0.680077f
C2034 a_9625_46129# a_10053_45546# 0.086776f
C2035 a_19862_44208# a_20365_43914# 0.075162f
C2036 a_18079_43940# a_15493_43940# 0.040279f
C2037 en_comp a_22400_42852# 0.721871f
C2038 a_11322_45546# a_11682_45822# 0.034435f
C2039 a_5066_45546# a_8953_45002# 0.013782f
C2040 a_19647_42308# VDD 0.227331f
C2041 a_16023_47582# a_15928_47570# 0.049827f
C2042 VDAC_Pi VDAC_Ni 3.18068f
C2043 a_n745_45366# a_n467_45028# 0.110406f
C2044 a_3877_44458# a_6755_46942# 0.388535f
C2045 VIN_N VREF 0.775904f
C2046 VIN_P VREF_GND 16.4969f
C2047 a_n2157_42858# a_n1991_42858# 0.905962f
C2048 a_14537_43396# a_14539_43914# 0.135541f
C2049 a_17719_45144# a_18315_45260# 0.017382f
C2050 a_16922_45042# a_19778_44110# 0.026041f
C2051 a_7499_43078# a_10729_43914# 0.23002f
C2052 a_19987_42826# a_20753_42852# 0.07365f
C2053 a_8333_44056# VDD 0.124235f
C2054 a_18479_47436# VDD 1.47669f
C2055 a_n1917_44484# a_n1899_43946# 0.012479f
C2056 a_17829_46910# VDD 0.37446f
C2057 a_n2129_43609# a_n1352_43396# 0.041828f
C2058 a_n1699_43638# a_n1917_43396# 0.209641f
C2059 a_n2267_43396# a_n1177_43370# 0.041762f
C2060 VDAC_P VCM 11.743501f
C2061 a_22725_38406# VDD 0.085997f
C2062 a_18597_46090# a_19466_46812# 0.074092f
C2063 a_n2497_47436# a_n1991_46122# 0.037858f
C2064 a_8128_46384# a_6755_46942# 0.01823f
C2065 a_9804_47204# a_10249_46116# 0.034717f
C2066 a_11309_47204# a_10467_46802# 0.023291f
C2067 a_1983_46706# a_1799_45572# 0.089984f
C2068 C8_P_btm C4_P_btm 0.145646f
C2069 C9_P_btm C3_P_btm 0.137552f
C2070 C10_P_btm C2_P_btm 0.327137f
C2071 C7_P_btm C5_P_btm 0.151416f
C2072 EN_VIN_BSTR_N C0_N_btm 0.12803f
C2073 a_16759_43396# a_16823_43084# 0.038761f
C2074 a_375_42282# VDD 0.591443f
C2075 a_19333_46634# a_19551_46910# 0.08213f
C2076 a_22165_42308# a_22223_42860# 0.171681f
C2077 a_16922_45042# a_20159_44458# 0.012027f
C2078 a_742_44458# a_556_44484# 0.044092f
C2079 a_6655_43762# VDD 0.132357f
C2080 a_10554_47026# VDD 0.205847f
C2081 a_n1761_44111# a_n1331_43914# 0.043168f
C2082 a_n2065_43946# a_n1549_44318# 0.110816f
C2083 a_n967_45348# a_n2157_42858# 0.02564f
C2084 a_15682_46116# a_16855_45546# 0.011741f
C2085 a_14635_42282# VDD 0.369964f
C2086 a_16855_45546# a_16680_45572# 0.233657f
C2087 a_15903_45785# a_16020_45572# 0.157972f
C2088 a_8199_44636# a_8975_43940# 0.028334f
C2089 a_9803_43646# a_9885_43646# 0.171361f
C2090 a_14579_43548# a_14205_43396# 0.066243f
C2091 a_4905_42826# a_4921_42308# 0.046918f
C2092 a_n967_45348# a_n1761_44111# 0.015839f
C2093 a_20202_43084# a_21356_42826# 0.011854f
C2094 a_n2129_44697# a_n1352_44484# 0.048248f
C2095 a_n1699_44726# a_n1917_44484# 0.209641f
C2096 a_n2267_44484# a_n1177_44458# 0.042415f
C2097 a_5807_45002# a_13249_42308# 0.725941f
C2098 a_18285_46348# a_18175_45572# 0.010439f
C2099 a_12891_46348# a_11827_44484# 0.020579f
C2100 a_11415_45002# a_15903_45785# 0.02962f
C2101 a_14543_43071# VDD 0.18866f
C2102 a_8199_44636# VDD 1.43837f
C2103 a_17973_43940# a_15493_43940# 0.028173f
C2104 a_19862_44208# a_20269_44172# 0.049487f
C2105 a_10490_45724# a_11682_45822# 0.014138f
C2106 a_19511_42282# VDD 0.244902f
C2107 a_7754_39964# VDAC_Ni 0.207118f
C2108 a_5343_44458# a_7963_42308# 0.108654f
C2109 SMPL_ON_N a_22591_46660# 0.011048f
C2110 VIN_P VREF 0.775904f
C2111 a_n2157_42858# a_n1853_43023# 0.290902f
C2112 a_16922_45042# a_18911_45144# 0.042178f
C2113 a_14537_43396# a_16112_44458# 0.093722f
C2114 a_7499_43078# a_10405_44172# 0.132405f
C2115 a_19987_42826# a_20356_42852# 0.014848f
C2116 a_18374_44850# a_18588_44850# 0.097745f
C2117 a_18443_44721# a_19006_44850# 0.049827f
C2118 a_18143_47464# VDD 0.388551f
C2119 a_1823_45246# a_3823_42558# 0.137565f
C2120 a_1823_45246# a_3503_45724# 0.295715f
C2121 a_14275_46494# a_14383_46116# 0.057222f
C2122 a_21259_43561# VDD 0.192954f
C2123 a_9223_42460# a_9377_42558# 0.010303f
C2124 a_8953_45546# a_5111_44636# 0.181796f
C2125 a_6511_45714# a_7227_45028# 0.213161f
C2126 a_6667_45809# a_6598_45938# 0.209641f
C2127 a_4921_42308# VDD 0.214995f
C2128 a_509_45822# VDD 0.190119f
C2129 a_n2129_43609# a_n1177_43370# 0.08445f
C2130 a_n2267_43396# a_n1917_43396# 0.227165f
C2131 a_n2433_43396# a_n1352_43396# 0.102325f
C2132 a_n1761_44111# a_n1853_43023# 0.019636f
C2133 VDAC_P VREF_GND 0.203715f
C2134 CAL_P RST_Z 0.551895f
C2135 a_22629_38406# VDD 0.315181f
C2136 a_n2497_47436# a_n1853_46287# 0.029452f
C2137 a_11309_47204# a_10428_46928# 0.025525f
C2138 a_948_46660# a_n2661_46098# 0.018472f
C2139 C9_P_btm C4_P_btm 0.154834f
C2140 C10_P_btm C3_P_btm 0.321945f
C2141 C8_P_btm C5_P_btm 0.145019f
C2142 C7_P_btm C6_P_btm 26.0771f
C2143 EN_VIN_BSTR_N C0_dummy_N_btm 0.026355f
C2144 a_16977_43638# a_16823_43084# 0.022663f
C2145 a_16751_45260# VDD 0.121848f
C2146 a_14180_45002# a_14309_45028# 0.062574f
C2147 a_19333_46634# a_19123_46287# 0.113955f
C2148 a_18287_44626# a_18989_43940# 0.193279f
C2149 a_18443_44721# a_18374_44850# 0.209641f
C2150 a_6452_43396# VDD 0.083252f
C2151 a_10623_46897# VDD 0.189083f
C2152 a_n2065_43946# a_n1331_43914# 0.053479f
C2153 a_n1761_44111# a_n1899_43946# 0.737653f
C2154 a_1239_47204# a_1431_47204# 0.219138f
C2155 a_1209_47178# a_2124_47436# 0.095065f
C2156 a_13291_42460# VDD 0.546706f
C2157 a_7845_44172# a_7287_43370# 0.011834f
C2158 a_15493_43940# a_20974_43370# 0.069596f
C2159 a_375_42282# a_196_42282# 0.165785f
C2160 a_15599_45572# a_16020_45572# 0.086708f
C2161 a_8199_44636# a_10057_43914# 0.113262f
C2162 a_n3690_38304# VDD 0.363068f
C2163 a_21513_45002# VDD 0.416919f
C2164 a_13667_43396# a_14205_43396# 0.076384f
C2165 a_14579_43548# a_14358_43442# 0.142377f
C2166 a_8953_45002# a_9482_43914# 0.010057f
C2167 a_2680_45002# a_2903_45348# 0.011458f
C2168 a_18479_45785# a_19113_45348# 0.013845f
C2169 a_9313_45822# a_5066_45546# 0.019449f
C2170 a_n2293_45010# a_1115_44172# 0.09282f
C2171 a_n2661_45010# a_1414_42308# 0.059385f
C2172 a_n967_45348# a_n2065_43946# 0.02253f
C2173 a_n2129_44697# a_n1177_44458# 0.027646f
C2174 a_n2267_44484# a_n1917_44484# 0.212549f
C2175 a_n2433_44484# a_n1352_44484# 0.102355f
C2176 a_n746_45260# a_n37_45144# 0.031257f
C2177 a_5807_45002# CLK 0.033646f
C2178 a_17339_46660# a_18341_45572# 0.015732f
C2179 a_8016_46348# a_8746_45002# 0.078716f
C2180 a_8953_45546# a_9049_44484# 0.03092f
C2181 a_8199_44636# a_10180_45724# 0.216999f
C2182 a_13460_43230# VDD 0.276534f
C2183 a_8349_46414# VDD 0.209819f
C2184 a_17737_43940# a_15493_43940# 0.037029f
C2185 a_10807_43548# a_11173_44260# 0.05223f
C2186 a_13249_42308# a_14495_45572# 0.027073f
C2187 a_11322_45546# a_10907_45822# 0.012408f
C2188 a_n2946_37984# a_n2946_37690# 0.050477f
C2189 a_22731_47423# a_22591_46660# 0.011433f
C2190 a_5807_45002# a_14035_46660# 0.025174f
C2191 a_22959_45036# VDD 0.30999f
C2192 a_17613_45144# a_17719_45144# 0.080654f
C2193 a_16922_45042# a_18587_45118# 0.021516f
C2194 a_14537_43396# a_15004_44636# 0.047224f
C2195 a_19987_42826# a_20256_42852# 0.015204f
C2196 a_18287_44626# a_19006_44850# 0.086658f
C2197 a_18443_44721# a_18588_44850# 0.057222f
C2198 en_comp a_n2267_43396# 0.028399f
C2199 a_1823_45246# a_3318_42354# 0.055532f
C2200 a_n967_45348# a_n2129_43609# 0.021282f
C2201 a_1823_45246# a_3316_45546# 0.099099f
C2202 a_14493_46090# a_14383_46116# 0.097745f
C2203 a_9223_42460# a_9293_42558# 0.011552f
C2204 a_22485_44484# a_15493_43940# 0.087012f
C2205 a_17339_46660# VDD 0.555596f
C2206 a_6511_45714# a_6598_45938# 0.06628f
C2207 a_6472_45840# a_7227_45028# 0.208286f
C2208 a_n2433_43396# a_n1177_43370# 0.043475f
C2209 a_n2129_43609# a_n1917_43396# 0.036131f
C2210 a_n2267_43396# a_n1699_43638# 0.179796f
C2211 VDAC_N VCM 11.7445f
C2212 CAL_P VDD 22.475801f
C2213 a_n2497_47436# a_n2157_46122# 0.034181f
C2214 a_1123_46634# a_n2661_46098# 0.041919f
C2215 C8_P_btm C6_P_btm 0.163943f
C2216 C10_P_btm C4_P_btm 0.703336f
C2217 C9_P_btm C5_P_btm 0.150576f
C2218 a_16409_43396# a_16823_43084# 0.020816f
C2219 a_16759_43396# a_16855_43396# 0.013793f
C2220 a_n967_45348# a_n2129_44697# 0.017689f
C2221 en_comp a_n2267_44484# 0.029536f
C2222 a_2905_45572# a_3175_45822# 0.046585f
C2223 a_14180_46812# a_14513_46634# 0.253235f
C2224 a_18579_44172# VDD 0.38178f
C2225 a_18287_44626# a_18374_44850# 0.053385f
C2226 a_18248_44752# a_18989_43940# 0.207562f
C2227 a_8103_44636# a_8375_44464# 0.13675f
C2228 a_5883_43914# a_6109_44484# 0.078113f
C2229 a_5111_44636# a_8333_44056# 0.280148f
C2230 a_11827_44484# a_14673_44172# 0.150125f
C2231 a_2123_42473# a_2351_42308# 0.084895f
C2232 a_9396_43370# VDD 0.288403f
C2233 a_10467_46802# VDD 0.401016f
C2234 a_n2065_43946# a_n1899_43946# 0.614122f
C2235 a_n863_45724# a_2713_42308# 0.044499f
C2236 en_comp a_n2472_42826# 0.019667f
C2237 a_15682_46116# a_16333_45814# 0.011944f
C2238 a_380_45546# a_997_45618# 0.070624f
C2239 a_n746_45260# a_175_44278# 0.159759f
C2240 a_1209_47178# a_1431_47204# 0.095209f
C2241 a_13003_42852# VDD 0.132655f
C2242 a_8034_45724# VDD 0.812726f
C2243 a_16333_45814# a_16680_45572# 0.051162f
C2244 a_15903_45785# a_15861_45028# 0.232345f
C2245 a_8016_46348# a_8975_43940# 0.01976f
C2246 a_11787_45002# a_11963_45334# 0.185422f
C2247 a_2680_45002# a_2809_45348# 0.010132f
C2248 a_n2104_46634# a_n2157_46122# 0.013135f
C2249 a_9127_43156# a_10083_42826# 0.011187f
C2250 a_20202_43084# a_19987_42826# 0.177726f
C2251 a_n2293_45010# a_644_44056# 0.014621f
C2252 a_11827_44484# a_12607_44458# 0.023193f
C2253 a_n2433_44484# a_n1177_44458# 0.043567f
C2254 a_n2129_44697# a_n1917_44484# 0.030172f
C2255 a_n2267_44484# a_n1699_44726# 0.172319f
C2256 a_n746_45260# a_n143_45144# 0.043399f
C2257 a_n2840_46634# VDD 0.306342f
C2258 a_20916_46384# SINGLE_ENDED 0.020511f
C2259 a_17339_46660# a_18479_45785# 0.027772f
C2260 a_8953_45546# a_7499_43078# 0.108436f
C2261 a_5807_45002# a_16922_45042# 0.030945f
C2262 a_8199_44636# a_10053_45546# 0.014322f
C2263 a_13635_43156# VDD 0.463701f
C2264 a_8016_46348# VDD 1.42798f
C2265 a_15682_43940# a_15493_43940# 0.067033f
C2266 a_10490_45724# a_10907_45822# 0.229517f
C2267 a_13059_46348# a_14539_43914# 0.05997f
C2268 a_8568_45546# a_9159_45572# 0.011449f
C2269 a_13904_45546# a_14495_45572# 0.092344f
C2270 a_n746_45260# a_n2661_46098# 0.049386f
C2271 a_15673_47210# a_15928_47570# 0.064178f
C2272 a_11682_45822# VDD 0.316586f
C2273 a_n745_45366# a_n967_45348# 0.010748f
C2274 a_n2661_45010# a_327_44734# 0.04375f
C2275 a_5807_45002# a_13885_46660# 0.014137f
C2276 a_22223_45036# VDD 0.300162f
C2277 a_n2472_42826# a_n2157_42858# 0.080495f
C2278 a_18479_45785# a_18579_44172# 0.045071f
C2279 a_16922_45042# a_18315_45260# 0.065907f
C2280 a_13556_45296# a_14539_43914# 0.025347f
C2281 a_12991_46634# a_13351_46090# 0.011685f
C2282 a_18248_44752# a_19006_44850# 0.056391f
C2283 a_17591_47464# VDD 0.421992f
C2284 a_n746_45260# a_742_44458# 0.0971f
C2285 a_167_45260# a_1848_45724# 0.359783f
C2286 a_13925_46122# a_14383_46116# 0.027606f
C2287 a_22485_44484# a_22223_43948# 0.016889f
C2288 a_20512_43084# a_15493_43940# 0.021257f
C2289 a_8199_44636# a_5111_44636# 0.024227f
C2290 a_13059_46348# a_14309_45028# 0.050896f
C2291 a_6511_45714# a_6667_45809# 0.113977f
C2292 a_6472_45840# a_6598_45938# 0.178024f
C2293 a_3905_42558# VDD 0.176395f
C2294 a_n2129_43609# a_n1699_43638# 0.022218f
C2295 a_n2433_43396# a_n1917_43396# 0.108815f
C2296 a_13163_45724# a_13159_45002# 0.010135f
C2297 VDAC_N VREF_GND 0.203821f
C2298 a_18597_46090# a_18834_46812# 0.010699f
C2299 a_1123_46634# a_1799_45572# 0.037438f
C2300 C8_P_btm C7_P_btm 31.072699f
C2301 C9_P_btm C6_P_btm 0.165353f
C2302 C10_P_btm C5_P_btm 0.51798f
C2303 a_16547_43609# a_16823_43084# 0.08061f
C2304 a_16019_45002# VDD 0.174085f
C2305 a_14797_45144# a_15060_45348# 0.010598f
C2306 a_18834_46812# a_19123_46287# 0.039405f
C2307 a_18287_44626# a_18443_44721# 0.10279f
C2308 a_8103_44636# a_7640_43914# 0.101633f
C2309 a_18248_44752# a_18374_44850# 0.170059f
C2310 a_8791_43396# VDD 0.191045f
C2311 a_10428_46928# VDD 0.278873f
C2312 a_n2065_43946# a_n1761_44111# 0.617556f
C2313 a_15682_46116# a_15765_45572# 0.015911f
C2314 a_1209_47178# a_1239_47204# 0.264529f
C2315 a_n2302_40160# a_n2216_40160# 0.011479f
C2316 a_n4334_40480# a_n4334_39616# 0.050585f
C2317 a_15493_43940# a_21381_43940# 0.02116f
C2318 a_15765_45572# a_16680_45572# 0.118759f
C2319 a_8016_46348# a_10057_43914# 0.09388f
C2320 a_6575_47204# a_8667_46634# 0.01088f
C2321 a_n4334_38304# VDD 0.385989f
C2322 a_8128_46384# a_8349_46414# 0.101217f
C2323 a_9127_43156# a_8952_43230# 0.234322f
C2324 a_n2293_45010# a_175_44278# 0.030523f
C2325 en_comp a_n2472_43914# 0.014244f
C2326 a_11827_44484# a_8975_43940# 0.076327f
C2327 a_n2129_44697# a_n1699_44726# 0.018607f
C2328 a_n2433_44484# a_n1917_44484# 0.113784f
C2329 a_n746_45260# a_n467_45028# 0.054826f
C2330 a_1823_45246# a_4704_46090# 0.164557f
C2331 a_2804_46116# a_3147_46376# 0.017019f
C2332 a_5111_44636# a_6452_43396# 0.024938f
C2333 a_17339_46660# a_18175_45572# 0.019286f
C2334 a_8016_46348# a_10180_45724# 0.259851f
C2335 a_8199_44636# a_9049_44484# 0.029722f
C2336 a_8953_45546# a_8568_45546# 0.136365f
C2337 a_12895_43230# VDD 0.212352f
C2338 a_7920_46348# VDD 0.100184f
C2339 a_14955_43940# a_15493_43940# 0.110232f
C2340 a_10949_43914# a_10555_44260# 0.034175f
C2341 a_10729_43914# a_11173_44260# 0.057346f
C2342 a_n1761_44111# a_n2129_43609# 0.029483f
C2343 a_13904_45546# a_13249_42308# 0.13587f
C2344 a_10490_45724# a_10210_45822# 0.014252f
C2345 a_8568_45546# a_8791_45572# 0.011458f
C2346 a_15811_47375# a_15928_47570# 0.161235f
C2347 a_22223_43948# a_22223_43396# 0.025171f
C2348 a_16147_45260# a_16751_45260# 0.054632f
C2349 a_11827_44484# VDD 0.615802f
C2350 a_16922_45042# a_17719_45144# 0.22253f
C2351 a_18248_44752# a_18588_44850# 0.027606f
C2352 a_16588_47582# VDD 0.282243f
C2353 en_comp a_n2433_43396# 0.036527f
C2354 a_n746_45260# a_n452_44636# 0.042999f
C2355 a_167_45260# a_997_45618# 0.052039f
C2356 a_6194_45824# a_6598_45938# 0.051162f
C2357 a_6472_45840# a_6667_45809# 0.215953f
C2358 a_1169_39043# a_1107_38525# 0.031327f
C2359 a_n2129_43609# a_n2267_43396# 0.230013f
C2360 a_n2433_43396# a_n1699_43638# 0.062578f
C2361 a_18780_47178# a_18834_46812# 0.010748f
C2362 VDAC_P VIN_P 0.255243f
C2363 C9_P_btm C7_P_btm 0.22201f
C2364 C10_P_btm C6_P_btm 0.895671f
C2365 a_19268_43646# a_19700_43370# 0.017165f
C2366 a_16243_43396# a_16823_43084# 0.05964f
C2367 a_15743_43084# a_16664_43396# 0.01372f
C2368 a_15595_45028# VDD 0.156299f
C2369 en_comp a_n2433_44484# 0.029809f
C2370 a_18834_46812# a_18285_46348# 0.144972f
C2371 a_13885_46660# a_14513_46634# 0.101344f
C2372 a_21195_42852# a_21671_42860# 0.177876f
C2373 a_6298_44484# a_7640_43914# 0.031665f
C2374 a_18248_44752# a_18443_44721# 0.206455f
C2375 a_17970_44736# a_18374_44850# 0.051162f
C2376 a_15015_46420# a_14840_46494# 0.233657f
C2377 a_1755_42282# a_2123_42473# 0.014573f
C2378 a_14635_42282# a_14113_42308# 0.052122f
C2379 a_8147_43396# VDD 0.393534f
C2380 a_10150_46912# VDD 0.284144f
C2381 a_n1099_45572# a_310_45028# 0.333219f
C2382 a_15682_46116# a_15903_45785# 0.011633f
C2383 a_n2497_47436# a_895_43940# 0.0309f
C2384 COMP_P a_22629_37990# 0.010153f
C2385 a_15493_43940# a_19741_43940# 0.027038f
C2386 a_15765_45572# a_16855_45546# 0.042415f
C2387 a_16333_45814# a_16115_45572# 0.209641f
C2388 a_8953_45546# a_5883_43914# 0.262126f
C2389 a_18479_45785# a_11827_44484# 0.03055f
C2390 a_2382_45260# a_2304_45348# 0.045704f
C2391 a_8128_46384# a_8016_46348# 0.09182f
C2392 a_22959_43396# a_22959_42860# 0.026152f
C2393 a_n2293_45010# a_n984_44318# 0.048428f
C2394 a_n2129_44697# a_n2267_44484# 0.698671f
C2395 a_n2433_44484# a_n1699_44726# 0.058433f
C2396 a_20411_46873# a_20708_46348# 0.081063f
C2397 a_n2497_47436# a_3065_45002# 0.022803f
C2398 a_1823_45246# a_4419_46090# 0.340207f
C2399 a_5883_43914# a_9028_43914# 0.05428f
C2400 a_5111_44636# a_9396_43370# 0.203348f
C2401 a_8199_44636# a_7499_43078# 0.859274f
C2402 a_8016_46348# a_10053_45546# 0.017312f
C2403 a_13113_42826# VDD 0.217254f
C2404 a_6419_46155# VDD 0.094119f
C2405 a_10729_43914# a_10555_44260# 0.038445f
C2406 a_8746_45002# a_10210_45822# 0.013725f
C2407 a_8568_45546# a_8697_45572# 0.010132f
C2408 a_18214_42558# VDD 0.295211f
C2409 a_15507_47210# a_15928_47570# 0.089677f
C2410 a_3754_39466# a_3754_39134# 0.296258f
C2411 a_10907_45822# VDD 0.352181f
C2412 a_12465_44636# a_11415_45002# 0.375509f
C2413 a_21359_45002# VDD 0.319372f
C2414 a_16922_45042# a_17613_45144# 0.10967f
C2415 a_13556_45296# a_15004_44636# 0.127354f
C2416 a_12251_46660# a_12594_46348# 0.011817f
C2417 a_16137_43396# a_18214_42558# 0.0459f
C2418 a_16763_47508# VDD 0.392885f
C2419 a_1823_45246# a_1848_45724# 0.028459f
C2420 a_16823_43084# VDD 0.159922f
C2421 a_8791_42308# a_9223_42460# 0.014257f
C2422 a_5663_43940# a_6101_44260# 0.013015f
C2423 a_6472_45840# a_6511_45714# 0.781352f
C2424 a_13381_47204# a_13487_47204# 0.152045f
C2425 a_n2433_43396# a_n2267_43396# 0.756435f
C2426 a_22537_39537# VDD 0.313136f
C2427 EN_VIN_BSTR_P C0_dummy_P_btm 0.026355f
C2428 C9_P_btm C8_P_btm 39.4538f
C2429 C10_P_btm C7_P_btm 1.39624f
C2430 VDAC_N VIN_N 0.256435f
C2431 a_6293_42852# a_5755_42852# 0.114235f
C2432 a_16137_43396# a_16823_43084# 0.038492f
C2433 a_15415_45028# VDD 0.191729f
C2434 a_n2661_45010# a_949_44458# 0.071688f
C2435 a_13885_46660# a_14180_46812# 0.150851f
C2436 a_17609_46634# a_18285_46348# 0.115413f
C2437 a_19279_43940# VDD 0.302681f
C2438 a_8387_43230# a_8495_42852# 0.057222f
C2439 a_21356_42826# a_21671_42860# 0.084365f
C2440 a_18248_44752# a_18287_44626# 0.633819f
C2441 a_6298_44484# a_6109_44484# 0.068396f
C2442 a_13291_42460# a_14113_42308# 0.025652f
C2443 a_7112_43396# VDD 0.273193f
C2444 a_9863_46634# VDD 0.411318f
C2445 a_n2472_43914# a_n2065_43946# 0.039807f
C2446 a_380_45546# a_310_45028# 0.057269f
C2447 a_11136_42852# VDD 0.132515f
C2448 a_15599_45572# a_16680_45572# 0.102355f
C2449 a_15765_45572# a_16115_45572# 0.20669f
C2450 a_8199_44636# a_9838_44484# 0.024921f
C2451 a_19862_44208# a_20922_43172# 0.164553f
C2452 a_20202_43084# a_20974_43370# 0.026132f
C2453 a_2274_45254# a_2304_45348# 0.062682f
C2454 a_8128_46384# a_7920_46348# 0.197919f
C2455 a_4905_42826# a_5379_42460# 0.077171f
C2456 a_8605_42826# a_8952_43230# 0.051162f
C2457 a_n2293_45010# a_n809_44244# 0.041966f
C2458 a_n2433_44484# a_n2267_44484# 0.730194f
C2459 a_14537_43396# a_14673_44172# 0.044194f
C2460 a_2698_46116# a_2804_46116# 0.313533f
C2461 a_9801_43940# VDD 0.19512f
C2462 a_5883_43914# a_8333_44056# 0.152643f
C2463 a_5111_44636# a_8791_43396# 0.05316f
C2464 a_20916_46384# VDD 0.302226f
C2465 a_8199_44636# a_8568_45546# 0.141772f
C2466 a_12545_42858# VDD 0.285703f
C2467 a_6165_46155# VDD 0.204296f
C2468 a_10405_44172# a_10555_44260# 0.085098f
C2469 a_19328_44172# a_19478_44306# 0.188181f
C2470 a_n2497_47436# a_n229_43646# 0.022782f
C2471 a_19332_42282# VDD 0.227361f
C2472 a_9313_45822# a_5807_45002# 0.031627f
C2473 a_n3690_38304# a_n3690_37440# 0.050585f
C2474 a_10210_45822# VDD 0.323342f
C2475 a_16147_45260# a_16019_45002# 0.186254f
C2476 a_22223_47212# a_22365_46825# 0.011422f
C2477 a_6545_47178# a_6419_46155# 0.080336f
C2478 a_21101_45002# VDD 0.2903f
C2479 a_18479_45785# a_19279_43940# 0.019159f
C2480 a_13556_45296# a_13720_44458# 0.212774f
C2481 a_16922_45042# a_17023_45118# 0.099834f
C2482 a_9482_43914# a_15004_44636# 0.34299f
C2483 a_3935_42891# a_3823_42558# 0.012124f
C2484 a_16023_47582# VDD 0.201413f
C2485 a_12891_46348# a_13777_45326# 0.03955f
C2486 a_n746_45260# a_n1177_44458# 0.064145f
C2487 a_8685_42308# a_9223_42460# 0.166964f
C2488 a_22223_46124# a_22223_45572# 0.025171f
C2489 a_6194_45824# a_6511_45714# 0.102325f
C2490 a_5379_42460# VDD 0.213136f
C2491 a_n23_45546# VDD 0.150941f
C2492 a_n2433_43396# a_n2129_43609# 0.283605f
C2493 a_22889_38993# VDD 0.495671f
C2494 a_9804_47204# a_9863_46634# 0.017882f
C2495 EN_VIN_BSTR_P C0_P_btm 0.12803f
C2496 a_383_46660# a_479_46660# 0.013793f
C2497 a_171_46873# a_n2661_46098# 0.168482f
C2498 C10_P_btm C8_P_btm 2.07867f
C2499 a_10775_45002# CLK 0.058141f
C2500 a_15743_43084# a_19268_43646# 0.010228f
C2501 a_14797_45144# VDD 0.124624f
C2502 a_n2661_45010# a_742_44458# 0.694478f
C2503 a_n2293_45010# a_n1352_44484# 0.020183f
C2504 a_13885_46660# a_14035_46660# 0.25868f
C2505 a_17609_46634# a_17829_46910# 0.111805f
C2506 a_20766_44850# VDD 0.197657f
C2507 a_21356_42826# a_21195_42852# 0.03853f
C2508 a_8605_42826# a_8495_42852# 0.097745f
C2509 a_626_44172# a_895_43940# 0.038336f
C2510 a_5518_44484# a_6109_44484# 0.050093f
C2511 a_17970_44736# a_18287_44626# 0.102355f
C2512 a_5343_44458# a_7640_43914# 0.152634f
C2513 a_19321_45002# a_19431_45546# 0.029441f
C2514 a_14493_46090# a_14840_46494# 0.051162f
C2515 a_13291_42460# a_13657_42558# 0.026223f
C2516 a_7287_43370# VDD 0.457521f
C2517 a_8492_46660# VDD 0.273866f
C2518 a_n863_45724# a_2351_42308# 0.038802f
C2519 a_380_45546# a_n1099_45572# 0.148825f
C2520 a_5807_45002# a_14539_43914# 0.066683f
C2521 a_21115_43940# a_21381_43940# 0.073198f
C2522 a_15599_45572# a_16855_45546# 0.043567f
C2523 a_15765_45572# a_16333_45814# 0.17072f
C2524 a_8016_46348# a_10157_44484# 0.016596f
C2525 a_7903_47542# a_8145_46902# 0.010369f
C2526 a_17715_44484# a_17737_43940# 0.289085f
C2527 a_10775_45002# a_10951_45334# 0.185422f
C2528 a_4905_42826# a_5267_42460# 0.146764f
C2529 a_8037_42858# a_8952_43230# 0.118759f
C2530 a_n23_44458# VDD 0.169093f
C2531 a_n2293_45010# a_n1549_44318# 0.014826f
C2532 a_n2433_44484# a_n2129_44697# 0.130072f
C2533 a_n2497_47436# a_2382_45260# 0.042349f
C2534 a_n746_45260# a_n967_45348# 0.028689f
C2535 a_626_44172# a_458_43396# 0.065365f
C2536 a_19594_46812# START 0.020669f
C2537 a_5111_44636# a_8147_43396# 0.08322f
C2538 a_8199_44636# a_8162_45546# 0.119979f
C2539 a_12089_42308# VDD 0.807892f
C2540 a_5497_46414# VDD 0.200657f
C2541 a_7542_44172# a_7499_43940# 0.157633f
C2542 a_8162_45546# a_8192_45572# 0.134163f
C2543 a_18907_42674# VDD 0.148872f
C2544 a_13487_47204# a_13569_47204# 0.014524f
C2545 a_1431_47204# a_1123_46634# 0.012069f
C2546 a_7754_39632# a_7754_39300# 0.296258f
C2547 a_n2661_45010# a_n467_45028# 0.227953f
C2548 a_12891_46348# a_13059_46348# 0.372745f
C2549 DATA[5] CLK 0.059607f
C2550 a_21005_45260# VDD 0.184261f
C2551 a_9482_43914# a_13720_44458# 0.188323f
C2552 a_22000_46634# a_20202_43084# 0.154237f
C2553 a_167_45260# a_310_45028# 0.035247f
C2554 a_12891_46348# a_13556_45296# 0.29495f
C2555 a_22400_42852# a_22485_38105# 0.198011f
C2556 a_8685_42308# a_8791_42308# 0.147376f
C2557 a_5907_45546# a_6511_45714# 0.043475f
C2558 a_6194_45824# a_6472_45840# 0.118423f
C2559 a_5267_42460# VDD 0.170631f
C2560 a_n356_45724# VDD 0.719282f
C2561 a_20202_43084# a_20512_43084# 0.130366f
C2562 a_22613_38993# VDD 0.533489f
C2563 EN_VIN_BSTR_P C1_P_btm 0.110046f
C2564 C10_P_btm C9_P_btm 53.3168f
C2565 a_8953_45002# CLK 0.310391f
C2566 a_14537_43396# VDD 0.779752f
C2567 a_n2661_45010# a_n452_44636# 0.020671f
C2568 a_14180_45002# a_14403_45348# 0.011458f
C2569 a_20835_44721# VDD 0.198384f
C2570 a_8037_42858# a_8495_42852# 0.027317f
C2571 a_20922_43172# a_21195_42852# 0.119168f
C2572 a_17767_44458# a_18287_44626# 0.043567f
C2573 a_17970_44736# a_18248_44752# 0.117156f
C2574 a_5343_44458# a_6109_44484# 0.285594f
C2575 a_5518_44484# a_5826_44734# 0.017351f
C2576 a_7499_43078# a_8791_43396# 0.04623f
C2577 a_2804_46116# a_2981_46116# 0.134298f
C2578 a_1138_42852# a_1337_46116# 0.039951f
C2579 a_13925_46122# a_14840_46494# 0.118759f
C2580 a_6547_43396# VDD 0.219105f
C2581 a_8667_46634# VDD 0.39254f
C2582 a_n863_45724# a_2123_42473# 0.036254f
C2583 a_n863_45724# a_310_45028# 0.033427f
C2584 a_n452_45724# a_n1099_45572# 0.053931f
C2585 a_n2497_47436# a_453_43940# 0.09742f
C2586 a_n785_47204# a_327_47204# 0.237391f
C2587 COMP_P CAL_P 0.037539f
C2588 a_2479_44172# a_2813_43396# 0.115852f
C2589 a_15493_43940# a_18533_43940# 0.052096f
C2590 a_15599_45572# a_16115_45572# 0.105995f
C2591 a_8199_44636# a_8701_44490# 0.25266f
C2592 VDAC_N VDAC_P 4.74149f
C2593 a_2684_37794# VDD 0.286899f
C2594 a_20731_45938# VDD 0.142103f
C2595 a_19431_45546# a_19778_44110# 0.010264f
C2596 a_20202_43084# a_21381_43940# 0.108097f
C2597 a_6755_46942# a_15368_46634# 0.033754f
C2598 a_n2472_46634# a_n2472_46090# 0.026152f
C2599 a_8605_42826# a_8387_43230# 0.209641f
C2600 a_8037_42858# a_9127_43156# 0.042737f
C2601 a_n2293_45010# a_n1331_43914# 0.02919f
C2602 a_2521_46116# a_2698_46116# 0.159555f
C2603 a_9165_43940# VDD 0.192035f
C2604 a_19321_45002# START 0.10793f
C2605 a_5111_44636# a_7112_43396# 0.041581f
C2606 a_20843_47204# VDD 0.188032f
C2607 a_12379_42858# VDD 0.484153f
C2608 a_5204_45822# VDD 0.359177f
C2609 a_7281_43914# a_7499_43940# 0.08213f
C2610 a_9672_43914# a_9895_44260# 0.011458f
C2611 a_13163_45724# a_13527_45546# 0.124682f
C2612 a_10053_45546# a_10210_45822# 0.18824f
C2613 a_18727_42674# VDD 0.181095f
C2614 VDAC_Pi a_3754_39134# 0.012307f
C2615 a_2113_38308# VDAC_Ni 0.318652f
C2616 a_3499_42826# a_3681_42891# 0.033957f
C2617 a_8697_45822# VDD 0.189893f
C2618 a_n2109_45247# en_comp 0.108653f
C2619 a_n2293_45010# a_n967_45348# 0.018659f
C2620 a_7499_43078# a_11827_44484# 0.104754f
C2621 a_5907_46634# a_5257_43370# 0.070316f
C2622 a_20567_45036# VDD 0.237324f
C2623 a_9482_43914# a_13076_44458# 0.103066f
C2624 a_19987_42826# a_20256_43172# 0.043356f
C2625 a_16241_47178# VDD 0.208959f
C2626 a_5205_44484# a_6671_43940# 0.049504f
C2627 a_16979_44734# a_17325_44484# 0.013377f
C2628 a_1176_45822# a_997_45618# 0.140567f
C2629 a_12891_46348# a_9482_43914# 0.314487f
C2630 a_14275_46494# a_14371_46494# 0.013793f
C2631 a_8325_42308# a_8791_42308# 0.173196f
C2632 a_16721_46634# VDD 0.186443f
C2633 a_5907_45546# a_6472_45840# 0.041762f
C2634 a_3823_42558# VDD 0.170296f
C2635 a_3503_45724# VDD 0.129733f
C2636 a_14955_43940# a_14955_43396# 0.012141f
C2637 en_comp a_22485_38105# 0.535686f
C2638 a_22581_37893# VDD 0.902719f
C2639 EN_VIN_BSTR_P C2_P_btm 0.118072f
C2640 a_18783_43370# a_15743_43084# 0.303966f
C2641 a_14180_45002# VDD 0.151315f
C2642 a_n2661_45010# a_n1352_44484# 0.051998f
C2643 a_14180_45002# a_14309_45348# 0.010132f
C2644 a_4955_46873# a_5068_46348# 0.081759f
C2645 a_17609_46634# a_17339_46660# 0.010277f
C2646 a_20679_44626# VDD 0.439119f
C2647 a_20922_43172# a_21356_42826# 0.017093f
C2648 a_17767_44458# a_18248_44752# 0.041822f
C2649 a_7499_43078# a_8147_43396# 0.227361f
C2650 a_1176_45822# a_1337_46116# 0.026848f
C2651 a_14493_46090# a_14275_46494# 0.209641f
C2652 a_13759_46122# a_14840_46494# 0.102325f
C2653 a_13925_46122# a_15015_46420# 0.042415f
C2654 a_14635_42282# a_14456_42282# 0.172313f
C2655 a_6765_43638# VDD 0.218204f
C2656 a_7927_46660# VDD 0.187888f
C2657 a_n863_45724# a_1755_42282# 0.050501f
C2658 a_8034_45724# a_8162_45546# 0.14162f
C2659 a_n863_45724# a_n1099_45572# 0.172847f
C2660 a_n23_47502# a_327_47204# 0.140943f
C2661 a_12800_43218# VDD 0.078978f
C2662 a_5111_44636# a_5379_42460# 0.118194f
C2663 a_15493_43940# a_19319_43548# 0.36082f
C2664 a_15599_45572# a_16333_45814# 0.053479f
C2665 a_15903_45785# a_15765_45572# 0.205788f
C2666 a_8199_44636# a_8103_44636# 0.256009f
C2667 a_13059_46348# a_14673_44172# 0.108306f
C2668 a_6886_37412# VDAC_P 0.062773f
C2669 a_1107_38525# VDD 0.374783f
C2670 a_20528_45572# VDD 0.08228f
C2671 a_n2840_43370# a_n2840_42826# 0.026152f
C2672 a_13249_42308# a_14539_43914# 0.032256f
C2673 a_18597_46090# a_19900_46494# 0.039688f
C2674 a_6755_46942# a_14976_45028# 0.029836f
C2675 a_8037_42858# a_8387_43230# 0.225358f
C2676 a_7871_42858# a_8952_43230# 0.102355f
C2677 a_n2293_45010# a_n1899_43946# 0.18948f
C2678 a_13556_45296# a_14673_44172# 0.137701f
C2679 a_167_45260# a_2698_46116# 0.019127f
C2680 a_375_42282# a_458_43396# 0.014454f
C2681 a_5111_44636# a_7287_43370# 0.104641f
C2682 a_19594_46812# VDD 0.349555f
C2683 a_10341_42308# VDD 0.931019f
C2684 a_5164_46348# VDD 0.717083f
C2685 a_9672_43914# a_9801_44260# 0.010132f
C2686 a_13059_46348# a_12607_44458# 0.033056f
C2687 a_18057_42282# VDD 0.130308f
C2688 a_n2293_45010# en_comp 0.066194f
C2689 a_18494_42460# VDD 0.73193f
C2690 a_10807_43548# a_11323_42473# 0.109765f
C2691 a_13556_45296# a_12607_44458# 0.01896f
C2692 a_11813_46116# a_12005_46116# 0.038046f
C2693 a_21363_46634# a_20202_43084# 0.048242f
C2694 a_16137_43396# a_18057_42282# 0.01884f
C2695 a_3499_42826# VDD 0.333472f
C2696 a_9313_45822# CLK 0.027301f
C2697 a_15673_47210# VDD 0.569224f
C2698 a_12891_46348# a_13348_45260# 0.097519f
C2699 a_14275_46494# a_14180_46482# 0.049827f
C2700 a_n2497_47436# a_n699_43396# 0.355158f
C2701 a_8325_42308# a_8685_42308# 0.141819f
C2702 a_18494_42460# a_16137_43396# 0.115144f
C2703 a_22315_44484# a_22223_43948# 0.012307f
C2704 a_16388_46812# VDD 0.797417f
C2705 a_5907_45546# a_6194_45824# 0.233657f
C2706 a_3318_42354# VDD 0.203036f
C2707 a_3316_45546# VDD 0.428912f
C2708 a_n2840_43370# a_n2433_43396# 0.039807f
C2709 a_17591_47464# a_17609_46634# 0.014668f
C2710 EN_VIN_BSTR_P C3_P_btm 0.100325f
C2711 a_383_46660# a_491_47026# 0.057222f
C2712 a_18525_43370# a_15743_43084# 0.058072f
C2713 a_16759_43396# a_16867_43762# 0.057222f
C2714 a_13777_45326# VDD 0.145151f
C2715 a_5257_43370# a_5111_42852# 0.013892f
C2716 a_n2661_45010# a_n1177_44458# 0.052759f
C2717 a_4955_46873# a_4704_46090# 0.109136f
C2718 a_20640_44752# VDD 0.246486f
C2719 a_17767_44458# a_17970_44736# 0.233657f
C2720 a_626_44172# a_453_43940# 0.163589f
C2721 a_7499_43078# a_7112_43396# 0.012965f
C2722 a_5807_45002# a_19256_45572# 0.015716f
C2723 a_18285_46348# a_18051_46116# 0.028958f
C2724 a_1208_46090# a_1337_46116# 0.062574f
C2725 a_13925_46122# a_14275_46494# 0.20669f
C2726 a_13759_46122# a_15015_46420# 0.043475f
C2727 a_1184_42692# a_2123_42473# 0.107417f
C2728 a_13291_42460# a_14456_42282# 0.015899f
C2729 a_6197_43396# VDD 0.408793f
C2730 a_8145_46902# VDD 0.199702f
C2731 a_n1079_45724# a_n1099_45572# 0.15766f
C2732 a_n2497_47436# a_1467_44172# 0.046456f
C2733 a_n23_47502# a_n785_47204# 0.031198f
C2734 a_5111_44636# a_5267_42460# 0.047489f
C2735 a_1414_42308# a_3457_43396# 0.094207f
C2736 a_19862_44208# a_20974_43370# 0.026213f
C2737 a_5066_45546# VDD 1.34058f
C2738 a_2277_45546# a_2274_45254# 0.011988f
C2739 a_15599_45572# a_15765_45572# 0.576512f
C2740 a_21188_45572# VDD 0.288663f
C2741 a_18597_46090# a_20075_46420# 0.073857f
C2742 a_18479_47436# a_20708_46348# 0.04299f
C2743 a_22223_43396# a_22223_42860# 0.026152f
C2744 a_8037_42858# a_8605_42826# 0.178024f
C2745 a_7871_42858# a_9127_43156# 0.043633f
C2746 a_n2293_45010# a_n1761_44111# 0.148418f
C2747 a_9482_43914# a_14673_44172# 0.42967f
C2748 a_167_45260# a_2521_46116# 0.328009f
C2749 a_5111_44636# a_6547_43396# 0.035842f
C2750 a_19321_45002# VDD 1.01574f
C2751 a_5257_43370# a_5205_44484# 0.021038f
C2752 a_10922_42852# VDD 0.216186f
C2753 a_5068_46348# VDD 0.085085f
C2754 a_6453_43914# a_6671_43940# 0.08213f
C2755 a_n2840_43914# a_n2840_43370# 0.025171f
C2756 a_17531_42308# VDD 0.262303f
C2757 a_n4334_38304# a_n4334_37440# 0.050585f
C2758 a_n746_45260# a_288_46660# 0.010226f
C2759 a_n2661_45010# a_n967_45348# 0.019427f
C2760 a_n2472_45002# en_comp 0.117861f
C2761 a_9482_43914# a_12607_44458# 0.151452f
C2762 a_15811_47375# VDD 0.979053f
C2763 a_11459_47204# DATA[5] 0.370451f
C2764 a_12891_46348# a_13159_45002# 0.031652f
C2765 a_n746_45260# a_n2129_44697# 0.17701f
C2766 a_13059_46348# VDD 0.955445f
C2767 a_5164_46348# a_4927_45028# 0.09665f
C2768 a_n2302_39072# a_n2302_38778# 0.050477f
C2769 a_2903_42308# VDD 0.22017f
C2770 a_3218_45724# VDD 0.133843f
C2771 a_22527_39145# VDD 0.626886f
C2772 EN_VIN_BSTR_P C4_P_btm 0.116925f
C2773 a_383_46660# a_288_46660# 0.049827f
C2774 a_601_46902# a_491_47026# 0.097745f
C2775 a_13556_45296# VDD 0.569056f
C2776 a_16759_43396# a_16664_43396# 0.049827f
C2777 a_18429_43548# a_15743_43084# 0.053516f
C2778 a_16977_43638# a_16867_43762# 0.097745f
C2779 a_18525_43370# a_18783_43370# 0.22264f
C2780 a_n2661_45010# a_n1917_44484# 0.015623f
C2781 a_n2293_45010# a_n2267_44484# 0.0118f
C2782 a_4651_46660# a_4704_46090# 0.013135f
C2783 a_20362_44736# VDD 0.275577f
C2784 a_7499_43078# a_7287_43370# 0.057949f
C2785 a_11827_44484# a_11541_44484# 0.0442f
C2786 a_19321_45002# a_18479_45785# 0.114441f
C2787 a_5807_45002# a_19431_45546# 0.01527f
C2788 a_13925_46122# a_14493_46090# 0.17072f
C2789 a_13759_46122# a_14275_46494# 0.105995f
C2790 a_6293_42852# VDD 0.401011f
C2791 a_13291_42460# a_13575_42558# 0.074792f
C2792 a_1184_42692# a_1755_42282# 0.016329f
C2793 a_7577_46660# VDD 0.249866f
C2794 a_n863_45724# a_n452_45724# 0.046903f
C2795 a_n2497_47436# a_1115_44172# 0.069778f
C2796 a_n746_45260# a_327_47204# 0.022743f
C2797 a_11554_42852# VDD 0.078978f
C2798 COMP_P a_22537_39537# 0.03695f
C2799 a_1609_45822# a_2274_45254# 0.11737f
C2800 a_15599_45572# a_15903_45785# 0.161702f
C2801 a_8530_39574# CAL_P 0.037066f
C2802 a_3726_37500# CAL_N 0.036205f
C2803 a_6886_37412# VDAC_N 0.067053f
C2804 a_12891_46348# a_5807_45002# 0.044188f
C2805 a_7227_47204# a_7411_46660# 0.011806f
C2806 a_21363_45546# VDD 0.36538f
C2807 a_8270_45546# a_9803_43646# 0.066865f
C2808 a_18597_46090# a_19335_46494# 0.036056f
C2809 a_6545_47178# a_5066_45546# 0.021464f
C2810 a_6755_46942# a_15009_46634# 0.012747f
C2811 a_15095_43370# a_15597_42852# 0.071983f
C2812 a_7871_42858# a_8387_43230# 0.106107f
C2813 a_n2293_45010# a_n2065_43946# 0.023134f
C2814 a_n2840_44458# a_n2433_44484# 0.039807f
C2815 a_n746_45260# a_n745_45366# 0.119822f
C2816 a_7499_43940# VDD 0.193884f
C2817 a_5343_44458# a_8333_44056# 0.092296f
C2818 a_5111_44636# a_6765_43638# 0.022146f
C2819 a_20202_43084# a_21613_42308# 0.07574f
C2820 a_19466_46812# a_20528_45572# 0.157758f
C2821 a_10991_42826# VDD 0.201891f
C2822 a_4704_46090# VDD 0.225404f
C2823 a_18326_43940# a_18451_43940# 0.145292f
C2824 a_14539_43914# a_15743_43084# 0.024623f
C2825 a_17303_42282# VDD 0.37938f
C2826 a_22731_47423# a_22959_47212# 0.08444f
C2827 a_n1557_42282# a_648_43396# 0.048175f
C2828 a_n2661_45010# en_comp 0.10363f
C2829 a_19594_46812# a_19466_46812# 0.100902f
C2830 a_5167_46660# a_5263_46660# 0.013793f
C2831 a_19778_44110# VDD 0.469922f
C2832 a_13017_45260# a_13076_44458# 0.011055f
C2833 a_9482_43914# a_8975_43940# 0.186623f
C2834 a_626_44172# a_n699_43396# 0.042617f
C2835 a_11813_46116# a_11387_46155# 0.080527f
C2836 a_15507_47210# VDD 0.441662f
C2837 a_9313_45822# DATA[5] 0.055804f
C2838 SMPL_ON_N a_21753_35474# 0.39912f
C2839 a_n2840_44458# a_n2840_43914# 0.026152f
C2840 a_13925_46122# a_14180_46482# 0.056391f
C2841 a_167_45260# a_n863_45724# 0.424358f
C2842 a_12891_46348# a_13017_45260# 0.210934f
C2843 a_5807_45002# a_6431_45366# 0.018543f
C2844 a_n2497_47436# a_2779_44458# 0.034441f
C2845 a_8337_42558# a_8325_42308# 0.01416f
C2846 a_15227_46910# VDD 0.229766f
C2847 a_20512_43084# a_19862_44208# 0.023947f
C2848 a_5164_46348# a_5111_44636# 0.024532f
C2849 a_2713_42308# VDD 0.208275f
C2850 a_2957_45546# VDD 0.192471f
C2851 a_11652_45724# a_11787_45002# 0.077604f
C2852 a_22589_40055# VDD 1.08898f
C2853 a_8128_46384# a_8145_46902# 0.012246f
C2854 EN_VIN_BSTR_P C5_P_btm 0.115337f
C2855 a_19998_34978# a_21753_35474# 0.150805f
C2856 a_33_46660# a_491_47026# 0.027606f
C2857 a_9482_43914# VDD 1.75061f
C2858 a_16409_43396# a_16867_43762# 0.027606f
C2859 a_17324_43396# a_15743_43084# 0.050725f
C2860 a_1823_45246# a_3539_42460# 0.678673f
C2861 a_n2661_45010# a_n1699_44726# 0.04137f
C2862 a_n2293_45010# a_n2129_44697# 0.021404f
C2863 a_8128_46384# a_5066_45546# 0.032968f
C2864 a_18597_46090# a_19240_46482# 0.025784f
C2865 a_20159_44458# VDD 0.345429f
C2866 a_16979_44734# a_17767_44458# 0.011457f
C2867 a_375_42282# a_453_43940# 0.021162f
C2868 a_19321_45002# a_18175_45572# 0.01259f
C2869 a_19123_46287# a_19240_46482# 0.157972f
C2870 a_13759_46122# a_14493_46090# 0.053479f
C2871 a_6031_43396# VDD 0.47547f
C2872 a_13291_42460# a_13070_42354# 0.155164f
C2873 a_1576_42282# a_1755_42282# 0.168925f
C2874 a_22959_42860# a_22775_42308# 0.019713f
C2875 a_7715_46873# VDD 0.414019f
C2876 a_n2497_47436# a_644_44056# 0.016428f
C2877 a_n746_45260# a_n785_47204# 0.198992f
C2878 a_3065_45002# a_3905_42558# 0.044632f
C2879 a_19862_44208# a_21381_43940# 0.113704f
C2880 a_11309_47204# a_5807_45002# 0.032739f
C2881 a_n2302_38778# VDD 0.35162f
C2882 a_20623_45572# VDD 0.200978f
C2883 a_327_44734# a_626_44172# 0.120093f
C2884 a_18597_46090# a_19553_46090# 0.021441f
C2885 a_18479_47436# a_20075_46420# 0.061108f
C2886 a_6755_46942# a_14084_46812# 0.052304f
C2887 a_n2840_46634# a_n2840_46090# 0.026152f
C2888 a_n1809_44850# VDD 0.132538f
C2889 a_7871_42858# a_8605_42826# 0.06628f
C2890 a_7765_42852# a_8037_42858# 0.309282f
C2891 a_2202_46116# a_167_45260# 0.159883f
C2892 a_6671_43940# VDD 0.227011f
C2893 a_5111_44636# a_6197_43396# 0.025934f
C2894 a_20202_43084# a_21887_42336# 0.082645f
C2895 a_n746_45260# a_556_44484# 0.045671f
C2896 a_10796_42968# VDD 0.270235f
C2897 a_15959_42545# a_16269_42308# 0.013793f
C2898 a_4419_46090# VDD 0.664887f
C2899 a_5663_43940# a_5829_43940# 0.143754f
C2900 a_8199_44636# a_8560_45348# 0.03862f
C2901 a_7499_43078# a_8697_45822# 0.038073f
C2902 a_18597_46090# a_15493_43940# 0.024181f
C2903 VDAC_Pi a_3754_39466# 0.308867f
C2904 a_19321_45002# a_19466_46812# 0.130025f
C2905 a_19594_46812# a_19333_46634# 0.060858f
C2906 VDD VCM 1.50561f
C2907 a_18911_45144# VDD 0.218047f
C2908 a_9482_43914# a_10057_43914# 0.401746f
C2909 a_18599_43230# a_18707_42852# 0.057222f
C2910 a_9313_45822# DATA[4] 0.0373f
C2911 SMPL_ON_N a_19998_34978# 0.01194f
C2912 a_n1853_46287# a_n356_45724# 0.011459f
C2913 a_13759_46122# a_14180_46482# 0.086708f
C2914 a_n2497_47436# a_949_44458# 0.127971f
C2915 a_5164_46348# a_5147_45002# 0.060833f
C2916 a_9313_45822# a_11459_47204# 0.210847f
C2917 a_1848_45724# VDD 0.100884f
C2918 a_11322_45546# a_11963_45334# 0.028732f
C2919 a_16375_45002# a_16237_45028# 0.035582f
C2920 a_8128_46384# a_7577_46660# 0.023306f
C2921 EN_VIN_BSTR_P C6_P_btm 0.118916f
C2922 a_1123_46634# a_948_46660# 0.234322f
C2923 a_33_46660# a_288_46660# 0.056391f
C2924 a_13348_45260# VDD 0.083657f
C2925 a_17499_43370# a_15743_43084# 0.049383f
C2926 a_16409_43396# a_16664_43396# 0.056391f
C2927 a_18429_43548# a_18525_43370# 0.419086f
C2928 a_n2661_45010# a_n2267_44484# 0.260289f
C2929 a_n2293_45010# a_n2433_44484# 0.016908f
C2930 a_18597_46090# a_16375_45002# 0.105669f
C2931 a_19615_44636# VDD 0.203841f
C2932 a_17339_46660# a_18051_46116# 0.040259f
C2933 a_13759_46122# a_13925_46122# 0.576786f
C2934 a_7411_46660# VDD 0.41059f
C2935 a_n863_45724# a_961_42354# 0.038222f
C2936 a_n1079_45724# a_n863_45724# 0.091159f
C2937 a_n2497_47436# a_175_44278# 0.05097f
C2938 a_n746_45260# a_n23_47502# 0.148631f
C2939 a_19862_44208# a_19741_43940# 0.038152f
C2940 a_5257_43370# a_5663_43940# 0.014098f
C2941 a_3726_37500# VDAC_P 0.059581f
C2942 a_20841_45814# VDD 0.209907f
C2943 a_20512_43084# a_20256_43172# 0.047194f
C2944 a_20974_43370# a_20749_43396# 0.0837f
C2945 a_18597_46090# a_18985_46122# 0.027318f
C2946 a_6755_46942# a_13607_46688# 0.129798f
C2947 a_n2012_44484# VDD 0.077632f
C2948 a_7871_42858# a_8037_42858# 0.772842f
C2949 a_1823_45246# a_167_45260# 0.155648f
C2950 a_19123_46287# a_18985_46122# 0.215692f
C2951 a_12891_46348# a_13249_42308# 0.166217f
C2952 SMPL_ON_P en_comp 0.034192f
C2953 a_5829_43940# VDD 0.156797f
C2954 a_20193_45348# a_15493_43940# 0.10893f
C2955 a_7499_43078# a_10341_42308# 0.42152f
C2956 a_5111_44636# a_6293_42852# 0.072755f
C2957 a_20202_43084# a_21335_42336# 0.227943f
C2958 a_10835_43094# VDD 0.43308f
C2959 a_5663_43940# a_5745_43940# 0.096132f
C2960 a_18079_43940# a_18326_43940# 0.152347f
C2961 a_11962_45724# a_13163_45724# 0.113317f
C2962 a_12427_45724# a_12791_45546# 0.124682f
C2963 a_8568_45546# a_8697_45822# 0.062574f
C2964 a_22731_47423# SMPL_ON_N 0.194951f
C2965 a_n2497_47436# a_n2661_46098# 0.026032f
C2966 a_5257_43370# a_4905_42826# 0.254437f
C2967 VDD VREF_GND 0.482759f
C2968 a_18587_45118# VDD 0.085535f
C2969 a_375_42282# a_n699_43396# 0.127058f
C2970 a_20623_46660# a_20719_46660# 0.013793f
C2971 a_18817_42826# a_18707_42852# 0.097745f
C2972 a_1847_42826# a_2713_42308# 0.015903f
C2973 a_14955_47212# VDD 0.301751f
C2974 a_16112_44458# a_16335_44484# 0.011458f
C2975 a_14311_47204# RST_Z 0.184572f
C2976 a_1823_45246# a_n863_45724# 0.207189f
C2977 a_n2497_47436# a_742_44458# 0.153038f
C2978 a_22400_42852# a_21613_42308# 0.02387f
C2979 a_8515_42308# a_8685_42308# 0.108744f
C2980 a_3600_43914# a_3499_42826# 0.125876f
C2981 a_19466_46812# a_19778_44110# 0.116901f
C2982 a_997_45618# VDD 0.12359f
C2983 a_11322_45546# a_11787_45002# 0.035999f
C2984 a_22537_40625# VDD 0.534319f
C2985 a_19250_34978# a_19998_34978# 0.08192f
C2986 EN_VIN_BSTR_P C7_P_btm 0.115875f
C2987 a_171_46873# a_288_46660# 0.159893f
C2988 a_13159_45002# VDD 0.321035f
C2989 a_21381_43940# a_21195_42852# 0.238789f
C2990 a_16759_43396# a_15743_43084# 0.033478f
C2991 a_16547_43609# a_16664_43396# 0.161376f
C2992 a_n2661_45010# a_n2129_44697# 0.18531f
C2993 a_14976_45028# a_15312_46660# 0.01024f
C2994 a_19339_43156# a_19987_42826# 0.016188f
C2995 a_14539_43914# a_16979_44734# 0.132799f
C2996 a_626_44172# a_644_44056# 0.126386f
C2997 a_5257_43370# VDD 0.922495f
C2998 a_n863_45724# a_1184_42692# 0.563857f
C2999 a_5883_43914# a_9165_43940# 0.019684f
C3000 a_11415_45002# a_22591_45572# 0.02488f
C3001 a_n452_47436# a_n785_47204# 0.03755f
C3002 a_1337_46116# VDD 0.20087f
C3003 a_2253_43940# a_2455_43940# 0.092725f
C3004 a_n2946_38778# VDD 0.383009f
C3005 a_6491_46660# a_5257_43370# 0.1719f
C3006 a_20273_45572# VDD 0.571099f
C3007 a_327_44734# a_375_42282# 0.067169f
C3008 a_18597_46090# a_18819_46122# 0.230891f
C3009 a_6755_46942# a_12816_46660# 0.061031f
C3010 a_18989_43940# VDD 0.342796f
C3011 a_7871_42858# a_7765_42852# 0.379881f
C3012 a_1138_42852# a_167_45260# 0.250282f
C3013 a_1823_45246# a_2202_46116# 0.25354f
C3014 a_19123_46287# a_18819_46122# 0.172712f
C3015 a_5745_43940# VDD 0.144352f
C3016 a_20193_45348# a_22223_43948# 0.041425f
C3017 a_5807_45002# VDD 1.75047f
C3018 a_5111_44636# a_6031_43396# 0.207345f
C3019 a_12379_46436# a_12638_46436# 0.093752f
C3020 a_10518_42984# VDD 0.273357f
C3021 a_5495_43940# a_5745_43940# 0.014406f
C3022 a_3699_46348# VDD 0.208984f
C3023 a_11962_45724# a_12791_45546# 0.124167f
C3024 a_n2497_47436# a_n447_43370# 0.192476f
C3025 a_18479_47436# a_15493_43940# 0.05409f
C3026 a_7754_39964# a_7754_39632# 0.296522f
C3027 a_6491_46660# a_5807_45002# 0.01567f
C3028 a_15143_45578# VDD 0.12071f
C3029 C10_N_btm VCM 10.5945f
C3030 VDD VREF 4.8299f
C3031 a_18315_45260# VDD 0.12623f
C3032 a_9482_43914# a_10334_44484# 0.015932f
C3033 a_20202_43084# a_21487_43396# 0.019942f
C3034 a_18249_42858# a_18707_42852# 0.027606f
C3035 a_14311_47204# VDD 0.241476f
C3036 a_16112_44458# a_16241_44484# 0.010132f
C3037 a_13487_47204# RST_Z 0.07884f
C3038 a_1138_42852# a_n863_45724# 0.135594f
C3039 a_5807_45002# a_5691_45260# 0.19412f
C3040 a_8515_42308# a_8325_42308# 0.134955f
C3041 a_16867_43762# VDD 0.132317f
C3042 a_2998_44172# a_3499_42826# 0.027036f
C3043 a_11031_47542# a_9313_45822# 0.063846f
C3044 a_n2946_39072# a_n2946_38778# 0.050477f
C3045 a_20193_45348# a_20753_42852# 0.04748f
C3046 a_18691_45572# a_18787_45572# 0.013793f
C3047 CAL_N RST_Z 0.058301f
C3048 a_22589_40599# VDD 0.821011f
C3049 a_8128_46384# a_7411_46660# 0.019875f
C3050 EN_VIN_BSTR_P C8_P_btm 0.090252f
C3051 a_601_46902# a_948_46660# 0.051162f
C3052 a_n133_46660# a_288_46660# 0.086708f
C3053 a_13017_45260# VDD 0.263701f
C3054 a_21381_43940# a_21356_42826# 0.196864f
C3055 a_16977_43638# a_15743_43084# 0.042866f
C3056 a_16243_43396# a_16664_43396# 0.090164f
C3057 a_n2661_45010# a_n2433_44484# 0.217176f
C3058 a_13249_42308# a_14673_44172# 0.026424f
C3059 a_20916_46384# a_21137_46414# 0.118131f
C3060 a_19339_43156# a_19164_43230# 0.233657f
C3061 a_7227_42852# a_7309_42852# 0.171361f
C3062 a_19006_44850# VDD 0.077608f
C3063 a_626_44172# a_175_44278# 0.017096f
C3064 a_5807_45002# a_18479_45785# 0.174313f
C3065 a_13351_46090# a_13759_46122# 0.043782f
C3066 a_1184_42692# a_961_42354# 0.100246f
C3067 a_22165_42308# a_21613_42308# 0.027246f
C3068 a_n863_45724# a_1576_42282# 0.05148f
C3069 a_5066_45546# a_8568_45546# 0.04527f
C3070 a_n2497_47436# a_n809_44244# 0.029871f
C3071 a_n815_47178# a_n785_47204# 0.123817f
C3072 a_3726_37500# VDAC_N 0.06247f
C3073 a_9804_47204# a_5807_45002# 0.039093f
C3074 a_20107_45572# VDD 0.458237f
C3075 a_6709_45028# a_7705_45326# 0.099282f
C3076 a_12465_44636# a_13925_46122# 0.018086f
C3077 a_18597_46090# a_17957_46116# 0.018356f
C3078 a_6755_46942# a_12991_46634# 0.077634f
C3079 a_18374_44850# VDD 0.203584f
C3080 a_7227_42852# a_7765_42852# 0.118623f
C3081 a_1176_45822# a_167_45260# 0.091673f
C3082 a_16131_47204# VDD 0.142103f
C3083 a_11309_47204# CLK 0.01087f
C3084 a_20202_43084# a_20712_42282# 0.028679f
C3085 a_10083_42826# VDD 0.461256f
C3086 a_17973_43940# a_18079_43940# 0.419086f
C3087 a_n2497_47436# a_n1352_43396# 0.061218f
C3088 a_18597_46090# a_21115_43940# 0.015966f
C3089 a_22223_47212# a_22731_47423# 0.011229f
C3090 a_6545_47178# a_5807_45002# 0.030195f
C3091 a_n746_45260# a_383_46660# 0.011439f
C3092 a_14495_45572# VDD 0.238674f
C3093 a_10490_45724# CLK 0.029352f
C3094 C10_N_btm VREF_GND 10.3207f
C3095 C9_N_btm VCM 6.06251f
C3096 a_18597_46090# a_11415_45002# 0.061694f
C3097 VDD VIN_N 1.51335f
C3098 a_5167_46660# a_5275_47026# 0.057222f
C3099 a_3877_44458# a_5257_43370# 0.142219f
C3100 a_17719_45144# VDD 0.1297f
C3101 a_9482_43914# a_10157_44484# 0.321004f
C3102 a_626_44172# a_742_44458# 0.022141f
C3103 a_n2661_45010# a_556_44484# 0.038106f
C3104 a_13487_47204# VDD 0.273369f
C3105 a_9067_47204# DATA[4] 0.354356f
C3106 a_12594_46348# a_12638_46436# 0.049443f
C3107 a_6755_46942# a_16020_45572# 0.010518f
C3108 a_16664_43396# VDD 0.077608f
C3109 a_14513_46634# VDD 0.223375f
C3110 a_5343_44458# a_8147_43396# 0.014327f
C3111 a_9863_47436# a_9313_45822# 0.049145f
C3112 a_2351_42308# VDD 0.188239f
C3113 a_7499_43078# a_9482_43914# 0.062333f
C3114 CAL_N VDD 26.0839f
C3115 EN_VIN_BSTR_N a_19998_34978# 0.573018f
C3116 EN_VIN_BSTR_P C9_P_btm 0.226529f
C3117 a_33_46660# a_948_46660# 0.117156f
C3118 a_5807_45002# a_3877_44458# 0.034811f
C3119 a_11963_45334# VDD 0.229584f
C3120 a_16409_43396# a_15743_43084# 0.586918f
C3121 a_17499_43370# a_18429_43548# 0.012474f
C3122 a_6755_46942# a_11415_45002# 0.02226f
C3123 a_3877_44458# a_3699_46348# 0.084544f
C3124 a_20916_46384# a_20708_46348# 0.189941f
C3125 a_8387_43230# a_8483_43230# 0.013793f
C3126 a_18588_44850# VDD 0.132317f
C3127 a_16112_44458# a_14539_43914# 0.13299f
C3128 a_11827_44484# a_14815_43914# 0.029578f
C3129 a_22165_42308# a_21887_42336# 0.110763f
C3130 a_n863_45724# a_1067_42314# 0.289393f
C3131 a_5066_45546# a_8162_45546# 0.025437f
C3132 a_14976_45028# a_15415_45028# 0.027906f
C3133 a_n2497_47436# a_n1549_44318# 0.018493f
C3134 COMP_P a_22527_39145# 0.033008f
C3135 a_19328_44172# a_19741_43940# 0.04732f
C3136 a_20269_44172# a_19319_43548# 0.12985f
C3137 a_16375_45002# a_16751_45260# 0.047561f
C3138 a_n3690_38528# VDD 0.363159f
C3139 a_3726_37500# a_6886_37412# 0.702909f
C3140 a_8128_46384# a_5807_45002# 0.023925f
C3141 a_7229_43940# a_7705_45326# 0.203098f
C3142 a_12465_44636# a_13759_46122# 0.018063f
C3143 a_6755_46942# a_12251_46660# 0.033714f
C3144 a_18443_44721# VDD 0.193515f
C3145 a_n746_45260# a_n2293_45010# 0.023201f
C3146 a_18285_46348# a_17957_46116# 0.12677f
C3147 a_7499_43078# a_10796_42968# 0.030705f
C3148 a_20193_45348# a_21115_43940# 0.01963f
C3149 a_19466_46812# a_20273_45572# 0.328586f
C3150 a_5257_43370# a_5111_44636# 0.22597f
C3151 a_8952_43230# VDD 0.273404f
C3152 a_3147_46376# VDD 0.341038f
C3153 a_11962_45724# a_12427_45724# 0.064229f
C3154 a_n2497_47436# a_n1177_43370# 0.062743f
C3155 a_13249_42308# VDD 0.653917f
C3156 a_20512_43084# a_19987_42826# 0.11919f
C3157 a_8746_45002# CLK 0.018523f
C3158 a_17339_46660# a_15493_43940# 0.020994f
C3159 a_n2293_45010# a_n2109_45247# 0.068458f
C3160 C10_N_btm VREF 14.773f
C3161 C8_N_btm VCM 2.61094f
C3162 C9_N_btm VREF_GND 5.18245f
C3163 RST_Z CLK 0.064624f
C3164 a_18597_46090# a_20202_43084# 0.04177f
C3165 VDD VIN_P 1.52779f
C3166 a_5167_46660# a_5072_46660# 0.049827f
C3167 a_5907_46634# a_6540_46812# 0.017547f
C3168 a_5385_46902# a_5275_47026# 0.097745f
C3169 a_5807_45002# a_19466_46812# 0.178376f
C3170 a_15095_43370# a_15567_42826# 0.167909f
C3171 a_17613_45144# VDD 0.094022f
C3172 a_9482_43914# a_9838_44484# 0.175591f
C3173 a_8953_45546# a_9885_43646# 0.011162f
C3174 a_n1441_43940# VDD 0.142719f
C3175 a_6575_47204# DATA[4] 0.15718f
C3176 a_5807_45002# a_5111_44636# 0.204193f
C3177 a_12594_46348# a_12379_46436# 0.04209f
C3178 a_19700_43370# VDD 0.28578f
C3179 a_18579_44172# a_15493_43940# 0.377126f
C3180 a_14180_46812# VDD 0.755623f
C3181 a_2675_43914# a_3499_42826# 0.010775f
C3182 a_9067_47204# a_9313_45822# 0.013659f
C3183 a_2123_42473# VDD 0.1936f
C3184 a_310_45028# VDD 0.360949f
C3185 EN_VIN_BSTR_N a_19250_34978# 0.651142f
C3186 EN_VIN_BSTR_P C10_P_btm 0.320569f
C3187 a_33_46660# a_1123_46634# 0.041798f
C3188 a_601_46902# a_383_46660# 0.209641f
C3189 VDAC_P RST_Z 0.158793f
C3190 a_11787_45002# VDD 0.153399f
C3191 a_16547_43609# a_15743_43084# 0.028834f
C3192 a_17499_43370# a_17324_43396# 0.234322f
C3193 a_16292_46812# a_16388_46812# 0.318472f
C3194 a_5755_42852# a_5837_42852# 0.171361f
C3195 a_8387_43230# a_8292_43218# 0.049827f
C3196 a_18817_42826# a_19164_43230# 0.051162f
C3197 a_1823_45246# a_4649_42852# 0.042816f
C3198 a_375_42282# a_175_44278# 0.017991f
C3199 a_17339_46660# a_16375_45002# 0.0296f
C3200 a_1208_46090# a_1431_46436# 0.011458f
C3201 a_n473_42460# a_n327_42308# 0.013377f
C3202 a_1067_42314# a_961_42354# 0.13675f
C3203 a_1576_42282# a_1184_42692# 0.033078f
C3204 a_5883_43914# a_7499_43940# 0.04798f
C3205 a_14976_45028# a_14797_45144# 0.137651f
C3206 a_11415_45002# a_22223_45572# 0.021019f
C3207 a_n452_47436# a_n746_45260# 0.187792f
C3208 a_8495_42852# VDD 0.132018f
C3209 a_19862_44208# a_19319_43548# 0.049274f
C3210 a_3065_45002# a_3823_42558# 0.198186f
C3211 a_5257_43370# a_3905_42865# 0.106385f
C3212 a_3316_45546# a_3429_45260# 0.142842f
C3213 a_20974_43370# a_22591_43396# 0.046632f
C3214 a_15861_45028# a_16237_45028# 0.062212f
C3215 a_7229_43940# a_6709_45028# 0.136786f
C3216 a_6755_46942# a_12469_46902# 0.042969f
C3217 a_18287_44626# VDD 0.389383f
C3218 a_n2497_47436# a_n967_45348# 0.021003f
C3219 a_1799_45572# a_1609_45822# 0.079527f
C3220 a_18285_46348# a_18189_46348# 0.118603f
C3221 a_12891_46348# a_12791_45546# 0.012918f
C3222 a_11309_47204# DATA[5] 0.080873f
C3223 a_7499_43078# a_10835_43094# 0.028158f
C3224 a_20193_45348# a_20935_43940# 0.016238f
C3225 a_19466_46812# a_20107_45572# 0.283769f
C3226 a_5257_43370# a_5147_45002# 0.836149f
C3227 a_9127_43156# VDD 0.468721f
C3228 a_15959_42545# a_16522_42674# 0.049827f
C3229 a_15890_42674# a_16104_42674# 0.097745f
C3230 a_17737_43940# a_17973_43940# 0.22264f
C3231 a_5013_44260# a_5025_43940# 0.011829f
C3232 a_2804_46116# VDD 0.159351f
C3233 a_14539_43914# a_16759_43396# 0.012597f
C3234 a_20202_43084# a_20193_45348# 0.116706f
C3235 a_n2497_47436# a_n1917_43396# 0.012526f
C3236 a_n746_45260# a_33_46660# 0.035747f
C3237 a_17124_42282# VDD 0.28176f
C3238 a_12465_44636# a_22223_47212# 0.175138f
C3239 a_13904_45546# VDD 0.135068f
C3240 C9_N_btm VREF 7.369471f
C3241 C10_N_btm VIN_N 3.66034f
C3242 RST_Z EN_OFFSET_CAL 0.044122f
C3243 C7_N_btm VCM 1.58335f
C3244 C8_N_btm VREF_GND 2.58605f
C3245 VDD CLK 0.49309f
C3246 a_18479_47436# a_11415_45002# 0.033153f
C3247 a_4817_46660# a_5275_47026# 0.031068f
C3248 a_5907_46634# a_5732_46660# 0.233657f
C3249 a_17023_45118# VDD 0.086861f
C3250 a_1847_42826# a_2351_42308# 0.120686f
C3251 a_16979_44734# a_17061_44734# 0.171361f
C3252 a_6575_47204# DATA[3] 0.055018f
C3253 a_n2497_47436# a_n1917_44484# 0.011319f
C3254 a_6755_46942# a_15861_45028# 0.033041f
C3255 a_5807_45002# a_5147_45002# 0.035651f
C3256 a_376_46348# a_380_45546# 0.011689f
C3257 a_12005_46116# a_12379_46436# 0.038694f
C3258 a_19268_43646# VDD 0.237793f
C3259 a_14035_46660# VDD 0.363878f
C3260 a_6575_47204# a_9313_45822# 0.017088f
C3261 a_1755_42282# VDD 0.215277f
C3262 a_22485_44484# a_22591_43396# 0.025074f
C3263 a_n1099_45572# VDD 0.89411f
C3264 VDAC_P VDD 5.18919f
C3265 a_15811_47375# a_16292_46812# 0.080078f
C3266 a_n133_46660# a_948_46660# 0.102355f
C3267 a_33_46660# a_383_46660# 0.20669f
C3268 a_10951_45334# VDD 0.226705f
C3269 a_16243_43396# a_15743_43084# 0.600668f
C3270 a_18479_45785# a_18287_44626# 0.024431f
C3271 a_18249_42858# a_19164_43230# 0.118759f
C3272 a_1208_46090# a_1337_46436# 0.010132f
C3273 a_1067_42314# a_1184_42692# 0.147283f
C3274 a_22485_44484# a_22591_44484# 0.15878f
C3275 a_5883_43914# a_6671_43940# 0.051304f
C3276 a_n2497_47436# a_n1899_43946# 0.040963f
C3277 a_14976_45028# a_14537_43396# 0.087031f
C3278 a_1241_43940# a_1443_43940# 0.092725f
C3279 a_3065_45002# a_3318_42354# 0.146272f
C3280 a_3316_45546# a_3065_45002# 0.141454f
C3281 a_16375_45002# a_16019_45002# 0.032313f
C3282 a_n4334_38528# VDD 0.385889f
C3283 a_7276_45260# a_6709_45028# 0.215102f
C3284 a_16147_45260# a_17719_45144# 0.049848f
C3285 a_6755_46942# a_11901_46660# 0.587021f
C3286 a_18248_44752# VDD 0.251171f
C3287 a_n863_45724# a_n1557_42282# 0.034373f
C3288 a_14537_43396# a_15433_44458# 0.018743f
C3289 a_n746_45260# a_n2661_45010# 0.400342f
C3290 a_1176_45822# a_1138_42852# 0.41217f
C3291 a_3737_43940# VDD 0.18423f
C3292 a_12089_42308# a_12563_42308# 0.03299f
C3293 a_18479_45785# a_19268_43646# 0.12682f
C3294 a_8953_45546# a_9885_42558# 0.024699f
C3295 a_7499_43078# a_10518_42984# 0.03265f
C3296 a_11827_44484# a_15493_43940# 0.010315f
C3297 a_20193_45348# a_20623_43914# 0.048456f
C3298 a_8387_43230# VDD 0.200672f
C3299 a_15959_42545# a_16104_42674# 0.057222f
C3300 a_15803_42450# a_16522_42674# 0.089677f
C3301 a_14539_43914# a_16977_43638# 0.013865f
C3302 a_22485_44484# a_20974_43370# 0.101193f
C3303 a_2698_46116# VDD 0.195879f
C3304 a_n2497_47436# a_n1699_43638# 0.038204f
C3305 a_18479_47436# a_20935_43940# 0.207572f
C3306 a_11415_45002# a_19113_45348# 0.012208f
C3307 a_n746_45260# a_171_46873# 0.120194f
C3308 a_16522_42674# VDD 0.077608f
C3309 a_11459_47204# a_11309_47204# 0.183357f
C3310 a_21811_47423# a_22223_47212# 0.031065f
C3311 a_13527_45546# VDD 0.1902f
C3312 a_10180_45724# CLK 0.095799f
C3313 a_n2661_45010# a_n2109_45247# 0.025907f
C3314 a_n2472_45002# a_n2293_45010# 0.177252f
C3315 C8_N_btm VREF 3.6701f
C3316 C9_N_btm VIN_N 1.82823f
C3317 C7_N_btm VREF_GND 1.61142f
C3318 C6_N_btm VCM 0.877241f
C3319 VDD EN_OFFSET_CAL 0.489629f
C3320 a_18479_47436# a_20202_43084# 0.040227f
C3321 a_4817_46660# a_5072_46660# 0.06121f
C3322 a_15095_43370# a_15279_43071# 0.105784f
C3323 a_12281_43396# a_12545_42858# 0.029151f
C3324 a_16922_45042# VDD 1.54713f
C3325 a_14539_43914# a_17061_44734# 0.020462f
C3326 a_7903_47542# DATA[3] 0.01066f
C3327 a_n2497_47436# a_n1699_44726# 0.012807f
C3328 a_15743_43084# VDD 0.572249f
C3329 a_13885_46660# VDD 0.499249f
C3330 a_1169_39043# comp_n 0.3874f
C3331 a_n3690_39392# a_n3690_38528# 0.050585f
C3332 a_10807_43548# a_10695_43548# 0.159782f
C3333 a_380_45546# VDD 0.154763f
C3334 a_8746_45002# a_8953_45002# 0.257529f
C3335 a_15811_47375# a_15559_46634# 0.018669f
C3336 a_n133_46660# a_1123_46634# 0.043619f
C3337 a_33_46660# a_601_46902# 0.17072f
C3338 VDAC_N RST_Z 0.154233f
C3339 a_10775_45002# VDD 0.148349f
C3340 a_16977_43638# a_17324_43396# 0.051162f
C3341 a_16137_43396# a_15743_43084# 0.029757f
C3342 a_n2840_45002# a_n2840_44458# 0.025171f
C3343 a_15559_46634# a_13059_46348# 0.167936f
C3344 a_8037_42858# a_8292_43218# 0.064178f
C3345 a_18817_42826# a_18599_43230# 0.209641f
C3346 a_18249_42858# a_19339_43156# 0.042415f
C3347 a_5111_42852# a_5193_42852# 0.171361f
C3348 a_12005_46116# a_12594_46348# 0.065075f
C3349 a_3539_42460# VDD 0.363092f
C3350 a_1067_42314# a_1576_42282# 0.017282f
C3351 a_n2497_47436# a_n1761_44111# 0.045728f
C3352 a_11415_45002# a_21513_45002# 0.050445f
C3353 COMP_P a_22537_40625# 0.120662f
C3354 a_2382_45260# a_3823_42558# 0.058499f
C3355 a_3316_45546# a_2680_45002# 0.050127f
C3356 a_20974_43370# a_22223_43396# 0.04256f
C3357 a_5205_44484# a_6709_45028# 0.095031f
C3358 a_7276_45260# a_7229_43940# 0.322065f
C3359 a_16147_45260# a_17613_45144# 0.028566f
C3360 a_18479_45785# a_16922_45042# 0.02321f
C3361 a_6755_46942# a_11813_46116# 0.028837f
C3362 a_17970_44736# VDD 0.27753f
C3363 a_10440_44484# CLK 0.013272f
C3364 a_1823_45246# a_4520_42826# 0.053569f
C3365 a_14537_43396# a_14815_43914# 0.015948f
C3366 a_17339_46660# a_17957_46116# 0.098952f
C3367 a_1208_46090# a_1138_42852# 0.043831f
C3368 a_20202_43084# a_19511_42282# 0.082529f
C3369 a_7499_43078# a_10083_42826# 0.375624f
C3370 a_20193_45348# a_20365_43914# 0.025746f
C3371 a_5204_45822# a_4880_45572# 0.046074f
C3372 a_8605_42826# VDD 0.204898f
C3373 a_15764_42576# a_16522_42674# 0.05936f
C3374 a_14539_43914# a_16409_43396# 0.031761f
C3375 a_20512_43084# a_20974_43370# 0.020132f
C3376 a_2521_46116# VDD 0.163553f
C3377 a_n2497_47436# a_n2267_43396# 0.222725f
C3378 a_18479_47436# a_20623_43914# 0.012705f
C3379 a_11322_45546# a_12427_45724# 0.010517f
C3380 a_11525_45546# a_11962_45724# 0.095856f
C3381 a_n746_45260# a_n133_46660# 0.042075f
C3382 a_16104_42674# VDD 0.134357f
C3383 a_9313_45822# a_11309_47204# 0.027145f
C3384 a_13163_45724# VDD 0.322298f
C3385 a_n2661_45010# a_n2293_45010# 0.400159f
C3386 C7_N_btm VREF 1.818f
C3387 C8_N_btm VIN_N 0.907642f
C3388 C6_N_btm VREF_GND 0.836236f
C3389 C5_N_btm VCM 0.719982f
C3390 VDD DATA[5] 0.504354f
C3391 a_5385_46902# a_5732_46660# 0.051162f
C3392 a_4955_46873# a_5072_46660# 0.17431f
C3393 a_12281_43396# a_12089_42308# 0.210903f
C3394 a_10775_45002# a_10057_43914# 0.010331f
C3395 a_17339_46660# a_11415_45002# 0.025523f
C3396 a_6755_46942# a_15682_46116# 0.116442f
C3397 a_13381_47204# VDD 0.130765f
C3398 a_9482_43914# a_11173_44260# 0.043729f
C3399 a_7227_47204# DATA[3] 0.357377f
C3400 a_n2497_47436# a_n2267_44484# 0.025633f
C3401 a_18783_43370# VDD 0.289099f
C3402 a_19279_43940# a_15493_43940# 0.019758f
C3403 a_5257_43370# a_5883_43914# 0.019234f
C3404 a_n2302_39072# a_n2216_39072# 0.011479f
C3405 a_20193_45348# a_22400_42852# 0.05078f
C3406 a_21381_43940# a_20974_43370# 0.02221f
C3407 a_n452_45724# VDD 0.112977f
C3408 a_10180_45724# a_10775_45002# 0.073185f
C3409 a_15507_47210# a_15559_46634# 0.011624f
C3410 VDAC_N VDD 4.61811f
C3411 a_n133_46660# a_383_46660# 0.105995f
C3412 a_6886_37412# RST_Z 0.031637f
C3413 a_8953_45002# VDD 1.24336f
C3414 a_16409_43396# a_17324_43396# 0.118759f
C3415 a_15368_46634# a_13059_46348# 0.101997f
C3416 a_18249_42858# a_18599_43230# 0.210876f
C3417 a_7765_42852# a_8292_43218# 0.157652f
C3418 a_18083_42858# a_19164_43230# 0.101963f
C3419 a_2382_45260# a_3499_42826# 0.040227f
C3420 a_7229_43940# a_7542_44172# 0.086946f
C3421 a_5275_47026# VDD 0.135766f
C3422 a_n2497_47436# a_n2065_43946# 0.036632f
C3423 a_20202_43084# a_21513_45002# 0.13666f
C3424 COMP_P a_22589_40599# 0.204694f
C3425 a_n815_47178# a_n452_47436# 0.107449f
C3426 a_2981_46116# VDD 0.111597f
C3427 a_18451_43940# a_18533_43940# 0.171361f
C3428 a_19328_44172# a_19319_43548# 0.033025f
C3429 a_2382_45260# a_3318_42354# 0.028613f
C3430 a_20193_45348# a_22223_42860# 0.017179f
C3431 a_3316_45546# a_2382_45260# 0.052075f
C3432 a_2112_39137# VDD 0.28506f
C3433 a_6431_45366# a_6709_45028# 0.112564f
C3434 a_16147_45260# a_17023_45118# 0.040001f
C3435 a_6755_46942# a_11735_46660# 0.61229f
C3436 a_17767_44458# VDD 0.348803f
C3437 a_21487_43396# a_21195_42852# 0.01192f
C3438 a_10334_44484# CLK 0.012484f
C3439 a_17339_46660# a_18189_46348# 0.170772f
C3440 a_1208_46090# a_1176_45822# 0.141891f
C3441 a_12089_42308# a_11551_42558# 0.109508f
C3442 a_7499_43078# a_8952_43230# 0.054554f
C3443 a_8037_42858# VDD 0.344922f
C3444 a_15764_42576# a_16104_42674# 0.029366f
C3445 a_167_45260# VDD 1.41955f
C3446 a_14539_43914# a_16547_43609# 0.01221f
C3447 a_n2497_47436# a_n2129_43609# 0.216536f
C3448 a_18597_46090# a_19862_44208# 0.536021f
C3449 a_11525_45546# a_11652_45724# 0.138143f
C3450 a_11322_45546# a_11962_45724# 0.270736f
C3451 a_10490_45724# a_12427_45724# 0.108721f
C3452 a_11415_45002# a_22223_45036# 0.011148f
C3453 a_11031_47542# a_11309_47204# 0.110775f
C3454 a_3754_39964# VDAC_Pi 0.296508f
C3455 a_12791_45546# VDD 0.205486f
C3456 a_4699_43561# a_3539_42460# 0.109444f
C3457 a_n2661_45010# a_n2472_45002# 0.065751f
C3458 a_15861_45028# a_16751_45260# 0.044248f
C3459 C6_N_btm VREF 1.41944f
C3460 C7_N_btm VIN_N 1.52449f
C3461 C5_N_btm VREF_GND 0.676559f
C3462 C4_N_btm VCM 0.716447f
C3463 VDD DATA[4] 0.326957f
C3464 a_4651_46660# a_5072_46660# 0.083408f
C3465 a_4817_46660# a_5732_46660# 0.118759f
C3466 a_12281_43396# a_12379_42858# 0.036584f
C3467 a_327_44734# a_n23_44458# 0.141544f
C3468 a_9482_43914# a_10555_44260# 0.088693f
C3469 a_n863_45724# a_2905_42968# 0.269475f
C3470 a_16112_44458# a_16241_44734# 0.062574f
C3471 a_14539_43914# a_14673_44172# 0.205935f
C3472 a_6851_47204# DATA[3] 0.146601f
C3473 a_11459_47204# VDD 0.34771f
C3474 a_n2497_47436# a_n2129_44697# 0.019202f
C3475 a_18525_43370# VDD 0.263553f
C3476 a_7542_44172# a_7845_44172# 0.137004f
C3477 a_19466_46812# a_16922_45042# 0.030378f
C3478 a_6575_47204# a_9067_47204# 0.210614f
C3479 a_n863_45724# VDD 1.89058f
C3480 a_18691_45572# a_18799_45938# 0.057222f
C3481 a_10180_45724# a_8953_45002# 0.107499f
C3482 a_6886_37412# VDD 0.235486f
C3483 a_171_46873# a_33_46660# 0.207108f
C3484 a_n133_46660# a_601_46902# 0.053479f
C3485 a_8191_45002# VDD 0.39677f
C3486 a_16977_43638# a_16759_43396# 0.209641f
C3487 a_16409_43396# a_17499_43370# 0.042737f
C3488 a_14976_45028# a_13059_46348# 0.209989f
C3489 a_15368_46634# a_15227_46910# 0.050747f
C3490 a_18249_42858# a_18817_42826# 0.16939f
C3491 a_18083_42858# a_19339_43156# 0.042271f
C3492 a_7871_42858# a_8292_43218# 0.086377f
C3493 a_4520_42826# a_4649_42852# 0.062574f
C3494 a_7229_43940# a_7281_43914# 0.164835f
C3495 a_3540_43646# VDD 0.209044f
C3496 a_5072_46660# VDD 0.081835f
C3497 a_5066_45546# a_4880_45572# 0.04794f
C3498 a_7309_42852# VDD 0.177437f
C3499 a_22775_42308# a_22485_38105# 0.330766f
C3500 a_20193_45348# a_22165_42308# 0.252856f
C3501 a_16147_45260# a_16922_45042# 0.016249f
C3502 a_6755_46942# a_11186_47026# 0.014167f
C3503 a_16979_44734# VDD 0.256327f
C3504 a_13556_45296# a_15433_44458# 0.1084f
C3505 a_17339_46660# a_17715_44484# 0.018672f
C3506 a_805_46414# a_1176_45822# 0.024739f
C3507 a_472_46348# a_1138_42852# 0.028956f
C3508 a_2455_43940# VDD 0.144352f
C3509 a_9804_47204# DATA[4] 0.015379f
C3510 a_7499_43078# a_9127_43156# 0.08498f
C3511 a_8953_45546# a_9803_42558# 0.031932f
C3512 a_20193_45348# a_19862_44208# 0.041264f
C3513 a_7765_42852# VDD 0.333322f
C3514 a_2202_46116# VDD 0.20904f
C3515 a_14539_43914# a_16243_43396# 0.029808f
C3516 a_20512_43084# a_21381_43940# 0.019564f
C3517 a_3600_43914# a_3992_43940# 0.016359f
C3518 a_n2497_47436# a_n2433_43396# 0.173242f
C3519 a_11322_45546# a_11652_45724# 0.26844f
C3520 a_10490_45724# a_11962_45724# 0.114064f
C3521 a_11415_45002# a_11827_44484# 0.169126f
C3522 C5_N_btm VREF 0.987144f
C3523 C6_N_btm VIN_N 0.391905f
C3524 VDD DATA[3] 0.309692f
C3525 C4_N_btm VREF_GND 0.671882f
C3526 C3_N_btm VCM 0.716273f
C3527 a_4817_46660# a_5907_46634# 0.042415f
C3528 a_5385_46902# a_5167_46660# 0.209641f
C3529 a_5807_45002# a_16292_46812# 0.202526f
C3530 a_14579_43548# a_15279_43071# 0.108607f
C3531 a_6755_46942# a_14840_46494# 0.021842f
C3532 a_20623_46660# a_20731_47026# 0.057222f
C3533 a_n1644_44306# VDD 0.082968f
C3534 a_16112_44458# a_14673_44172# 0.077293f
C3535 a_6491_46660# DATA[3] 0.011549f
C3536 a_9313_45822# VDD 0.5747f
C3537 a_n2497_47436# a_n2433_44484# 0.027254f
C3538 a_18429_43548# VDD 0.163446f
C3539 a_2127_44172# a_2253_44260# 0.013015f
C3540 a_1414_42308# a_3499_42826# 0.023314f
C3541 a_961_42354# VDD 0.091526f
C3542 a_n1079_45724# VDD 0.172275f
C3543 a_18691_45572# a_18596_45572# 0.049827f
C3544 a_18909_45814# a_18799_45938# 0.097745f
C3545 a_19431_45546# a_19256_45572# 0.233657f
C3546 VDAC_N C10_N_btm 0.883474p
C3547 a_n133_46660# a_33_46660# 0.580914f
C3548 a_7705_45326# VDD 0.211554f
C3549 a_16409_43396# a_16759_43396# 0.20669f
C3550 a_16243_43396# a_17324_43396# 0.102355f
C3551 a_1823_45246# a_4905_42826# 0.110836f
C3552 a_14976_45028# a_15227_46910# 0.060892f
C3553 a_18083_42858# a_18599_43230# 0.113784f
C3554 a_6540_46812# VDD 0.084698f
C3555 a_5837_42852# VDD 0.1774f
C3556 a_21613_42308# a_22485_38105# 0.026117f
C3557 a_3905_42865# a_3539_42460# 0.022817f
C3558 a_6491_46660# a_6540_46812# 0.079263f
C3559 a_20974_43370# a_21855_43396# 0.029556f
C3560 a_18597_46090# a_21195_42852# 0.01512f
C3561 a_10249_46116# a_11186_47026# 0.172467f
C3562 a_14539_43914# VDD 0.873589f
C3563 a_4520_42826# a_5111_42852# 0.047152f
C3564 a_13556_45296# a_14815_43914# 0.378519f
C3565 a_9482_43914# a_15433_44458# 0.20244f
C3566 a_472_46348# a_1176_45822# 0.146555f
C3567 a_2253_43940# VDD 0.156797f
C3568 a_8953_45546# a_9223_42460# 0.166987f
C3569 a_11415_45002# a_10907_45822# 0.050963f
C3570 a_7871_42858# VDD 0.395222f
C3571 a_14113_42308# a_16522_42674# 0.183181f
C3572 a_1823_45246# VDD 1.7584f
C3573 a_3600_43914# a_3737_43940# 0.126609f
C3574 a_18479_47436# a_19862_44208# 0.138185f
C3575 a_11322_45546# a_11525_45546# 0.055031f
C3576 a_10490_45724# a_11652_45724# 0.044431f
C3577 a_20202_43084# a_11827_44484# 0.032881f
C3578 a_11415_45002# a_21359_45002# 0.015551f
C3579 a_9313_45822# a_9804_47204# 0.171044f
C3580 a_12427_45724# VDD 0.33808f
C3581 a_458_43396# a_648_43396# 0.045837f
C3582 a_15861_45028# a_16019_45002# 0.04712f
C3583 a_n2840_45002# a_n2661_45010# 0.189331f
C3584 VDD DATA[2] 0.3216f
C3585 C4_N_btm VREF 0.98728f
C3586 C5_N_btm VIN_N 0.502041f
C3587 C3_N_btm VREF_GND 0.67174f
C3588 C2_N_btm VCM 0.716172f
C3589 a_21811_47423# a_21363_46634# 0.010128f
C3590 a_3877_44458# a_5072_46660# 0.021873f
C3591 a_4651_46660# a_5732_46660# 0.102355f
C3592 a_4817_46660# a_5167_46660# 0.218775f
C3593 a_14309_45028# VDD 0.189806f
C3594 a_4905_42826# a_5193_42852# 0.016389f
C3595 a_20556_43646# a_20749_43396# 0.018955f
C3596 a_6755_46942# a_15015_46420# 0.133517f
C3597 a_20841_46902# a_20731_47026# 0.097745f
C3598 a_21363_46634# a_22000_46634# 0.017308f
C3599 a_20623_46660# a_20528_46660# 0.049827f
C3600 a_17595_43084# a_17749_42852# 0.010303f
C3601 a_n863_45724# a_1847_42826# 0.216819f
C3602 a_15004_44636# a_14673_44172# 0.039287f
C3603 a_6545_47178# DATA[3] 0.178561f
C3604 a_11031_47542# VDD 0.214104f
C3605 a_n1853_46287# a_n1099_45572# 0.067343f
C3606 a_17324_43396# VDD 0.274722f
C3607 a_7281_43914# a_7542_44172# 0.060549f
C3608 a_1184_42692# VDD 0.813074f
C3609 a_n2946_39072# a_n2860_39072# 0.011479f
C3610 a_n4334_39392# a_n4334_38528# 0.050585f
C3611 a_7903_47542# a_6575_47204# 0.046223f
C3612 a_18341_45572# a_18799_45938# 0.027606f
C3613 a_9049_44484# a_8953_45002# 0.031391f
C3614 VDAC_N C9_N_btm 0.44188p
C3615 a_n133_46660# a_171_46873# 0.163873f
C3616 a_6709_45028# VDD 0.390566f
C3617 a_16243_43396# a_17499_43370# 0.043633f
C3618 a_16409_43396# a_16977_43638# 0.17072f
C3619 a_15781_43660# a_15743_43084# 0.050751f
C3620 a_15009_46634# a_13059_46348# 0.054389f
C3621 a_17333_42852# a_18249_42858# 0.311255f
C3622 a_18083_42858# a_18817_42826# 0.0532f
C3623 a_7227_42852# a_7573_43172# 0.013377f
C3624 a_2896_43646# VDD 0.208317f
C3625 a_5732_46660# VDD 0.277366f
C3626 a_12891_46348# a_13076_44458# 0.182315f
C3627 a_5193_42852# VDD 0.187605f
C3628 a_18451_43940# a_18797_44260# 0.013377f
C3629 a_17715_44484# a_11827_44484# 0.037803f
C3630 comp_n VDD 0.504807f
C3631 a_6545_47178# a_6540_46812# 0.013617f
C3632 a_18799_45938# VDD 0.132317f
C3633 a_6431_45366# a_5205_44484# 0.018787f
C3634 a_10249_46116# a_10768_47026# 0.027091f
C3635 a_16112_44458# VDD 0.182397f
C3636 a_14579_43548# a_14635_42282# 0.124652f
C3637 a_9482_43914# a_14815_43914# 0.024524f
C3638 a_472_46348# a_1208_46090# 0.088629f
C3639 a_1443_43940# VDD 0.144342f
C3640 a_15928_47570# VDD 0.08228f
C3641 a_7499_43078# a_8605_42826# 0.026478f
C3642 a_8199_44636# a_9803_42558# 0.036259f
C3643 a_18494_42460# a_15493_43940# 0.02195f
C3644 a_4419_46090# a_4880_45572# 0.032829f
C3645 a_7227_42852# VDD 0.254613f
C3646 a_1138_42852# VDD 0.397518f
C3647 a_10490_45724# a_11525_45546# 0.06936f
C3648 a_11415_45002# a_21101_45002# 0.018873f
C3649 a_2113_38308# VDAC_Pi 0.170941f
C3650 a_9313_45822# a_8128_46384# 0.013269f
C3651 a_11962_45724# VDD 0.210594f
C3652 a_15861_45028# a_15595_45028# 0.072432f
C3653 C3_N_btm VREF 0.984942f
C3654 C4_N_btm VIN_N 0.50261f
C3655 C2_N_btm VREF_GND 0.671742f
C3656 C1_N_btm VCM 0.716121f
C3657 a_4817_46660# a_5385_46902# 0.170485f
C3658 a_4651_46660# a_5907_46634# 0.043482f
C3659 a_3877_44458# a_6540_46812# 0.244975f
C3660 a_5807_45002# a_15368_46634# 0.029781f
C3661 VDD DATA[1] 0.321585f
C3662 a_14579_43548# a_14543_43071# 0.032593f
C3663 a_21363_46634# a_21188_46660# 0.233657f
C3664 a_20273_46660# a_20731_47026# 0.027606f
C3665 a_17595_43084# a_17665_42852# 0.011552f
C3666 a_n863_45724# a_791_42968# 0.338631f
C3667 a_9863_47436# VDD 0.207794f
C3668 a_6755_46942# a_15765_45572# 0.026052f
C3669 a_15368_46634# a_15143_45578# 0.105334f
C3670 a_17499_43370# VDD 0.453381f
C3671 a_11415_45002# a_14797_45144# 0.021281f
C3672 a_5257_43370# a_5518_44484# 0.095452f
C3673 a_7227_47204# a_6575_47204# 0.028925f
C3674 a_1576_42282# VDD 0.26017f
C3675 a_20512_43084# a_21855_43396# 0.013929f
C3676 a_20202_43084# a_19279_43940# 0.020761f
C3677 a_18909_45814# a_19256_45572# 0.051162f
C3678 a_18341_45572# a_18596_45572# 0.056391f
C3679 VDAC_N C8_N_btm 0.220913p
C3680 EN_VIN_BSTR_P a_n217_35014# 0.651142f
C3681 a_3726_37500# RST_Z 1.60318f
C3682 a_7229_43940# VDD 0.821851f
C3683 a_16243_43396# a_16759_43396# 0.106647f
C3684 a_15009_46634# a_15227_46910# 0.08213f
C3685 a_3877_44458# a_1823_45246# 0.231164f
C3686 a_18083_42858# a_18249_42858# 0.699797f
C3687 a_12607_44458# a_13720_44458# 0.122704f
C3688 a_12883_44458# a_13076_44458# 0.142643f
C3689 a_16388_46812# a_16375_45002# 0.039999f
C3690 a_5907_46634# VDD 0.341121f
C3691 a_12891_46348# a_12883_44458# 0.018059f
C3692 a_4649_42852# VDD 0.194775f
C3693 SMPL_ON_P a_n1605_47204# 0.194856f
C3694 a_19321_45002# a_15493_43940# 0.050579f
C3695 a_8530_39574# CAL_N 0.644218f
C3696 a_18596_45572# VDD 0.077608f
C3697 a_18597_46090# a_20922_43172# 0.021228f
C3698 a_20916_46384# a_20202_43084# 0.181561f
C3699 a_10467_46802# a_11735_46660# 0.096658f
C3700 a_10554_47026# a_10768_47026# 0.097745f
C3701 a_10623_46897# a_11186_47026# 0.049827f
C3702 a_15004_44636# VDD 0.090175f
C3703 a_3935_42891# a_4520_42826# 0.017436f
C3704 a_13556_45296# a_13857_44734# 0.01375f
C3705 a_472_46348# a_805_46414# 0.360492f
C3706 a_1241_43940# VDD 0.162129f
C3707 a_8199_44636# a_9223_42460# 0.065156f
C3708 a_8953_45546# a_8685_42308# 0.250058f
C3709 a_7499_43078# a_8037_42858# 0.160087f
C3710 a_5755_42852# VDD 0.179985f
C3711 a_1176_45822# VDD 0.781481f
C3712 a_10490_45724# a_11322_45546# 0.246478f
C3713 a_11415_45002# a_21005_45260# 0.01592f
C3714 a_9863_47436# a_9804_47204# 0.109361f
C3715 a_11652_45724# VDD 0.155048f
C3716 C2_N_btm VREF 0.987884f
C3717 C1_N_btm VREF_GND 0.673422f
C3718 C0_N_btm VCM 0.717064f
C3719 a_4651_46660# a_5167_46660# 0.102946f
C3720 a_3877_44458# a_5732_46660# 0.040487f
C3721 a_5807_45002# a_14976_45028# 0.026261f
C3722 VDD DATA[0] 1.05526f
C3723 C3_N_btm VIN_N 0.455045f
C3724 a_8953_45546# a_9803_43646# 0.091141f
C3725 a_n467_45028# a_n23_44458# 0.038286f
C3726 a_8953_45002# a_9838_44484# 0.013986f
C3727 a_9313_45822# a_9049_44484# 0.119007f
C3728 a_18285_46348# a_18280_46660# 0.089884f
C3729 a_20273_46660# a_20528_46660# 0.056391f
C3730 a_7845_44172# VDD 0.11772f
C3731 a_18599_43230# a_18695_43230# 0.013793f
C3732 a_n863_45724# a_685_42968# 0.052365f
C3733 a_9067_47204# VDD 0.47483f
C3734 a_6755_46942# a_15903_45785# 0.192397f
C3735 a_n1853_46287# a_n452_45724# 0.080546f
C3736 a_16759_43396# VDD 0.191873f
C3737 a_18579_44172# a_19862_44208# 0.091151f
C3738 a_11415_45002# a_14537_43396# 0.04406f
C3739 a_5257_43370# a_5343_44458# 0.063407f
C3740 a_3218_45724# a_3260_45572# 0.010055f
C3741 a_6851_47204# a_6575_47204# 0.027563f
C3742 a_1067_42314# VDD 0.128996f
C3743 a_n2472_45546# VDD 0.290266f
C3744 a_18341_45572# a_19256_45572# 0.116691f
C3745 a_18479_45785# a_18596_45572# 0.183223f
C3746 a_3726_37500# VDD 0.341303f
C3747 VDAC_N C7_N_btm 0.11042p
C3748 a_7276_45260# VDD 0.093163f
C3749 a_16547_43609# a_16409_43396# 0.206231f
C3750 a_16243_43396# a_16977_43638# 0.053479f
C3751 a_4905_42826# a_5111_42852# 0.105155f
C3752 a_1823_45246# a_4235_43370# 0.029154f
C3753 a_19321_45002# a_18985_46122# 0.019556f
C3754 a_18083_42858# a_17333_42852# 0.284837f
C3755 a_12607_44458# a_13076_44458# 0.200168f
C3756 a_22315_44484# a_22485_44484# 0.109468f
C3757 a_5167_46660# VDD 0.203378f
C3758 a_7499_43078# a_7309_42852# 0.011818f
C3759 a_12891_46348# a_12607_44458# 0.067773f
C3760 a_n2497_47436# a_n746_45260# 0.046973f
C3761 a_22223_46124# EN_OFFSET_CAL 0.011048f
C3762 a_13904_45546# a_14127_45572# 0.011458f
C3763 a_1169_39043# VDD 0.505762f
C3764 a_19256_45572# VDD 0.27151f
C3765 a_10467_46802# a_11186_47026# 0.082642f
C3766 a_10623_46897# a_10768_47026# 0.057222f
C3767 a_13720_44458# VDD 0.202097f
C3768 a_9482_43914# a_13857_44734# 0.011887f
C3769 a_10341_42308# a_10723_42308# 0.024028f
C3770 a_19778_44110# a_15493_43940# 0.033844f
C3771 a_5111_42852# VDD 0.178652f
C3772 a_1208_46090# VDD 0.178097f
C3773 a_5111_44636# a_5193_42852# 0.018763f
C3774 a_13249_42308# a_13575_42558# 0.088907f
C3775 a_11415_45002# a_20567_45036# 0.011165f
C3776 a_11525_45546# VDD 0.133093f
C3777 a_1823_45246# a_3905_42865# 0.218008f
C3778 C0_N_btm VREF_GND 0.350401f
C3779 C0_dummy_N_btm VCM 0.311452f
C3780 RST_Z SINGLE_ENDED 0.0318f
C3781 a_4651_46660# a_5385_46902# 0.053479f
C3782 a_4955_46873# a_4817_46660# 0.318259f
C3783 a_3877_44458# a_5907_46634# 0.073504f
C3784 VDD CLK_DATA 0.422202f
C3785 C2_N_btm VIN_N 0.502408f
C3786 C1_N_btm VREF 0.98698f
C3787 a_20411_46873# a_20528_46660# 0.170785f
C3788 a_20841_46902# a_21188_46660# 0.051162f
C3789 a_7542_44172# VDD 0.412456f
C3790 a_18599_43230# a_18504_43218# 0.049827f
C3791 a_16795_42852# a_16877_42852# 0.171361f
C3792 a_6575_47204# VDD 1.32036f
C3793 a_6755_46942# a_15599_45572# 0.024601f
C3794 a_n1853_46287# a_n863_45724# 0.019522f
C3795 a_16977_43638# VDD 0.206333f
C3796 a_18579_44172# a_19478_44306# 0.040429f
C3797 a_11415_45002# a_14180_45002# 0.025987f
C3798 a_6491_46660# a_6575_47204# 0.029984f
C3799 a_18494_42460# a_20356_42852# 0.014237f
C3800 a_18479_45785# a_19256_45572# 0.044595f
C3801 a_18909_45814# a_18691_45572# 0.209641f
C3802 a_18341_45572# a_19431_45546# 0.041762f
C3803 a_18175_45572# a_18596_45572# 0.086708f
C3804 VDAC_N C6_N_btm 55.2142f
C3805 a_5205_44484# VDD 0.508148f
C3806 a_4905_42826# a_4520_42826# 0.147708f
C3807 a_16243_43396# a_16409_43396# 0.575934f
C3808 a_1823_45246# a_4093_43548# 0.17443f
C3809 a_2905_45572# a_3218_45724# 0.021505f
C3810 a_19321_45002# a_18819_46122# 0.018323f
C3811 a_17701_42308# a_17333_42852# 0.061051f
C3812 a_5755_42852# a_6101_43172# 0.013377f
C3813 a_17061_44734# VDD 0.17647f
C3814 a_12607_44458# a_12883_44458# 0.11453f
C3815 a_11189_46129# a_11387_46155# 0.320331f
C3816 a_1427_43646# VDD 0.19291f
C3817 a_5385_46902# VDD 0.203316f
C3818 a_14537_43396# a_14955_43396# 0.027267f
C3819 a_22400_42852# a_22537_39537# 0.019618f
C3820 a_n1920_47178# a_n1605_47204# 0.08571f
C3821 a_n1533_46116# VDD 0.143145f
C3822 a_13904_45546# a_14033_45572# 0.010132f
C3823 a_8530_39574# VDAC_P 0.064895f
C3824 a_20974_43370# a_21487_43396# 0.03755f
C3825 a_19431_45546# VDD 0.342308f
C3826 a_6755_46942# a_8270_45546# 0.045608f
C3827 a_10428_46928# a_11186_47026# 0.055625f
C3828 a_13076_44458# VDD 0.180665f
C3829 a_n863_45724# a_1568_43370# 0.202455f
C3830 a_1138_42852# a_791_42968# 0.100783f
C3831 a_n2497_47436# a_n2293_45010# 0.233882f
C3832 a_16388_46812# a_17957_46116# 0.140894f
C3833 a_376_46348# a_472_46348# 0.318161f
C3834 a_10341_42308# a_10533_42308# 0.035479f
C3835 a_12891_46348# VDD 1.01428f
C3836 a_8199_44636# a_8685_42308# 0.114007f
C3837 a_7499_43078# a_7871_42858# 0.146369f
C3838 a_11827_44484# a_19862_44208# 0.015537f
C3839 a_4520_42826# VDD 0.142755f
C3840 a_15959_42545# a_15890_42674# 0.209641f
C3841 a_2675_43914# a_3353_43940# 0.011812f
C3842 a_805_46414# VDD 0.154663f
C3843 a_13249_42308# a_13070_42354# 0.141799f
C3844 a_8746_45002# a_10490_45724# 0.116339f
C3845 a_11322_45546# VDD 0.370908f
C3846 a_1823_45246# a_3600_43914# 0.016141f
C3847 C0_dummy_P_btm VCM 0.311452f
C3848 RST_Z START 0.033428f
C3849 VDD SINGLE_ENDED 0.210835f
C3850 a_4651_46660# a_4817_46660# 0.57393f
C3851 a_3877_44458# a_5167_46660# 0.032716f
C3852 C1_N_btm VIN_N 0.39234f
C3853 C0_N_btm VREF 0.443884f
C3854 a_8270_45546# a_8953_45546# 1.06716f
C3855 a_20273_46660# a_21188_46660# 0.118759f
C3856 a_20107_46660# a_20528_46660# 0.083408f
C3857 a_7281_43914# VDD 0.198809f
C3858 a_7903_47542# VDD 0.202868f
C3859 a_n1853_46287# a_n1079_45724# 0.02186f
C3860 a_16409_43396# VDD 0.250832f
C3861 a_12359_47026# VDD 0.142103f
C3862 a_5663_43940# a_6453_43914# 0.017005f
C3863 a_11415_45002# a_13777_45326# 0.021087f
C3864 a_6851_47204# a_7227_47204# 0.241208f
C3865 a_6545_47178# a_6575_47204# 0.11927f
C3866 a_564_42282# VDD 0.293756f
C3867 a_20202_43084# a_20679_44626# 0.035147f
C3868 a_8270_45546# a_9028_43914# 0.233359f
C3869 a_18341_45572# a_18691_45572# 0.206455f
C3870 a_18175_45572# a_19256_45572# 0.102355f
C3871 a_n1550_35448# a_n217_35014# 0.08192f
C3872 VDAC_N C5_N_btm 27.606901f
C3873 a_6431_45366# VDD 0.203167f
C3874 a_16137_43396# a_16409_43396# 0.011989f
C3875 a_16243_43396# a_16547_43609# 0.165289f
C3876 a_2905_45572# a_2957_45546# 0.137248f
C3877 a_17595_43084# a_17333_42852# 0.057438f
C3878 a_16241_44734# VDD 0.189894f
C3879 a_5111_44636# a_7845_44172# 0.063408f
C3880 a_n746_45260# a_626_44172# 0.011647f
C3881 a_11189_46129# a_11133_46155# 0.203074f
C3882 a_n1557_42282# VDD 0.355513f
C3883 a_4817_46660# VDD 0.370615f
C3884 a_14537_43396# a_15095_43370# 0.019641f
C3885 a_21613_42308# a_22775_42308# 0.225363f
C3886 a_22400_42852# a_22889_38993# 0.13715f
C3887 a_7754_38470# VDAC_P 0.063714f
C3888 a_20974_43370# a_20556_43646# 0.076332f
C3889 a_3905_42865# a_4649_42852# 0.04156f
C3890 a_18691_45572# VDD 0.191893f
C3891 a_19321_45002# a_11415_45002# 0.065361f
C3892 a_10428_46928# a_10768_47026# 0.027606f
C3893 a_12883_44458# VDD 0.263743f
C3894 a_11309_47204# VDD 0.358104f
C3895 a_3065_45002# a_3539_42460# 0.300764f
C3896 a_7499_43078# a_7227_42852# 0.126148f
C3897 a_19466_46812# a_19256_45572# 0.041135f
C3898 a_3935_42891# VDD 0.096403f
C3899 a_15803_42450# a_15890_42674# 0.07009f
C3900 a_472_46348# VDD 0.706547f
C3901 a_20202_43084# a_18494_42460# 0.166633f
C3902 a_15890_42674# VDD 0.203548f
C3903 a_6575_47204# a_8128_46384# 0.105633f
C3904 a_10490_45724# VDD 0.162001f
C3905 a_1823_45246# a_2998_44172# 0.062531f
C3906 C0_P_btm VCM 0.717283f
C3907 VDD START 0.114358f
C3908 a_4651_46660# a_4955_46873# 0.140348f
C3909 a_3877_44458# a_5385_46902# 0.021989f
C3910 C0_N_btm VIN_N 0.529671f
C3911 a_20841_46902# a_20623_46660# 0.209641f
C3912 a_20273_46660# a_21363_46634# 0.042415f
C3913 a_13059_46348# a_11415_45002# 0.225168f
C3914 a_6453_43914# VDD 0.194953f
C3915 a_16414_43172# a_16245_42852# 0.08213f
C3916 a_18249_42858# a_18504_43218# 0.05936f
C3917 a_7227_47204# VDD 0.430714f
C3918 a_11189_46129# a_10586_45546# 0.028266f
C3919 a_6761_42308# a_7227_42308# 0.173849f
C3920 a_16547_43609# VDD 0.31275f
C3921 a_18579_44172# a_19328_44172# 0.053539f
C3922 a_19279_43940# a_19862_44208# 0.012567f
C3923 a_12156_46660# VDD 0.082428f
C3924 a_1115_44172# a_1241_44260# 0.013015f
C3925 a_5111_44636# a_5111_42852# 0.148196f
C3926 a_11415_45002# a_13556_45296# 0.16025f
C3927 a_3503_45724# a_3775_45552# 0.13675f
C3928 a_19319_43548# a_19741_43940# 0.048788f
C3929 a_n2840_45546# VDD 0.302566f
C3930 a_20202_43084# a_20640_44752# 0.027593f
C3931 a_18175_45572# a_19431_45546# 0.043567f
C3932 a_18479_45785# a_18691_45572# 0.036486f
C3933 a_18341_45572# a_18909_45814# 0.170692f
C3934 a_n1550_35448# EN_VIN_BSTR_P 0.573018f
C3935 VDAC_N C4_N_btm 13.8047f
C3936 a_16137_43396# a_16547_43609# 0.151161f
C3937 a_16795_42852# a_17333_42852# 0.108694f
C3938 a_17595_43084# a_18083_42858# 0.046381f
C3939 a_14673_44172# VDD 0.381917f
C3940 SMPL_ON_P a_n1550_35448# 0.012033f
C3941 a_5111_44636# a_7542_44172# 0.039468f
C3942 a_n1641_46494# a_n1533_46116# 0.057222f
C3943 a_18989_43940# a_15493_43940# 0.025737f
C3944 a_14537_43396# a_14205_43396# 0.080783f
C3945 a_4955_46873# VDD 0.467566f
C3946 a_11415_45002# a_21363_45546# 0.011178f
C3947 a_20202_43084# a_21188_45572# 0.013137f
C3948 a_11189_46129# a_11136_45572# 0.042798f
C3949 a_22400_42852# a_22613_38993# 0.038807f
C3950 a_8292_43218# VDD 0.08228f
C3951 a_18597_46090# a_20974_43370# 0.025672f
C3952 a_n2302_39072# VDD 0.355374f
C3953 a_n2302_37690# a_n2216_37690# 0.011479f
C3954 a_8530_39574# VDAC_N 0.06498f
C3955 a_3499_42826# a_n2293_42282# 0.058548f
C3956 a_18909_45814# VDD 0.205795f
C3957 a_5111_44636# a_5205_44484# 0.200189f
C3958 a_8746_45002# a_8975_43940# 0.016889f
C3959 a_n2293_45010# a_626_44172# 0.024201f
C3960 a_12607_44458# VDD 0.188171f
C3961 a_n1557_42282# a_196_42282# 0.031105f
C3962 a_n2497_47436# a_n2661_45010# 0.281004f
C3963 a_16388_46812# a_17715_44484# 0.032772f
C3964 a_n2293_42282# a_3318_42354# 0.01699f
C3965 a_19466_46812# a_19431_45546# 0.038922f
C3966 a_3681_42891# VDD 0.223661f
C3967 COMP_P comp_n 0.032515f
C3968 a_15764_42576# a_15890_42674# 0.181217f
C3969 a_15803_42450# a_15959_42545# 0.110532f
C3970 a_376_46348# VDD 0.116284f
C3971 a_11415_45002# a_19778_44110# 0.030651f
C3972 a_7903_47542# a_8128_46384# 0.109077f
C3973 a_15959_42545# VDD 0.19373f
C3974 a_8746_45002# VDD 0.970181f
C3975 a_3905_42865# a_5111_42852# 0.079376f
C3976 a_17339_46660# a_18451_43940# 0.012866f
C3977 a_15599_45572# a_16751_45260# 0.012353f
C3978 C0_P_btm VREF_GND 0.350485f
C3979 C1_P_btm VCM 0.716121f
C3980 VDD RST_Z 4.72787f
C3981 a_3160_47472# a_3699_46348# 0.109505f
C3982 a_3877_44458# a_4817_46660# 0.017126f
C3983 C0_dummy_N_btm VIN_N 0.544204f
C3984 a_7499_43078# a_7845_44172# 0.112307f
C3985 a_8270_45546# a_8199_44636# 0.95539f
C3986 a_5807_45002# a_16375_45002# 0.042941f
C3987 a_17339_46660# a_17639_46660# 0.081726f
C3988 a_20273_46660# a_20623_46660# 0.20669f
C3989 a_20107_46660# a_21188_46660# 0.102355f
C3990 a_5663_43940# VDD 0.133666f
C3991 a_15567_42826# a_16245_42852# 0.03084f
C3992 a_17333_42852# a_18504_43218# 0.157683f
C3993 a_2382_45260# a_3737_43940# 0.027805f
C3994 a_6851_47204# VDD 0.287724f
C3995 a_8270_45546# a_8192_45572# 0.048422f
C3996 a_16243_43396# VDD 0.39865f
C3997 a_19279_43940# a_19478_44306# 0.03583f
C3998 a_18579_44172# a_18451_43940# 0.147572f
C3999 a_5495_43940# a_5663_43940# 0.227135f
C4000 a_11415_45002# a_9482_43914# 0.309633f
C4001 a_6491_46660# a_6851_47204# 0.132946f
C4002 a_n327_42558# VDD 0.198414f
C4003 a_18479_45785# a_18909_45814# 0.023226f
C4004 a_18175_45572# a_18691_45572# 0.105995f
C4005 VDAC_N C3_N_btm 6.907279f
C4006 a_12465_44636# a_6755_46942# 0.021176f
C4007 a_13487_47204# a_14084_46812# 0.012167f
C4008 a_16137_43396# a_16243_43396# 0.182209f
C4009 a_n863_45724# a_895_43940# 0.015488f
C4010 a_15009_46634# a_14180_46812# 0.123843f
C4011 a_2959_46660# a_3147_46376# 0.010696f
C4012 a_5807_45002# a_18985_46122# 0.017912f
C4013 a_17595_43084# a_17701_42308# 0.141211f
C4014 a_5111_42852# a_5457_43172# 0.013377f
C4015 SMPL_ON_P a_n2002_35448# 0.399437f
C4016 a_n746_45260# a_375_42282# 0.41439f
C4017 a_n1423_46090# a_n1533_46116# 0.097745f
C4018 a_4905_42826# VDD 0.439034f
C4019 a_14537_43396# a_14358_43442# 0.1418f
C4020 a_20193_45348# a_20974_43370# 0.026944f
C4021 a_4651_46660# VDD 0.457722f
C4022 a_20202_43084# a_21363_45546# 0.029873f
C4023 a_21887_42336# a_21613_42308# 0.071168f
C4024 a_22400_42852# a_22581_37893# 0.031385f
C4025 a_n2497_47436# a_n1605_47204# 0.0417f
C4026 a_19321_45002# a_20623_43914# 0.294126f
C4027 a_8530_39574# a_6886_37412# 0.616015f
C4028 a_7754_38470# VDAC_N 0.110605f
C4029 a_18341_45572# VDD 0.2432f
C4030 a_5147_45002# a_5205_44484# 0.018671f
C4031 a_8975_43940# VDD 0.257588f
C4032 a_n1557_42282# a_n473_42460# 0.077371f
C4033 a_n863_45724# a_458_43396# 0.122956f
C4034 a_16721_46634# a_15682_46116# 0.010175f
C4035 a_16388_46812# a_17583_46090# 0.033313f
C4036 a_2382_45260# a_3539_42460# 0.110439f
C4037 a_2905_42968# VDD 0.142081f
C4038 a_15486_42560# a_15890_42674# 0.051162f
C4039 a_13575_42558# a_13921_42308# 0.013377f
C4040 a_15764_42576# a_15959_42545# 0.21686f
C4041 a_895_43940# a_2455_43940# 0.01899f
C4042 a_10949_43914# a_12429_44172# 0.156922f
C4043 a_n1076_46494# VDD 0.294742f
C4044 a_10180_45724# a_8746_45002# 0.304016f
C4045 a_10053_45546# a_10490_45724# 0.084842f
C4046 a_20990_47178# a_21177_47436# 0.159555f
C4047 a_15803_42450# VDD 0.448709f
C4048 a_3905_42865# a_4520_42826# 0.054799f
C4049 a_15903_45785# a_16019_45002# 0.139976f
C4050 C1_P_btm VREF_GND 0.673422f
C4051 C2_P_btm VCM 0.716172f
C4052 a_3877_44458# a_4955_46873# 0.029242f
C4053 C0_P_btm VREF 0.443926f
C4054 a_7499_43078# a_7542_44172# 0.069089f
C4055 a_7229_43940# a_5883_43914# 0.026061f
C4056 a_20107_46660# a_21363_46634# 0.043567f
C4057 a_20273_46660# a_20841_46902# 0.17072f
C4058 a_5495_43940# VDD 0.173477f
C4059 a_18083_42858# a_18504_43218# 0.088127f
C4060 a_22959_45036# a_22959_44484# 0.025171f
C4061 a_20193_45348# a_22485_44484# 0.027057f
C4062 a_6491_46660# VDD 0.436756f
C4063 a_10355_46116# a_10586_45546# 0.012906f
C4064 a_6773_42558# a_6761_42308# 0.01129f
C4065 a_16137_43396# VDD 0.483673f
C4066 a_18579_44172# a_18326_43940# 0.096332f
C4067 a_5013_44260# a_5663_43940# 0.083171f
C4068 a_1823_45246# a_3429_45260# 0.047931f
C4069 a_11415_45002# a_13348_45260# 0.036052f
C4070 a_18597_46090# a_20512_43084# 0.023158f
C4071 a_6545_47178# a_6851_47204# 0.134581f
C4072 a_6755_46942# a_15682_43940# 0.028635f
C4073 a_18479_45785# a_18341_45572# 0.21997f
C4074 a_18175_45572# a_18909_45814# 0.053479f
C4075 a_16375_45002# a_17719_45144# 0.201099f
C4076 VDAC_N C2_N_btm 3.46253f
C4077 a_n2302_37690# VDD 0.350119f
C4078 a_5691_45260# VDD 0.205518f
C4079 a_4093_43548# a_4520_42826# 0.077799f
C4080 a_4235_43370# a_3935_42891# 0.082011f
C4081 a_1138_42852# a_1049_43396# 0.022078f
C4082 a_n863_45724# a_2479_44172# 0.047943f
C4083 a_14084_46812# a_14180_46812# 0.318161f
C4084 a_5807_45002# a_18819_46122# 0.012467f
C4085 a_10057_43914# a_8975_43940# 0.069663f
C4086 a_n1991_46122# a_n1533_46116# 0.034619f
C4087 a_14537_43396# a_14579_43548# 0.046172f
C4088 a_21335_42336# a_21613_42308# 0.110671f
C4089 a_n2497_47436# SMPL_ON_P 0.131317f
C4090 a_n863_45724# a_2680_45002# 0.024737f
C4091 a_18597_46090# a_21381_43940# 0.080234f
C4092 a_n2946_39072# VDD 0.383374f
C4093 a_7754_38470# a_6886_37412# 0.181496f
C4094 a_18479_45785# VDD 0.536075f
C4095 a_n2293_45010# a_375_42282# 0.021456f
C4096 a_n2661_45010# a_626_44172# 0.0195f
C4097 a_8746_45002# a_10440_44484# 0.027688f
C4098 a_10057_43914# VDD 0.399284f
C4099 a_2075_43172# a_2905_42968# 0.023236f
C4100 a_n1557_42282# a_n961_42308# 0.041329f
C4101 a_20193_45348# a_20205_45028# 0.012189f
C4102 a_1799_45572# a_1848_45724# 0.080562f
C4103 a_16388_46812# a_15682_46116# 0.044769f
C4104 a_8270_45546# a_8034_45724# 0.031124f
C4105 a_n901_46420# a_n1076_46494# 0.234322f
C4106 a_9804_47204# VDD 0.410522f
C4107 a_5883_43914# a_7845_44172# 0.02286f
C4108 a_18494_42460# a_20269_44172# 0.017863f
C4109 a_15764_42576# a_15803_42450# 0.901878f
C4110 a_20193_45348# a_22223_43396# 0.020364f
C4111 a_2479_44172# a_2455_43940# 0.025354f
C4112 a_895_43940# a_2253_43940# 0.053882f
C4113 a_10949_43914# a_11750_44172# 0.05299f
C4114 a_n901_46420# VDD 0.518805f
C4115 a_10053_45546# a_8746_45002# 0.075884f
C4116 a_22485_38105# a_22629_38406# 0.206945f
C4117 a_15764_42576# VDD 0.258303f
C4118 a_10180_45724# VDD 0.336512f
C4119 a_3905_42865# a_3935_42891# 0.240349f
C4120 en_comp a_1107_38525# 0.206093f
C4121 C2_P_btm VREF_GND 0.671742f
C4122 C3_P_btm VCM 0.716273f
C4123 C0_dummy_P_btm VIN_P 0.544204f
C4124 C1_P_btm VREF 0.98698f
C4125 a_3160_47472# a_3147_46376# 0.208295f
C4126 a_3877_44458# a_4651_46660# 0.032518f
C4127 a_8270_45546# a_8016_46348# 0.036831f
C4128 a_20107_46660# a_20623_46660# 0.105914f
C4129 a_5013_44260# VDD 0.198233f
C4130 a_15567_42826# a_15597_42852# 0.025037f
C4131 a_20193_45348# a_20512_43084# 0.160912f
C4132 a_6545_47178# VDD 0.386368f
C4133 a_19279_43940# a_19328_44172# 0.120319f
C4134 a_20362_44736# a_20365_43914# 0.012553f
C4135 a_5013_44260# a_5495_43940# 0.251039f
C4136 a_11415_45002# a_13159_45002# 0.141106f
C4137 a_1823_45246# a_3065_45002# 0.607468f
C4138 a_6545_47178# a_6491_46660# 0.181574f
C4139 a_196_42282# VDD 0.291844f
C4140 a_18175_45572# a_18341_45572# 0.577068f
C4141 a_16375_45002# a_17613_45144# 0.040514f
C4142 VDAC_N C1_N_btm 1.7375f
C4143 a_4927_45028# VDD 0.159822f
C4144 a_1138_42852# a_1209_43370# 0.01435f
C4145 a_13059_46348# a_14205_43396# 0.049915f
C4146 a_14084_46812# a_14035_46660# 0.086342f
C4147 a_16795_42852# a_17595_43084# 0.010079f
C4148 a_n1917_44484# a_n1821_44484# 0.013793f
C4149 a_10440_44484# a_8975_43940# 0.045841f
C4150 a_4699_43561# VDD 0.262218f
C4151 a_n473_42460# a_n327_42558# 0.171361f
C4152 a_13556_45296# a_14205_43396# 0.012255f
C4153 a_20193_45348# a_21381_43940# 0.01388f
C4154 a_3877_44458# VDD 0.786903f
C4155 a_11415_45002# a_20273_45572# 0.01364f
C4156 a_22400_42852# a_22527_39145# 0.228292f
C4157 a_n1736_46482# VDD 0.083417f
C4158 a_14955_43940# a_15037_43940# 0.171361f
C4159 a_5343_44458# a_8037_42858# 0.019942f
C4160 a_n863_45724# a_2382_45260# 0.119625f
C4161 a_6491_46660# a_3877_44458# 0.02519f
C4162 a_n2946_37690# a_n2860_37690# 0.011479f
C4163 a_20974_43370# a_21259_43561# 0.049502f
C4164 a_18175_45572# VDD 0.38478f
C4165 a_4927_45028# a_5691_45260# 0.018415f
C4166 a_8746_45002# a_10334_44484# 0.019787f
C4167 a_5807_45002# a_11415_45002# 0.05094f
C4168 a_10440_44484# VDD 0.159539f
C4169 a_n1557_42282# a_n1329_42308# 0.075734f
C4170 a_1847_42826# a_2905_42968# 0.097535f
C4171 a_10341_42308# a_9803_42558# 0.108853f
C4172 a_8128_46384# VDD 0.403575f
C4173 a_5111_44636# a_4905_42826# 0.128918f
C4174 a_5883_43914# a_7542_44172# 0.187537f
C4175 a_18494_42460# a_19862_44208# 0.019692f
C4176 a_19466_46812# a_18341_45572# 0.02497f
C4177 a_1847_42826# VDD 0.527555f
C4178 a_14113_42308# a_15890_42674# 0.022182f
C4179 a_15486_42560# a_15803_42450# 0.102355f
C4180 a_2479_44172# a_2253_43940# 0.010537f
C4181 a_10729_43914# a_11750_44172# 0.144893f
C4182 a_10949_43914# a_10807_43548# 0.034945f
C4183 a_2127_44172# a_2455_43940# 0.096132f
C4184 a_895_43940# a_1443_43940# 0.016028f
C4185 a_22959_46660# EN_OFFSET_CAL 0.050989f
C4186 a_n1641_46494# VDD 0.226065f
C4187 a_9049_44484# a_8746_45002# 0.025877f
C4188 a_22485_38105# CAL_P 0.026856f
C4189 a_20894_47436# a_20990_47178# 0.313533f
C4190 a_15486_42560# VDD 0.275297f
C4191 a_10053_45546# VDD 0.150582f
C4192 a_3905_42865# a_3681_42891# 0.101054f
C4193 a_1568_43370# a_1427_43646# 0.046825f
C4194 a_1138_42852# a_895_43940# 0.017458f
C4195 C3_P_btm VREF_GND 0.67174f
C4196 C4_P_btm VCM 0.716447f
C4197 a_2905_45572# a_3147_46376# 0.02017f
C4198 C10_N_btm VDD 2.40001f
C4199 C0_P_btm VIN_P 0.529671f
C4200 C2_P_btm VREF 0.987884f
C4201 a_20411_46873# a_20273_46660# 0.219954f
C4202 a_20107_46660# a_20841_46902# 0.053479f
C4203 a_5244_44056# VDD 0.146618f
C4204 a_4007_47204# DATA[2] 0.337596f
C4205 a_19466_46812# VDD 0.664497f
C4206 a_5244_44056# a_5495_43940# 0.107037f
C4207 a_11415_45002# a_13017_45260# 0.100288f
C4208 a_1823_45246# a_2680_45002# 0.073588f
C4209 a_n473_42460# VDD 0.27195f
C4210 a_18175_45572# a_18479_45785# 0.280208f
C4211 a_16375_45002# a_17023_45118# 0.014031f
C4212 VDAC_N C0_N_btm 0.901121f
C4213 VDAC_P C0_dummy_P_btm 0.88451f
C4214 a_n2002_35448# a_n1550_35448# 0.150805f
C4215 a_n2946_37690# VDD 0.38221f
C4216 a_5111_44636# VDD 1.28013f
C4217 a_8191_45002# a_8560_45348# 0.03364f
C4218 a_n863_45724# a_453_43940# 0.02533f
C4219 a_13059_46348# a_14358_43442# 0.041731f
C4220 a_14084_46812# a_13885_46660# 0.237373f
C4221 a_5807_45002# a_18189_46348# 0.033239f
C4222 a_4520_42826# a_4743_43172# 0.011458f
C4223 a_5147_45002# a_5663_43940# 0.019985f
C4224 a_5111_44636# a_5495_43940# 0.037006f
C4225 a_10334_44484# a_8975_43940# 0.044798f
C4226 a_10440_44484# a_10057_43914# 0.026774f
C4227 a_n1641_46494# a_n1545_46494# 0.013793f
C4228 a_4235_43370# VDD 0.229422f
C4229 a_11415_45002# a_20107_45572# 0.019157f
C4230 a_22400_42852# a_22589_40055# 0.663766f
C4231 a_n2497_47436# a_n1920_47178# 0.049461f
C4232 a_2479_44172# a_2896_43646# 0.026857f
C4233 a_3905_42865# a_4905_42826# 0.404829f
C4234 a_5343_44458# a_7765_42852# 0.010279f
C4235 a_18189_46348# a_18315_45260# 0.101775f
C4236 a_310_45028# a_n37_45144# 0.112458f
C4237 a_n863_45724# a_2274_45254# 0.17549f
C4238 a_19321_45002# a_19862_44208# 0.090113f
C4239 a_6545_47178# a_3877_44458# 0.026367f
C4240 a_n3690_39392# VDD 0.363068f
C4241 en_comp a_22527_39145# 0.393507f
C4242 a_16147_45260# VDD 0.197706f
C4243 a_5111_44636# a_5691_45260# 0.130044f
C4244 a_n2661_45010# a_375_42282# 0.017053f
C4245 a_10334_44484# VDD 0.19332f
C4246 a_n1557_42282# COMP_P 0.123881f
C4247 a_1847_42826# a_2075_43172# 0.103349f
C4248 a_n1423_46090# a_n1076_46494# 0.051162f
C4249 a_5883_43914# a_7281_43914# 0.029594f
C4250 a_16922_45042# a_15493_43940# 0.019907f
C4251 a_791_42968# VDD 0.128737f
C4252 a_14113_42308# a_15959_42545# 0.036113f
C4253 a_15486_42560# a_15764_42576# 0.118759f
C4254 a_15051_42282# a_15803_42450# 0.043619f
C4255 a_10729_43914# a_10807_43548# 0.238591f
C4256 a_2127_44172# a_2253_43940# 0.143754f
C4257 a_895_43940# a_1241_43940# 0.054548f
C4258 a_n1423_46090# VDD 0.227012f
C4259 a_6667_45809# a_6977_45572# 0.013793f
C4260 a_10053_45546# a_10180_45724# 0.144403f
C4261 a_7499_43078# a_8746_45002# 0.153858f
C4262 a_n2302_37984# a_n2216_37984# 0.011479f
C4263 a_15051_42282# VDD 0.461307f
C4264 a_9049_44484# VDD 0.680993f
C4265 a_1049_43396# a_1427_43646# 0.010711f
C4266 a_15493_43940# a_15743_43084# 0.206331f
C4267 C4_P_btm VREF_GND 0.671882f
C4268 C5_P_btm VCM 0.719982f
C4269 C9_N_btm VDD 0.345685f
C4270 C1_P_btm VIN_P 0.39234f
C4271 C3_P_btm VREF 0.984942f
C4272 a_7229_43940# a_6298_44484# 0.028942f
C4273 a_20107_46660# a_20273_46660# 0.608339f
C4274 a_3905_42865# VDD 0.788273f
C4275 a_3815_47204# DATA[2] 0.022461f
C4276 a_5815_47464# VDD 0.399354f
C4277 a_n2472_46090# a_n2472_45546# 0.025171f
C4278 a_19333_46634# VDD 0.199048f
C4279 a_5244_44056# a_5013_44260# 0.094334f
C4280 a_11415_45002# a_11963_45334# 0.031636f
C4281 a_1823_45246# a_2382_45260# 0.801932f
C4282 a_167_45260# a_1667_45002# 0.05322f
C4283 a_n961_42308# VDD 0.24416f
C4284 a_18494_42460# a_20256_43172# 0.052522f
C4285 a_16375_45002# a_16922_45042# 0.170835f
C4286 VDAC_N C0_dummy_N_btm 0.885361f
C4287 VDAC_P C0_P_btm 0.901219f
C4288 CAL_P EN_VIN_BSTR_N 0.040136f
C4289 a_5147_45002# VDD 0.574918f
C4290 a_n863_45724# a_1414_42308# 0.711805f
C4291 a_13059_46348# a_14579_43548# 0.171744f
C4292 a_13607_46688# a_13885_46660# 0.11044f
C4293 a_5807_45002# a_17715_44484# 0.045558f
C4294 a_4520_42826# a_4649_43172# 0.010132f
C4295 a_5147_45002# a_5495_43940# 0.086203f
C4296 a_5111_44636# a_5013_44260# 0.029412f
C4297 a_n1917_44484# a_n1809_44850# 0.057222f
C4298 a_10157_44484# a_8975_43940# 0.045547f
C4299 a_n1641_46494# a_n1736_46482# 0.049827f
C4300 a_13059_46348# a_12839_46116# 0.098052f
C4301 a_4093_43548# VDD 0.216874f
C4302 a_22165_42308# a_17303_42282# 0.095988f
C4303 a_19511_42282# a_21125_42558# 0.01129f
C4304 a_13483_43940# a_13565_43940# 0.171361f
C4305 a_1414_42308# a_3540_43646# 0.022584f
C4306 a_5343_44458# a_7871_42858# 0.020081f
C4307 a_n863_45724# a_1667_45002# 0.20954f
C4308 a_8530_39574# a_3726_37500# 1.35509f
C4309 en_comp a_22589_40055# 0.260977f
C4310 a_21381_43940# a_21259_43561# 0.013931f
C4311 a_5147_45002# a_5691_45260# 0.035185f
C4312 a_5111_44636# a_4927_45028# 0.134309f
C4313 a_7499_43078# a_8975_43940# 0.519621f
C4314 a_6755_46942# a_7832_46660# 0.025487f
C4315 a_10157_44484# VDD 0.174233f
C4316 a_13059_46348# a_14840_46494# 0.031849f
C4317 a_n1991_46122# a_n1076_46494# 0.124988f
C4318 a_5883_43914# a_6453_43914# 0.051468f
C4319 a_19778_44110# a_19862_44208# 0.213467f
C4320 a_11415_45002# a_13249_42308# 0.071546f
C4321 a_685_42968# VDD 0.088446f
C4322 a_14113_42308# a_15803_42450# 0.289859f
C4323 a_15051_42282# a_15764_42576# 0.042737f
C4324 a_10729_43914# a_10949_43914# 0.418928f
C4325 a_n1991_46122# VDD 0.581018f
C4326 a_2112_39137# VDAC_Ni 0.018095f
C4327 a_14113_42308# VDD 0.365578f
C4328 a_7499_43078# VDD 1.87959f
C4329 a_1209_43370# a_1427_43646# 0.08213f
C4330 a_1049_43396# a_n1557_42282# 0.211757f
C4331 a_n863_45724# a_n699_43396# 0.23135f
C4332 a_8270_45546# a_9801_43940# 0.014887f
C4333 C5_P_btm VREF_GND 0.676559f
C4334 C6_P_btm VCM 0.877162f
C4335 C8_N_btm VDD 0.19922f
C4336 C2_P_btm VIN_P 0.502408f
C4337 C4_P_btm VREF 0.98728f
C4338 a_20107_46660# a_20411_46873# 0.316529f
C4339 a_3600_43914# VDD 0.22716f
C4340 a_16795_42852# a_17141_43172# 0.013377f
C4341 a_3785_47178# DATA[2] 0.119025f
C4342 a_14539_43914# a_14815_43914# 0.099149f
C4343 a_5129_47502# VDD 0.20906f
C4344 a_15781_43660# VDD 0.196099f
C4345 a_3905_42865# a_5013_44260# 0.182997f
C4346 a_11415_45002# a_11787_45002# 0.072246f
C4347 a_1823_45246# a_2274_45254# 0.255985f
C4348 a_167_45260# a_327_44734# 0.199136f
C4349 COMP_P RST_Z 0.03403f
C4350 a_n1329_42308# VDD 0.237697f
C4351 a_16147_45260# a_18175_45572# 0.108647f
C4352 VDAC_P C1_P_btm 1.74268f
C4353 a_n3690_37440# VDD 0.363068f
C4354 a_4558_45348# VDD 0.25277f
C4355 a_15781_43660# a_16137_43396# 0.089942f
C4356 a_n863_45724# a_1467_44172# 0.021736f
C4357 a_5147_45002# a_5013_44260# 0.189328f
C4358 a_5111_44636# a_5244_44056# 0.01138f
C4359 a_n1917_44484# a_n2012_44484# 0.049827f
C4360 a_9838_44484# a_8975_43940# 0.055678f
C4361 a_n1699_44726# a_n1809_44850# 0.097745f
C4362 a_10334_44484# a_10440_44484# 0.313533f
C4363 a_1756_43548# VDD 0.138878f
C4364 a_22400_42852# a_22537_40625# 0.93502f
C4365 a_n2497_47436# a_n2288_47178# 0.067981f
C4366 a_22959_46124# VDD 0.309939f
C4367 a_n863_45724# a_327_44734# 0.353745f
C4368 a_n4334_39392# VDD 0.385989f
C4369 a_7754_38470# a_3726_37500# 0.124796f
C4370 VDAC_Ni a_6886_37412# 0.178275f
C4371 a_20193_45348# a_21613_42308# 0.137559f
C4372 a_5147_45002# a_4927_45028# 0.168157f
C4373 a_7499_43078# a_10057_43914# 0.262644f
C4374 a_9838_44484# VDD 0.242131f
C4375 a_n1557_42282# a_n1736_42282# 0.170341f
C4376 a_n1423_46090# a_n1641_46494# 0.209641f
C4377 a_n1991_46122# a_n901_46420# 0.041816f
C4378 a_n1853_46287# a_n1076_46494# 0.056078f
C4379 a_5883_43914# a_5663_43940# 0.153361f
C4380 a_19778_44110# a_19478_44306# 0.099524f
C4381 a_6298_44484# a_7542_44172# 0.014735f
C4382 a_12465_44636# a_11827_44484# 0.785011f
C4383 a_14113_42308# a_15764_42576# 0.229529f
C4384 a_15051_42282# a_15486_42560# 0.234322f
C4385 a_n1853_46287# VDD 0.645231f
C4386 a_22591_46660# EN_OFFSET_CAL 0.047938f
C4387 a_10405_44172# a_10949_43914# 0.05348f
C4388 a_13657_42558# VDD 0.195727f
C4389 a_22485_38105# a_22537_39537# 0.559814f
C4390 a_8568_45546# VDD 0.182812f
C4391 a_1209_43370# a_n1557_42282# 0.113851f
C4392 a_742_44458# a_1755_42282# 0.013027f
C4393 a_1138_42852# a_453_43940# 0.018298f
C4394 C7_N_btm VDD 0.121904f
C4395 a_5807_45002# a_11813_46116# 0.037525f
C4396 C3_P_btm VIN_P 0.455045f
C4397 C9_N_btm C10_N_btm 53.3168f
C4398 C5_P_btm VREF 0.987144f
C4399 C6_P_btm VREF_GND 0.836236f
C4400 C7_P_btm VCM 1.58335f
C4401 a_7229_43940# a_5343_44458# 0.196399f
C4402 a_5205_44484# a_6298_44484# 0.085118f
C4403 a_2998_44172# VDD 0.362233f
C4404 a_11827_44484# a_22485_44484# 0.015798f
C4405 a_15681_43442# VDD 0.159054f
C4406 a_18834_46812# VDD 0.116625f
C4407 a_1823_45246# a_1667_45002# 0.24808f
C4408 COMP_P VDD 3.52636f
C4409 a_16375_45002# a_16405_45348# 0.012425f
C4410 VDAC_P C2_P_btm 3.46245f
C4411 a_4574_45260# VDD 0.122256f
C4412 a_1414_42308# a_1184_42692# 0.115223f
C4413 a_19333_46634# a_19466_46812# 0.167526f
C4414 a_5807_45002# a_15682_46116# 0.062679f
C4415 a_5147_45002# a_5244_44056# 0.122327f
C4416 a_n2267_44484# a_n1809_44850# 0.027606f
C4417 a_5883_43914# a_8975_43940# 0.50976f
C4418 a_n1991_46122# a_n1736_46482# 0.06121f
C4419 a_1568_43370# VDD 0.433732f
C4420 a_n961_42308# a_n473_42460# 0.011409f
C4421 a_22400_42852# a_22589_40599# 0.135364f
C4422 a_3905_42865# a_4235_43370# 0.041971f
C4423 a_1823_45246# a_n699_43396# 0.08003f
C4424 a_17715_44484# a_17613_45144# 0.012898f
C4425 a_20193_45348# a_21887_42336# 0.169001f
C4426 en_comp a_22537_40625# 0.021487f
C4427 a_4558_45348# a_4927_45028# 0.123258f
C4428 a_5147_45002# a_5111_44636# 0.562127f
C4429 a_15861_45028# a_17613_45144# 0.016666f
C4430 a_8667_46634# a_8270_45546# 0.046604f
C4431 a_5883_43914# VDD 0.859221f
C4432 a_13059_46348# a_14275_46494# 0.036863f
C4433 a_n1991_46122# a_n1641_46494# 0.219633f
C4434 a_n2157_46122# a_n1076_46494# 0.102355f
C4435 a_n1853_46287# a_n901_46420# 0.049679f
C4436 a_14635_42282# a_14853_42852# 0.01129f
C4437 a_5343_44458# a_7845_44172# 0.103601f
C4438 a_5883_43914# a_5495_43940# 0.09813f
C4439 a_6298_44484# a_7281_43914# 0.010383f
C4440 a_5204_45822# a_5263_45724# 0.109078f
C4441 a_3877_44458# a_4558_45348# 0.028316f
C4442 a_n746_45260# a_n23_44458# 0.046452f
C4443 a_11551_42558# a_11897_42308# 0.013377f
C4444 a_14113_42308# a_15486_42560# 0.039784f
C4445 a_n2157_46122# VDD 0.42567f
C4446 a_11415_45002# EN_OFFSET_CAL 0.14622f
C4447 a_10405_44172# a_10729_43914# 0.083277f
C4448 a_1414_42308# a_1443_43940# 0.018064f
C4449 a_11415_45002# a_16922_45042# 0.012903f
C4450 a_n2946_37984# a_n2860_37984# 0.011479f
C4451 a_22485_38105# a_22889_38993# 0.089418f
C4452 a_8162_45546# VDD 0.266272f
C4453 a_458_43396# a_n1557_42282# 0.027865f
C4454 a_4093_43548# a_4235_43370# 0.515101f
C4455 a_8270_45546# a_9165_43940# 0.063297f
C4456 a_18597_46090# a_20411_46873# 0.070431f
C4457 C6_N_btm VDD 0.210613f
C4458 C4_P_btm VIN_P 0.50261f
C4459 C8_N_btm C10_N_btm 2.07867f
C4460 C6_P_btm VREF 1.41944f
C4461 C8_P_btm VCM 2.61094f
C4462 C7_P_btm VREF_GND 1.61142f
C4463 a_5205_44484# a_5518_44484# 0.135771f
C4464 a_2889_44172# VDD 0.1447f
C4465 a_11827_44484# a_20512_43084# 0.030456f
C4466 a_n863_45724# a_n13_43084# 0.041588f
C4467 a_15004_44636# a_14815_43914# 0.078606f
C4468 a_8975_43940# a_11541_44484# 0.028558f
C4469 a_8199_44636# a_10586_45546# 0.057648f
C4470 a_17609_46634# VDD 0.501057f
C4471 a_n1549_44318# a_n1441_43940# 0.057222f
C4472 a_3065_45002# a_3935_42891# 0.01149f
C4473 a_167_45260# a_n37_45144# 0.277898f
C4474 a_1169_39587# a_1169_39043# 0.054961f
C4475 a_19443_46116# VDD 0.132317f
C4476 a_7499_43078# a_5111_44636# 0.753731f
C4477 VDAC_P C3_P_btm 6.90991f
C4478 a_n4334_37440# VDD 0.385859f
C4479 a_n746_45260# a_n356_45724# 0.030083f
C4480 a_2443_46660# a_167_45260# 0.012819f
C4481 a_5147_45002# a_3905_42865# 0.048808f
C4482 a_n2129_44697# a_n1809_44850# 0.026556f
C4483 a_n2267_44484# a_n2012_44484# 0.05936f
C4484 a_10157_44484# a_10334_44484# 0.159555f
C4485 a_n1853_46287# a_n1736_46482# 0.170096f
C4486 a_9625_46129# a_9823_46155# 0.321686f
C4487 a_1049_43396# VDD 0.196328f
C4488 a_14539_43914# a_15493_43940# 0.625897f
C4489 a_n2833_47464# a_n2497_47436# 0.217831f
C4490 a_22223_46124# VDD 0.300745f
C4491 a_3905_42865# a_4093_43548# 0.032751f
C4492 a_18494_42460# a_19987_42826# 0.098055f
C4493 a_167_45260# a_949_44458# 0.021626f
C4494 a_1138_42852# a_n699_43396# 0.024181f
C4495 a_18189_46348# a_16922_45042# 0.015824f
C4496 a_n863_45724# a_n37_45144# 0.056531f
C4497 en_comp a_22589_40599# 0.021612f
C4498 a_4574_45260# a_4927_45028# 0.047624f
C4499 a_15861_45028# a_17023_45118# 0.076138f
C4500 a_8701_44490# VDD 0.164475f
C4501 a_685_42968# a_791_42968# 0.13675f
C4502 a_n863_45724# a_104_43370# 0.046664f
C4503 a_13059_46348# a_14493_46090# 0.029059f
C4504 a_n1991_46122# a_n1423_46090# 0.175891f
C4505 a_n2157_46122# a_n901_46420# 0.043559f
C4506 a_n1853_46287# a_n1641_46494# 0.033696f
C4507 a_n2293_42282# a_1755_42282# 0.875855f
C4508 a_19778_44110# a_19328_44172# 0.064774f
C4509 a_5343_44458# a_7542_44172# 0.014194f
C4510 a_3877_44458# a_4574_45260# 0.010367f
C4511 a_n1533_42852# VDD 0.142813f
C4512 a_14113_42308# a_15051_42282# 0.077852f
C4513 a_1467_44172# a_1443_43940# 0.011516f
C4514 a_5257_43370# a_5708_44484# 0.056224f
C4515 a_22485_38105# a_22613_38993# 0.253409f
C4516 a_2684_37794# VDAC_Pi 0.133177f
C4517 a_7230_45938# VDD 0.077608f
C4518 a_458_43396# a_766_43646# 0.017351f
C4519 a_n863_45724# a_949_44458# 0.034335f
C4520 a_1138_42852# a_1467_44172# 0.034446f
C4521 a_18479_47436# a_20273_46660# 0.018124f
C4522 C5_N_btm VDD 0.267489f
C4523 C5_P_btm VIN_P 0.502041f
C4524 C8_N_btm C9_N_btm 39.4538f
C4525 C7_N_btm C10_N_btm 1.39624f
C4526 C7_P_btm VREF 1.818f
C4527 C9_P_btm VCM 6.06251f
C4528 C8_P_btm VREF_GND 2.58605f
C4529 a_20202_43084# a_15743_43084# 0.021267f
C4530 a_5205_44484# a_5343_44458# 0.129692f
C4531 a_10249_46116# a_10355_46116# 0.182836f
C4532 a_2675_43914# VDD 0.200923f
C4533 a_n2840_46090# a_n2840_45546# 0.025171f
C4534 a_3823_42558# a_4169_42308# 0.013377f
C4535 a_16292_46812# VDD 0.123916f
C4536 a_n1331_43914# a_n1441_43940# 0.097745f
C4537 a_167_45260# a_n143_45144# 0.03701f
C4538 a_n1736_42282# VDD 0.227152f
C4539 a_17478_45572# a_17668_45572# 0.045837f
C4540 VDAC_P C4_P_btm 13.8049f
C4541 a_8530_39574# RST_Z 0.431385f
C4542 a_3429_45260# VDD 0.142923f
C4543 a_1414_42308# a_1067_42314# 0.100434f
C4544 a_1568_43370# a_1847_42826# 0.153113f
C4545 a_n863_45724# a_175_44278# 0.113317f
C4546 a_n2129_44697# a_n2012_44484# 0.172424f
C4547 a_n2157_46122# a_n1736_46482# 0.086708f
C4548 a_9625_46129# a_9569_46155# 0.204034f
C4549 a_13059_46348# a_14180_46482# 0.025233f
C4550 a_n2497_47436# a_626_44172# 0.249352f
C4551 a_1209_43370# VDD 0.191694f
C4552 a_5066_45546# a_5263_45724# 0.022243f
C4553 a_10807_43548# a_11257_43940# 0.013221f
C4554 a_17715_44484# a_16922_45042# 0.039816f
C4555 a_n863_45724# a_n143_45144# 0.033306f
C4556 a_21811_47423# a_20916_46384# 0.109084f
C4557 en_comp CAL_N 0.023818f
C4558 a_4558_45348# a_5147_45002# 0.09356f
C4559 a_15861_45028# a_16922_45042# 0.259169f
C4560 a_8103_44636# VDD 0.124028f
C4561 a_13059_46348# a_13925_46122# 0.056739f
C4562 a_5807_45002# a_6511_45714# 0.012932f
C4563 a_8270_45546# a_5066_45546# 0.189476f
C4564 a_n2157_46122# a_n1641_46494# 0.105995f
C4565 a_n1853_46287# a_n1423_46090# 0.043126f
C4566 a_n2472_46090# VDD 0.224658f
C4567 a_22365_46825# EN_OFFSET_CAL 0.195393f
C4568 a_1115_44172# a_1443_43940# 0.096132f
C4569 a_1467_44172# a_1241_43940# 0.011879f
C4570 a_18479_47436# a_20894_47436# 0.032517f
C4571 a_14456_42282# VDD 0.265543f
C4572 a_22485_38105# a_22581_37893# 0.902394f
C4573 a_6812_45938# VDD 0.132317f
C4574 a_n863_45724# a_742_44458# 0.629795f
C4575 a_1138_42852# a_1115_44172# 0.012127f
C4576 C4_N_btm VDD 0.265463f
C4577 a_18479_47436# a_20411_46873# 0.192791f
C4578 C6_P_btm VIN_P 0.391898f
C4579 C7_N_btm C9_N_btm 0.22201f
C4580 C6_N_btm C10_N_btm 0.895671f
C4581 C8_P_btm VREF 3.6701f
C4582 C10_P_btm VCM 10.5945f
C4583 C9_P_btm VREF_GND 5.18245f
C4584 a_3539_42460# a_n2293_42282# 0.010651f
C4585 a_5111_44636# a_5883_43914# 0.281106f
C4586 a_10249_46116# a_9823_46155# 0.082191f
C4587 a_895_43940# VDD 0.318652f
C4588 a_13720_44458# a_14112_44734# 0.016359f
C4589 a_4700_47436# VDD 0.086132f
C4590 a_12465_44636# a_14537_43396# 0.031033f
C4591 a_5755_42308# a_6171_42473# 0.017801f
C4592 a_15559_46634# VDD 0.301657f
C4593 a_n1899_43946# a_n1441_43940# 0.03441f
C4594 a_2382_45260# a_3935_42891# 0.061675f
C4595 a_10586_45546# a_11682_45822# 0.014019f
C4596 a_15861_45028# a_17668_45572# 0.065471f
C4597 a_8199_44636# a_8375_44464# 0.043989f
C4598 a_7754_38470# RST_Z 0.034995f
C4599 a_8530_39574# VDD 0.346613f
C4600 a_22629_37990# a_22737_36887# 0.08947f
C4601 VDAC_P C5_P_btm 27.6071f
C4602 a_3065_45002# VDD 0.501045f
C4603 a_15095_43370# a_15743_43084# 0.022008f
C4604 a_1799_45572# a_167_45260# 0.061186f
C4605 a_n2433_44484# a_n2012_44484# 0.093133f
C4606 a_8199_44636# a_10355_46116# 0.176325f
C4607 a_8953_45546# a_9569_46155# 0.014447f
C4608 a_13059_46348# a_12638_46436# 0.053952f
C4609 a_5257_43370# a_6472_45840# 0.012073f
C4610 a_458_43396# VDD 0.431902f
C4611 a_3067_47026# VDD 0.132018f
C4612 a_15015_46420# a_15143_45578# 0.011172f
C4613 a_19511_42282# a_21335_42336# 0.011904f
C4614 a_10807_43548# a_11173_43940# 0.013678f
C4615 a_21137_46414# VDD 0.219745f
C4616 a_n863_45724# a_n467_45028# 0.037721f
C4617 VDAC_Ni a_3726_37500# 1.5261f
C4618 a_20193_45348# a_20712_42282# 0.010791f
C4619 a_2813_43396# a_3457_43396# 0.026697f
C4620 a_9049_44484# a_5883_43914# 0.025986f
C4621 a_7927_46660# a_8023_46660# 0.013793f
C4622 a_6755_46942# a_6969_46634# 0.085936f
C4623 a_6298_44484# VDD 1.21616f
C4624 a_13059_46348# a_13759_46122# 0.249771f
C4625 a_5807_45002# a_6472_45840# 0.016039f
C4626 a_n1853_46287# a_n1991_46122# 0.737461f
C4627 a_n2157_46122# a_n1423_46090# 0.053479f
C4628 a_15433_44458# a_14673_44172# 0.027789f
C4629 a_16922_45042# a_20365_43914# 0.021687f
C4630 a_3877_44458# a_3429_45260# 0.02987f
C4631 a_18579_44172# a_18533_43940# 0.011624f
C4632 a_n2840_46090# VDD 0.295278f
C4633 a_1115_44172# a_1241_43940# 0.143754f
C4634 a_8568_45546# a_7499_43078# 0.070368f
C4635 a_18479_47436# a_19787_47423# 0.029306f
C4636 a_13575_42558# VDD 0.182133f
C4637 VCM VSS 63.4818f
C4638 VREF_GND VSS 60.3924f
C4639 VREF VSS 43.355f
C4640 VIN_N VSS 17.425707f
C4641 VIN_P VSS 17.402405f
C4642 CLK VSS 3.412422f
C4643 EN_OFFSET_CAL VSS 0.505642f
C4644 DATA[5] VSS 0.561058f
C4645 DATA[4] VSS 0.755679f
C4646 DATA[3] VSS 1.01838f
C4647 DATA[2] VSS 0.536983f
C4648 DATA[1] VSS 0.550109f
C4649 DATA[0] VSS 0.616231f
C4650 CLK_DATA VSS 0.488979f
C4651 SINGLE_ENDED VSS 0.60168f
C4652 START VSS 0.991673f
C4653 RST_Z VSS 16.923779f
C4654 VDD VSS 0.589169p
C4655 C10_N_btm VSS 0.213734p
C4656 C9_N_btm VSS 82.96518f
C4657 C8_N_btm VSS 48.225792f
C4658 C7_N_btm VSS 0.183895p
C4659 C6_N_btm VSS 0.110285p
C4660 C5_N_btm VSS 68.25825f
C4661 C4_N_btm VSS 47.407547f
C4662 C3_N_btm VSS 27.93639f
C4663 C2_N_btm VSS 21.322378f
C4664 C1_N_btm VSS 16.07949f
C4665 C0_N_btm VSS 14.840141f
C4666 C0_dummy_N_btm VSS 13.25974f
C4667 C0_dummy_P_btm VSS 13.247499f
C4668 C0_P_btm VSS 14.833541f
C4669 C1_P_btm VSS 16.090279f
C4670 C2_P_btm VSS 21.349722f
C4671 C3_P_btm VSS 27.92746f
C4672 C4_P_btm VSS 47.39849f
C4673 C5_P_btm VSS 68.252174f
C4674 C6_P_btm VSS 0.110274p
C4675 C7_P_btm VSS 0.183882p
C4676 C8_P_btm VSS 48.210182f
C4677 C9_P_btm VSS 82.93767f
C4678 C10_P_btm VSS 0.213718p
C4679 a_21753_35474# VSS 0.730911f
C4680 a_19998_34978# VSS 1.75018f
C4681 a_19250_34978# VSS 1.69804f
C4682 EN_VIN_BSTR_N VSS 9.35845f
C4683 a_n217_35014# VSS 1.73445f
C4684 EN_VIN_BSTR_P VSS 9.590905f
C4685 a_n1550_35448# VSS 1.7497f
C4686 a_n2002_35448# VSS 0.735333f
C4687 a_22737_36887# VSS 0.092029f
C4688 a_22737_37285# VSS 0.095943f
C4689 a_22629_37990# VSS 0.468764f
C4690 a_22725_38406# VSS 0.010928f
C4691 a_22629_38406# VSS 0.583873f
C4692 CAL_P VSS 11.759019f
C4693 a_22537_39537# VSS 2.61801f
C4694 a_22889_38993# VSS 0.497542f
C4695 a_22613_38993# VSS 0.357645f
C4696 a_22581_37893# VSS 1.83807f
C4697 a_22527_39145# VSS 2.28699f
C4698 a_22589_40055# VSS 1.23689f
C4699 a_22537_40625# VSS 1.58437f
C4700 a_22589_40599# VSS 1.83268f
C4701 CAL_N VSS 9.176875f
C4702 VDAC_P VSS 1.825184p
C4703 VDAC_N VSS 1.823233p
C4704 a_6886_37412# VSS 3.84933f
C4705 a_3726_37500# VSS 4.51772f
C4706 a_n2302_37690# VSS 0.514517f
C4707 a_n2946_37690# VSS 0.517242f
C4708 a_n3690_37440# VSS 0.548488f
C4709 a_n4334_37440# VSS 0.561497f
C4710 a_8530_39574# VSS 2.76298f
C4711 a_7754_38470# VSS 3.2456f
C4712 VDAC_Ni VSS 3.07545f
C4713 a_7754_38636# VSS 0.353706f
C4714 a_3754_38802# VSS 0.390074f
C4715 a_7754_38968# VSS 0.330037f
C4716 a_3754_39134# VSS 0.401983f
C4717 a_7754_39300# VSS 0.330682f
C4718 a_3754_39466# VSS 0.401172f
C4719 a_7754_39632# VSS 0.340942f
C4720 VDAC_Pi VSS 3.946555f
C4721 a_7754_39964# VSS 2.62481f
C4722 a_3754_39964# VSS 0.671366f
C4723 a_2113_38308# VSS 2.6473f
C4724 a_n2302_37984# VSS 0.483504f
C4725 a_n2946_37984# VSS 0.485942f
C4726 a_n3690_38304# VSS 0.517812f
C4727 a_n4334_38304# VSS 0.529531f
C4728 a_2684_37794# VSS 0.414596f
C4729 a_1107_38525# VSS 0.6415f
C4730 a_n2302_38778# VSS 0.483515f
C4731 a_n2946_38778# VSS 0.485895f
C4732 a_n3690_38528# VSS 0.516979f
C4733 a_n4334_38528# VSS 0.529888f
C4734 a_2112_39137# VSS 0.414404f
C4735 comp_n VSS 0.572075f
C4736 a_1169_39043# VSS 0.615041f
C4737 a_n2302_39072# VSS 0.483504f
C4738 a_n2946_39072# VSS 0.486447f
C4739 a_n3690_39392# VSS 0.517965f
C4740 a_n4334_39392# VSS 0.529516f
C4741 a_1169_39587# VSS 0.633906f
C4742 a_n2302_39866# VSS 0.483537f
C4743 a_n2946_39866# VSS 0.527929f
C4744 a_n3690_39616# VSS 0.574329f
C4745 a_n4334_39616# VSS 0.529903f
C4746 a_n2302_40160# VSS 0.522244f
C4747 a_n4334_40480# VSS 0.578721f
C4748 a_22485_38105# VSS 1.90993f
C4749 a_22775_42308# VSS 0.602116f
C4750 a_21613_42308# VSS 0.725532f
C4751 a_21887_42336# VSS 0.234022f
C4752 a_21335_42336# VSS 0.259392f
C4753 a_20712_42282# VSS 0.349662f
C4754 a_20107_42308# VSS 0.344464f
C4755 a_19647_42308# VSS 0.313304f
C4756 a_19511_42282# VSS 0.751141f
C4757 a_19332_42282# VSS 0.31505f
C4758 a_18907_42674# VSS 0.209311f
C4759 a_18727_42674# VSS 0.233526f
C4760 a_18057_42282# VSS 0.370712f
C4761 a_17531_42308# VSS 0.253358f
C4762 a_17303_42282# VSS 1.19776f
C4763 a_17124_42282# VSS 0.332693f
C4764 a_16522_42674# VSS 0.073862f
C4765 a_15890_42674# VSS 0.180637f
C4766 a_15959_42545# VSS 0.263128f
C4767 a_15803_42450# VSS 0.566963f
C4768 a_15764_42576# VSS 0.298494f
C4769 a_15486_42560# VSS 0.263746f
C4770 a_15051_42282# VSS 0.790649f
C4771 a_14113_42308# VSS 1.42448f
C4772 a_14456_42282# VSS 0.33927f
C4773 a_13575_42558# VSS 0.370369f
C4774 a_13070_42354# VSS 0.222095f
C4775 a_12563_42308# VSS 0.330976f
C4776 a_11551_42558# VSS 0.372919f
C4777 a_11323_42473# VSS 0.253445f
C4778 a_10723_42308# VSS 0.342975f
C4779 a_10533_42308# VSS 0.310658f
C4780 a_9803_42558# VSS 0.370474f
C4781 a_9223_42460# VSS 0.236204f
C4782 a_8791_42308# VSS 0.301f
C4783 a_8685_42308# VSS 0.163732f
C4784 a_8325_42308# VSS 0.316205f
C4785 a_8515_42308# VSS 0.250762f
C4786 a_7963_42308# VSS 0.256292f
C4787 a_7227_42308# VSS 0.359705f
C4788 a_6761_42308# VSS 0.447596f
C4789 a_6171_42473# VSS 0.257988f
C4790 a_5755_42308# VSS 0.314735f
C4791 a_4921_42308# VSS 0.511258f
C4792 a_5379_42460# VSS 0.564806f
C4793 a_5267_42460# VSS 0.204309f
C4794 a_3823_42558# VSS 0.381485f
C4795 a_3318_42354# VSS 0.238394f
C4796 a_2903_42308# VSS 0.340659f
C4797 a_2713_42308# VSS 0.31991f
C4798 a_2351_42308# VSS 0.210162f
C4799 a_2123_42473# VSS 0.21778f
C4800 a_1755_42282# VSS 3.17706f
C4801 a_961_42354# VSS 0.215753f
C4802 a_1184_42692# VSS 0.222827f
C4803 a_1576_42282# VSS 0.327109f
C4804 a_1067_42314# VSS 0.32917f
C4805 a_564_42282# VSS 0.36802f
C4806 a_196_42282# VSS 0.343186f
C4807 a_n473_42460# VSS 0.366068f
C4808 a_n961_42308# VSS 0.328065f
C4809 a_n1329_42308# VSS 0.30898f
C4810 COMP_P VSS 11.200387f
C4811 a_n1736_42282# VSS 0.320711f
C4812 a_n2104_42282# VSS 0.346472f
C4813 a_n2472_42282# VSS 0.335792f
C4814 a_n2840_42282# VSS 0.343361f
C4815 a_22400_42852# VSS 1.97851f
C4816 a_20256_43172# VSS 0.192089f
C4817 a_18504_43218# VSS 0.078212f
C4818 a_14635_42282# VSS 0.336817f
C4819 a_13291_42460# VSS 0.197331f
C4820 a_12800_43218# VSS 0.073862f
C4821 a_11554_42852# VSS 0.073028f
C4822 a_8292_43218# VSS 0.073862f
C4823 a_n2293_42282# VSS 2.62914f
C4824 a_22959_42860# VSS 0.34332f
C4825 a_22223_42860# VSS 0.328988f
C4826 a_22165_42308# VSS 0.354098f
C4827 a_21671_42860# VSS 0.316857f
C4828 a_21195_42852# VSS 0.277519f
C4829 a_21356_42826# VSS 0.304166f
C4830 a_20922_43172# VSS 0.266814f
C4831 a_19987_42826# VSS 0.378798f
C4832 a_19164_43230# VSS 0.264863f
C4833 a_19339_43156# VSS 0.471496f
C4834 a_18599_43230# VSS 0.266382f
C4835 a_18817_42826# VSS 0.182139f
C4836 a_18249_42858# VSS 0.302863f
C4837 a_17333_42852# VSS 0.29982f
C4838 a_18083_42858# VSS 0.578693f
C4839 a_17701_42308# VSS 0.179963f
C4840 a_17595_43084# VSS 0.205109f
C4841 a_16795_42852# VSS 0.362281f
C4842 a_16414_43172# VSS 0.270304f
C4843 a_15567_42826# VSS 0.316627f
C4844 a_15279_43071# VSS 0.248252f
C4845 a_14543_43071# VSS 0.246071f
C4846 a_13460_43230# VSS 0.259861f
C4847 a_13635_43156# VSS 0.7696f
C4848 a_12895_43230# VSS 0.250159f
C4849 a_13113_42826# VSS 0.174096f
C4850 a_12545_42858# VSS 0.287468f
C4851 a_12089_42308# VSS 0.283874f
C4852 a_12379_42858# VSS 0.549229f
C4853 a_10341_42308# VSS 0.317389f
C4854 a_10922_42852# VSS 0.176112f
C4855 a_10991_42826# VSS 0.261283f
C4856 a_10796_42968# VSS 0.29877f
C4857 a_10835_43094# VSS 0.59174f
C4858 a_10518_42984# VSS 0.260322f
C4859 a_10083_42826# VSS 0.762957f
C4860 a_8952_43230# VSS 0.261046f
C4861 a_9127_43156# VSS 0.77314f
C4862 a_8387_43230# VSS 0.255573f
C4863 a_8605_42826# VSS 0.181157f
C4864 a_8037_42858# VSS 0.293593f
C4865 a_7765_42852# VSS 0.252651f
C4866 a_7871_42858# VSS 0.503534f
C4867 a_7227_42852# VSS 0.36607f
C4868 a_5755_42852# VSS 0.383967f
C4869 a_5111_42852# VSS 0.354197f
C4870 a_4520_42826# VSS 0.334784f
C4871 a_3935_42891# VSS 0.26911f
C4872 a_3681_42891# VSS 0.301094f
C4873 a_2905_42968# VSS 0.305424f
C4874 a_2075_43172# VSS 0.537699f
C4875 a_1847_42826# VSS 0.670072f
C4876 a_791_42968# VSS 0.335942f
C4877 a_685_42968# VSS 0.220885f
C4878 a_n1736_43218# VSS 0.073862f
C4879 a_n13_43084# VSS 0.368998f
C4880 a_n1076_43230# VSS 0.263204f
C4881 a_n901_43156# VSS 0.76245f
C4882 a_n1641_43230# VSS 0.256397f
C4883 a_n1423_42826# VSS 0.1805f
C4884 a_n1991_42858# VSS 0.295941f
C4885 a_n1853_43023# VSS 1.30078f
C4886 a_n2157_42858# VSS 0.556569f
C4887 a_n2472_42826# VSS 0.301801f
C4888 a_n2840_42826# VSS 0.327636f
C4889 a_20749_43396# VSS 0.253248f
C4890 a_22959_43396# VSS 0.345439f
C4891 a_22591_43396# VSS 0.335697f
C4892 a_22223_43396# VSS 0.333609f
C4893 a_21855_43396# VSS 0.334538f
C4894 a_19095_43396# VSS 0.132304f
C4895 a_21487_43396# VSS 0.293844f
C4896 a_21259_43561# VSS 0.217667f
C4897 a_16823_43084# VSS 1.23251f
C4898 a_16664_43396# VSS 0.080001f
C4899 a_19700_43370# VSS 0.335707f
C4900 a_19268_43646# VSS 0.242693f
C4901 a_15743_43084# VSS 1.49489f
C4902 a_18783_43370# VSS 0.360096f
C4903 a_18525_43370# VSS 0.361236f
C4904 a_18429_43548# VSS 0.222219f
C4905 a_17324_43396# VSS 0.258017f
C4906 a_17499_43370# VSS 0.762886f
C4907 a_16759_43396# VSS 0.252915f
C4908 a_16977_43638# VSS 0.178776f
C4909 a_16409_43396# VSS 0.290743f
C4910 a_16547_43609# VSS 0.561468f
C4911 a_16243_43396# VSS 0.562369f
C4912 a_16137_43396# VSS 0.635905f
C4913 a_15781_43660# VSS 0.234761f
C4914 a_15681_43442# VSS 0.20154f
C4915 a_12281_43396# VSS 0.691406f
C4916 a_14955_43396# VSS 0.266041f
C4917 a_15095_43370# VSS 0.436411f
C4918 a_14205_43396# VSS 0.2933f
C4919 a_14358_43442# VSS 0.198188f
C4920 a_14579_43548# VSS 0.293668f
C4921 a_13667_43396# VSS 0.265557f
C4922 a_10695_43548# VSS 0.279385f
C4923 a_9803_43646# VSS 0.371929f
C4924 a_3457_43396# VSS 0.379621f
C4925 a_2813_43396# VSS 0.412407f
C4926 a_6452_43396# VSS 0.073862f
C4927 a_9396_43370# VSS 0.338475f
C4928 a_8791_43396# VSS 0.235222f
C4929 a_8147_43396# VSS 0.256103f
C4930 a_7112_43396# VSS 0.256956f
C4931 a_7287_43370# VSS 0.754599f
C4932 a_6547_43396# VSS 0.253718f
C4933 a_6765_43638# VSS 0.174622f
C4934 a_6197_43396# VSS 0.290517f
C4935 a_6293_42852# VSS 0.473619f
C4936 a_6031_43396# VSS 0.541083f
C4937 a_648_43396# VSS 0.231254f
C4938 a_3539_42460# VSS 0.337918f
C4939 a_n1557_42282# VSS 0.870257f
C4940 a_4905_42826# VSS 0.781685f
C4941 a_4699_43561# VSS 0.267684f
C4942 a_4235_43370# VSS 0.33553f
C4943 a_4093_43548# VSS 0.320586f
C4944 a_1756_43548# VSS 0.322408f
C4945 a_1568_43370# VSS 0.63594f
C4946 a_1049_43396# VSS 0.216408f
C4947 a_1209_43370# VSS 0.281234f
C4948 a_458_43396# VSS 0.252302f
C4949 a_n2012_43396# VSS 0.073862f
C4950 a_104_43370# VSS 0.297328f
C4951 a_n447_43370# VSS 0.269574f
C4952 a_n1352_43396# VSS 0.260107f
C4953 a_n1177_43370# VSS 0.478516f
C4954 a_n1917_43396# VSS 0.258245f
C4955 a_n1699_43638# VSS 0.175452f
C4956 a_n2267_43396# VSS 0.297246f
C4957 a_n2129_43609# VSS 1.07965f
C4958 a_n2433_43396# VSS 0.56533f
C4959 a_n2840_43370# VSS 0.316787f
C4960 a_20974_43370# VSS 0.458091f
C4961 a_21381_43940# VSS 0.358332f
C4962 a_19319_43548# VSS 0.229395f
C4963 a_11173_44260# VSS 0.219946f
C4964 a_10555_44260# VSS 0.346315f
C4965 a_22959_43948# VSS 0.341565f
C4966 a_15493_43940# VSS 0.460801f
C4967 a_22223_43948# VSS 0.31992f
C4968 a_21115_43940# VSS 0.204633f
C4969 a_20935_43940# VSS 0.222887f
C4970 a_20623_43914# VSS 0.371294f
C4971 a_20365_43914# VSS 0.359455f
C4972 a_20269_44172# VSS 0.225063f
C4973 a_19862_44208# VSS 0.562087f
C4974 a_19478_44306# VSS 0.278384f
C4975 a_19328_44172# VSS 0.2031f
C4976 a_18451_43940# VSS 0.377396f
C4977 a_18326_43940# VSS 0.276559f
C4978 a_18079_43940# VSS 0.21121f
C4979 a_17973_43940# VSS 0.359917f
C4980 a_17737_43940# VSS 0.386318f
C4981 a_15682_43940# VSS 1.9643f
C4982 a_14955_43940# VSS 0.365393f
C4983 a_13483_43940# VSS 0.376442f
C4984 a_12429_44172# VSS 0.389129f
C4985 a_11750_44172# VSS 0.221782f
C4986 a_10807_43548# VSS 0.451031f
C4987 a_10949_43914# VSS 0.257331f
C4988 a_10729_43914# VSS 0.34307f
C4989 a_10405_44172# VSS 0.142993f
C4990 a_9672_43914# VSS 0.323006f
C4991 a_9028_43914# VSS 0.398016f
C4992 a_8333_44056# VSS 0.331632f
C4993 a_3499_42826# VSS 0.380221f
C4994 a_n1644_44306# VSS 0.080042f
C4995 a_7845_44172# VSS 0.239173f
C4996 a_7542_44172# VSS 0.283767f
C4997 a_7281_43914# VSS 0.271121f
C4998 a_6453_43914# VSS 0.26639f
C4999 a_5663_43940# VSS 0.488325f
C5000 a_5495_43940# VSS 0.212229f
C5001 a_5013_44260# VSS 0.279924f
C5002 a_5244_44056# VSS 0.216368f
C5003 a_3905_42865# VSS 0.9893f
C5004 a_3600_43914# VSS 0.422049f
C5005 a_2998_44172# VSS 0.503048f
C5006 a_2889_44172# VSS 0.217034f
C5007 a_2675_43914# VSS 0.2974f
C5008 a_895_43940# VSS 0.237723f
C5009 a_2479_44172# VSS 0.817462f
C5010 a_2127_44172# VSS 0.517911f
C5011 a_453_43940# VSS 0.285192f
C5012 a_1414_42308# VSS 1.07452f
C5013 a_1467_44172# VSS 0.187431f
C5014 a_1115_44172# VSS 0.52592f
C5015 a_644_44056# VSS 0.227493f
C5016 a_175_44278# VSS 0.226801f
C5017 a_n984_44318# VSS 0.27358f
C5018 a_n809_44244# VSS 0.785904f
C5019 a_n1549_44318# VSS 0.264547f
C5020 a_n1331_43914# VSS 0.185087f
C5021 a_n1899_43946# VSS 0.299008f
C5022 a_n1761_44111# VSS 0.392075f
C5023 a_n2065_43946# VSS 0.658803f
C5024 a_n2472_43914# VSS 0.3103f
C5025 a_n2840_43914# VSS 0.345355f
C5026 a_22959_44484# VSS 0.343897f
C5027 a_22591_44484# VSS 0.315361f
C5028 a_22485_44484# VSS 0.590119f
C5029 a_20512_43084# VSS 0.561552f
C5030 a_22315_44484# VSS 0.238239f
C5031 a_21398_44850# VSS 0.073862f
C5032 a_18579_44172# VSS 0.812679f
C5033 a_19279_43940# VSS 1.69633f
C5034 a_20766_44850# VSS 0.177656f
C5035 a_20835_44721# VSS 0.260406f
C5036 a_20679_44626# VSS 0.58931f
C5037 a_20640_44752# VSS 0.296084f
C5038 a_20362_44736# VSS 0.255907f
C5039 a_20159_44458# VSS 0.483669f
C5040 a_19615_44636# VSS 0.238459f
C5041 a_19006_44850# VSS 0.073862f
C5042 a_14673_44172# VSS 0.290001f
C5043 a_11541_44484# VSS 0.139071f
C5044 a_15433_44458# VSS 0.301508f
C5045 a_14815_43914# VSS 0.445698f
C5046 a_9159_44484# VSS 0.158168f
C5047 a_10617_44484# VSS 0.119149f
C5048 a_5708_44484# VSS 0.231649f
C5049 a_3363_44484# VSS 0.27629f
C5050 a_556_44484# VSS 0.201935f
C5051 a_8375_44464# VSS 0.211867f
C5052 a_7640_43914# VSS 0.542377f
C5053 a_6109_44484# VSS 0.648821f
C5054 a_n23_44458# VSS 0.278255f
C5055 a_n2012_44484# VSS 0.080001f
C5056 a_18989_43940# VSS 0.423174f
C5057 a_18374_44850# VSS 0.179731f
C5058 a_18443_44721# VSS 0.253971f
C5059 a_18287_44626# VSS 0.507939f
C5060 a_18248_44752# VSS 0.294917f
C5061 a_17970_44736# VSS 0.26161f
C5062 a_17767_44458# VSS 0.474097f
C5063 a_16979_44734# VSS 0.363013f
C5064 a_14539_43914# VSS 1.18088f
C5065 a_16112_44458# VSS 0.326339f
C5066 a_15004_44636# VSS 0.254778f
C5067 a_13720_44458# VSS 0.403209f
C5068 a_13076_44458# VSS 0.38829f
C5069 a_12883_44458# VSS 0.287544f
C5070 a_12607_44458# VSS 0.499331f
C5071 a_8975_43940# VSS 0.652857f
C5072 a_10057_43914# VSS 0.654189f
C5073 a_10440_44484# VSS 0.210149f
C5074 a_10334_44484# VSS 0.210217f
C5075 a_10157_44484# VSS 0.208916f
C5076 a_9838_44484# VSS 0.276258f
C5077 a_5883_43914# VSS 0.792825f
C5078 a_8701_44490# VSS 0.358059f
C5079 a_8103_44636# VSS 0.340824f
C5080 a_6298_44484# VSS 1.93814f
C5081 a_5518_44484# VSS 0.242995f
C5082 a_5343_44458# VSS 1.28071f
C5083 a_4743_44484# VSS 0.327178f
C5084 a_n699_43396# VSS 1.82142f
C5085 a_2779_44458# VSS 0.532137f
C5086 a_949_44458# VSS 1.97734f
C5087 a_742_44458# VSS 1.02263f
C5088 a_n452_44636# VSS 0.254732f
C5089 a_n1352_44484# VSS 0.269853f
C5090 a_n1177_44458# VSS 0.493891f
C5091 a_n1917_44484# VSS 0.280038f
C5092 a_n1699_44726# VSS 0.197478f
C5093 a_n2267_44484# VSS 0.308908f
C5094 a_n2129_44697# VSS 0.307327f
C5095 a_n2433_44484# VSS 0.679598f
C5096 a_n2840_44458# VSS 0.316322f
C5097 a_16237_45028# VSS 0.017944f
C5098 a_20193_45348# VSS 1.70015f
C5099 a_19113_45348# VSS 0.367248f
C5100 a_22959_45036# VSS 0.345334f
C5101 a_22223_45036# VSS 0.354178f
C5102 a_11827_44484# VSS 1.28091f
C5103 a_21359_45002# VSS 0.397791f
C5104 a_21101_45002# VSS 0.35202f
C5105 a_21005_45260# VSS 0.212992f
C5106 a_20567_45036# VSS 0.31908f
C5107 a_18494_42460# VSS 1.15626f
C5108 a_19778_44110# VSS 0.599421f
C5109 a_18911_45144# VSS 0.307008f
C5110 a_18587_45118# VSS 0.214925f
C5111 a_18315_45260# VSS 0.334834f
C5112 a_17719_45144# VSS 0.331229f
C5113 a_17613_45144# VSS 0.244364f
C5114 a_17023_45118# VSS 0.20885f
C5115 a_16922_45042# VSS 0.818675f
C5116 a_8560_45348# VSS 0.185033f
C5117 a_2304_45348# VSS 0.182367f
C5118 a_626_44172# VSS 0.67926f
C5119 a_375_42282# VSS 0.447027f
C5120 a_16751_45260# VSS 0.316547f
C5121 a_16019_45002# VSS 0.25377f
C5122 a_15595_45028# VSS 0.214111f
C5123 a_15415_45028# VSS 0.221991f
C5124 a_14797_45144# VSS 0.249222f
C5125 a_14537_43396# VSS 1.73146f
C5126 a_14180_45002# VSS 0.327485f
C5127 a_13777_45326# VSS 0.272936f
C5128 a_13556_45296# VSS 1.01916f
C5129 a_9482_43914# VSS 3.42654f
C5130 a_13348_45260# VSS 0.243533f
C5131 a_13159_45002# VSS 0.265737f
C5132 a_13017_45260# VSS 0.362048f
C5133 a_11963_45334# VSS 0.226884f
C5134 a_11787_45002# VSS 0.212512f
C5135 a_10951_45334# VSS 0.228638f
C5136 a_10775_45002# VSS 0.204487f
C5137 a_8953_45002# VSS 1.94941f
C5138 a_8191_45002# VSS 0.325964f
C5139 a_7705_45326# VSS 0.273009f
C5140 a_6709_45028# VSS 0.354418f
C5141 a_7229_43940# VSS 0.786182f
C5142 a_7276_45260# VSS 0.251523f
C5143 a_5205_44484# VSS 0.546179f
C5144 a_6431_45366# VSS 0.233718f
C5145 a_5691_45260# VSS 0.370273f
C5146 a_4927_45028# VSS 0.520892f
C5147 a_5111_44636# VSS 3.44603f
C5148 a_5147_45002# VSS 0.803306f
C5149 a_4558_45348# VSS 0.446148f
C5150 a_4574_45260# VSS 0.208274f
C5151 a_3429_45260# VSS 0.274034f
C5152 a_3065_45002# VSS 0.864786f
C5153 a_2680_45002# VSS 0.321351f
C5154 a_2382_45260# VSS 1.03422f
C5155 a_2274_45254# VSS 0.187307f
C5156 a_1667_45002# VSS 0.345429f
C5157 a_327_44734# VSS 0.419171f
C5158 a_n37_45144# VSS 0.321746f
C5159 a_n143_45144# VSS 0.209896f
C5160 a_n467_45028# VSS 0.311181f
C5161 a_n967_45348# VSS 0.453992f
C5162 en_comp VSS 7.84057f
C5163 a_n745_45366# VSS 0.257282f
C5164 a_n2109_45247# VSS 0.252392f
C5165 a_n2293_45010# VSS 0.614925f
C5166 a_n2472_45002# VSS 0.298945f
C5167 a_n2661_45010# VSS 0.839496f
C5168 a_n2840_45002# VSS 0.340687f
C5169 a_22959_45572# VSS 0.34535f
C5170 a_22591_45572# VSS 0.363695f
C5171 a_22223_45572# VSS 0.334964f
C5172 a_21513_45002# VSS 0.669089f
C5173 a_20528_45572# VSS 0.073082f
C5174 a_21188_45572# VSS 0.284872f
C5175 a_21363_45546# VSS 0.515994f
C5176 a_20623_45572# VSS 0.256236f
C5177 a_20841_45814# VSS 0.180037f
C5178 a_20273_45572# VSS 0.288513f
C5179 a_20107_45572# VSS 0.541125f
C5180 a_17668_45572# VSS 0.217142f
C5181 a_18596_45572# VSS 0.073862f
C5182 a_19256_45572# VSS 0.257674f
C5183 a_19431_45546# VSS 0.487121f
C5184 a_18691_45572# VSS 0.255356f
C5185 a_18909_45814# VSS 0.178658f
C5186 a_18341_45572# VSS 0.291608f
C5187 a_18479_45785# VSS 1.15946f
C5188 a_18175_45572# VSS 0.516981f
C5189 a_16147_45260# VSS 0.506229f
C5190 a_16020_45572# VSS 0.073862f
C5191 a_17478_45572# VSS 0.232341f
C5192 a_15861_45028# VSS 0.449058f
C5193 a_16680_45572# VSS 0.258674f
C5194 a_16855_45546# VSS 0.471485f
C5195 a_16115_45572# VSS 0.253972f
C5196 a_16333_45814# VSS 0.178165f
C5197 a_15765_45572# VSS 0.291326f
C5198 a_15903_45785# VSS 0.4164f
C5199 a_15599_45572# VSS 0.50233f
C5200 a_15037_45618# VSS 0.209713f
C5201 a_11136_45572# VSS 0.17156f
C5202 a_9159_45572# VSS 0.151638f
C5203 a_8192_45572# VSS 0.17002f
C5204 a_11682_45822# VSS 0.010374f
C5205 a_10907_45822# VSS 0.547001f
C5206 a_10210_45822# VSS 0.012573f
C5207 a_15143_45578# VSS 0.315994f
C5208 a_14495_45572# VSS 0.325874f
C5209 a_13249_42308# VSS 1.08648f
C5210 a_13904_45546# VSS 0.327907f
C5211 a_13527_45546# VSS 0.245514f
C5212 a_13163_45724# VSS 0.180841f
C5213 a_12791_45546# VSS 0.237787f
C5214 a_12427_45724# VSS 0.190531f
C5215 a_11962_45724# VSS 0.218739f
C5216 a_11652_45724# VSS 0.258015f
C5217 a_11525_45546# VSS 0.346102f
C5218 a_11322_45546# VSS 0.62914f
C5219 a_10490_45724# VSS 0.972668f
C5220 a_8746_45002# VSS 0.547616f
C5221 a_10180_45724# VSS 0.281135f
C5222 a_10053_45546# VSS 0.373668f
C5223 a_9049_44484# VSS 0.249658f
C5224 a_7499_43078# VSS 3.22587f
C5225 a_8568_45546# VSS 0.317032f
C5226 a_8162_45546# VSS 0.376225f
C5227 a_7230_45938# VSS 0.078992f
C5228 a_4880_45572# VSS 0.182839f
C5229 a_3775_45552# VSS 0.209244f
C5230 a_7227_45028# VSS 0.439395f
C5231 a_6598_45938# VSS 0.185967f
C5232 a_6667_45809# VSS 0.264656f
C5233 a_6511_45714# VSS 0.647716f
C5234 a_6472_45840# VSS 0.310105f
C5235 a_6194_45824# VSS 0.2717f
C5236 a_5907_45546# VSS 0.592148f
C5237 a_5263_45724# VSS 0.250928f
C5238 a_4099_45572# VSS 0.33915f
C5239 a_2277_45546# VSS 0.303704f
C5240 a_1609_45822# VSS 0.5528f
C5241 a_509_45822# VSS 0.010571f
C5242 a_n23_45546# VSS 0.281189f
C5243 a_n356_45724# VSS 0.32306f
C5244 a_3503_45724# VSS 0.322319f
C5245 a_3316_45546# VSS 0.336134f
C5246 a_3218_45724# VSS 0.379893f
C5247 a_2957_45546# VSS 0.276358f
C5248 a_1848_45724# VSS 0.245258f
C5249 a_997_45618# VSS 0.248122f
C5250 a_310_45028# VSS 0.207165f
C5251 a_n1099_45572# VSS 0.339525f
C5252 a_380_45546# VSS 0.337145f
C5253 a_n452_45724# VSS 0.253614f
C5254 a_n863_45724# VSS 3.49288f
C5255 a_n1079_45724# VSS 0.289271f
C5256 a_n2472_45546# VSS 0.340801f
C5257 a_n2840_45546# VSS 0.344757f
C5258 a_19240_46482# VSS 0.073862f
C5259 a_16375_45002# VSS 1.44161f
C5260 a_14180_46482# VSS 0.073862f
C5261 a_12638_46436# VSS 0.162178f
C5262 a_12379_46436# VSS 0.275423f
C5263 a_10586_45546# VSS 0.542658f
C5264 a_8034_45724# VSS 0.299594f
C5265 a_5066_45546# VSS 0.436834f
C5266 a_2981_46116# VSS 0.091491f
C5267 a_n1736_46482# VSS 0.07565f
C5268 a_22959_46124# VSS 0.345245f
C5269 a_22223_46124# VSS 0.354467f
C5270 a_21137_46414# VSS 0.340736f
C5271 a_20708_46348# VSS 0.268156f
C5272 a_19900_46494# VSS 0.26164f
C5273 a_20075_46420# VSS 0.475201f
C5274 a_19335_46494# VSS 0.260378f
C5275 a_19553_46090# VSS 0.179968f
C5276 a_18985_46122# VSS 0.297132f
C5277 a_18819_46122# VSS 0.545109f
C5278 a_17957_46116# VSS 0.309446f
C5279 a_18189_46348# VSS 0.296366f
C5280 a_17715_44484# VSS 0.55862f
C5281 a_17583_46090# VSS 0.307562f
C5282 a_15682_46116# VSS 1.96743f
C5283 a_14840_46494# VSS 0.263367f
C5284 a_15015_46420# VSS 0.472948f
C5285 a_14275_46494# VSS 0.258968f
C5286 a_14493_46090# VSS 0.176122f
C5287 a_13925_46122# VSS 0.294602f
C5288 a_13759_46122# VSS 0.518292f
C5289 a_13351_46090# VSS 0.304427f
C5290 a_12594_46348# VSS 0.284494f
C5291 a_12005_46116# VSS 0.381711f
C5292 a_11387_46155# VSS 0.260117f
C5293 a_11133_46155# VSS 0.299642f
C5294 a_11189_46129# VSS 0.32558f
C5295 a_10355_46116# VSS 0.290668f
C5296 a_9823_46155# VSS 0.261206f
C5297 a_9569_46155# VSS 0.304755f
C5298 a_9625_46129# VSS 0.369694f
C5299 a_8953_45546# VSS 1.00397f
C5300 a_8199_44636# VSS 2.29742f
C5301 a_8349_46414# VSS 0.273442f
C5302 a_8016_46348# VSS 0.539696f
C5303 a_7920_46348# VSS 0.269852f
C5304 a_6419_46155# VSS 0.273686f
C5305 a_6165_46155# VSS 0.303989f
C5306 a_5497_46414# VSS 0.304684f
C5307 a_5204_45822# VSS 0.338817f
C5308 a_5164_46348# VSS 0.419282f
C5309 a_5068_46348# VSS 0.25855f
C5310 a_4704_46090# VSS 0.296767f
C5311 a_4419_46090# VSS 0.357571f
C5312 a_3699_46348# VSS 0.226584f
C5313 a_3147_46376# VSS 0.52775f
C5314 a_2804_46116# VSS 0.222855f
C5315 a_2698_46116# VSS 0.215567f
C5316 a_2521_46116# VSS 0.220999f
C5317 a_167_45260# VSS 1.32487f
C5318 a_2202_46116# VSS 0.273578f
C5319 a_1823_45246# VSS 2.36307f
C5320 a_1138_42852# VSS 0.456566f
C5321 a_1176_45822# VSS 0.278365f
C5322 a_1208_46090# VSS 0.348206f
C5323 a_805_46414# VSS 0.27506f
C5324 a_472_46348# VSS 0.32751f
C5325 a_376_46348# VSS 0.285607f
C5326 a_n1076_46494# VSS 0.262147f
C5327 a_n901_46420# VSS 0.762523f
C5328 a_n1641_46494# VSS 0.256945f
C5329 a_n1423_46090# VSS 0.176189f
C5330 a_n1991_46122# VSS 0.305274f
C5331 a_n1853_46287# VSS 0.341802f
C5332 a_n2157_46122# VSS 0.525314f
C5333 a_n2472_46090# VSS 0.290925f
C5334 a_n2840_46090# VSS 0.340313f
C5335 a_22959_46660# VSS 0.338967f
C5336 a_22591_46660# VSS 0.292786f
C5337 a_11415_45002# VSS 1.63684f
C5338 a_20202_43084# VSS 1.05073f
C5339 a_22365_46825# VSS 0.208388f
C5340 a_18280_46660# VSS 0.29316f
C5341 a_17639_46660# VSS 0.308795f
C5342 a_20528_46660# VSS 0.07565f
C5343 a_22000_46634# VSS 0.295895f
C5344 a_21188_46660# VSS 0.261124f
C5345 a_21363_46634# VSS 0.488515f
C5346 a_20623_46660# VSS 0.258464f
C5347 a_20841_46902# VSS 0.180869f
C5348 a_20273_46660# VSS 0.309206f
C5349 a_20411_46873# VSS 0.393328f
C5350 a_20107_46660# VSS 0.575208f
C5351 a_19123_46287# VSS 0.477642f
C5352 a_18285_46348# VSS 0.577053f
C5353 a_17339_46660# VSS 0.927636f
C5354 a_16721_46634# VSS 0.305539f
C5355 a_16388_46812# VSS 1.42609f
C5356 a_13059_46348# VSS 2.36107f
C5357 a_14513_46634# VSS 0.29862f
C5358 a_14180_46812# VSS 0.368158f
C5359 a_14035_46660# VSS 0.322858f
C5360 a_13885_46660# VSS 0.297377f
C5361 a_12156_46660# VSS 0.074642f
C5362 a_19466_46812# VSS 0.675335f
C5363 a_19333_46634# VSS 0.289568f
C5364 a_18834_46812# VSS 0.198054f
C5365 a_17609_46634# VSS 0.205547f
C5366 a_16292_46812# VSS 0.271203f
C5367 a_15559_46634# VSS 0.394779f
C5368 a_15368_46634# VSS 0.278142f
C5369 a_14976_45028# VSS 0.479565f
C5370 a_15009_46634# VSS 0.270859f
C5371 a_14084_46812# VSS 0.251005f
C5372 a_13607_46688# VSS 0.218935f
C5373 a_12816_46660# VSS 0.260317f
C5374 a_12991_46634# VSS 0.475827f
C5375 a_12251_46660# VSS 0.270927f
C5376 a_12469_46902# VSS 0.193369f
C5377 a_11901_46660# VSS 0.303844f
C5378 a_11813_46116# VSS 0.563718f
C5379 a_11735_46660# VSS 0.520568f
C5380 a_11186_47026# VSS 0.078586f
C5381 a_8270_45546# VSS 0.779033f
C5382 a_7832_46660# VSS 0.073862f
C5383 a_6969_46634# VSS 0.289597f
C5384 a_6755_46942# VSS 3.33348f
C5385 a_10249_46116# VSS 0.414443f
C5386 a_10554_47026# VSS 0.191251f
C5387 a_10623_46897# VSS 0.283572f
C5388 a_10467_46802# VSS 0.523954f
C5389 a_10428_46928# VSS 0.314538f
C5390 a_10150_46912# VSS 0.276624f
C5391 a_9863_46634# VSS 0.607398f
C5392 a_8492_46660# VSS 0.283316f
C5393 a_8667_46634# VSS 0.596387f
C5394 a_7927_46660# VSS 0.269867f
C5395 a_8145_46902# VSS 0.179735f
C5396 a_7577_46660# VSS 0.314978f
C5397 a_7715_46873# VSS 0.546182f
C5398 a_7411_46660# VSS 0.532412f
C5399 a_5257_43370# VSS 1.42323f
C5400 a_5072_46660# VSS 0.073862f
C5401 a_6540_46812# VSS 0.248814f
C5402 a_5732_46660# VSS 0.260482f
C5403 a_5907_46634# VSS 0.473347f
C5404 a_5167_46660# VSS 0.263586f
C5405 a_5385_46902# VSS 0.17737f
C5406 a_4817_46660# VSS 0.296797f
C5407 a_4955_46873# VSS 0.365781f
C5408 a_4651_46660# VSS 0.548065f
C5409 a_3877_44458# VSS 2.8543f
C5410 a_2864_46660# VSS 0.080001f
C5411 a_3524_46660# VSS 0.267612f
C5412 a_3699_46634# VSS 0.499647f
C5413 a_2959_46660# VSS 0.261026f
C5414 a_3177_46902# VSS 0.184239f
C5415 a_2609_46660# VSS 0.302878f
C5416 a_2443_46660# VSS 0.657702f
C5417 a_n2661_46098# VSS 2.05975f
C5418 a_1799_45572# VSS 0.30194f
C5419 a_491_47026# VSS 0.010533f
C5420 a_288_46660# VSS 0.075217f
C5421 a_1983_46706# VSS 0.205951f
C5422 a_948_46660# VSS 0.263413f
C5423 a_1123_46634# VSS 0.776627f
C5424 a_383_46660# VSS 0.269735f
C5425 a_601_46902# VSS 0.192316f
C5426 a_33_46660# VSS 0.309712f
C5427 a_171_46873# VSS 0.579977f
C5428 a_n133_46660# VSS 0.576523f
C5429 a_n1021_46688# VSS 0.271211f
C5430 a_n2104_46634# VSS 0.340006f
C5431 a_n2472_46634# VSS 0.323981f
C5432 a_n2840_46634# VSS 0.328049f
C5433 a_20916_46384# VSS 0.827544f
C5434 a_20843_47204# VSS 0.121976f
C5435 a_19594_46812# VSS 0.277274f
C5436 a_19321_45002# VSS 1.15234f
C5437 a_5807_45002# VSS 2.5828f
C5438 a_15928_47570# VSS 0.075455f
C5439 a_12891_46348# VSS 1.22195f
C5440 a_11309_47204# VSS 0.423399f
C5441 a_9804_47204# VSS 0.528639f
C5442 a_8128_46384# VSS 0.573494f
C5443 a_2747_46873# VSS 0.287894f
C5444 a_22959_47212# VSS 0.322938f
C5445 SMPL_ON_N VSS 7.32671f
C5446 a_22731_47423# VSS 0.227778f
C5447 a_22223_47212# VSS 0.332189f
C5448 a_12465_44636# VSS 5.61685f
C5449 a_21811_47423# VSS 0.23358f
C5450 a_21496_47436# VSS 0.249536f
C5451 a_21177_47436# VSS 0.223524f
C5452 a_20990_47178# VSS 0.224581f
C5453 a_20894_47436# VSS 0.233111f
C5454 a_19787_47423# VSS 0.258015f
C5455 a_19386_47436# VSS 0.209882f
C5456 a_18597_46090# VSS 2.82344f
C5457 a_18780_47178# VSS 0.319719f
C5458 a_18479_47436# VSS 1.19826f
C5459 a_18143_47464# VSS 0.579061f
C5460 a_17591_47464# VSS 0.576556f
C5461 a_16588_47582# VSS 0.263715f
C5462 a_16763_47508# VSS 0.587861f
C5463 a_16023_47582# VSS 0.264352f
C5464 a_16241_47178# VSS 0.18232f
C5465 a_15673_47210# VSS 0.315684f
C5466 a_15811_47375# VSS 0.349499f
C5467 a_15507_47210# VSS 0.556554f
C5468 a_14955_47212# VSS 0.358339f
C5469 a_14311_47204# VSS 0.248858f
C5470 a_13487_47204# VSS 0.643275f
C5471 a_13381_47204# VSS 0.225132f
C5472 a_11459_47204# VSS 0.553679f
C5473 a_9313_45822# VSS 1.04727f
C5474 a_11031_47542# VSS 0.247302f
C5475 a_9863_47436# VSS 0.265619f
C5476 a_9067_47204# VSS 0.606182f
C5477 a_6575_47204# VSS 0.798434f
C5478 a_7903_47542# VSS 0.258657f
C5479 a_7227_47204# VSS 0.610401f
C5480 a_6851_47204# VSS 0.346433f
C5481 a_6491_46660# VSS 0.343406f
C5482 a_6545_47178# VSS 0.597936f
C5483 a_5815_47464# VSS 0.594449f
C5484 a_5129_47502# VSS 0.361487f
C5485 a_4700_47436# VSS 0.271201f
C5486 a_4007_47204# VSS 0.628996f
C5487 a_3815_47204# VSS 0.440491f
C5488 a_3785_47178# VSS 0.541893f
C5489 a_3381_47502# VSS 0.320926f
C5490 a_3160_47472# VSS 0.607125f
C5491 a_2905_45572# VSS 0.47073f
C5492 a_2952_47436# VSS 0.275026f
C5493 a_2553_47502# VSS 0.294118f
C5494 a_2124_47436# VSS 0.276508f
C5495 a_1431_47204# VSS 0.595895f
C5496 a_1239_47204# VSS 0.33333f
C5497 a_1209_47178# VSS 0.474725f
C5498 a_327_47204# VSS 0.581187f
C5499 a_n785_47204# VSS 0.361759f
C5500 a_n23_47502# VSS 0.278861f
C5501 a_n746_45260# VSS 0.993718f
C5502 a_n452_47436# VSS 0.28781f
C5503 a_n815_47178# VSS 0.513835f
C5504 a_n1605_47204# VSS 0.250546f
C5505 SMPL_ON_P VSS 12.32981f
C5506 a_n1920_47178# VSS 0.310881f
C5507 a_n2288_47178# VSS 0.346995f
C5508 a_n2497_47436# VSS 2.31207f
C5509 a_n2833_47464# VSS 0.602779f
C5510 a_5342_30871.t0 VSS 0.051002f
C5511 a_5342_30871.t7 VSS 0.04948f
C5512 a_5342_30871.t8 VSS 0.079338f
C5513 a_5342_30871.n0 VSS 0.18907f
C5514 a_5342_30871.t4 VSS 0.671533f
C5515 a_5342_30871.t5 VSS 0.691556f
C5516 a_5342_30871.n1 VSS 0.865919f
C5517 a_5342_30871.t9 VSS 0.671533f
C5518 a_5342_30871.t6 VSS 0.691556f
C5519 a_5342_30871.n2 VSS 0.901731f
C5520 a_5342_30871.n3 VSS 10.8884f
C5521 a_5342_30871.n4 VSS 5.4481f
C5522 a_5342_30871.t3 VSS 0.033152f
C5523 a_5342_30871.t2 VSS 0.033152f
C5524 a_5342_30871.n5 VSS 0.066303f
C5525 a_5342_30871.n6 VSS 0.464133f
C5526 a_5342_30871.n7 VSS 0.153042f
C5527 a_5342_30871.t1 VSS 0.051002f
C5528 C8_P_btm.t0 VSS 0.1469f
C5529 C8_P_btm.t1 VSS 0.1469f
C5530 C8_P_btm.n0 VSS 0.453952f
C5531 C8_P_btm.t2 VSS 0.1469f
C5532 C8_P_btm.t3 VSS 0.1469f
C5533 C8_P_btm.n1 VSS 0.468327f
C5534 C8_P_btm.n2 VSS 1.81139f
C5535 C8_P_btm.t6 VSS 0.167162f
C5536 C8_P_btm.t7 VSS 0.167162f
C5537 C8_P_btm.n3 VSS 0.847137f
C5538 C8_P_btm.n4 VSS 1.20098f
C5539 C8_P_btm.t9 VSS 0.167162f
C5540 C8_P_btm.t8 VSS 0.167162f
C5541 C8_P_btm.n5 VSS 0.853379f
C5542 C8_P_btm.n6 VSS 0.927507f
C5543 C8_P_btm.t5 VSS 0.041791f
C5544 C8_P_btm.t4 VSS 0.041791f
C5545 C8_P_btm.n7 VSS 0.156641f
C5546 C8_P_btm.n8 VSS 2.62073f
C5547 C8_P_btm.n9 VSS 2.45049f
C5548 C8_P_btm.n10 VSS 1.08519f
C5549 C8_P_btm.n11 VSS 1.08899f
C5550 C8_P_btm.n12 VSS 1.08899f
C5551 C8_P_btm.n13 VSS 1.08519f
C5552 C8_P_btm.n14 VSS 1.08899f
C5553 C8_P_btm.n15 VSS 1.08899f
C5554 C8_P_btm.n16 VSS 1.08899f
C5555 C8_P_btm.n17 VSS 1.08899f
C5556 C8_P_btm.n18 VSS 1.08519f
C5557 C8_P_btm.n19 VSS 1.08899f
C5558 C8_P_btm.n20 VSS 1.08899f
C5559 C8_P_btm.n21 VSS 1.08519f
C5560 C8_P_btm.n22 VSS 1.08899f
C5561 C8_P_btm.n23 VSS 1.08899f
C5562 C8_P_btm.n24 VSS 1.08899f
C5563 C8_P_btm.n25 VSS 1.05133f
C5564 C8_P_btm.n26 VSS 1.08899f
C5565 C8_P_btm.n27 VSS 1.08899f
C5566 C8_P_btm.n28 VSS 1.08899f
C5567 C8_P_btm.n29 VSS 1.08899f
C5568 C8_P_btm.n30 VSS 1.08899f
C5569 C8_P_btm.n31 VSS 1.48645f
C5570 C8_P_btm.n32 VSS 1.08899f
C5571 C8_P_btm.n33 VSS 0.801269f
C5572 C8_P_btm.n34 VSS 1.08899f
C5573 C8_P_btm.n35 VSS 1.08899f
C5574 C8_P_btm.n36 VSS 1.08899f
C5575 C8_P_btm.n37 VSS 1.08899f
C5576 C8_P_btm.n38 VSS 1.08899f
C5577 C8_P_btm.n39 VSS 1.55314f
C5578 C8_P_btm.n40 VSS 1.70585f
C5579 C8_P_btm.n41 VSS 1.3116f
C5580 C8_P_btm.n42 VSS 1.08519f
C5581 C8_P_btm.n43 VSS 1.08519f
C5582 C8_P_btm.n44 VSS 1.08899f
C5583 C8_P_btm.n45 VSS 1.08519f
C5584 C8_P_btm.n46 VSS 1.08519f
C5585 C8_P_btm.n47 VSS 1.08519f
C5586 C8_P_btm.n48 VSS 1.08519f
C5587 C8_P_btm.n49 VSS 1.08519f
C5588 C8_P_btm.n50 VSS 1.08519f
C5589 C8_P_btm.n51 VSS 1.39409f
C5590 C8_P_btm.n52 VSS 4.75265f
C5591 C8_P_btm.n53 VSS 3.37111f
C5592 C8_P_btm.n54 VSS 1.08899f
C5593 C8_P_btm.n55 VSS 1.08899f
C5594 C8_P_btm.n56 VSS 1.08899f
C5595 C8_P_btm.n57 VSS 1.08899f
C5596 C8_P_btm.n58 VSS 1.08899f
C5597 C8_P_btm.n59 VSS 1.08899f
C5598 C8_P_btm.n60 VSS 1.08899f
C5599 C8_P_btm.n61 VSS 1.08899f
C5600 C8_P_btm.n62 VSS 1.08899f
C5601 C8_P_btm.n63 VSS 1.08899f
C5602 C8_P_btm.n64 VSS 1.08899f
C5603 C8_P_btm.n65 VSS 1.08519f
C5604 C8_P_btm.n66 VSS 1.08519f
C5605 C8_P_btm.n67 VSS 1.08519f
C5606 C8_P_btm.n68 VSS 1.08899f
C5607 C8_P_btm.n69 VSS 1.08899f
C5608 C8_P_btm.n70 VSS 1.08899f
C5609 C8_P_btm.n71 VSS 1.08899f
C5610 C8_P_btm.n72 VSS 1.08899f
C5611 C8_P_btm.n73 VSS 1.08899f
C5612 C8_P_btm.n74 VSS 1.08899f
C5613 C8_P_btm.n75 VSS 1.08899f
C5614 C8_P_btm.n76 VSS 0.801269f
C5615 C8_P_btm.n77 VSS 0.801269f
C5616 C8_P_btm.n78 VSS 1.08899f
C5617 C8_P_btm.n79 VSS 0.801269f
C5618 C8_P_btm.n80 VSS 1.08899f
C5619 C8_P_btm.n81 VSS 1.08899f
C5620 C8_P_btm.n82 VSS 1.08899f
C5621 C8_P_btm.n83 VSS 1.3691f
C5622 C8_P_btm.n84 VSS 1.08899f
C5623 C8_P_btm.n85 VSS 1.08899f
C5624 C8_P_btm.n86 VSS 0.801269f
C5625 C8_P_btm.n87 VSS 1.08899f
C5626 C8_P_btm.n88 VSS 0.801269f
C5627 C8_P_btm.n89 VSS 1.08899f
C5628 C8_P_btm.n90 VSS 1.08899f
C5629 C8_P_btm.n91 VSS 1.08899f
C5630 C8_P_btm.n92 VSS 1.3691f
C5631 C8_P_btm.n93 VSS 1.08899f
C5632 C8_P_btm.n94 VSS 1.08899f
C5633 C8_P_btm.n95 VSS 0.801269f
C5634 C8_P_btm.n96 VSS 1.08899f
C5635 C8_P_btm.n97 VSS 0.801269f
C5636 C8_P_btm.n98 VSS 1.08899f
C5637 C8_P_btm.n99 VSS 1.08899f
C5638 C8_P_btm.n100 VSS 1.08899f
C5639 C8_P_btm.n101 VSS 1.08899f
C5640 C8_P_btm.n102 VSS 1.08899f
C5641 C8_P_btm.n103 VSS 1.08519f
C5642 C8_P_btm.n104 VSS 1.08899f
C5643 C8_P_btm.n105 VSS 1.08899f
C5644 C8_P_btm.n106 VSS 1.08899f
C5645 C8_P_btm.n107 VSS 1.08899f
C5646 C8_P_btm.n108 VSS 0.801269f
C5647 C8_P_btm.n109 VSS 0.801269f
C5648 C8_P_btm.n110 VSS 1.08899f
C5649 C8_P_btm.n111 VSS 1.08899f
C5650 C8_P_btm.n112 VSS 1.08899f
C5651 C8_P_btm.n113 VSS 0.801269f
C5652 C8_P_btm.n114 VSS 0.801269f
C5653 C8_P_btm.n115 VSS 1.55307f
C5654 C8_P_btm.n116 VSS 1.08519f
C5655 C8_P_btm.n117 VSS 1.08899f
C5656 C8_P_btm.n118 VSS 1.08519f
C5657 C8_P_btm.n119 VSS 1.08899f
C5658 C8_P_btm.n120 VSS 1.08899f
C5659 C8_P_btm.n121 VSS 1.08899f
C5660 C8_P_btm.n122 VSS 1.08519f
C5661 C8_P_btm.n123 VSS 1.08899f
C5662 C8_P_btm.n124 VSS 1.08899f
C5663 C8_P_btm.n125 VSS 1.08519f
C5664 C8_P_btm.n126 VSS 1.08899f
C5665 C8_P_btm.n127 VSS 1.08899f
C5666 C8_P_btm.n128 VSS 1.08899f
C5667 C8_P_btm.n129 VSS 1.08899f
C5668 C8_P_btm.n130 VSS 3.37122f
C5669 C8_P_btm.n131 VSS 1.08899f
C5670 C8_P_btm.n132 VSS 1.08899f
C5671 C8_P_btm.n133 VSS 1.08899f
C5672 C8_P_btm.n134 VSS 1.08519f
C5673 C8_P_btm.n135 VSS 1.08899f
C5674 C8_P_btm.n136 VSS 1.08899f
C5675 C8_P_btm.n137 VSS 1.08519f
C5676 C8_P_btm.n138 VSS 1.08899f
C5677 C8_P_btm.n139 VSS 1.08899f
C5678 C8_P_btm.n140 VSS 1.08899f
C5679 C8_P_btm.n141 VSS 1.08899f
C5680 C8_P_btm.n142 VSS 1.08899f
C5681 C8_P_btm.n143 VSS 1.08899f
C5682 C8_P_btm.n144 VSS 1.08519f
C5683 C8_P_btm.n145 VSS 1.08519f
C5684 C8_P_btm.n146 VSS 1.08519f
C5685 C8_P_btm.n147 VSS 1.08519f
C5686 C8_P_btm.n148 VSS 1.08519f
C5687 C8_P_btm.n149 VSS 1.08899f
C5688 C8_P_btm.n150 VSS 1.08899f
C5689 C8_P_btm.n151 VSS 1.08899f
C5690 C8_P_btm.n152 VSS 1.08899f
C5691 C8_P_btm.n153 VSS 1.08519f
C5692 C8_P_btm.n154 VSS 1.39409f
C5693 C8_P_btm.n155 VSS 3.37111f
C5694 C8_P_btm.n156 VSS 7.05489f
C5695 C8_P_btm.n157 VSS 1.08899f
C5696 C8_P_btm.n158 VSS 1.08899f
C5697 C8_P_btm.n159 VSS 1.08899f
C5698 C8_P_btm.n160 VSS 1.3941f
C5699 C8_P_btm.n161 VSS 1.08519f
C5700 C8_P_btm.n162 VSS 1.08519f
C5701 C8_P_btm.n163 VSS 1.08519f
C5702 C8_P_btm.n164 VSS 1.08899f
C5703 C8_P_btm.n165 VSS 1.08899f
C5704 C8_P_btm.n166 VSS 1.08899f
C5705 C8_P_btm.n167 VSS 1.08899f
C5706 C8_P_btm.n168 VSS 1.08519f
C5707 C8_P_btm.n169 VSS 1.08519f
C5708 C8_P_btm.n170 VSS 1.08519f
C5709 C8_P_btm.n171 VSS 1.08899f
C5710 C8_P_btm.n172 VSS 1.08899f
C5711 C8_P_btm.n173 VSS 1.08899f
C5712 C8_P_btm.n174 VSS 1.08899f
C5713 C8_P_btm.n175 VSS 1.08519f
C5714 C8_P_btm.n176 VSS 1.31159f
C5715 C8_P_btm.n177 VSS 1.70573f
C5716 C8_P_btm.n178 VSS 1.08899f
C5717 C8_P_btm.n179 VSS 1.08899f
C5718 C8_P_btm.n180 VSS 1.08899f
C5719 C8_P_btm.n181 VSS 1.08899f
C5720 C8_P_btm.n182 VSS 1.08899f
C5721 C8_P_btm.n183 VSS 1.08899f
C5722 C8_P_btm.n184 VSS 2.37473f
C5723 C8_P_btm.n185 VSS 1.05126f
C5724 C8_P_btm.n186 VSS 1.48659f
C5725 C8_P_btm.n187 VSS 1.08899f
C5726 C8_P_btm.n188 VSS 1.3691f
C5727 C8_P_btm.n189 VSS 1.3691f
C5728 C8_P_btm.n190 VSS 1.3691f
C5729 C8_P_btm.n191 VSS 1.08899f
C5730 C8_P_btm.n192 VSS 1.08899f
C5731 C8_P_btm.n193 VSS 1.08899f
C5732 C8_P_btm.n194 VSS 0.801269f
C5733 C8_P_btm.n195 VSS 0.801269f
C5734 C8_P_btm.n196 VSS 0.801269f
C5735 C8_P_btm.n197 VSS 0.801269f
C5736 C8_P_btm.n198 VSS 1.08899f
C5737 C8_P_btm.n199 VSS 1.08899f
C5738 C8_P_btm.n200 VSS 1.3691f
C5739 C8_P_btm.n201 VSS 1.3691f
C5740 C8_P_btm.n202 VSS 1.08899f
C5741 C8_P_btm.n203 VSS 1.3691f
C5742 C8_P_btm.n204 VSS 1.3691f
C5743 C8_P_btm.n205 VSS 1.3691f
C5744 C8_P_btm.n206 VSS 1.08899f
C5745 C8_P_btm.n207 VSS 1.08899f
C5746 C8_P_btm.n208 VSS 1.08899f
C5747 C8_P_btm.n209 VSS 1.87981f
C5748 C8_P_btm.n210 VSS 1.8931f
C5749 C8_P_btm.n211 VSS 0.801269f
C5750 C8_P_btm.n212 VSS 0.801269f
C5751 C8_P_btm.n213 VSS 1.08899f
C5752 C8_P_btm.n214 VSS 1.08899f
C5753 C8_P_btm.n215 VSS 1.3691f
C5754 C8_P_btm.n216 VSS 1.3691f
C5755 C8_P_btm.n217 VSS 1.08899f
C5756 C8_P_btm.n218 VSS 1.3691f
C5757 C8_P_btm.n219 VSS 1.3691f
C5758 C8_P_btm.n220 VSS 1.3691f
C5759 C8_P_btm.n221 VSS 1.3691f
C5760 C8_P_btm.n222 VSS 1.08899f
C5761 C8_P_btm.n223 VSS 1.08899f
C5762 C8_P_btm.n224 VSS 1.08899f
C5763 C8_P_btm.n225 VSS 0.801269f
C5764 C8_P_btm.n226 VSS 0.801269f
C5765 C8_P_btm.n227 VSS 0.801269f
C5766 C8_P_btm.n228 VSS 0.801269f
C5767 C8_P_btm.n229 VSS 1.08899f
C5768 C8_P_btm.n230 VSS 1.08899f
C5769 C8_P_btm.n231 VSS 1.08899f
C5770 C8_P_btm.n232 VSS 1.08899f
C5771 C8_P_btm.n233 VSS 1.08899f
C5772 C8_P_btm.n234 VSS 2.37461f
C5773 C8_P_btm.n235 VSS 1.08519f
C5774 C8_P_btm.n236 VSS 1.08519f
C5775 C8_P_btm.n237 VSS 1.08899f
C5776 C8_P_btm.n238 VSS 1.08899f
C5777 C8_P_btm.n239 VSS 1.08899f
C5778 C8_P_btm.n240 VSS 1.08899f
C5779 C8_P_btm.n241 VSS 1.08519f
C5780 C8_P_btm.n242 VSS 1.08519f
C5781 C8_P_btm.n243 VSS 1.08519f
C5782 C8_P_btm.n244 VSS 1.08519f
C5783 C8_P_btm.n245 VSS 1.08899f
C5784 C8_P_btm.n246 VSS 1.08899f
C5785 C8_P_btm.n247 VSS 1.08899f
C5786 C8_P_btm.n248 VSS 1.08899f
C5787 C8_P_btm.n249 VSS 1.08519f
C5788 C8_P_btm.n250 VSS 2.45777f
C5789 C0_dummy_P_btm.t1 VSS 0.580759f
C5790 C0_dummy_P_btm.t0 VSS 0.30854f
C5791 C0_dummy_P_btm.n0 VSS 5.98126f
C5792 a_n2661_42282.t1 VSS 0.091035f
C5793 a_n2661_42282.t3 VSS 0.044507f
C5794 a_n2661_42282.t2 VSS 0.028401f
C5795 a_n2661_42282.n0 VSS 0.867409f
C5796 a_n2661_42282.n1 VSS 3.66259f
C5797 a_n2661_42282.t0 VSS 0.106053f
C5798 a_n4318_38680.t0 VSS 0.040452f
C5799 a_n4318_38680.t4 VSS 0.067578f
C5800 a_n4318_38680.t5 VSS 0.042323f
C5801 a_n4318_38680.n0 VSS 0.901461f
C5802 a_n4318_38680.t2 VSS 0.026294f
C5803 a_n4318_38680.t3 VSS 0.026294f
C5804 a_n4318_38680.n1 VSS 0.052587f
C5805 a_n4318_38680.n2 VSS 4.58118f
C5806 a_n4318_38680.n3 VSS 0.121382f
C5807 a_n4318_38680.t1 VSS 0.040452f
C5808 C2_P_btm.t3 VSS 1.57745f
C5809 C2_P_btm.t2 VSS 0.479134f
C5810 C2_P_btm.t0 VSS 0.321405f
C5811 C2_P_btm.n0 VSS 2.53294f
C5812 C2_P_btm.n1 VSS 3.886f
C5813 C2_P_btm.t1 VSS 0.219545f
C5814 C2_P_btm.n2 VSS 4.60349f
C5815 a_n2109_47186.t1 VSS 0.047239f
C5816 a_n2109_47186.t2 VSS 0.018723f
C5817 a_n2109_47186.t3 VSS 0.02934f
C5818 a_n2109_47186.n0 VSS 0.473524f
C5819 a_n2109_47186.n1 VSS 2.02574f
C5820 a_n2109_47186.t0 VSS 0.105439f
C5821 a_n2312_38680.t0 VSS 0.056936f
C5822 a_n2312_38680.t5 VSS 0.094012f
C5823 a_n2312_38680.t4 VSS 0.058647f
C5824 a_n2312_38680.n0 VSS 2.32091f
C5825 a_n2312_38680.t2 VSS 0.037008f
C5826 a_n2312_38680.t3 VSS 0.037008f
C5827 a_n2312_38680.n1 VSS 0.074016f
C5828 a_n2312_38680.n2 VSS 9.39369f
C5829 a_n2312_38680.n3 VSS 0.170845f
C5830 a_n2312_38680.t1 VSS 0.056936f
C5831 a_n356_44636.t2 VSS 0.031631f
C5832 a_n356_44636.t4 VSS 0.025547f
C5833 a_n356_44636.n0 VSS 0.180344f
C5834 a_n356_44636.t3 VSS 0.020365f
C5835 a_n356_44636.t5 VSS 0.037044f
C5836 a_n356_44636.n1 VSS 0.069187f
C5837 a_n356_44636.n2 VSS 3.30191f
C5838 a_n356_44636.t1 VSS 0.070506f
C5839 a_n356_44636.n3 VSS 3.51112f
C5840 a_n356_44636.t0 VSS 0.152343f
C5841 a_8685_43396.t3 VSS 0.03388f
C5842 a_8685_43396.t2 VSS 0.023031f
C5843 a_8685_43396.n0 VSS 0.512976f
C5844 a_8685_43396.t1 VSS 0.049789f
C5845 a_8685_43396.n1 VSS 3.76267f
C5846 a_8685_43396.t0 VSS 0.117656f
C5847 C0_dummy_N_btm.t1 VSS 0.580759f
C5848 C0_dummy_N_btm.t0 VSS 0.30854f
C5849 C0_dummy_N_btm.n0 VSS 5.98126f
C5850 a_13678_32519.t4 VSS 2.33335f
C5851 a_13678_32519.t3 VSS 0.038955f
C5852 a_13678_32519.t2 VSS 0.038955f
C5853 a_13678_32519.n0 VSS 0.07791f
C5854 a_13678_32519.n1 VSS 19.011099f
C5855 a_13678_32519.t0 VSS 0.059931f
C5856 a_13678_32519.n2 VSS 0.179832f
C5857 a_13678_32519.t1 VSS 0.059931f
C5858 a_11341_43940.t2 VSS 0.09126f
C5859 a_11341_43940.t1 VSS 0.106349f
C5860 a_11341_43940.t3 VSS 0.01717f
C5861 a_11341_43940.t4 VSS 0.026906f
C5862 a_11341_43940.n0 VSS 0.928043f
C5863 a_11341_43940.n1 VSS 4.09928f
C5864 a_11341_43940.n2 VSS 0.111184f
C5865 a_11341_43940.t0 VSS 0.019808f
C5866 a_n2293_46098.t1 VSS 0.041602f
C5867 a_n2293_46098.t2 VSS 0.011145f
C5868 a_n2293_46098.t3 VSS 0.017465f
C5869 a_n2293_46098.n0 VSS 0.566037f
C5870 a_n2293_46098.n1 VSS 2.3181f
C5871 a_n2293_46098.t0 VSS 0.045647f
C5872 a_n2293_46634.t2 VSS 0.014897f
C5873 a_n2293_46634.t1 VSS 0.07098f
C5874 a_n2293_46634.t3 VSS 0.020984f
C5875 a_n2293_46634.t4 VSS 0.01339f
C5876 a_n2293_46634.n0 VSS 1.16322f
C5877 a_n2293_46634.n1 VSS 5.37172f
C5878 a_n2293_46634.n2 VSS 0.029911f
C5879 a_n2293_46634.t0 VSS 0.014897f
C5880 a_19963_31679.t3 VSS 0.038709f
C5881 a_19963_31679.t2 VSS 0.038709f
C5882 a_19963_31679.n0 VSS 0.134606f
C5883 a_19963_31679.t4 VSS 2.72762f
C5884 a_19963_31679.n1 VSS 14.819401f
C5885 a_19963_31679.t0 VSS 0.059552f
C5886 a_19963_31679.n2 VSS 0.12186f
C5887 a_19963_31679.t1 VSS 0.059552f
C5888 C5_N_btm.t2 VSS 1.10875f
C5889 C5_N_btm.t3 VSS 0.344593f
C5890 C5_N_btm.t1 VSS 0.231154f
C5891 C5_N_btm.n0 VSS 1.75362f
C5892 C5_N_btm.n1 VSS 2.74079f
C5893 C5_N_btm.t0 VSS 0.148423f
C5894 C5_N_btm.n2 VSS 3.53899f
C5895 CAL_P.n0 VSS 1.89859f
C5896 CAL_P.t4 VSS 5.35363f
C5897 CAL_P.n1 VSS 3.77122f
C5898 CAL_P.t3 VSS 4.80383f
C5899 CAL_P.n2 VSS 3.86937f
C5900 CAL_P.t6 VSS 5.34448f
C5901 CAL_P.n3 VSS 2.01614f
C5902 CAL_P.t1 VSS 0.011104f
C5903 CAL_P.n5 VSS 0.341163f
C5904 CAL_P.n6 VSS 0.520365f
C5905 CAL_P.t5 VSS 0.103479f
C5906 RST_Z.t5 VSS 0.088732f
C5907 RST_Z.t3 VSS 0.318957f
C5908 RST_Z.n0 VSS 2.83283f
C5909 RST_Z.t0 VSS 0.04971f
C5910 RST_Z.t4 VSS 0.031045f
C5911 RST_Z.n1 VSS 0.097381f
C5912 RST_Z.n2 VSS 6.84398f
C5913 RST_Z.t2 VSS 0.029113f
C5914 RST_Z.t1 VSS 0.04668f
C5915 RST_Z.n3 VSS 0.110098f
C5916 a_4338_37500.t5 VSS 0.099543f
C5917 a_4338_37500.t3 VSS 0.025975f
C5918 a_4338_37500.t4 VSS 0.025975f
C5919 a_4338_37500.n0 VSS 0.071898f
C5920 a_4338_37500.n1 VSS 0.347491f
C5921 a_4338_37500.t2 VSS 0.098471f
C5922 a_4338_37500.n2 VSS 0.476562f
C5923 a_4338_37500.t6 VSS 0.024676f
C5924 a_4338_37500.t1 VSS 0.024676f
C5925 a_4338_37500.n3 VSS 0.110266f
C5926 a_4338_37500.n4 VSS 1.30834f
C5927 a_4338_37500.t0 VSS 0.086124f
C5928 a_n2661_43922.t2 VSS 0.017685f
C5929 a_n2661_43922.t4 VSS 0.015897f
C5930 a_n2661_43922.t3 VSS 0.024912f
C5931 a_n2661_43922.n0 VSS 0.832411f
C5932 a_n2661_43922.t1 VSS 0.034907f
C5933 a_n2661_43922.n1 VSS 5.59707f
C5934 a_n2661_43922.n2 VSS 0.059431f
C5935 a_n2661_43922.t0 VSS 0.017685f
C5936 a_n2810_45572.t3 VSS 0.038905f
C5937 a_n2810_45572.t2 VSS 0.038905f
C5938 a_n2810_45572.n0 VSS 0.135289f
C5939 a_n2810_45572.t4 VSS 0.061654f
C5940 a_n2810_45572.t5 VSS 0.098832f
C5941 a_n2810_45572.n1 VSS 2.1946f
C5942 a_n2810_45572.n2 VSS 9.08962f
C5943 a_n2810_45572.t0 VSS 0.059855f
C5944 a_n2810_45572.n3 VSS 0.122478f
C5945 a_n2810_45572.t1 VSS 0.059855f
C5946 a_n3420_37440.t0 VSS 0.038822f
C5947 a_n3420_37440.t6 VSS 0.025234f
C5948 a_n3420_37440.t5 VSS 0.025234f
C5949 a_n3420_37440.n0 VSS 0.052302f
C5950 a_n3420_37440.t7 VSS 0.025234f
C5951 a_n3420_37440.t4 VSS 0.025234f
C5952 a_n3420_37440.n1 VSS 0.062067f
C5953 a_n3420_37440.n2 VSS 0.231597f
C5954 a_n3420_37440.t8 VSS 0.063087f
C5955 a_n3420_37440.t10 VSS 0.039615f
C5956 a_n3420_37440.n3 VSS 0.091296f
C5957 a_n3420_37440.t9 VSS 0.826046f
C5958 a_n3420_37440.n4 VSS 8.277861f
C5959 a_n3420_37440.n5 VSS 0.149475f
C5960 a_n3420_37440.t1 VSS 0.038822f
C5961 a_n3420_37440.t2 VSS 0.038822f
C5962 a_n3420_37440.n6 VSS 0.100045f
C5963 a_n3420_37440.n7 VSS 0.268793f
C5964 a_n3420_37440.n8 VSS 0.081597f
C5965 a_n3420_37440.t3 VSS 0.038822f
C5966 C4_P_btm.t0 VSS 1.26438f
C5967 C4_P_btm.t3 VSS 0.389904f
C5968 C4_P_btm.t1 VSS 0.261549f
C5969 C4_P_btm.n0 VSS 2.01038f
C5970 C4_P_btm.n1 VSS 3.13259f
C5971 C4_P_btm.t2 VSS 0.171423f
C5972 C4_P_btm.n2 VSS 3.85704f
C5973 a_9145_43396.t1 VSS 0.161715f
C5974 a_9145_43396.t2 VSS 0.066775f
C5975 a_9145_43396.t3 VSS 0.045494f
C5976 a_9145_43396.n0 VSS 0.652408f
C5977 a_9145_43396.n1 VSS 3.59257f
C5978 a_9145_43396.t0 VSS 0.181042f
C5979 a_9313_44734.t4 VSS 0.01997f
C5980 a_9313_44734.t3 VSS 0.031295f
C5981 a_9313_44734.n0 VSS 1.20515f
C5982 a_9313_44734.t1 VSS 0.050734f
C5983 a_9313_44734.n1 VSS 5.94398f
C5984 a_9313_44734.t2 VSS 0.035269f
C5985 a_9313_44734.n2 VSS 0.094597f
C5986 a_9313_44734.t0 VSS 0.019007f
C5987 CLK.t0 VSS 0.014189f
C5988 CLK.t1 VSS 0.030339f
C5989 CLK.t6 VSS 0.014189f
C5990 CLK.t7 VSS 0.030339f
C5991 CLK.t3 VSS 0.014189f
C5992 CLK.t5 VSS 0.030339f
C5993 CLK.t4 VSS 0.014189f
C5994 CLK.t2 VSS 0.030339f
C5995 CLK.n0 VSS 0.069262f
C5996 CLK.n1 VSS 0.091226f
C5997 CLK.n2 VSS 0.091226f
C5998 CLK.n3 VSS 0.315718f
C5999 a_14209_32519.t4 VSS 2.20549f
C6000 a_14209_32519.t3 VSS 0.042182f
C6001 a_14209_32519.t2 VSS 0.042182f
C6002 a_14209_32519.n0 VSS 0.084365f
C6003 a_14209_32519.n1 VSS 18.9013f
C6004 a_14209_32519.t0 VSS 0.064896f
C6005 a_14209_32519.n2 VSS 0.194731f
C6006 a_14209_32519.t1 VSS 0.064896f
C6007 a_n2293_45546.t3 VSS 0.027578f
C6008 a_n2293_45546.t2 VSS 0.14257f
C6009 a_n2293_45546.t4 VSS 0.027602f
C6010 a_n2293_45546.t5 VSS 0.017614f
C6011 a_n2293_45546.n0 VSS 0.198188f
C6012 a_n2293_45546.n1 VSS 1.20435f
C6013 a_n2293_45546.t1 VSS 0.142802f
C6014 a_n2293_45546.n2 VSS 0.23154f
C6015 a_n2293_45546.n3 VSS 0.078731f
C6016 a_n2293_45546.t0 VSS 0.029029f
C6017 a_n2956_38216.t0 VSS 0.055071f
C6018 a_n2956_38216.t4 VSS 0.056727f
C6019 a_n2956_38216.t5 VSS 0.090934f
C6020 a_n2956_38216.n0 VSS 2.19941f
C6021 a_n2956_38216.t2 VSS 0.035796f
C6022 a_n2956_38216.t3 VSS 0.035796f
C6023 a_n2956_38216.n1 VSS 0.071593f
C6024 a_n2956_38216.n2 VSS 9.13435f
C6025 a_n2956_38216.n3 VSS 0.165251f
C6026 a_n2956_38216.t1 VSS 0.055071f
C6027 a_n3420_38528.t0 VSS 0.057935f
C6028 a_n3420_38528.t6 VSS 0.037658f
C6029 a_n3420_38528.t5 VSS 0.037658f
C6030 a_n3420_38528.n0 VSS 0.078052f
C6031 a_n3420_38528.t7 VSS 0.037658f
C6032 a_n3420_38528.t4 VSS 0.037658f
C6033 a_n3420_38528.n1 VSS 0.092624f
C6034 a_n3420_38528.n2 VSS 0.345621f
C6035 a_n3420_38528.t9 VSS 0.094147f
C6036 a_n3420_38528.t10 VSS 0.059119f
C6037 a_n3420_38528.n3 VSS 0.136244f
C6038 a_n3420_38528.t8 VSS 1.22451f
C6039 a_n3420_38528.n4 VSS 12.292f
C6040 a_n3420_38528.n5 VSS 0.223067f
C6041 a_n3420_38528.t1 VSS 0.057935f
C6042 a_n3420_38528.t2 VSS 0.057935f
C6043 a_n3420_38528.n6 VSS 0.1493f
C6044 a_n3420_38528.n7 VSS 0.40113f
C6045 a_n3420_38528.n8 VSS 0.12177f
C6046 a_n3420_38528.t3 VSS 0.057935f
C6047 a_14401_32519.t0 VSS 0.052319f
C6048 a_14401_32519.t2 VSS 0.034007f
C6049 a_14401_32519.t3 VSS 0.034007f
C6050 a_14401_32519.n0 VSS 0.125944f
C6051 a_14401_32519.t4 VSS 0.165676f
C6052 a_14401_32519.t5 VSS 0.190508f
C6053 a_14401_32519.n1 VSS 4.55239f
C6054 a_14401_32519.n2 VSS 12.9882f
C6055 a_14401_32519.n3 VSS 0.10468f
C6056 a_14401_32519.t1 VSS 0.052319f
C6057 a_n3674_38216.t0 VSS 0.036091f
C6058 a_n3674_38216.t5 VSS 0.03776f
C6059 a_n3674_38216.t4 VSS 0.060293f
C6060 a_n3674_38216.n0 VSS 0.943199f
C6061 a_n3674_38216.t2 VSS 0.023459f
C6062 a_n3674_38216.t3 VSS 0.023459f
C6063 a_n3674_38216.n1 VSS 0.046918f
C6064 a_n3674_38216.n2 VSS 4.284431f
C6065 a_n3674_38216.n3 VSS 0.108298f
C6066 a_n3674_38216.t1 VSS 0.036091f
C6067 a_n2661_45546.t2 VSS 0.013372f
C6068 a_n2661_45546.t3 VSS 0.018836f
C6069 a_n2661_45546.t4 VSS 0.01202f
C6070 a_n2661_45546.n0 VSS 0.45609f
C6071 a_n2661_45546.t1 VSS 0.026392f
C6072 a_n2661_45546.n1 VSS 2.41498f
C6073 a_n2661_45546.n2 VSS 0.044935f
C6074 a_n2661_45546.t0 VSS 0.013372f
C6075 C7_N_btm.t2 VSS 0.15694f
C6076 C7_N_btm.t3 VSS 0.15694f
C6077 C7_N_btm.n0 VSS 0.933237f
C6078 C7_N_btm.t4 VSS 1.12025f
C6079 C7_N_btm.n1 VSS 2.0822f
C6080 C7_N_btm.t1 VSS 1.12621f
C6081 C7_N_btm.n2 VSS 1.11461f
C6082 C7_N_btm.t0 VSS 0.21231f
C6083 C7_N_btm.n3 VSS 2.68842f
C6084 a_n2956_37592.t0 VSS 0.042448f
C6085 a_n2956_37592.t2 VSS 0.027591f
C6086 a_n2956_37592.t3 VSS 0.027591f
C6087 a_n2956_37592.n0 VSS 0.102183f
C6088 a_n2956_37592.t4 VSS 0.07009f
C6089 a_n2956_37592.t5 VSS 0.043724f
C6090 a_n2956_37592.n1 VSS 1.92651f
C6091 a_n2956_37592.n2 VSS 6.43248f
C6092 a_n2956_37592.n3 VSS 0.08493f
C6093 a_n2956_37592.t1 VSS 0.042448f
C6094 a_n4064_37440.t2 VSS 0.056069f
C6095 a_n4064_37440.t5 VSS 0.036445f
C6096 a_n4064_37440.t4 VSS 0.036445f
C6097 a_n4064_37440.n0 VSS 0.075538f
C6098 a_n4064_37440.t7 VSS 0.036445f
C6099 a_n4064_37440.t6 VSS 0.036445f
C6100 a_n4064_37440.n1 VSS 0.089641f
C6101 a_n4064_37440.n2 VSS 0.337923f
C6102 a_n4064_37440.t10 VSS 0.091114f
C6103 a_n4064_37440.t8 VSS 0.057215f
C6104 a_n4064_37440.n3 VSS 0.163695f
C6105 a_n4064_37440.t9 VSS 1.11699f
C6106 a_n4064_37440.n4 VSS 12.434799f
C6107 a_n4064_37440.n5 VSS 0.216361f
C6108 a_n4064_37440.t1 VSS 0.056069f
C6109 a_n4064_37440.t0 VSS 0.056069f
C6110 a_n4064_37440.n6 VSS 0.144491f
C6111 a_n4064_37440.n7 VSS 0.384297f
C6112 a_n4064_37440.n8 VSS 0.117848f
C6113 a_n4064_37440.t3 VSS 0.056069f
C6114 a_6945_45028.t2 VSS 0.025062f
C6115 a_6945_45028.t1 VSS 0.053493f
C6116 a_6945_45028.t3 VSS 0.022528f
C6117 a_6945_45028.t4 VSS 0.035304f
C6118 a_6945_45028.n0 VSS 1.45092f
C6119 a_6945_45028.n1 VSS 8.10634f
C6120 a_6945_45028.n2 VSS 0.081286f
C6121 a_6945_45028.t0 VSS 0.025062f
C6122 a_5649_42852.t1 VSS 0.112596f
C6123 a_5649_42852.t3 VSS 0.04889f
C6124 a_5649_42852.t2 VSS 0.031198f
C6125 a_5649_42852.n0 VSS 1.89654f
C6126 a_5649_42852.n1 VSS 5.7852f
C6127 a_5649_42852.t0 VSS 0.125581f
C6128 a_2982_43646.t0 VSS 0.014708f
C6129 a_2982_43646.n0 VSS 0.019387f
C6130 a_2982_43646.t7 VSS 0.019978f
C6131 a_2982_43646.t6 VSS 0.012748f
C6132 a_2982_43646.n1 VSS 0.980887f
C6133 a_2982_43646.n2 VSS 5.3119f
C6134 a_2982_43646.t5 VSS 0.014708f
C6135 a_2982_43646.t4 VSS 0.014708f
C6136 a_2982_43646.n3 VSS 0.03557f
C6137 a_2982_43646.n4 VSS 0.111694f
C6138 a_2982_43646.n5 VSS 0.029883f
C6139 a_2982_43646.t1 VSS 0.014708f
C6140 C3_P_btm.t0 VSS 1.36935f
C6141 C3_P_btm.t1 VSS 0.419015f
C6142 C3_P_btm.t3 VSS 0.281077f
C6143 C3_P_btm.n0 VSS 2.18805f
C6144 C3_P_btm.n1 VSS 3.46981f
C6145 C3_P_btm.t2 VSS 0.213431f
C6146 C3_P_btm.n2 VSS 4.00802f
C6147 a_1666_39587.t2 VSS 0.089771f
C6148 a_1666_39587.t1 VSS 0.077332f
C6149 a_1666_39587.t6 VSS 0.128406f
C6150 a_1666_39587.t5 VSS 0.06994f
C6151 a_1666_39587.n0 VSS 0.787042f
C6152 a_1666_39587.t4 VSS 0.03269f
C6153 a_1666_39587.t3 VSS 0.020416f
C6154 a_1666_39587.n1 VSS 0.076534f
C6155 a_1666_39587.n2 VSS 0.593943f
C6156 a_1666_39587.n3 VSS 0.314727f
C6157 a_1666_39587.n4 VSS 0.596985f
C6158 a_1666_39587.t0 VSS 0.312213f
C6159 a_3357_43084.t2 VSS 0.028174f
C6160 a_3357_43084.t3 VSS 0.039686f
C6161 a_3357_43084.t4 VSS 0.025325f
C6162 a_3357_43084.n0 VSS 1.58232f
C6163 a_3357_43084.t5 VSS 0.02912f
C6164 a_3357_43084.t6 VSS 0.046638f
C6165 a_3357_43084.n1 VSS 0.126276f
C6166 a_3357_43084.n2 VSS 7.36849f
C6167 a_3357_43084.t1 VSS 0.055608f
C6168 a_3357_43084.n3 VSS 0.37551f
C6169 a_3357_43084.n4 VSS 0.094676f
C6170 a_3357_43084.t0 VSS 0.028174f
C6171 C5_P_btm.t2 VSS 1.10875f
C6172 C5_P_btm.t3 VSS 0.344593f
C6173 C5_P_btm.t1 VSS 0.231154f
C6174 C5_P_btm.n0 VSS 1.75362f
C6175 C5_P_btm.n1 VSS 2.74079f
C6176 C5_P_btm.t0 VSS 0.148423f
C6177 C5_P_btm.n2 VSS 3.53531f
C6178 a_n4064_38528.t0 VSS 0.056191f
C6179 a_n4064_38528.t6 VSS 0.036524f
C6180 a_n4064_38528.t7 VSS 0.036524f
C6181 a_n4064_38528.n0 VSS 0.075703f
C6182 a_n4064_38528.t4 VSS 0.036524f
C6183 a_n4064_38528.t5 VSS 0.036524f
C6184 a_n4064_38528.n1 VSS 0.089836f
C6185 a_n4064_38528.n2 VSS 0.338658f
C6186 a_n4064_38528.t10 VSS 0.091313f
C6187 a_n4064_38528.t9 VSS 0.057339f
C6188 a_n4064_38528.n3 VSS 0.164051f
C6189 a_n4064_38528.t8 VSS 1.07833f
C6190 a_n4064_38528.n4 VSS 12.569f
C6191 a_n4064_38528.n5 VSS 0.216831f
C6192 a_n4064_38528.t1 VSS 0.056191f
C6193 a_n4064_38528.t2 VSS 0.056191f
C6194 a_n4064_38528.n6 VSS 0.144806f
C6195 a_n4064_38528.n7 VSS 0.385132f
C6196 a_n4064_38528.n8 VSS 0.118104f
C6197 a_n4064_38528.t3 VSS 0.056191f
C6198 C2_N_btm.t3 VSS 1.57745f
C6199 C2_N_btm.t2 VSS 0.479134f
C6200 C2_N_btm.t0 VSS 0.321405f
C6201 C2_N_btm.n0 VSS 2.53294f
C6202 C2_N_btm.n1 VSS 3.886f
C6203 C2_N_btm.t1 VSS 0.219545f
C6204 C2_N_btm.n2 VSS 4.6214f
C6205 a_19721_31679.t4 VSS 2.76161f
C6206 a_19721_31679.t2 VSS 0.039317f
C6207 a_19721_31679.t3 VSS 0.039317f
C6208 a_19721_31679.n0 VSS 0.078634f
C6209 a_19721_31679.n1 VSS 14.778599f
C6210 a_19721_31679.t0 VSS 0.060487f
C6211 a_19721_31679.n2 VSS 0.181503f
C6212 a_19721_31679.t1 VSS 0.060487f
C6213 a_n4318_37592.t3 VSS 0.023524f
C6214 a_n4318_37592.t2 VSS 0.023524f
C6215 a_n4318_37592.n0 VSS 0.081801f
C6216 a_n4318_37592.t4 VSS 0.060459f
C6217 a_n4318_37592.t5 VSS 0.037864f
C6218 a_n4318_37592.n1 VSS 0.93849f
C6219 a_n4318_37592.n2 VSS 4.4879f
C6220 a_n4318_37592.t0 VSS 0.03619f
C6221 a_n4318_37592.n3 VSS 0.074055f
C6222 a_n4318_37592.t1 VSS 0.03619f
C6223 a_n357_42282.t0 VSS 0.024977f
C6224 a_n357_42282.t8 VSS 0.035183f
C6225 a_n357_42282.t7 VSS 0.022451f
C6226 a_n357_42282.n0 VSS 0.089445f
C6227 a_n357_42282.t9 VSS 0.042092f
C6228 a_n357_42282.t4 VSS 0.026431f
C6229 a_n357_42282.n1 VSS 0.195409f
C6230 a_n357_42282.t10 VSS 0.026458f
C6231 a_n357_42282.t14 VSS 0.052239f
C6232 a_n357_42282.n2 VSS 0.056361f
C6233 a_n357_42282.n3 VSS 1.91332f
C6234 a_n357_42282.t17 VSS 0.052239f
C6235 a_n357_42282.t16 VSS 0.026458f
C6236 a_n357_42282.n4 VSS 0.081682f
C6237 a_n357_42282.n5 VSS 2.40747f
C6238 a_n357_42282.t5 VSS 0.026458f
C6239 a_n357_42282.t13 VSS 0.052239f
C6240 a_n357_42282.n6 VSS 0.057633f
C6241 a_n357_42282.n7 VSS 2.09016f
C6242 a_n357_42282.t12 VSS 0.026458f
C6243 a_n357_42282.t11 VSS 0.052239f
C6244 a_n357_42282.n8 VSS 0.057633f
C6245 a_n357_42282.n9 VSS 3.21356f
C6246 a_n357_42282.t6 VSS 0.026458f
C6247 a_n357_42282.t15 VSS 0.052239f
C6248 a_n357_42282.n10 VSS 0.057633f
C6249 a_n357_42282.n11 VSS 4.42489f
C6250 a_n357_42282.n12 VSS 0.926356f
C6251 a_n357_42282.t3 VSS 0.016235f
C6252 a_n357_42282.t2 VSS 0.016235f
C6253 a_n357_42282.n13 VSS 0.03247f
C6254 a_n357_42282.n14 VSS 0.218959f
C6255 a_n357_42282.n15 VSS 0.074947f
C6256 a_n357_42282.t1 VSS 0.024977f
C6257 a_20447_31679.t0 VSS 0.060321f
C6258 a_20447_31679.t3 VSS 0.039209f
C6259 a_20447_31679.t2 VSS 0.039209f
C6260 a_20447_31679.n0 VSS 0.145208f
C6261 a_20447_31679.t4 VSS 2.97925f
C6262 a_20447_31679.n1 VSS 14.5558f
C6263 a_20447_31679.n2 VSS 0.120691f
C6264 a_20447_31679.t1 VSS 0.060321f
C6265 a_7174_31319.t0 VSS 0.062239f
C6266 a_7174_31319.t4 VSS 0.360616f
C6267 a_7174_31319.t5 VSS 0.342606f
C6268 a_7174_31319.n0 VSS 22.9714f
C6269 a_7174_31319.t3 VSS 0.040455f
C6270 a_7174_31319.t2 VSS 0.040455f
C6271 a_7174_31319.n1 VSS 0.08091f
C6272 a_7174_31319.n2 VSS 13.1523f
C6273 a_7174_31319.n3 VSS 0.186758f
C6274 a_7174_31319.t1 VSS 0.062239f
C6275 VDAC_Pi.t3 VSS 0.042772f
C6276 VDAC_Pi.t0 VSS 0.042772f
C6277 VDAC_Pi.n0 VSS 0.095084f
C6278 VDAC_Pi.t2 VSS 0.042772f
C6279 VDAC_Pi.t1 VSS 0.042772f
C6280 VDAC_Pi.n1 VSS 0.09446f
C6281 VDAC_Pi.n2 VSS 0.665943f
C6282 VDAC_Pi.t8 VSS 0.180328f
C6283 VDAC_Pi.t10 VSS 0.150409f
C6284 VDAC_Pi.n3 VSS 2.14996f
C6285 VDAC_Pi.n4 VSS 0.329095f
C6286 VDAC_Pi.t4 VSS 0.042772f
C6287 VDAC_Pi.t5 VSS 0.042772f
C6288 VDAC_Pi.n5 VSS 0.109636f
C6289 VDAC_Pi.n6 VSS 0.242751f
C6290 VDAC_Pi.t6 VSS 0.042772f
C6291 VDAC_Pi.t7 VSS 0.042772f
C6292 VDAC_Pi.n7 VSS 0.109636f
C6293 VDAC_Pi.n8 VSS 0.442463f
C6294 VDAC_Pi.t9 VSS 0.046473f
C6295 a_413_45260.t3 VSS 0.041164f
C6296 a_413_45260.t4 VSS 0.026268f
C6297 a_413_45260.n0 VSS 1.88871f
C6298 a_413_45260.t5 VSS 0.030204f
C6299 a_413_45260.t2 VSS 0.048374f
C6300 a_413_45260.n1 VSS 0.154616f
C6301 a_413_45260.n2 VSS 8.684461f
C6302 a_413_45260.t1 VSS 0.057637f
C6303 a_413_45260.n3 VSS 0.504089f
C6304 a_413_45260.t0 VSS 0.164481f
C6305 a_n2661_46634.t2 VSS 0.018393f
C6306 a_n2661_46634.t3 VSS 0.025909f
C6307 a_n2661_46634.t4 VSS 0.016533f
C6308 a_n2661_46634.n0 VSS 1.16528f
C6309 a_n2661_46634.t1 VSS 0.082955f
C6310 a_n2661_46634.n1 VSS 5.63437f
C6311 a_n2661_46634.n2 VSS 0.03816f
C6312 a_n2661_46634.t0 VSS 0.018393f
C6313 a_n4318_40392.t2 VSS 0.028084f
C6314 a_n4318_40392.t3 VSS 0.028084f
C6315 a_n4318_40392.n0 VSS 0.09766f
C6316 a_n4318_40392.t5 VSS 0.045205f
C6317 a_n4318_40392.t4 VSS 0.07218f
C6318 a_n4318_40392.n1 VSS 0.822403f
C6319 a_n4318_40392.n2 VSS 4.13156f
C6320 a_n4318_40392.t0 VSS 0.043207f
C6321 a_n4318_40392.n3 VSS 0.088412f
C6322 a_n4318_40392.t1 VSS 0.043207f
C6323 a_4361_42308.t1 VSS 0.068622f
C6324 a_4361_42308.t3 VSS 0.042621f
C6325 a_4361_42308.t2 VSS 0.027198f
C6326 a_4361_42308.n0 VSS 1.58022f
C6327 a_4361_42308.n1 VSS 11.0282f
C6328 a_4361_42308.t0 VSS 0.153167f
C6329 a_11453_44696.t1 VSS 0.075872f
C6330 a_11453_44696.n0 VSS 0.122039f
C6331 a_11453_44696.t3 VSS 0.021486f
C6332 a_11453_44696.t4 VSS 0.033671f
C6333 a_11453_44696.n1 VSS 0.282188f
C6334 a_11453_44696.t5 VSS 0.027854f
C6335 a_11453_44696.t2 VSS 0.03218f
C6336 a_11453_44696.n2 VSS 0.219214f
C6337 a_11453_44696.n3 VSS 5.53396f
C6338 a_11453_44696.n4 VSS 0.067948f
C6339 a_11453_44696.t0 VSS 0.083591f
C6340 C3_N_btm.t2 VSS 1.36935f
C6341 C3_N_btm.t1 VSS 0.419015f
C6342 C3_N_btm.t3 VSS 0.281077f
C6343 C3_N_btm.n0 VSS 2.18805f
C6344 C3_N_btm.n1 VSS 3.46981f
C6345 C3_N_btm.t0 VSS 0.213431f
C6346 C3_N_btm.n2 VSS 4.00579f
C6347 a_5932_42308.t5 VSS 0.081492f
C6348 a_5932_42308.t7 VSS 0.050824f
C6349 a_5932_42308.n0 VSS 0.224341f
C6350 a_5932_42308.t4 VSS 0.360472f
C6351 a_5932_42308.t6 VSS 0.346979f
C6352 a_5932_42308.n1 VSS 15.369901f
C6353 a_5932_42308.n2 VSS 9.56684f
C6354 a_5932_42308.t3 VSS 0.034052f
C6355 a_5932_42308.t2 VSS 0.034052f
C6356 a_5932_42308.n3 VSS 0.068103f
C6357 a_5932_42308.n4 VSS 0.600938f
C6358 a_5932_42308.t0 VSS 0.052387f
C6359 a_5932_42308.n5 VSS 0.157196f
C6360 a_5932_42308.t1 VSS 0.052387f
C6361 C1_P_btm.t2 VSS 1.54443f
C6362 C1_P_btm.t3 VSS 0.46356f
C6363 C1_P_btm.t1 VSS 0.312474f
C6364 C1_P_btm.n0 VSS 2.48776f
C6365 C1_P_btm.n1 VSS 3.86765f
C6366 C1_P_btm.t0 VSS 0.279285f
C6367 C1_P_btm.n2 VSS 4.72888f
C6368 a_n1435_47204.t2 VSS 0.011955f
C6369 a_n1435_47204.t3 VSS 0.019038f
C6370 a_n1435_47204.n0 VSS 0.39724f
C6371 a_n1435_47204.t1 VSS 0.020213f
C6372 a_n1435_47204.n1 VSS 1.71165f
C6373 a_n1435_47204.t0 VSS 0.039902f
C6374 a_n4318_38216.t0 VSS 0.037409f
C6375 a_n4318_38216.t2 VSS 0.024316f
C6376 a_n4318_38216.t3 VSS 0.024316f
C6377 a_n4318_38216.n0 VSS 0.090053f
C6378 a_n4318_38216.t5 VSS 0.03914f
C6379 a_n4318_38216.t4 VSS 0.062495f
C6380 a_n4318_38216.n1 VSS 1.01125f
C6381 a_n4318_38216.n2 VSS 4.29876f
C6382 a_n4318_38216.n3 VSS 0.074849f
C6383 a_n4318_38216.t1 VSS 0.037409f
C6384 C1_N_btm.t2 VSS 1.54443f
C6385 C1_N_btm.t1 VSS 0.46356f
C6386 C1_N_btm.t3 VSS 0.312474f
C6387 C1_N_btm.n0 VSS 2.48776f
C6388 C1_N_btm.n1 VSS 3.86765f
C6389 C1_N_btm.t0 VSS 0.279285f
C6390 C1_N_btm.n2 VSS 4.72639f
C6391 a_5700_37509.t2 VSS 0.087988f
C6392 a_5700_37509.t9 VSS 0.231968f
C6393 a_5700_37509.t12 VSS 0.231968f
C6394 a_5700_37509.n0 VSS 0.462462f
C6395 a_5700_37509.t6 VSS 0.231968f
C6396 a_5700_37509.t13 VSS 0.231968f
C6397 a_5700_37509.n1 VSS 0.462027f
C6398 a_5700_37509.n2 VSS 0.180212f
C6399 a_5700_37509.t7 VSS 0.231968f
C6400 a_5700_37509.t14 VSS 0.231968f
C6401 a_5700_37509.n3 VSS 0.462027f
C6402 a_5700_37509.n4 VSS 0.127652f
C6403 a_5700_37509.t18 VSS 0.231968f
C6404 a_5700_37509.t10 VSS 0.231968f
C6405 a_5700_37509.n5 VSS 0.462027f
C6406 a_5700_37509.n6 VSS 0.692908f
C6407 a_5700_37509.t5 VSS 0.231968f
C6408 a_5700_37509.t19 VSS 0.231968f
C6409 a_5700_37509.n7 VSS 0.561806f
C6410 a_5700_37509.t8 VSS 0.231968f
C6411 a_5700_37509.t4 VSS 0.231968f
C6412 a_5700_37509.n8 VSS 0.556177f
C6413 a_5700_37509.n9 VSS 1.57381f
C6414 a_5700_37509.t16 VSS 0.231968f
C6415 a_5700_37509.t17 VSS 0.231968f
C6416 a_5700_37509.n10 VSS 0.556177f
C6417 a_5700_37509.n11 VSS 0.827046f
C6418 a_5700_37509.t15 VSS 0.231968f
C6419 a_5700_37509.t11 VSS 0.231968f
C6420 a_5700_37509.n12 VSS 0.556177f
C6421 a_5700_37509.n13 VSS 1.34054f
C6422 a_5700_37509.n14 VSS 3.49156f
C6423 a_5700_37509.t3 VSS 0.319458f
C6424 a_5700_37509.n15 VSS 1.6989f
C6425 a_5700_37509.t1 VSS 0.321046f
C6426 a_5700_37509.n16 VSS 1.25965f
C6427 a_5700_37509.n17 VSS 0.200876f
C6428 a_5700_37509.t0 VSS 0.087988f
C6429 VDAC_N.t20 VSS 0.506181f
C6430 VDAC_N.t16 VSS 0.505972f
C6431 VDAC_N.n0 VSS 0.565755f
C6432 VDAC_N.t12 VSS 0.505972f
C6433 VDAC_N.n1 VSS 0.296463f
C6434 VDAC_N.t15 VSS 0.505972f
C6435 VDAC_N.n2 VSS 0.396124f
C6436 VDAC_N.t9 VSS 0.506181f
C6437 VDAC_N.t14 VSS 0.505972f
C6438 VDAC_N.n3 VSS 0.565755f
C6439 VDAC_N.t18 VSS 0.505972f
C6440 VDAC_N.n4 VSS 0.296463f
C6441 VDAC_N.t8 VSS 0.505972f
C6442 VDAC_N.n5 VSS 0.589481f
C6443 VDAC_N.t10 VSS 0.505972f
C6444 VDAC_N.n6 VSS 0.588782f
C6445 VDAC_N.t11 VSS 0.505972f
C6446 VDAC_N.n7 VSS 0.296463f
C6447 VDAC_N.t13 VSS 0.505972f
C6448 VDAC_N.n8 VSS 0.296463f
C6449 VDAC_N.t19 VSS 0.505972f
C6450 VDAC_N.n9 VSS 0.315895f
C6451 VDAC_N.t23 VSS 0.506181f
C6452 VDAC_N.t21 VSS 0.505972f
C6453 VDAC_N.n10 VSS 0.565755f
C6454 VDAC_N.t17 VSS 0.505972f
C6455 VDAC_N.n11 VSS 0.296463f
C6456 VDAC_N.t22 VSS 0.505972f
C6457 VDAC_N.n12 VSS 0.305239f
C6458 VDAC_N.n13 VSS 0.242053f
C6459 VDAC_N.n14 VSS 0.39001f
C6460 VDAC_N.t0 VSS 0.343856f
C6461 VDAC_N.t3 VSS 0.343856f
C6462 VDAC_N.n15 VSS 1.31693f
C6463 VDAC_N.t2 VSS 0.343856f
C6464 VDAC_N.t5 VSS 0.343856f
C6465 VDAC_N.n16 VSS 1.28614f
C6466 VDAC_N.n17 VSS 1.81413f
C6467 VDAC_N.t1 VSS 0.343856f
C6468 VDAC_N.t7 VSS 0.343856f
C6469 VDAC_N.n18 VSS 1.31693f
C6470 VDAC_N.t4 VSS 0.343856f
C6471 VDAC_N.t6 VSS 0.343856f
C6472 VDAC_N.n19 VSS 1.28614f
C6473 VDAC_N.n20 VSS 1.81153f
C6474 VDAC_N.n21 VSS 1.67456f
C6475 VDAC_N.n22 VSS 45.5905f
C6476 a_17364_32525.t2 VSS 0.035856f
C6477 a_17364_32525.t3 VSS 0.035856f
C6478 a_17364_32525.n0 VSS 0.13279f
C6479 a_17364_32525.t4 VSS 1.46122f
C6480 a_17364_32525.n1 VSS 15.213599f
C6481 a_17364_32525.t0 VSS 0.055162f
C6482 a_17364_32525.n2 VSS 0.11037f
C6483 a_17364_32525.t1 VSS 0.055162f
C6484 w_10694_33990.n0 VSS 0.03242f
C6485 w_10694_33990.n1 VSS 0.034459f
C6486 w_10694_33990.n2 VSS 0.063869f
C6487 w_10694_33990.n3 VSS 0.074218f
C6488 w_10694_33990.n4 VSS 0.010162f
C6489 w_10694_33990.n5 VSS 0.147702f
C6490 w_10694_33990.n6 VSS 0.035533f
C6491 w_10694_33990.n7 VSS 0.285954f
C6492 w_10694_33990.n8 VSS 0.57917f
C6493 w_10694_33990.n9 VSS 0.255268f
C6494 w_10694_33990.n10 VSS 0.186992f
C6495 w_10694_33990.n11 VSS 1.44388f
C6496 w_10694_33990.t8 VSS 0.087008f
C6497 w_10694_33990.t5 VSS 0.018651f
C6498 w_10694_33990.n12 VSS 0.03807f
C6499 w_10694_33990.n13 VSS 2.76283f
C6500 w_10694_33990.t6 VSS 0.068357f
C6501 w_10694_33990.n14 VSS 1.4451f
C6502 w_10694_33990.n15 VSS 0.112291f
C6503 w_10694_33990.n16 VSS 0.66405f
C6504 w_10694_33990.n17 VSS 0.670596f
C6505 w_10694_33990.t17 VSS 0.086193f
C6506 w_10694_33990.n18 VSS 0.165131f
C6507 w_10694_33990.n19 VSS 0.157894f
C6508 w_10694_33990.n20 VSS 0.027781f
C6509 w_10694_33990.n21 VSS 0.027078f
C6510 w_10694_33990.n22 VSS 0.339416f
C6511 w_10694_33990.n23 VSS 0.028432f
C6512 w_10694_33990.t12 VSS 0.332239f
C6513 w_10694_33990.t10 VSS 0.168607f
C6514 w_10694_33990.t16 VSS 0.227151f
C6515 w_10694_33990.t14 VSS 0.168607f
C6516 w_10694_33990.n24 VSS 0.030935f
C6517 w_10694_33990.n25 VSS 0.027157f
C6518 w_10694_33990.t11 VSS 0.024969f
C6519 w_10694_33990.t15 VSS 0.024969f
C6520 w_10694_33990.n26 VSS 0.05604f
C6521 w_10694_33990.t13 VSS 0.091524f
C6522 w_10694_33990.n27 VSS 0.293976f
C6523 w_10694_33990.n28 VSS 0.039757f
C6524 w_10694_33990.n29 VSS 0.195444f
C6525 w_10694_33990.n30 VSS 0.074292f
C6526 w_10694_33990.n31 VSS 0.103874f
C6527 w_10694_33990.n32 VSS 0.026372f
C6528 w_10694_33990.n33 VSS 0.133386f
C6529 w_10694_33990.n34 VSS 0.022735f
C6530 w_10694_33990.n35 VSS 0.010162f
C6531 w_10694_33990.n36 VSS 0.088242f
C6532 w_10694_33990.t0 VSS 0.167665f
C6533 w_10694_33990.n37 VSS 0.108398f
C6534 w_10694_33990.n38 VSS 0.010162f
C6535 w_10694_33990.n39 VSS 0.022735f
C6536 w_10694_33990.n40 VSS 0.030935f
C6537 w_10694_33990.n41 VSS 0.011287f
C6538 w_10694_33990.n42 VSS 0.038036f
C6539 w_10694_33990.n43 VSS 0.112405f
C6540 w_10694_33990.n44 VSS 0.056392f
C6541 w_10694_33990.n45 VSS 0.037579f
C6542 w_10694_33990.n46 VSS 0.03779f
C6543 w_10694_33990.n47 VSS 0.081873f
C6544 w_10694_33990.n48 VSS 0.127359f
C6545 w_10694_33990.n49 VSS 0.088323f
C6546 w_10694_33990.n50 VSS 0.278854f
C6547 w_10694_33990.n51 VSS 1.44514f
C6548 w_10694_33990.t9 VSS 0.087008f
C6549 w_10694_33990.t3 VSS 0.018651f
C6550 w_10694_33990.n52 VSS 0.03807f
C6551 w_10694_33990.n53 VSS 2.76283f
C6552 w_10694_33990.t4 VSS 0.068357f
C6553 w_10694_33990.n54 VSS 1.44713f
C6554 w_10694_33990.n55 VSS 0.65106f
C6555 w_10694_33990.n56 VSS 0.614609f
C6556 w_10694_33990.n57 VSS 0.047876f
C6557 w_10694_33990.n58 VSS 0.145098f
C6558 w_10694_33990.n59 VSS 0.20272f
C6559 w_10694_33990.n60 VSS 0.158546f
C6560 w_10694_33990.n61 VSS 3.92883f
C6561 w_10694_33990.t2 VSS 6.74843f
C6562 w_10694_33990.n62 VSS 6.49835f
C6563 w_10694_33990.t7 VSS 6.71766f
C6564 w_10694_33990.n63 VSS 3.64426f
C6565 w_10694_33990.n64 VSS 0.156949f
C6566 w_10694_33990.n65 VSS 0.098091f
C6567 w_10694_33990.n66 VSS 0.035533f
C6568 w_10694_33990.n67 VSS 0.01988f
C6569 w_10694_33990.n68 VSS 0.024428f
C6570 w_10694_33990.n69 VSS 0.021603f
C6571 w_10694_33990.t1 VSS 0.020155f
C6572 a_n2661_44458.t1 VSS 0.059422f
C6573 a_n2661_44458.t3 VSS 0.026806f
C6574 a_n2661_44458.t4 VSS 0.017105f
C6575 a_n2661_44458.n0 VSS 0.77788f
C6576 a_n2661_44458.n1 VSS 5.61926f
C6577 a_n2661_44458.t2 VSS 0.016281f
C6578 a_n2661_44458.n2 VSS 0.027569f
C6579 a_n2661_44458.n3 VSS 0.034535f
C6580 a_n2661_44458.n4 VSS 0.015858f
C6581 a_5742_30871.t0 VSS 0.03516f
C6582 a_5742_30871.t5 VSS 0.111338f
C6583 a_5742_30871.t8 VSS 0.128026f
C6584 a_5742_30871.n0 VSS 0.49678f
C6585 a_5742_30871.t4 VSS 0.111338f
C6586 a_5742_30871.t6 VSS 0.128026f
C6587 a_5742_30871.n1 VSS 0.430179f
C6588 a_5742_30871.n2 VSS 11.229099f
C6589 a_5742_30871.t9 VSS 0.054693f
C6590 a_5742_30871.t7 VSS 0.03411f
C6591 a_5742_30871.n3 VSS 0.127149f
C6592 a_5742_30871.n4 VSS 6.79781f
C6593 a_5742_30871.t3 VSS 0.022854f
C6594 a_5742_30871.t2 VSS 0.022854f
C6595 a_5742_30871.n5 VSS 0.045707f
C6596 a_5742_30871.n6 VSS 0.28425f
C6597 a_5742_30871.n7 VSS 0.105502f
C6598 a_5742_30871.t1 VSS 0.03516f
C6599 SMPL_ON_P.t9 VSS 0.040546f
C6600 SMPL_ON_P.t8 VSS 0.065013f
C6601 SMPL_ON_P.n0 VSS 0.277894f
C6602 SMPL_ON_P.t5 VSS 0.027166f
C6603 SMPL_ON_P.t7 VSS 0.027166f
C6604 SMPL_ON_P.n1 VSS 0.083843f
C6605 SMPL_ON_P.t4 VSS 0.027166f
C6606 SMPL_ON_P.t6 VSS 0.027166f
C6607 SMPL_ON_P.n2 VSS 0.059996f
C6608 SMPL_ON_P.n3 VSS 0.324651f
C6609 SMPL_ON_P.t0 VSS 0.041793f
C6610 SMPL_ON_P.t2 VSS 0.041793f
C6611 SMPL_ON_P.n4 VSS 0.127258f
C6612 SMPL_ON_P.t3 VSS 0.041793f
C6613 SMPL_ON_P.t1 VSS 0.041793f
C6614 SMPL_ON_P.n5 VSS 0.092582f
C6615 SMPL_ON_P.n6 VSS 0.44185f
C6616 SMPL_ON_P.n7 VSS 5.77296f
C6617 COMP_P.t1 VSS 0.030382f
C6618 COMP_P.t0 VSS 0.030382f
C6619 COMP_P.n0 VSS 0.067302f
C6620 COMP_P.t3 VSS 0.030382f
C6621 COMP_P.t2 VSS 0.030382f
C6622 COMP_P.n1 VSS 0.09251f
C6623 COMP_P.n2 VSS 0.322778f
C6624 COMP_P.t4 VSS 0.019748f
C6625 COMP_P.t7 VSS 0.019748f
C6626 COMP_P.n3 VSS 0.06095f
C6627 COMP_P.t6 VSS 0.019748f
C6628 COMP_P.t5 VSS 0.019748f
C6629 COMP_P.n4 VSS 0.043614f
C6630 COMP_P.n5 VSS 0.237297f
C6631 COMP_P.n6 VSS 0.119216f
C6632 COMP_P.t10 VSS 0.050694f
C6633 COMP_P.t9 VSS 0.027786f
C6634 COMP_P.n7 VSS 0.210023f
C6635 COMP_P.t8 VSS 0.031402f
C6636 COMP_P.t11 VSS 0.050293f
C6637 COMP_P.n8 VSS 2.91043f
C6638 COMP_P.n9 VSS 10.529799f
C6639 a_n1741_47186.t4 VSS 0.018856f
C6640 a_n1741_47186.t5 VSS 0.018856f
C6641 a_n1741_47186.n0 VSS 0.038054f
C6642 a_n1741_47186.t8 VSS 0.025145f
C6643 a_n1741_47186.t9 VSS 0.039404f
C6644 a_n1741_47186.n1 VSS 1.34953f
C6645 a_n1741_47186.n2 VSS 8.13925f
C6646 a_n1741_47186.t3 VSS 0.029009f
C6647 a_n1741_47186.t2 VSS 0.029009f
C6648 a_n1741_47186.n3 VSS 0.061932f
C6649 a_n1741_47186.n4 VSS 0.163192f
C6650 a_n1741_47186.t7 VSS 0.029009f
C6651 a_n1741_47186.t6 VSS 0.029009f
C6652 a_n1741_47186.n5 VSS 0.062191f
C6653 a_n1741_47186.n6 VSS 0.223111f
C6654 a_n1741_47186.t0 VSS 0.029009f
C6655 a_n1741_47186.n7 VSS 0.086432f
C6656 a_n1741_47186.t1 VSS 0.029009f
C6657 a_n443_42852.t1 VSS 0.019211f
C6658 a_n443_42852.t4 VSS 0.012487f
C6659 a_n443_42852.t6 VSS 0.012487f
C6660 a_n443_42852.n0 VSS 0.048023f
C6661 a_n443_42852.t7 VSS 0.012487f
C6662 a_n443_42852.t5 VSS 0.012487f
C6663 a_n443_42852.n1 VSS 0.028533f
C6664 a_n443_42852.n2 VSS 0.15892f
C6665 a_n443_42852.t17 VSS 0.01395f
C6666 a_n443_42852.t13 VSS 0.013014f
C6667 a_n443_42852.n3 VSS 0.065551f
C6668 a_n443_42852.t14 VSS 0.03167f
C6669 a_n443_42852.t12 VSS 0.065775f
C6670 a_n443_42852.n4 VSS 1.41345f
C6671 a_n443_42852.t20 VSS 0.01414f
C6672 a_n443_42852.t22 VSS 0.017129f
C6673 a_n443_42852.n5 VSS 0.353441f
C6674 a_n443_42852.t21 VSS 0.026036f
C6675 a_n443_42852.t11 VSS 0.017738f
C6676 a_n443_42852.n6 VSS 0.064904f
C6677 a_n443_42852.n7 VSS 2.30852f
C6678 a_n443_42852.t19 VSS 0.031994f
C6679 a_n443_42852.t24 VSS 0.019821f
C6680 a_n443_42852.n8 VSS 0.075058f
C6681 a_n443_42852.n9 VSS 2.90642f
C6682 a_n443_42852.t8 VSS 0.01761f
C6683 a_n443_42852.t25 VSS 0.029884f
C6684 a_n443_42852.t9 VSS 0.01761f
C6685 a_n443_42852.t10 VSS 0.029884f
C6686 a_n443_42852.n10 VSS 0.050141f
C6687 a_n443_42852.n11 VSS 0.075573f
C6688 a_n443_42852.n12 VSS 0.524192f
C6689 a_n443_42852.n13 VSS 0.832394f
C6690 a_n443_42852.t16 VSS 0.012818f
C6691 a_n443_42852.t18 VSS 0.013727f
C6692 a_n443_42852.n14 VSS 0.052066f
C6693 a_n443_42852.n15 VSS 0.102646f
C6694 a_n443_42852.t23 VSS 0.02033f
C6695 a_n443_42852.t15 VSS 0.032375f
C6696 a_n443_42852.n16 VSS 0.04599f
C6697 a_n443_42852.n17 VSS 0.178545f
C6698 a_n443_42852.n18 VSS 0.098927f
C6699 a_n443_42852.t2 VSS 0.019211f
C6700 a_n443_42852.t0 VSS 0.019211f
C6701 a_n443_42852.n19 VSS 0.042906f
C6702 a_n443_42852.n20 VSS 0.16317f
C6703 a_n443_42852.n21 VSS 0.058337f
C6704 a_n443_42852.t3 VSS 0.019211f
C6705 a_8696_44636.t4 VSS 0.029695f
C6706 a_8696_44636.t3 VSS 0.017499f
C6707 a_8696_44636.n0 VSS 0.079251f
C6708 a_8696_44636.t5 VSS 0.019335f
C6709 a_8696_44636.t6 VSS 0.014051f
C6710 a_8696_44636.n1 VSS 0.042181f
C6711 a_8696_44636.t7 VSS 0.01364f
C6712 a_8696_44636.t9 VSS 0.016512f
C6713 a_8696_44636.n2 VSS 0.226971f
C6714 a_8696_44636.n3 VSS 3.69645f
C6715 a_8696_44636.t2 VSS 0.016502f
C6716 a_8696_44636.t8 VSS 0.013632f
C6717 a_8696_44636.n4 VSS 0.062351f
C6718 a_8696_44636.n5 VSS 0.200459f
C6719 a_8696_44636.n6 VSS 0.191216f
C6720 a_8696_44636.t1 VSS 0.043594f
C6721 a_8696_44636.n7 VSS 0.139889f
C6722 a_8696_44636.t0 VSS 0.076774f
C6723 a_n1057_35014.t0 VSS 0.036613f
C6724 a_n1057_35014.n0 VSS 1.87506f
C6725 a_n1057_35014.n1 VSS 1.90362f
C6726 a_n1057_35014.n2 VSS 0.577258f
C6727 a_n1057_35014.n3 VSS 1.73867f
C6728 a_n1057_35014.n4 VSS 0.445111f
C6729 a_n1057_35014.t5 VSS 5.31306f
C6730 a_n1057_35014.n5 VSS 4.34405f
C6731 a_n1057_35014.t6 VSS 5.31306f
C6732 a_n1057_35014.n6 VSS 1.81069f
C6733 a_n1057_35014.n7 VSS 0.484f
C6734 a_n1057_35014.n8 VSS 0.21532f
C6735 a_n1057_35014.n9 VSS 0.174526f
C6736 a_n1057_35014.n10 VSS 0.420322f
C6737 a_n1057_35014.n11 VSS 0.445839f
C6738 a_n1057_35014.t4 VSS 5.31306f
C6739 a_n1057_35014.t7 VSS 5.31306f
C6740 a_n1057_35014.n12 VSS 4.14858f
C6741 a_n1057_35014.n13 VSS 0.472991f
C6742 a_n1057_35014.n14 VSS 0.492963f
C6743 a_n1057_35014.t2 VSS 0.036613f
C6744 a_n1057_35014.t3 VSS 0.036613f
C6745 a_n1057_35014.n15 VSS 0.093314f
C6746 a_n1057_35014.n16 VSS 0.559196f
C6747 a_n1057_35014.n17 VSS 0.099788f
C6748 a_n1057_35014.t1 VSS 0.036613f
C6749 a_2711_45572.n0 VSS 0.014123f
C6750 a_2711_45572.t4 VSS 0.013151f
C6751 a_2711_45572.n1 VSS 0.109517f
C6752 a_2711_45572.t7 VSS 0.015734f
C6753 a_2711_45572.n2 VSS 0.021444f
C6754 a_2711_45572.n3 VSS 1.0594f
C6755 a_2711_45572.t11 VSS 0.015734f
C6756 a_2711_45572.n4 VSS 0.029102f
C6757 a_2711_45572.n5 VSS 2.17871f
C6758 a_2711_45572.t8 VSS 0.013151f
C6759 a_2711_45572.n6 VSS 0.031902f
C6760 a_2711_45572.n7 VSS 0.689222f
C6761 a_2711_45572.n8 VSS 0.112965f
C6762 a_2711_45572.n9 VSS 0.028492f
C6763 VIN_P.t9 VSS 0.268837f
C6764 VIN_P.t10 VSS 0.265605f
C6765 VIN_P.n0 VSS 1.60998f
C6766 VIN_P.t0 VSS 0.144996f
C6767 VIN_P.t5 VSS 0.144996f
C6768 VIN_P.n1 VSS 0.513004f
C6769 VIN_P.t12 VSS 0.062178f
C6770 VIN_P.t11 VSS 0.060662f
C6771 VIN_P.n2 VSS 0.20897f
C6772 VIN_P.t7 VSS 0.06066f
C6773 VIN_P.n3 VSS 0.113566f
C6774 VIN_P.t2 VSS 0.064106f
C6775 VIN_P.n4 VSS 0.172747f
C6776 VIN_P.t15 VSS 0.063671f
C6777 VIN_P.n5 VSS 0.140791f
C6778 VIN_P.t6 VSS 0.063671f
C6779 VIN_P.n6 VSS 0.152702f
C6780 VIN_P.t8 VSS 0.063671f
C6781 VIN_P.n7 VSS 0.152702f
C6782 VIN_P.t1 VSS 0.063671f
C6783 VIN_P.n8 VSS 0.163687f
C6784 VIN_P.t3 VSS 0.036249f
C6785 VIN_P.t14 VSS 0.036249f
C6786 VIN_P.n9 VSS 0.098859f
C6787 VIN_P.n10 VSS 0.216413f
C6788 VIN_P.t13 VSS 0.136218f
C6789 VIN_P.n11 VSS 0.814626f
C6790 VIN_P.n12 VSS 0.960503f
C6791 VIN_P.t4 VSS 0.674566f
C6792 VIN_P.n13 VSS 1.45115f
C6793 VIN_P.n14 VSS 6.8455f
C6794 a_3754_38470.t7 VSS 0.029992f
C6795 a_3754_38470.t10 VSS 0.029993f
C6796 a_3754_38470.t6 VSS 0.02996f
C6797 a_3754_38470.n0 VSS 0.086396f
C6798 a_3754_38470.t8 VSS 0.029993f
C6799 a_3754_38470.t3 VSS 0.02996f
C6800 a_3754_38470.n1 VSS 0.083014f
C6801 a_3754_38470.n2 VSS 0.053306f
C6802 a_3754_38470.t9 VSS 0.029992f
C6803 a_3754_38470.t4 VSS 0.02996f
C6804 a_3754_38470.n3 VSS 0.088448f
C6805 a_3754_38470.n4 VSS 0.053306f
C6806 a_3754_38470.t5 VSS 0.02996f
C6807 a_3754_38470.n5 VSS 0.029854f
C6808 a_3754_38470.n6 VSS 0.071966f
C6809 a_3754_38470.t2 VSS 0.034572f
C6810 a_3754_38470.n7 VSS 0.413441f
C6811 a_3754_38470.t1 VSS 0.044659f
C6812 a_3754_38470.n8 VSS 0.933763f
C6813 a_3754_38470.t0 VSS 0.367463f
C6814 a_13717_47436.t3 VSS 0.068802f
C6815 a_13717_47436.t2 VSS 0.109568f
C6816 a_13717_47436.n0 VSS 1.43054f
C6817 a_13717_47436.t1 VSS 0.116329f
C6818 a_13717_47436.n1 VSS 6.94383f
C6819 a_13717_47436.t0 VSS 0.230934f
C6820 a_1273_38525.t1 VSS 0.016522f
C6821 a_1273_38525.t2 VSS 0.016522f
C6822 a_1273_38525.t0 VSS 0.016522f
C6823 a_1273_38525.n0 VSS 0.039533f
C6824 a_1273_38525.t7 VSS 0.010739f
C6825 a_1273_38525.t5 VSS 0.010739f
C6826 a_1273_38525.n1 VSS 0.02697f
C6827 a_1273_38525.t4 VSS 0.010739f
C6828 a_1273_38525.t6 VSS 0.010739f
C6829 a_1273_38525.n2 VSS 0.022828f
C6830 a_1273_38525.n3 VSS 0.085426f
C6831 a_1273_38525.t11 VSS 0.060909f
C6832 a_1273_38525.t8 VSS 0.058644f
C6833 a_1273_38525.n4 VSS 0.525844f
C6834 a_1273_38525.n5 VSS 0.234962f
C6835 a_1273_38525.t13 VSS 0.060841f
C6836 a_1273_38525.t10 VSS 0.058639f
C6837 a_1273_38525.n6 VSS 0.634717f
C6838 a_1273_38525.t12 VSS 0.071684f
C6839 a_1273_38525.n7 VSS 0.290078f
C6840 a_1273_38525.t9 VSS 0.071685f
C6841 a_1273_38525.n8 VSS 0.252398f
C6842 a_1273_38525.n9 VSS 0.32433f
C6843 a_1273_38525.n10 VSS 0.120033f
C6844 a_1273_38525.n11 VSS 0.115928f
C6845 a_1273_38525.n12 VSS 0.035505f
C6846 a_1273_38525.t3 VSS 0.016522f
C6847 a_19479_31679.t0 VSS 0.056919f
C6848 a_19479_31679.t4 VSS 2.66617f
C6849 a_19479_31679.t2 VSS 0.036998f
C6850 a_19479_31679.t3 VSS 0.036998f
C6851 a_19479_31679.n0 VSS 0.073995f
C6852 a_19479_31679.n1 VSS 14.9012f
C6853 a_19479_31679.n2 VSS 0.170796f
C6854 a_19479_31679.t1 VSS 0.056919f
C6855 a_15227_44166.t14 VSS 0.015806f
C6856 a_15227_44166.n0 VSS 0.02596f
C6857 a_15227_44166.n1 VSS 0.019901f
C6858 a_15227_44166.t10 VSS 0.010006f
C6859 a_15227_44166.t7 VSS 0.015935f
C6860 a_15227_44166.n2 VSS 0.036323f
C6861 a_15227_44166.t15 VSS 0.016379f
C6862 a_15227_44166.n3 VSS 0.029978f
C6863 a_15227_44166.n4 VSS 0.294522f
C6864 a_15227_44166.t12 VSS 0.015935f
C6865 a_15227_44166.t4 VSS 0.010006f
C6866 a_15227_44166.n5 VSS 0.024086f
C6867 a_15227_44166.t9 VSS 0.012634f
C6868 a_15227_44166.n6 VSS 0.039462f
C6869 a_15227_44166.t16 VSS 0.014709f
C6870 a_15227_44166.n7 VSS 0.018786f
C6871 a_15227_44166.t5 VSS 0.014709f
C6872 a_15227_44166.n8 VSS 0.020866f
C6873 a_15227_44166.n9 VSS 0.014304f
C6874 a_15227_44166.t25 VSS 0.016377f
C6875 a_15227_44166.n10 VSS 0.033317f
C6876 a_15227_44166.n11 VSS 0.306929f
C6877 a_15227_44166.n12 VSS 0.190119f
C6878 a_15227_44166.n13 VSS 0.145795f
C6879 a_15227_44166.n14 VSS 0.115162f
C6880 a_15227_44166.n15 VSS 0.020473f
C6881 a_15227_44166.n16 VSS 0.10391f
C6882 a_15227_44166.n17 VSS 0.162159f
C6883 a_15227_44166.n18 VSS 0.295897f
C6884 a_15227_44166.t13 VSS 0.019131f
C6885 a_15227_44166.n19 VSS 0.032293f
C6886 a_15227_44166.n20 VSS 0.347652f
C6887 a_15227_44166.n21 VSS 0.012293f
C6888 a_15227_44166.n22 VSS 0.094211f
C6889 a_15227_44166.n23 VSS 0.028374f
C6890 a_19692_46634.t1 VSS 0.01118f
C6891 a_19692_46634.t2 VSS 0.061503f
C6892 a_19692_46634.t11 VSS 0.028513f
C6893 a_19692_46634.t10 VSS 0.017812f
C6894 a_19692_46634.n0 VSS 0.084119f
C6895 a_19692_46634.t4 VSS 0.023029f
C6896 a_19692_46634.t3 VSS 0.01266f
C6897 a_19692_46634.n1 VSS 0.04558f
C6898 a_19692_46634.t12 VSS 0.015881f
C6899 a_19692_46634.t7 VSS 0.019663f
C6900 a_19692_46634.n2 VSS 0.10453f
C6901 a_19692_46634.n3 VSS 0.147521f
C6902 a_19692_46634.n4 VSS 0.697911f
C6903 a_19692_46634.t8 VSS 0.026756f
C6904 a_19692_46634.t9 VSS 0.015767f
C6905 a_19692_46634.n5 VSS 0.036273f
C6906 a_19692_46634.t6 VSS 0.026756f
C6907 a_19692_46634.t5 VSS 0.015767f
C6908 a_19692_46634.n6 VSS 0.036273f
C6909 a_19692_46634.n7 VSS 0.045244f
C6910 a_19692_46634.n8 VSS 0.805821f
C6911 a_19692_46634.n9 VSS 0.152509f
C6912 a_19692_46634.n10 VSS 0.057753f
C6913 a_19692_46634.t0 VSS 0.01118f
C6914 a_n4318_39304.t3 VSS 0.027585f
C6915 a_n4318_39304.t2 VSS 0.027585f
C6916 a_n4318_39304.n0 VSS 0.102161f
C6917 a_n4318_39304.t4 VSS 0.044402f
C6918 a_n4318_39304.t5 VSS 0.070898f
C6919 a_n4318_39304.n1 VSS 1.03911f
C6920 a_n4318_39304.n2 VSS 4.31847f
C6921 a_n4318_39304.t0 VSS 0.042439f
C6922 a_n4318_39304.n3 VSS 0.084912f
C6923 a_n4318_39304.t1 VSS 0.042439f
C6924 a_n2956_39304.t4 VSS 0.060807f
C6925 a_n2956_39304.t5 VSS 0.097476f
C6926 a_n2956_39304.n0 VSS 2.37214f
C6927 a_n2956_39304.t3 VSS 0.038371f
C6928 a_n2956_39304.t2 VSS 0.038371f
C6929 a_n2956_39304.n1 VSS 0.076743f
C6930 a_n2956_39304.n2 VSS 9.420889f
C6931 a_n2956_39304.t0 VSS 0.059033f
C6932 a_n2956_39304.n3 VSS 0.177139f
C6933 a_n2956_39304.t1 VSS 0.059033f
C6934 a_5934_30871.t0 VSS 0.059171f
C6935 a_5934_30871.t4 VSS 0.443837f
C6936 a_5934_30871.t6 VSS 0.412182f
C6937 a_5934_30871.n0 VSS 19.026999f
C6938 a_5934_30871.t7 VSS 0.092045f
C6939 a_5934_30871.t5 VSS 0.057405f
C6940 a_5934_30871.n1 VSS 0.269364f
C6941 a_5934_30871.n2 VSS 11.3934f
C6942 a_5934_30871.t3 VSS 0.038461f
C6943 a_5934_30871.t2 VSS 0.038461f
C6944 a_5934_30871.n3 VSS 0.076922f
C6945 a_5934_30871.n4 VSS 0.455085f
C6946 a_5934_30871.n5 VSS 0.177553f
C6947 a_5934_30871.t1 VSS 0.059171f
C6948 a_13507_46334.t1 VSS 0.027351f
C6949 a_13507_46334.t4 VSS 0.013373f
C6950 a_13507_46334.n0 VSS 0.037272f
C6951 a_13507_46334.n1 VSS 0.117224f
C6952 a_13507_46334.t11 VSS 0.010429f
C6953 a_13507_46334.t3 VSS 0.016833f
C6954 a_13507_46334.n2 VSS 0.035028f
C6955 a_13507_46334.t13 VSS 0.015344f
C6956 a_13507_46334.n3 VSS 0.118627f
C6957 a_13507_46334.n4 VSS 0.812176f
C6958 a_13507_46334.t2 VSS 0.014238f
C6959 a_13507_46334.n5 VSS 0.035768f
C6960 a_13507_46334.n6 VSS 0.352271f
C6961 a_13507_46334.t6 VSS 0.016865f
C6962 a_13507_46334.n7 VSS 0.038933f
C6963 a_13507_46334.t5 VSS 0.016865f
C6964 a_13507_46334.n8 VSS 0.036322f
C6965 a_13507_46334.n9 VSS 1.29738f
C6966 a_13507_46334.n10 VSS 0.90886f
C6967 a_13507_46334.n11 VSS 0.095082f
C6968 a_13507_46334.t0 VSS 0.039857f
C6969 a_n3420_37984.t1 VSS 0.057946f
C6970 a_n3420_37984.t6 VSS 0.037665f
C6971 a_n3420_37984.t5 VSS 0.037665f
C6972 a_n3420_37984.n0 VSS 0.078068f
C6973 a_n3420_37984.t7 VSS 0.037665f
C6974 a_n3420_37984.t4 VSS 0.037665f
C6975 a_n3420_37984.n1 VSS 0.092642f
C6976 a_n3420_37984.n2 VSS 0.34569f
C6977 a_n3420_37984.t9 VSS 1.22031f
C6978 a_n3420_37984.t8 VSS 0.059131f
C6979 a_n3420_37984.t10 VSS 0.094166f
C6980 a_n3420_37984.n3 VSS 0.136687f
C6981 a_n3420_37984.n4 VSS 12.295401f
C6982 a_n3420_37984.n5 VSS 0.223115f
C6983 a_n3420_37984.t2 VSS 0.057946f
C6984 a_n3420_37984.t0 VSS 0.057946f
C6985 a_n3420_37984.n6 VSS 0.14933f
C6986 a_n3420_37984.n7 VSS 0.40121f
C6987 a_n3420_37984.n8 VSS 0.121794f
C6988 a_n3420_37984.t3 VSS 0.057946f
C6989 a_n4315_30879.n0 VSS 0.030923f
C6990 a_n4315_30879.n1 VSS 0.018381f
C6991 a_n4315_30879.n2 VSS 0.099492f
C6992 a_n4315_30879.t18 VSS 0.013186f
C6993 a_n4315_30879.t19 VSS 0.020998f
C6994 a_n4315_30879.n3 VSS 0.04468f
C6995 a_n4315_30879.t12 VSS 0.421831f
C6996 a_n4315_30879.t13 VSS 0.421766f
C6997 a_n4315_30879.n4 VSS 0.311515f
C6998 a_n4315_30879.t14 VSS 0.421766f
C6999 a_n4315_30879.n5 VSS 0.158559f
C7000 a_n4315_30879.t9 VSS 0.421766f
C7001 a_n4315_30879.n6 VSS 0.158559f
C7002 a_n4315_30879.t24 VSS 0.421766f
C7003 a_n4315_30879.n7 VSS 0.158559f
C7004 a_n4315_30879.t11 VSS 0.421766f
C7005 a_n4315_30879.n8 VSS 0.158559f
C7006 a_n4315_30879.t25 VSS 0.421766f
C7007 a_n4315_30879.n9 VSS 0.158559f
C7008 a_n4315_30879.t21 VSS 0.421766f
C7009 a_n4315_30879.n10 VSS 0.158559f
C7010 a_n4315_30879.t15 VSS 0.421766f
C7011 a_n4315_30879.n11 VSS 0.158559f
C7012 a_n4315_30879.t23 VSS 0.421766f
C7013 a_n4315_30879.n12 VSS 0.158559f
C7014 a_n4315_30879.t17 VSS 0.421766f
C7015 a_n4315_30879.n13 VSS 0.158559f
C7016 a_n4315_30879.t10 VSS 0.421766f
C7017 a_n4315_30879.n14 VSS 0.158559f
C7018 a_n4315_30879.t16 VSS 0.421766f
C7019 a_n4315_30879.n15 VSS 0.158559f
C7020 a_n4315_30879.t22 VSS 0.421766f
C7021 a_n4315_30879.n16 VSS 0.158559f
C7022 a_n4315_30879.t20 VSS 0.421766f
C7023 a_n4315_30879.n17 VSS 0.158254f
C7024 a_n4315_30879.t8 VSS 0.421766f
C7025 a_n4315_30879.n18 VSS 1.17914f
C7026 a_n4315_30879.n19 VSS 1.27875f
C7027 a_n4315_30879.n20 VSS 0.050661f
C7028 a_n4315_30879.t2 VSS 0.01246f
C7029 a_n4315_30879.t1 VSS 0.01246f
C7030 a_n4315_30879.n21 VSS 0.025632f
C7031 a_n4315_30879.n22 VSS 0.103414f
C7032 a_n4315_30879.t0 VSS 0.01246f
C7033 a_n4315_30879.n23 VSS 0.031712f
C7034 a_n4315_30879.t3 VSS 0.01246f
C7035 a_n3674_39304.t0 VSS 0.039449f
C7036 a_n3674_39304.t3 VSS 0.025642f
C7037 a_n3674_39304.t2 VSS 0.025642f
C7038 a_n3674_39304.n0 VSS 0.089167f
C7039 a_n3674_39304.t4 VSS 0.041274f
C7040 a_n3674_39304.t5 VSS 0.065904f
C7041 a_n3674_39304.n1 VSS 0.966541f
C7042 a_n3674_39304.n2 VSS 4.52621f
C7043 a_n3674_39304.n3 VSS 0.080724f
C7044 a_n3674_39304.t1 VSS 0.039449f
C7045 a_n1925_46634.t1 VSS 0.022876f
C7046 a_n1925_46634.t4 VSS 0.022897f
C7047 a_n1925_46634.t5 VSS 0.014611f
C7048 a_n1925_46634.n0 VSS 0.65448f
C7049 a_n1925_46634.t3 VSS 0.122746f
C7050 a_n1925_46634.t2 VSS 0.118458f
C7051 a_n1925_46634.n1 VSS 0.283321f
C7052 a_n1925_46634.n2 VSS 3.48918f
C7053 a_n1925_46634.n3 VSS 0.047354f
C7054 a_n1925_46634.t0 VSS 0.024081f
C7055 a_n3420_39616.t0 VSS 0.047804f
C7056 a_n3420_39616.t6 VSS 0.031072f
C7057 a_n3420_39616.t5 VSS 0.031072f
C7058 a_n3420_39616.n0 VSS 0.064403f
C7059 a_n3420_39616.t7 VSS 0.031072f
C7060 a_n3420_39616.t4 VSS 0.031072f
C7061 a_n3420_39616.n1 VSS 0.076426f
C7062 a_n3420_39616.n2 VSS 0.28518f
C7063 a_n3420_39616.t9 VSS 0.077683f
C7064 a_n3420_39616.t8 VSS 0.04878f
C7065 a_n3420_39616.n3 VSS 0.112418f
C7066 a_n3420_39616.t10 VSS 0.606935f
C7067 a_n3420_39616.t11 VSS 0.624337f
C7068 a_n3420_39616.n4 VSS 2.16864f
C7069 a_n3420_39616.n5 VSS 7.88099f
C7070 a_n3420_39616.n6 VSS 0.184059f
C7071 a_n3420_39616.t2 VSS 0.047804f
C7072 a_n3420_39616.t1 VSS 0.047804f
C7073 a_n3420_39616.n7 VSS 0.123191f
C7074 a_n3420_39616.n8 VSS 0.330982f
C7075 a_n3420_39616.n9 VSS 0.100476f
C7076 a_n3420_39616.t3 VSS 0.047804f
C7077 a_20205_31679.t0 VSS 0.058088f
C7078 a_20205_31679.t2 VSS 0.037757f
C7079 a_20205_31679.t3 VSS 0.037757f
C7080 a_20205_31679.n0 VSS 0.139831f
C7081 a_20205_31679.t4 VSS 2.88037f
C7082 a_20205_31679.n1 VSS 14.6719f
C7083 a_20205_31679.n2 VSS 0.116222f
C7084 a_20205_31679.t1 VSS 0.058088f
C7085 a_17538_32519.t0 VSS 0.057897f
C7086 a_17538_32519.t2 VSS 0.037633f
C7087 a_17538_32519.t3 VSS 0.037633f
C7088 a_17538_32519.n0 VSS 0.130863f
C7089 a_17538_32519.t5 VSS 0.762306f
C7090 a_17538_32519.t4 VSS 0.784162f
C7091 a_17538_32519.n1 VSS 4.32327f
C7092 a_17538_32519.n2 VSS 12.6899f
C7093 a_17538_32519.n3 VSS 0.118472f
C7094 a_17538_32519.t1 VSS 0.057897f
C7095 C9_N_btm.t9 VSS 0.137574f
C7096 C9_N_btm.t10 VSS 0.137574f
C7097 C9_N_btm.n0 VSS 0.439559f
C7098 C9_N_btm.t14 VSS 0.137574f
C7099 C9_N_btm.t16 VSS 0.137574f
C7100 C9_N_btm.n1 VSS 0.425131f
C7101 C9_N_btm.n2 VSS 1.33616f
C7102 C9_N_btm.t15 VSS 0.137574f
C7103 C9_N_btm.t13 VSS 0.137574f
C7104 C9_N_btm.n3 VSS 0.425131f
C7105 C9_N_btm.n4 VSS 0.684407f
C7106 C9_N_btm.t11 VSS 0.137574f
C7107 C9_N_btm.t12 VSS 0.137574f
C7108 C9_N_btm.n5 VSS 0.425131f
C7109 C9_N_btm.n6 VSS 1.08525f
C7110 C9_N_btm.t5 VSS 0.156549f
C7111 C9_N_btm.t6 VSS 0.156549f
C7112 C9_N_btm.n7 VSS 0.645454f
C7113 C9_N_btm.t4 VSS 0.156549f
C7114 C9_N_btm.t7 VSS 0.156549f
C7115 C9_N_btm.n8 VSS 0.630592f
C7116 C9_N_btm.n9 VSS 1.02683f
C7117 C9_N_btm.n10 VSS 0.61298f
C7118 C9_N_btm.t8 VSS 0.961787f
C7119 C9_N_btm.n11 VSS 0.767348f
C7120 C9_N_btm.t0 VSS 0.156549f
C7121 C9_N_btm.t2 VSS 0.156549f
C7122 C9_N_btm.n12 VSS 0.63781f
C7123 C9_N_btm.t3 VSS 0.156549f
C7124 C9_N_btm.t1 VSS 0.156549f
C7125 C9_N_btm.n13 VSS 0.651901f
C7126 C9_N_btm.n14 VSS 1.03801f
C7127 C9_N_btm.n15 VSS 2.51129f
C7128 C9_N_btm.n16 VSS 2.29472f
C7129 C9_N_btm.n17 VSS 1.01629f
C7130 C9_N_btm.n18 VSS 1.01985f
C7131 C9_N_btm.n19 VSS 1.01985f
C7132 C9_N_btm.n20 VSS 1.01629f
C7133 C9_N_btm.n21 VSS 1.01985f
C7134 C9_N_btm.n22 VSS 1.01985f
C7135 C9_N_btm.n23 VSS 1.01985f
C7136 C9_N_btm.n24 VSS 1.01985f
C7137 C9_N_btm.n25 VSS 1.01629f
C7138 C9_N_btm.n26 VSS 1.01985f
C7139 C9_N_btm.n27 VSS 1.01985f
C7140 C9_N_btm.n28 VSS 1.01629f
C7141 C9_N_btm.n29 VSS 1.01985f
C7142 C9_N_btm.n30 VSS 1.01985f
C7143 C9_N_btm.n31 VSS 1.01985f
C7144 C9_N_btm.n32 VSS 1.01985f
C7145 C9_N_btm.n33 VSS 1.01629f
C7146 C9_N_btm.n34 VSS 1.01985f
C7147 C9_N_btm.n35 VSS 1.01985f
C7148 C9_N_btm.n36 VSS 1.01629f
C7149 C9_N_btm.n37 VSS 1.01985f
C7150 C9_N_btm.n38 VSS 1.01985f
C7151 C9_N_btm.n39 VSS 1.01985f
C7152 C9_N_btm.n40 VSS 1.28199f
C7153 C9_N_btm.n41 VSS 1.01985f
C7154 C9_N_btm.n42 VSS 1.01985f
C7155 C9_N_btm.n43 VSS 1.01985f
C7156 C9_N_btm.n44 VSS 1.01985f
C7157 C9_N_btm.n45 VSS 1.01985f
C7158 C9_N_btm.n46 VSS 1.01985f
C7159 C9_N_btm.n47 VSS 1.01985f
C7160 C9_N_btm.n48 VSS 1.02004f
C7161 C9_N_btm.n49 VSS 1.01985f
C7162 C9_N_btm.n50 VSS 0.750397f
C7163 C9_N_btm.n51 VSS 1.02004f
C7164 C9_N_btm.n52 VSS 1.01985f
C7165 C9_N_btm.n53 VSS 1.01985f
C7166 C9_N_btm.n54 VSS 1.01985f
C7167 C9_N_btm.n55 VSS 1.01985f
C7168 C9_N_btm.n56 VSS 1.01985f
C7169 C9_N_btm.n57 VSS 1.01985f
C7170 C9_N_btm.n58 VSS 1.01629f
C7171 C9_N_btm.n59 VSS 1.01629f
C7172 C9_N_btm.n60 VSS 1.01985f
C7173 C9_N_btm.n61 VSS 1.02004f
C7174 C9_N_btm.n62 VSS 0.750397f
C7175 C9_N_btm.n63 VSS 0.750397f
C7176 C9_N_btm.n64 VSS 1.02004f
C7177 C9_N_btm.n65 VSS 1.02004f
C7178 C9_N_btm.n66 VSS 1.45446f
C7179 C9_N_btm.n67 VSS 1.59744f
C7180 C9_N_btm.n68 VSS 1.22831f
C7181 C9_N_btm.n69 VSS 1.01985f
C7182 C9_N_btm.n70 VSS 1.01985f
C7183 C9_N_btm.n71 VSS 1.01985f
C7184 C9_N_btm.n72 VSS 1.01985f
C7185 C9_N_btm.n73 VSS 1.01629f
C7186 C9_N_btm.n74 VSS 1.01629f
C7187 C9_N_btm.n75 VSS 1.01629f
C7188 C9_N_btm.n76 VSS 1.01629f
C7189 C9_N_btm.n77 VSS 1.01985f
C7190 C9_N_btm.n78 VSS 1.01629f
C7191 C9_N_btm.n79 VSS 1.01985f
C7192 C9_N_btm.n80 VSS 1.01985f
C7193 C9_N_btm.n81 VSS 1.01985f
C7194 C9_N_btm.n82 VSS 1.01629f
C7195 C9_N_btm.n83 VSS 1.01985f
C7196 C9_N_btm.n84 VSS 1.01985f
C7197 C9_N_btm.n85 VSS 1.01985f
C7198 C9_N_btm.n86 VSS 1.01985f
C7199 C9_N_btm.n87 VSS 1.01985f
C7200 C9_N_btm.n88 VSS 1.01985f
C7201 C9_N_btm.n89 VSS 1.01985f
C7202 C9_N_btm.n90 VSS 1.01629f
C7203 C9_N_btm.n91 VSS 1.01629f
C7204 C9_N_btm.n92 VSS 1.01985f
C7205 C9_N_btm.n93 VSS 1.01985f
C7206 C9_N_btm.n94 VSS 1.01985f
C7207 C9_N_btm.n95 VSS 1.01629f
C7208 C9_N_btm.n96 VSS 1.01629f
C7209 C9_N_btm.n97 VSS 1.01629f
C7210 C9_N_btm.n98 VSS 1.01629f
C7211 C9_N_btm.n99 VSS 1.01985f
C7212 C9_N_btm.n100 VSS 1.30559f
C7213 C9_N_btm.n101 VSS 1.01985f
C7214 C9_N_btm.n102 VSS 2.29472f
C7215 C9_N_btm.n103 VSS 4.45069f
C7216 C9_N_btm.n104 VSS 3.1571f
C7217 C9_N_btm.n105 VSS 1.01985f
C7218 C9_N_btm.n106 VSS 1.01985f
C7219 C9_N_btm.n107 VSS 1.01985f
C7220 C9_N_btm.n108 VSS 1.01985f
C7221 C9_N_btm.n109 VSS 1.01985f
C7222 C9_N_btm.n110 VSS 1.01985f
C7223 C9_N_btm.n111 VSS 1.01985f
C7224 C9_N_btm.n112 VSS 1.01985f
C7225 C9_N_btm.n113 VSS 1.01985f
C7226 C9_N_btm.n114 VSS 1.01985f
C7227 C9_N_btm.n115 VSS 1.01985f
C7228 C9_N_btm.n116 VSS 1.01985f
C7229 C9_N_btm.n117 VSS 1.01985f
C7230 C9_N_btm.n118 VSS 1.01985f
C7231 C9_N_btm.n119 VSS 1.01629f
C7232 C9_N_btm.n120 VSS 1.01629f
C7233 C9_N_btm.n121 VSS 1.01629f
C7234 C9_N_btm.n122 VSS 1.01629f
C7235 C9_N_btm.n123 VSS 1.01985f
C7236 C9_N_btm.n124 VSS 1.01985f
C7237 C9_N_btm.n125 VSS 1.01985f
C7238 C9_N_btm.n126 VSS 1.01985f
C7239 C9_N_btm.n127 VSS 1.01985f
C7240 C9_N_btm.n128 VSS 1.01985f
C7241 C9_N_btm.n129 VSS 1.01985f
C7242 C9_N_btm.n130 VSS 1.01985f
C7243 C9_N_btm.n131 VSS 1.01985f
C7244 C9_N_btm.n132 VSS 1.01985f
C7245 C9_N_btm.n133 VSS 1.01985f
C7246 C9_N_btm.n134 VSS 1.01985f
C7247 C9_N_btm.n135 VSS 1.01985f
C7248 C9_N_btm.n136 VSS 1.02004f
C7249 C9_N_btm.n137 VSS 1.02004f
C7250 C9_N_btm.n138 VSS 0.750397f
C7251 C9_N_btm.n139 VSS 0.750397f
C7252 C9_N_btm.n140 VSS 0.750397f
C7253 C9_N_btm.n141 VSS 1.02004f
C7254 C9_N_btm.n142 VSS 0.750397f
C7255 C9_N_btm.n143 VSS 1.02004f
C7256 C9_N_btm.n144 VSS 1.01985f
C7257 C9_N_btm.n145 VSS 1.01985f
C7258 C9_N_btm.n146 VSS 1.01985f
C7259 C9_N_btm.n147 VSS 1.01985f
C7260 C9_N_btm.n148 VSS 1.01985f
C7261 C9_N_btm.n149 VSS 1.01985f
C7262 C9_N_btm.n150 VSS 1.01985f
C7263 C9_N_btm.n151 VSS 1.01985f
C7264 C9_N_btm.n152 VSS 1.01985f
C7265 C9_N_btm.n153 VSS 1.28199f
C7266 C9_N_btm.n154 VSS 1.01985f
C7267 C9_N_btm.n155 VSS 1.01985f
C7268 C9_N_btm.n156 VSS 1.01985f
C7269 C9_N_btm.n157 VSS 1.01985f
C7270 C9_N_btm.n158 VSS 1.01985f
C7271 C9_N_btm.n159 VSS 1.01985f
C7272 C9_N_btm.n160 VSS 1.01985f
C7273 C9_N_btm.n161 VSS 1.01985f
C7274 C9_N_btm.n162 VSS 1.01985f
C7275 C9_N_btm.n163 VSS 1.02004f
C7276 C9_N_btm.n164 VSS 1.01985f
C7277 C9_N_btm.n165 VSS 1.02004f
C7278 C9_N_btm.n166 VSS 0.750397f
C7279 C9_N_btm.n167 VSS 1.02004f
C7280 C9_N_btm.n168 VSS 1.01985f
C7281 C9_N_btm.n169 VSS 1.01985f
C7282 C9_N_btm.n170 VSS 1.01985f
C7283 C9_N_btm.n171 VSS 1.01985f
C7284 C9_N_btm.n172 VSS 1.01985f
C7285 C9_N_btm.n173 VSS 1.01985f
C7286 C9_N_btm.n174 VSS 1.01985f
C7287 C9_N_btm.n175 VSS 1.01985f
C7288 C9_N_btm.n176 VSS 1.28199f
C7289 C9_N_btm.n177 VSS 1.28199f
C7290 C9_N_btm.n178 VSS 1.01985f
C7291 C9_N_btm.n179 VSS 1.01985f
C7292 C9_N_btm.n180 VSS 1.01985f
C7293 C9_N_btm.n181 VSS 1.01985f
C7294 C9_N_btm.n182 VSS 1.01985f
C7295 C9_N_btm.n183 VSS 1.01985f
C7296 C9_N_btm.n184 VSS 2.48581f
C7297 C9_N_btm.n185 VSS 0.984432f
C7298 C9_N_btm.n186 VSS 1.01985f
C7299 C9_N_btm.n187 VSS 1.01985f
C7300 C9_N_btm.n188 VSS 2.48581f
C7301 C9_N_btm.n189 VSS 1.01985f
C7302 C9_N_btm.n190 VSS 1.01985f
C7303 C9_N_btm.n191 VSS 1.01985f
C7304 C9_N_btm.n192 VSS 1.01985f
C7305 C9_N_btm.n193 VSS 1.01985f
C7306 C9_N_btm.n194 VSS 1.01985f
C7307 C9_N_btm.n195 VSS 1.01985f
C7308 C9_N_btm.n196 VSS 1.01985f
C7309 C9_N_btm.n197 VSS 1.02004f
C7310 C9_N_btm.n198 VSS 1.01985f
C7311 C9_N_btm.n199 VSS 1.02004f
C7312 C9_N_btm.n200 VSS 0.750397f
C7313 C9_N_btm.n201 VSS 1.01985f
C7314 C9_N_btm.n202 VSS 1.02004f
C7315 C9_N_btm.n203 VSS 1.01985f
C7316 C9_N_btm.n204 VSS 1.01985f
C7317 C9_N_btm.n205 VSS 1.01985f
C7318 C9_N_btm.n206 VSS 1.01985f
C7319 C9_N_btm.n207 VSS 1.01985f
C7320 C9_N_btm.n208 VSS 1.01985f
C7321 C9_N_btm.n209 VSS 1.01985f
C7322 C9_N_btm.n210 VSS 1.28199f
C7323 C9_N_btm.n211 VSS 1.01985f
C7324 C9_N_btm.n212 VSS 1.28199f
C7325 C9_N_btm.n213 VSS 1.28199f
C7326 C9_N_btm.n214 VSS 1.01985f
C7327 C9_N_btm.n215 VSS 1.01985f
C7328 C9_N_btm.n216 VSS 1.01985f
C7329 C9_N_btm.n217 VSS 1.01985f
C7330 C9_N_btm.n218 VSS 1.01985f
C7331 C9_N_btm.n219 VSS 1.01985f
C7332 C9_N_btm.n220 VSS 1.01985f
C7333 C9_N_btm.n221 VSS 1.01985f
C7334 C9_N_btm.n222 VSS 1.28199f
C7335 C9_N_btm.n223 VSS 1.28199f
C7336 C9_N_btm.n224 VSS 1.01985f
C7337 C9_N_btm.n225 VSS 1.01985f
C7338 C9_N_btm.n226 VSS 1.01985f
C7339 C9_N_btm.n227 VSS 1.01985f
C7340 C9_N_btm.n228 VSS 1.01985f
C7341 C9_N_btm.n229 VSS 1.01985f
C7342 C9_N_btm.n230 VSS 1.01985f
C7343 C9_N_btm.n231 VSS 1.01985f
C7344 C9_N_btm.n232 VSS 1.01985f
C7345 C9_N_btm.n233 VSS 1.01985f
C7346 C9_N_btm.n234 VSS 1.01985f
C7347 C9_N_btm.n235 VSS 1.02004f
C7348 C9_N_btm.n236 VSS 1.45446f
C7349 C9_N_btm.n237 VSS 1.02004f
C7350 C9_N_btm.n238 VSS 1.01985f
C7351 C9_N_btm.n239 VSS 1.01985f
C7352 C9_N_btm.n240 VSS 1.01985f
C7353 C9_N_btm.n241 VSS 1.01985f
C7354 C9_N_btm.n242 VSS 1.01985f
C7355 C9_N_btm.n243 VSS 1.01985f
C7356 C9_N_btm.n244 VSS 1.01985f
C7357 C9_N_btm.n245 VSS 1.01985f
C7358 C9_N_btm.n246 VSS 1.01985f
C7359 C9_N_btm.n247 VSS 1.01985f
C7360 C9_N_btm.n248 VSS 1.01985f
C7361 C9_N_btm.n249 VSS 1.01985f
C7362 C9_N_btm.n250 VSS 1.01985f
C7363 C9_N_btm.n251 VSS 1.01985f
C7364 C9_N_btm.n252 VSS 1.01985f
C7365 C9_N_btm.n253 VSS 1.01985f
C7366 C9_N_btm.n254 VSS 1.01985f
C7367 C9_N_btm.n255 VSS 1.01985f
C7368 C9_N_btm.n256 VSS 1.01985f
C7369 C9_N_btm.n257 VSS 1.01985f
C7370 C9_N_btm.n258 VSS 1.01985f
C7371 C9_N_btm.n259 VSS 1.01985f
C7372 C9_N_btm.n260 VSS 1.01985f
C7373 C9_N_btm.n261 VSS 1.01985f
C7374 C9_N_btm.n262 VSS 1.01985f
C7375 C9_N_btm.n263 VSS 1.01985f
C7376 C9_N_btm.n264 VSS 1.01985f
C7377 C9_N_btm.n265 VSS 1.01985f
C7378 C9_N_btm.n266 VSS 1.01985f
C7379 C9_N_btm.n267 VSS 1.01985f
C7380 C9_N_btm.n268 VSS 1.01985f
C7381 C9_N_btm.n269 VSS 1.01985f
C7382 C9_N_btm.n270 VSS 1.01985f
C7383 C9_N_btm.n271 VSS 1.01985f
C7384 C9_N_btm.n272 VSS 1.01985f
C7385 C9_N_btm.n273 VSS 1.01985f
C7386 C9_N_btm.n274 VSS 1.01985f
C7387 C9_N_btm.n275 VSS 1.01985f
C7388 C9_N_btm.n276 VSS 1.01985f
C7389 C9_N_btm.n277 VSS 1.01985f
C7390 C9_N_btm.n278 VSS 1.01985f
C7391 C9_N_btm.n279 VSS 1.01985f
C7392 C9_N_btm.n280 VSS 1.0161f
C7393 C9_N_btm.n281 VSS 1.01629f
C7394 C9_N_btm.n282 VSS 1.01629f
C7395 C9_N_btm.n283 VSS 1.01985f
C7396 C9_N_btm.n284 VSS 1.01985f
C7397 C9_N_btm.n285 VSS 1.01629f
C7398 C9_N_btm.n286 VSS 1.01629f
C7399 C9_N_btm.n287 VSS 1.01629f
C7400 C9_N_btm.n288 VSS 1.01629f
C7401 C9_N_btm.n289 VSS 1.01629f
C7402 C9_N_btm.n290 VSS 1.01629f
C7403 C9_N_btm.n291 VSS 1.01985f
C7404 C9_N_btm.n292 VSS 1.01985f
C7405 C9_N_btm.n293 VSS 1.01629f
C7406 C9_N_btm.n294 VSS 1.01629f
C7407 C9_N_btm.n295 VSS 1.01629f
C7408 C9_N_btm.n296 VSS 1.01629f
C7409 C9_N_btm.n297 VSS 1.01629f
C7410 C9_N_btm.n298 VSS 1.30559f
C7411 C9_N_btm.n299 VSS 1.01985f
C7412 C9_N_btm.n300 VSS 1.01985f
C7413 C9_N_btm.n301 VSS 3.1571f
C7414 C9_N_btm.n302 VSS 4.45069f
C7415 C9_N_btm.n303 VSS 1.02004f
C7416 C9_N_btm.n304 VSS 1.59759f
C7417 C9_N_btm.n305 VSS 1.22835f
C7418 C9_N_btm.n306 VSS 1.01629f
C7419 C9_N_btm.n307 VSS 1.01629f
C7420 C9_N_btm.n308 VSS 1.01629f
C7421 C9_N_btm.n309 VSS 1.01629f
C7422 C9_N_btm.n310 VSS 1.01985f
C7423 C9_N_btm.n311 VSS 1.01985f
C7424 C9_N_btm.n312 VSS 1.01629f
C7425 C9_N_btm.n313 VSS 1.01629f
C7426 C9_N_btm.n314 VSS 1.01629f
C7427 C9_N_btm.n315 VSS 1.01629f
C7428 C9_N_btm.n316 VSS 1.01629f
C7429 C9_N_btm.n317 VSS 1.01629f
C7430 C9_N_btm.n318 VSS 1.01985f
C7431 C9_N_btm.n319 VSS 1.01985f
C7432 C9_N_btm.n320 VSS 1.01629f
C7433 C9_N_btm.n321 VSS 1.01629f
C7434 C9_N_btm.n322 VSS 1.01629f
C7435 C9_N_btm.n323 VSS 1.01629f
C7436 C9_N_btm.n324 VSS 1.01629f
C7437 C9_N_btm.n325 VSS 1.01629f
C7438 C9_N_btm.n326 VSS 1.01985f
C7439 C9_N_btm.n327 VSS 1.01985f
C7440 C9_N_btm.n328 VSS 1.01629f
C7441 C9_N_btm.n329 VSS 1.01629f
C7442 C9_N_btm.n330 VSS 1.30558f
C7443 C9_N_btm.n331 VSS 3.157f
C7444 C9_N_btm.n332 VSS 4.45062f
C7445 C9_N_btm.n333 VSS 1.01985f
C7446 C9_N_btm.n334 VSS 1.01985f
C7447 C9_N_btm.n335 VSS 1.01985f
C7448 C9_N_btm.n336 VSS 1.01985f
C7449 C9_N_btm.n337 VSS 1.01985f
C7450 C9_N_btm.n338 VSS 1.01985f
C7451 C9_N_btm.n339 VSS 1.01985f
C7452 C9_N_btm.n340 VSS 1.01985f
C7453 C9_N_btm.n341 VSS 1.01985f
C7454 C9_N_btm.n342 VSS 1.01985f
C7455 C9_N_btm.n343 VSS 1.01985f
C7456 C9_N_btm.n344 VSS 1.01985f
C7457 C9_N_btm.n345 VSS 1.01985f
C7458 C9_N_btm.n346 VSS 1.01985f
C7459 C9_N_btm.n347 VSS 1.01985f
C7460 C9_N_btm.n348 VSS 1.01985f
C7461 C9_N_btm.n349 VSS 1.01985f
C7462 C9_N_btm.n350 VSS 1.01985f
C7463 C9_N_btm.n351 VSS 1.01985f
C7464 C9_N_btm.n352 VSS 1.01985f
C7465 C9_N_btm.n353 VSS 1.01985f
C7466 C9_N_btm.n354 VSS 1.01985f
C7467 C9_N_btm.n355 VSS 1.01985f
C7468 C9_N_btm.n356 VSS 1.01985f
C7469 C9_N_btm.n357 VSS 1.01985f
C7470 C9_N_btm.n358 VSS 1.01985f
C7471 C9_N_btm.n359 VSS 1.01985f
C7472 C9_N_btm.n360 VSS 1.01985f
C7473 C9_N_btm.n361 VSS 1.02004f
C7474 C9_N_btm.n362 VSS 0.750397f
C7475 C9_N_btm.n363 VSS 0.750397f
C7476 C9_N_btm.n364 VSS 0.750397f
C7477 C9_N_btm.n365 VSS 1.02004f
C7478 C9_N_btm.n366 VSS 1.02004f
C7479 C9_N_btm.n367 VSS 0.750397f
C7480 C9_N_btm.n368 VSS 0.750397f
C7481 C9_N_btm.n369 VSS 1.01985f
C7482 C9_N_btm.n370 VSS 1.01985f
C7483 C9_N_btm.n371 VSS 1.01985f
C7484 C9_N_btm.n372 VSS 1.01985f
C7485 C9_N_btm.n373 VSS 1.01985f
C7486 C9_N_btm.n374 VSS 1.01985f
C7487 C9_N_btm.n375 VSS 1.01985f
C7488 C9_N_btm.n376 VSS 1.01985f
C7489 C9_N_btm.n377 VSS 1.02004f
C7490 C9_N_btm.n378 VSS 1.02004f
C7491 C9_N_btm.n379 VSS 0.750397f
C7492 C9_N_btm.n380 VSS 0.750397f
C7493 C9_N_btm.n381 VSS 0.750397f
C7494 C9_N_btm.n382 VSS 0.750397f
C7495 C9_N_btm.n383 VSS 1.02004f
C7496 C9_N_btm.n384 VSS 1.02004f
C7497 C9_N_btm.n385 VSS 1.01985f
C7498 C9_N_btm.n386 VSS 1.01985f
C7499 C9_N_btm.n387 VSS 1.01985f
C7500 C9_N_btm.n388 VSS 1.01985f
C7501 C9_N_btm.n389 VSS 1.01985f
C7502 C9_N_btm.n390 VSS 1.28199f
C7503 C9_N_btm.n391 VSS 1.28199f
C7504 C9_N_btm.n392 VSS 1.28199f
C7505 C9_N_btm.n393 VSS 1.28199f
C7506 C9_N_btm.n394 VSS 1.28199f
C7507 C9_N_btm.n395 VSS 1.28199f
C7508 C9_N_btm.n396 VSS 1.01985f
C7509 C9_N_btm.n397 VSS 1.01985f
C7510 C9_N_btm.n398 VSS 1.01985f
C7511 C9_N_btm.n399 VSS 1.01985f
C7512 C9_N_btm.n400 VSS 1.01985f
C7513 C9_N_btm.n401 VSS 1.02004f
C7514 C9_N_btm.n402 VSS 1.01985f
C7515 C9_N_btm.n403 VSS 1.23745f
C7516 C9_N_btm.n404 VSS 0.575754f
C7517 C9_N_btm.n405 VSS 1.02004f
C7518 C9_N_btm.n406 VSS 0.750397f
C7519 C9_N_btm.n407 VSS 1.01985f
C7520 C9_N_btm.n408 VSS 1.02004f
C7521 C9_N_btm.n409 VSS 0.750397f
C7522 C9_N_btm.n410 VSS 0.750397f
C7523 C9_N_btm.n411 VSS 1.02004f
C7524 C9_N_btm.n412 VSS 1.01985f
C7525 C9_N_btm.n413 VSS 1.01985f
C7526 C9_N_btm.n414 VSS 1.01985f
C7527 C9_N_btm.n415 VSS 1.01985f
C7528 C9_N_btm.n416 VSS 1.01985f
C7529 C9_N_btm.n417 VSS 1.01985f
C7530 C9_N_btm.n418 VSS 1.01985f
C7531 C9_N_btm.n419 VSS 1.02004f
C7532 C9_N_btm.n420 VSS 1.02004f
C7533 C9_N_btm.n421 VSS 0.750397f
C7534 C9_N_btm.n422 VSS 0.750397f
C7535 C9_N_btm.n423 VSS 0.750397f
C7536 C9_N_btm.n424 VSS 1.45446f
C7537 C9_N_btm.n425 VSS 1.02004f
C7538 C9_N_btm.n426 VSS 1.01985f
C7539 C9_N_btm.n427 VSS 1.01985f
C7540 C9_N_btm.n428 VSS 1.01985f
C7541 C9_N_btm.n429 VSS 1.01985f
C7542 C9_N_btm.n430 VSS 1.01985f
C7543 C9_N_btm.n431 VSS 1.01985f
C7544 C9_N_btm.n432 VSS 1.01985f
C7545 C9_N_btm.n433 VSS 1.01985f
C7546 C9_N_btm.n434 VSS 0.984432f
C7547 C9_N_btm.n435 VSS 1.39202f
C7548 C9_N_btm.n436 VSS 1.28199f
C7549 C9_N_btm.n437 VSS 1.28199f
C7550 C9_N_btm.n438 VSS 1.39202f
C7551 C9_N_btm.n439 VSS 1.01985f
C7552 C9_N_btm.n440 VSS 1.01985f
C7553 C9_N_btm.n441 VSS 1.01985f
C7554 C9_N_btm.n442 VSS 1.01985f
C7555 C9_N_btm.n443 VSS 1.01985f
C7556 C9_N_btm.n444 VSS 1.02004f
C7557 C9_N_btm.n445 VSS 0.750397f
C7558 C9_N_btm.n446 VSS 0.750397f
C7559 C9_N_btm.n447 VSS 1.02004f
C7560 C9_N_btm.n448 VSS 1.02004f
C7561 C9_N_btm.n449 VSS 1.23727f
C7562 C9_N_btm.n450 VSS 0.575754f
C7563 C9_N_btm.n451 VSS 1.45446f
C7564 C9_N_btm.n452 VSS 0.750397f
C7565 C9_N_btm.n453 VSS 1.02004f
C7566 C9_N_btm.n454 VSS 1.01985f
C7567 C9_N_btm.n455 VSS 1.01985f
C7568 C9_N_btm.n456 VSS 1.01985f
C7569 C9_N_btm.n457 VSS 1.01985f
C7570 C9_N_btm.n458 VSS 1.01985f
C7571 C9_N_btm.n459 VSS 1.01985f
C7572 C9_N_btm.n460 VSS 1.01985f
C7573 C9_N_btm.n461 VSS 1.01985f
C7574 C9_N_btm.n462 VSS 1.28199f
C7575 C9_N_btm.n463 VSS 1.28199f
C7576 C9_N_btm.n464 VSS 1.28199f
C7577 C9_N_btm.n465 VSS 1.28199f
C7578 C9_N_btm.n466 VSS 1.01985f
C7579 C9_N_btm.n467 VSS 1.01985f
C7580 C9_N_btm.n468 VSS 1.01985f
C7581 C9_N_btm.n469 VSS 1.28199f
C7582 C9_N_btm.n470 VSS 1.28199f
C7583 C9_N_btm.n471 VSS 1.28199f
C7584 C9_N_btm.n472 VSS 1.01985f
C7585 C9_N_btm.n473 VSS 1.01985f
C7586 C9_N_btm.n474 VSS 1.01985f
C7587 C9_N_btm.n475 VSS 1.01985f
C7588 C9_N_btm.n476 VSS 1.01985f
C7589 C9_N_btm.n477 VSS 1.02004f
C7590 C9_N_btm.n478 VSS 0.750397f
C7591 C9_N_btm.n479 VSS 0.750397f
C7592 C9_N_btm.n480 VSS 0.750398f
C7593 C9_N_btm.n481 VSS 1.02004f
C7594 C9_N_btm.n482 VSS 1.02004f
C7595 C9_N_btm.n483 VSS 1.01985f
C7596 C9_N_btm.n484 VSS 1.01985f
C7597 C9_N_btm.n485 VSS 1.01985f
C7598 C9_N_btm.n486 VSS 1.01985f
C7599 C9_N_btm.n487 VSS 1.01985f
C7600 C9_N_btm.n488 VSS 1.01985f
C7601 C9_N_btm.n489 VSS 1.01985f
C7602 C9_N_btm.n490 VSS 1.01985f
C7603 C9_N_btm.n491 VSS 1.01629f
C7604 C9_N_btm.n492 VSS 1.01985f
C7605 C9_N_btm.n493 VSS 1.01985f
C7606 C9_N_btm.n494 VSS 1.01985f
C7607 C9_N_btm.n495 VSS 1.01985f
C7608 C9_N_btm.n496 VSS 1.01629f
C7609 C9_N_btm.n497 VSS 1.01629f
C7610 C9_N_btm.n498 VSS 1.01629f
C7611 C9_N_btm.n499 VSS 1.01629f
C7612 C9_N_btm.n500 VSS 1.01985f
C7613 C9_N_btm.n501 VSS 1.01985f
C7614 C9_N_btm.n502 VSS 1.01985f
C7615 C9_N_btm.n503 VSS 1.01985f
C7616 C9_N_btm.n504 VSS 1.01629f
C7617 C9_N_btm.n505 VSS 1.01629f
C7618 C9_N_btm.n506 VSS 1.01629f
C7619 C9_N_btm.n507 VSS 1.01629f
C7620 C9_N_btm.n508 VSS 1.01985f
C7621 C9_N_btm.n509 VSS 1.01985f
C7622 C9_N_btm.n510 VSS 1.01985f
C7623 C9_N_btm.n511 VSS 1.01985f
C7624 C9_N_btm.n512 VSS 1.01629f
C7625 C9_N_btm.n513 VSS 2.2847f
C7626 a_21588_30879.t0 VSS 0.024382f
C7627 a_21588_30879.t6 VSS 0.825305f
C7628 a_21588_30879.t8 VSS 0.825432f
C7629 a_21588_30879.t4 VSS 0.825304f
C7630 a_21588_30879.n0 VSS 0.612275f
C7631 a_21588_30879.t11 VSS 0.825304f
C7632 a_21588_30879.n1 VSS 0.310265f
C7633 a_21588_30879.t7 VSS 0.825304f
C7634 a_21588_30879.n2 VSS 0.310265f
C7635 a_21588_30879.t9 VSS 0.825304f
C7636 a_21588_30879.n3 VSS 0.310265f
C7637 a_21588_30879.t10 VSS 0.825304f
C7638 a_21588_30879.n4 VSS 0.310265f
C7639 a_21588_30879.t5 VSS 0.825304f
C7640 a_21588_30879.n5 VSS 0.309233f
C7641 a_21588_30879.n6 VSS 3.61172f
C7642 a_21588_30879.t3 VSS 0.015848f
C7643 a_21588_30879.t2 VSS 0.015848f
C7644 a_21588_30879.n7 VSS 0.031697f
C7645 a_21588_30879.n8 VSS 3.13783f
C7646 a_21588_30879.n9 VSS 0.073162f
C7647 a_21588_30879.t1 VSS 0.024382f
C7648 a_n2293_42834.t2 VSS 0.014014f
C7649 a_n2293_42834.t1 VSS 0.029912f
C7650 a_n2293_42834.t4 VSS 0.012597f
C7651 a_n2293_42834.t3 VSS 0.01974f
C7652 a_n2293_42834.n0 VSS 0.604238f
C7653 a_n2293_42834.n1 VSS 3.36003f
C7654 a_n2293_42834.n2 VSS 0.045452f
C7655 a_n2293_42834.t0 VSS 0.014014f
C7656 C6_N_btm.t1 VSS 1.67804f
C7657 C6_N_btm.t3 VSS 0.051941f
C7658 C6_N_btm.t2 VSS 0.051941f
C7659 C6_N_btm.n0 VSS 0.247039f
C7660 C6_N_btm.t5 VSS 0.051941f
C7661 C6_N_btm.t4 VSS 0.051941f
C7662 C6_N_btm.n1 VSS 0.138138f
C7663 C6_N_btm.n2 VSS 1.35068f
C7664 C6_N_btm.n3 VSS 2.10571f
C7665 C6_N_btm.t0 VSS 0.120999f
C7666 C6_N_btm.n4 VSS 2.99373f
C7667 a_20692_30879.t4 VSS 3.0248f
C7668 a_20692_30879.t3 VSS 0.037079f
C7669 a_20692_30879.t2 VSS 0.037079f
C7670 a_20692_30879.n0 VSS 0.074157f
C7671 a_20692_30879.n1 VSS 14.541599f
C7672 a_20692_30879.t0 VSS 0.057044f
C7673 a_20692_30879.n2 VSS 0.171171f
C7674 a_20692_30879.t1 VSS 0.057044f
C7675 C4_N_btm.t3 VSS 1.26438f
C7676 C4_N_btm.t2 VSS 0.389904f
C7677 C4_N_btm.t1 VSS 0.261549f
C7678 C4_N_btm.n0 VSS 2.01038f
C7679 C4_N_btm.n1 VSS 3.13259f
C7680 C4_N_btm.t0 VSS 0.171423f
C7681 C4_N_btm.n2 VSS 3.85704f
C7682 a_14097_32519.t0 VSS 0.065966f
C7683 a_14097_32519.t4 VSS 2.34954f
C7684 a_14097_32519.t3 VSS 0.042878f
C7685 a_14097_32519.t2 VSS 0.042878f
C7686 a_14097_32519.n0 VSS 0.085756f
C7687 a_14097_32519.n1 VSS 18.5491f
C7688 a_14097_32519.n2 VSS 0.197942f
C7689 a_14097_32519.t1 VSS 0.065966f
C7690 a_n2956_38680.t0 VSS 0.056669f
C7691 a_n2956_38680.t2 VSS 0.036835f
C7692 a_n2956_38680.t3 VSS 0.036835f
C7693 a_n2956_38680.n0 VSS 0.128088f
C7694 a_n2956_38680.t4 VSS 0.093572f
C7695 a_n2956_38680.t5 VSS 0.058372f
C7696 a_n2956_38680.n1 VSS 2.33493f
C7697 a_n2956_38680.n2 VSS 9.08207f
C7698 a_n2956_38680.n3 VSS 0.115959f
C7699 a_n2956_38680.t1 VSS 0.056669f
C7700 a_n4209_39304.t1 VSS 0.036477f
C7701 a_n4209_39304.t6 VSS 0.02371f
C7702 a_n4209_39304.t7 VSS 0.02371f
C7703 a_n4209_39304.n0 VSS 0.090526f
C7704 a_n4209_39304.t5 VSS 0.02371f
C7705 a_n4209_39304.t4 VSS 0.02371f
C7706 a_n4209_39304.n1 VSS 0.05381f
C7707 a_n4209_39304.n2 VSS 0.291258f
C7708 a_n4209_39304.t9 VSS 0.038601f
C7709 a_n4209_39304.t10 VSS 0.061472f
C7710 a_n4209_39304.n3 VSS 0.1308f
C7711 a_n4209_39304.t11 VSS 1.23487f
C7712 a_n4209_39304.t8 VSS 1.23471f
C7713 a_n4209_39304.n4 VSS 4.17954f
C7714 a_n4209_39304.n5 VSS 4.12475f
C7715 a_n4209_39304.n6 VSS 0.148307f
C7716 a_n4209_39304.t2 VSS 0.036477f
C7717 a_n4209_39304.t0 VSS 0.036477f
C7718 a_n4209_39304.n7 VSS 0.075037f
C7719 a_n4209_39304.n8 VSS 0.302739f
C7720 a_n4209_39304.n9 VSS 0.092834f
C7721 a_n4209_39304.t3 VSS 0.036477f
C7722 a_768_44030.t1 VSS 0.010205f
C7723 a_768_44030.t0 VSS 0.010205f
C7724 a_768_44030.t2 VSS 0.010205f
C7725 a_768_44030.n0 VSS 0.03041f
C7726 a_768_44030.n1 VSS 0.019124f
C7727 a_768_44030.n2 VSS 0.015105f
C7728 a_768_44030.n3 VSS 0.086126f
C7729 a_768_44030.n4 VSS 0.078f
C7730 a_768_44030.t8 VSS 0.017198f
C7731 a_768_44030.t22 VSS 0.010799f
C7732 a_768_44030.n5 VSS 0.025728f
C7733 a_768_44030.n6 VSS 0.027156f
C7734 a_768_44030.n7 VSS 0.033472f
C7735 a_768_44030.n8 VSS 0.550196f
C7736 a_768_44030.t23 VSS 0.015875f
C7737 a_768_44030.t13 VSS 0.015875f
C7738 a_768_44030.n9 VSS 0.026635f
C7739 a_768_44030.n10 VSS 0.052106f
C7740 a_768_44030.n11 VSS 0.606757f
C7741 a_768_44030.t25 VSS 0.010799f
C7742 a_768_44030.t14 VSS 0.017198f
C7743 a_768_44030.n12 VSS 0.028066f
C7744 a_768_44030.n13 VSS 0.217952f
C7745 a_768_44030.n14 VSS 0.024903f
C7746 a_768_44030.n15 VSS 0.810065f
C7747 a_768_44030.t18 VSS 0.010799f
C7748 a_768_44030.t16 VSS 0.017198f
C7749 a_768_44030.n16 VSS 0.027124f
C7750 a_768_44030.n17 VSS 1.25227f
C7751 a_768_44030.n18 VSS 0.340801f
C7752 a_768_44030.t19 VSS 0.017198f
C7753 a_768_44030.t9 VSS 0.010799f
C7754 a_768_44030.n19 VSS 0.025596f
C7755 a_768_44030.n20 VSS 0.356559f
C7756 a_768_44030.n21 VSS 0.065592f
C7757 a_768_44030.n22 VSS 0.020472f
C7758 a_768_44030.t3 VSS 0.010205f
C7759 a_n4209_37414.t1 VSS 0.048411f
C7760 a_n4209_37414.t4 VSS 0.031467f
C7761 a_n4209_37414.t6 VSS 0.031467f
C7762 a_n4209_37414.n0 VSS 0.120144f
C7763 a_n4209_37414.t5 VSS 0.031467f
C7764 a_n4209_37414.t7 VSS 0.031467f
C7765 a_n4209_37414.n1 VSS 0.071416f
C7766 a_n4209_37414.n2 VSS 0.351271f
C7767 a_n4209_37414.t8 VSS 0.081584f
C7768 a_n4209_37414.t10 VSS 0.05123f
C7769 a_n4209_37414.n3 VSS 0.171345f
C7770 a_n4209_37414.t9 VSS 1.46067f
C7771 a_n4209_37414.n4 VSS 9.31613f
C7772 a_n4209_37414.n5 VSS 0.199599f
C7773 a_n4209_37414.t2 VSS 0.048411f
C7774 a_n4209_37414.t0 VSS 0.048411f
C7775 a_n4209_37414.n6 VSS 0.123208f
C7776 a_n4209_37414.n7 VSS 0.434301f
C7777 a_n4209_37414.n8 VSS 0.099587f
C7778 a_n4209_37414.t3 VSS 0.048411f
C7779 a_20820_30879.t5 VSS 1.61926f
C7780 a_20820_30879.t4 VSS 1.61947f
C7781 a_20820_30879.n0 VSS 7.88484f
C7782 a_20820_30879.t3 VSS 0.031094f
C7783 a_20820_30879.t2 VSS 0.031094f
C7784 a_20820_30879.n1 VSS 0.062189f
C7785 a_20820_30879.n2 VSS 6.21284f
C7786 a_20820_30879.t0 VSS 0.047838f
C7787 a_20820_30879.n3 VSS 0.143545f
C7788 a_20820_30879.t1 VSS 0.047838f
C7789 a_4915_47217.t11 VSS 0.012274f
C7790 a_4915_47217.t4 VSS 0.033738f
C7791 a_4915_47217.n0 VSS 0.171274f
C7792 a_4915_47217.t7 VSS 0.012567f
C7793 a_4915_47217.t2 VSS 0.018288f
C7794 a_4915_47217.n1 VSS 0.062818f
C7795 a_4915_47217.n2 VSS 1.37164f
C7796 a_4915_47217.t3 VSS 0.015286f
C7797 a_4915_47217.t5 VSS 0.02594f
C7798 a_4915_47217.t8 VSS 0.015286f
C7799 a_4915_47217.t6 VSS 0.02594f
C7800 a_4915_47217.n3 VSS 0.043524f
C7801 a_4915_47217.n4 VSS 0.065599f
C7802 a_4915_47217.n5 VSS 0.414469f
C7803 a_4915_47217.t10 VSS 0.027605f
C7804 a_4915_47217.t9 VSS 0.017236f
C7805 a_4915_47217.n6 VSS 0.100243f
C7806 a_4915_47217.n7 VSS 0.73963f
C7807 a_4915_47217.n8 VSS 0.024126f
C7808 a_4915_47217.t1 VSS 0.052375f
C7809 a_4915_47217.n9 VSS 0.09553f
C7810 a_4915_47217.t0 VSS 0.054615f
C7811 a_17517_44484.t1 VSS 0.120389f
C7812 a_17517_44484.t2 VSS 0.054492f
C7813 a_17517_44484.t3 VSS 0.034773f
C7814 a_17517_44484.n0 VSS 0.380383f
C7815 a_17517_44484.n1 VSS 2.26754f
C7816 a_17517_44484.t0 VSS 0.142418f
C7817 a_765_45546.t0 VSS 0.026757f
C7818 a_765_45546.t2 VSS 0.021248f
C7819 a_765_45546.t3 VSS 0.021248f
C7820 a_765_45546.n0 VSS 0.042608f
C7821 a_765_45546.t6 VSS 0.035808f
C7822 a_765_45546.t11 VSS 0.022485f
C7823 a_765_45546.n1 VSS 0.067065f
C7824 a_765_45546.t7 VSS 0.022485f
C7825 a_765_45546.t8 VSS 0.035808f
C7826 a_765_45546.n2 VSS 0.053245f
C7827 a_765_45546.n3 VSS 4.06584f
C7828 a_765_45546.t10 VSS 0.022485f
C7829 a_765_45546.t9 VSS 0.035808f
C7830 a_765_45546.n4 VSS 0.062716f
C7831 a_765_45546.n5 VSS 4.61854f
C7832 a_765_45546.t4 VSS 0.054982f
C7833 a_765_45546.t5 VSS 0.041499f
C7834 a_765_45546.n6 VSS 0.146724f
C7835 a_765_45546.n7 VSS 0.102399f
C7836 a_765_45546.n8 VSS 0.123476f
C7837 a_765_45546.n9 VSS 0.055519f
C7838 a_765_45546.t1 VSS 0.021248f
C7839 a_n3565_38216.t4 VSS 0.031524f
C7840 a_n3565_38216.t7 VSS 0.031524f
C7841 a_n3565_38216.n0 VSS 0.120358f
C7842 a_n3565_38216.t5 VSS 0.031524f
C7843 a_n3565_38216.t6 VSS 0.031524f
C7844 a_n3565_38216.n1 VSS 0.071544f
C7845 a_n3565_38216.n2 VSS 0.346162f
C7846 a_n3565_38216.t9 VSS 0.051322f
C7847 a_n3565_38216.t8 VSS 0.08173f
C7848 a_n3565_38216.n3 VSS 0.1309f
C7849 a_n3565_38216.t10 VSS 1.52735f
C7850 a_n3565_38216.n4 VSS 9.186629f
C7851 a_n3565_38216.n5 VSS 0.199965f
C7852 a_n3565_38216.t2 VSS 0.048498f
C7853 a_n3565_38216.t0 VSS 0.048498f
C7854 a_n3565_38216.n6 VSS 0.099765f
C7855 a_n3565_38216.n7 VSS 0.440761f
C7856 a_n3565_38216.t1 VSS 0.048498f
C7857 a_n3565_38216.n8 VSS 0.123428f
C7858 a_n3565_38216.t3 VSS 0.048498f
C7859 a_12741_44636.t2 VSS 0.036748f
C7860 a_12741_44636.t4 VSS 0.011477f
C7861 a_12741_44636.n0 VSS 0.100961f
C7862 a_12741_44636.t3 VSS 0.013488f
C7863 a_12741_44636.n1 VSS 0.050629f
C7864 a_12741_44636.n2 VSS 1.8523f
C7865 a_12741_44636.n3 VSS 0.085454f
C7866 a_12741_44636.n4 VSS 0.016904f
C7867 a_1423_45028.t0 VSS 0.028842f
C7868 a_1423_45028.t3 VSS 0.018747f
C7869 a_1423_45028.t2 VSS 0.018747f
C7870 a_1423_45028.n0 VSS 0.090336f
C7871 a_1423_45028.t7 VSS 0.038158f
C7872 a_1423_45028.t5 VSS 0.025843f
C7873 a_1423_45028.n1 VSS 0.352783f
C7874 a_1423_45028.t4 VSS 0.048391f
C7875 a_1423_45028.t6 VSS 0.026432f
C7876 a_1423_45028.n2 VSS 0.089285f
C7877 a_1423_45028.n3 VSS 2.94577f
C7878 a_1423_45028.n4 VSS 0.329914f
C7879 a_1423_45028.n5 VSS 0.057913f
C7880 a_1423_45028.t1 VSS 0.028842f
C7881 a_18194_34908.n0 VSS 0.022699f
C7882 a_18194_34908.n1 VSS 0.016243f
C7883 a_18194_34908.n2 VSS 0.088729f
C7884 a_18194_34908.t15 VSS 0.073797f
C7885 a_18194_34908.t11 VSS 0.077755f
C7886 a_18194_34908.n3 VSS 0.097484f
C7887 a_18194_34908.t13 VSS 0.073797f
C7888 a_18194_34908.t14 VSS 0.073797f
C7889 a_18194_34908.n4 VSS 0.055342f
C7890 a_18194_34908.n5 VSS 0.051459f
C7891 a_18194_34908.n6 VSS 0.240972f
C7892 a_18194_34908.t10 VSS 0.073546f
C7893 a_18194_34908.t12 VSS 0.077665f
C7894 a_18194_34908.n7 VSS 0.090055f
C7895 a_18194_34908.n8 VSS 0.378189f
C7896 a_18194_34908.t8 VSS 0.073546f
C7897 a_18194_34908.t9 VSS 0.077665f
C7898 a_18194_34908.n9 VSS 0.090055f
C7899 a_18194_34908.n10 VSS 0.243257f
C7900 a_18194_34908.n11 VSS 0.070983f
C7901 a_18194_34908.t1 VSS 0.011315f
C7902 a_18194_34908.t0 VSS 0.011315f
C7903 a_18194_34908.n12 VSS 0.034453f
C7904 a_18194_34908.n13 VSS 0.11877f
C7905 a_18194_34908.t2 VSS 0.011315f
C7906 a_18194_34908.n14 VSS 0.025065f
C7907 a_18194_34908.t3 VSS 0.011315f
C7908 C0_N_btm.t0 VSS 1.3641f
C7909 C0_N_btm.t2 VSS 0.406352f
C7910 C0_N_btm.t3 VSS 0.273912f
C7911 C0_N_btm.n0 VSS 2.20629f
C7912 C0_N_btm.n1 VSS 3.34443f
C7913 C0_N_btm.t1 VSS 0.195052f
C7914 C0_N_btm.n2 VSS 3.77254f
C7915 a_1606_42308.t3 VSS 0.035276f
C7916 a_1606_42308.t2 VSS 0.035276f
C7917 a_1606_42308.n0 VSS 0.130642f
C7918 a_1606_42308.t4 VSS 0.084422f
C7919 a_1606_42308.t6 VSS 0.052651f
C7920 a_1606_42308.n1 VSS 0.183637f
C7921 a_1606_42308.t7 VSS 0.351678f
C7922 a_1606_42308.t5 VSS 0.349599f
C7923 a_1606_42308.n2 VSS 16.647598f
C7924 a_1606_42308.n3 VSS 9.93149f
C7925 a_1606_42308.n4 VSS 0.480587f
C7926 a_1606_42308.t0 VSS 0.05427f
C7927 a_1606_42308.n5 VSS 0.108585f
C7928 a_1606_42308.t1 VSS 0.05427f
C7929 a_n743_46660.t1 VSS 0.038866f
C7930 a_n743_46660.t8 VSS 0.031818f
C7931 a_n743_46660.t2 VSS 0.011575f
C7932 a_n743_46660.n0 VSS 0.061379f
C7933 a_n743_46660.t11 VSS 0.016255f
C7934 a_n743_46660.t9 VSS 0.026034f
C7935 a_n743_46660.n1 VSS 0.056914f
C7936 a_n743_46660.n2 VSS 1.13789f
C7937 a_n743_46660.t5 VSS 0.045933f
C7938 a_n743_46660.t7 VSS 0.024182f
C7939 a_n743_46660.n3 VSS 0.154076f
C7940 a_n743_46660.n4 VSS 3.74127f
C7941 a_n743_46660.t3 VSS 0.031818f
C7942 a_n743_46660.t10 VSS 0.011575f
C7943 a_n743_46660.n5 VSS 0.07926f
C7944 a_n743_46660.t6 VSS 0.011575f
C7945 a_n743_46660.t4 VSS 0.031818f
C7946 a_n743_46660.n6 VSS 0.058074f
C7947 a_n743_46660.n7 VSS 0.538399f
C7948 a_n743_46660.n8 VSS 1.24634f
C7949 a_n743_46660.n9 VSS 0.325871f
C7950 a_n743_46660.t0 VSS 0.119075f
C7951 a_n2661_42834.t4 VSS 0.019831f
C7952 a_n2661_42834.t3 VSS 0.031077f
C7953 a_n2661_42834.n0 VSS 1.08426f
C7954 a_n2661_42834.t1 VSS 0.043545f
C7955 a_n2661_42834.n1 VSS 7.10303f
C7956 a_n2661_42834.t2 VSS 0.022062f
C7957 a_n2661_42834.n2 VSS 0.074138f
C7958 a_n2661_42834.t0 VSS 0.022062f
C7959 a_10809_44734.t1 VSS 0.021966f
C7960 a_10809_44734.t2 VSS 0.090351f
C7961 a_10809_44734.t6 VSS 0.019745f
C7962 a_10809_44734.t4 VSS 0.030942f
C7963 a_10809_44734.n0 VSS 0.746529f
C7964 a_10809_44734.t5 VSS 0.036362f
C7965 a_10809_44734.t3 VSS 0.022704f
C7966 a_10809_44734.n1 VSS 0.07098f
C7967 a_10809_44734.n2 VSS 5.92306f
C7968 a_10809_44734.n3 VSS 0.465697f
C7969 a_10809_44734.n4 VSS 0.049698f
C7970 a_10809_44734.t0 VSS 0.021966f
C7971 a_n3674_39768.t0 VSS 0.038961f
C7972 a_n3674_39768.t2 VSS 0.025325f
C7973 a_n3674_39768.t3 VSS 0.025325f
C7974 a_n3674_39768.n0 VSS 0.088064f
C7975 a_n3674_39768.t5 VSS 0.065088f
C7976 a_n3674_39768.t4 VSS 0.040763f
C7977 a_n3674_39768.n1 VSS 0.896286f
C7978 a_n3674_39768.n2 VSS 4.6015f
C7979 a_n3674_39768.n3 VSS 0.079725f
C7980 a_n3674_39768.t1 VSS 0.038961f
C7981 a_4791_45118.t0 VSS 0.011828f
C7982 a_4791_45118.n0 VSS 0.022208f
C7983 a_4791_45118.t21 VSS 0.010922f
C7984 a_4791_45118.t20 VSS 0.013522f
C7985 a_4791_45118.n1 VSS 0.0771f
C7986 a_4791_45118.t17 VSS 0.015837f
C7987 a_4791_45118.n2 VSS 0.029578f
C7988 a_4791_45118.n3 VSS 0.125163f
C7989 a_4791_45118.t13 VSS 0.010843f
C7990 a_4791_45118.t12 VSS 0.0184f
C7991 a_4791_45118.t23 VSS 0.010843f
C7992 a_4791_45118.t16 VSS 0.0184f
C7993 a_4791_45118.n4 VSS 0.030872f
C7994 a_4791_45118.n5 VSS 0.046558f
C7995 a_4791_45118.t14 VSS 0.0195f
C7996 a_4791_45118.t5 VSS 0.064581f
C7997 a_4791_45118.t22 VSS 0.010922f
C7998 a_4791_45118.t8 VSS 0.013522f
C7999 a_4791_45118.n6 VSS 0.0771f
C8000 a_4791_45118.t9 VSS 0.015837f
C8001 a_4791_45118.n7 VSS 0.029578f
C8002 a_4791_45118.n8 VSS 0.110676f
C8003 a_4791_45118.n9 VSS 0.662852f
C8004 a_4791_45118.n10 VSS 0.104858f
C8005 a_4791_45118.n11 VSS 0.269169f
C8006 a_4791_45118.n12 VSS 0.033804f
C8007 a_4791_45118.n13 VSS 0.293538f
C8008 a_4791_45118.t7 VSS 0.010734f
C8009 a_4791_45118.n14 VSS 0.028899f
C8010 a_4791_45118.t11 VSS 0.019699f
C8011 a_4791_45118.t15 VSS 0.012204f
C8012 a_4791_45118.n15 VSS 0.044442f
C8013 a_4791_45118.n16 VSS 0.366829f
C8014 a_4791_45118.n17 VSS 0.250733f
C8015 a_4791_45118.n18 VSS 0.130292f
C8016 a_4791_45118.n19 VSS 0.024526f
C8017 a_4791_45118.t1 VSS 0.011828f
C8018 a_n881_46662.t19 VSS 0.011174f
C8019 a_n881_46662.n1 VSS 0.024996f
C8020 a_n881_46662.n2 VSS 0.018098f
C8021 a_n881_46662.n3 VSS 0.019454f
C8022 a_n881_46662.n4 VSS 0.018098f
C8023 a_n881_46662.n5 VSS 0.020208f
C8024 a_n881_46662.n6 VSS 0.022278f
C8025 a_n881_46662.n7 VSS 0.509844f
C8026 a_n881_46662.t21 VSS 0.011208f
C8027 a_n881_46662.n8 VSS 0.016873f
C8028 a_n881_46662.n9 VSS 0.141885f
C8029 a_n881_46662.n10 VSS 0.196598f
C8030 a_n881_46662.n11 VSS 0.018098f
C8031 a_n881_46662.n12 VSS 0.195897f
C8032 a_n881_46662.n13 VSS 0.230733f
C8033 a_n881_46662.n14 VSS 0.018098f
C8034 a_n881_46662.n15 VSS 0.188146f
C8035 a_n881_46662.n16 VSS 0.018098f
C8036 a_n881_46662.n17 VSS 0.118203f
C8037 a_n881_46662.n18 VSS 0.287638f
C8038 a_n881_46662.n19 VSS 0.389663f
C8039 a_n881_46662.n20 VSS 0.068829f
C8040 a_n881_46662.n21 VSS 0.015826f
C8041 a_13887_32519.t0 VSS 0.061798f
C8042 a_13887_32519.t4 VSS 2.31163f
C8043 a_13887_32519.t2 VSS 0.040168f
C8044 a_13887_32519.t3 VSS 0.040168f
C8045 a_13887_32519.n0 VSS 0.080337f
C8046 a_13887_32519.n1 VSS 18.618698f
C8047 a_13887_32519.n2 VSS 0.185435f
C8048 a_13887_32519.t1 VSS 0.061798f
C8049 a_n4209_38502.t0 VSS 0.046968f
C8050 a_n4209_38502.t7 VSS 0.030529f
C8051 a_n4209_38502.t4 VSS 0.030529f
C8052 a_n4209_38502.n0 VSS 0.116562f
C8053 a_n4209_38502.t6 VSS 0.030529f
C8054 a_n4209_38502.t5 VSS 0.030529f
C8055 a_n4209_38502.n1 VSS 0.069287f
C8056 a_n4209_38502.n2 VSS 0.340799f
C8057 a_n4209_38502.t8 VSS 0.079152f
C8058 a_n4209_38502.t10 VSS 0.049703f
C8059 a_n4209_38502.n3 VSS 0.166236f
C8060 a_n4209_38502.t9 VSS 1.43874f
C8061 a_n4209_38502.n4 VSS 9.19838f
C8062 a_n4209_38502.n5 VSS 0.193648f
C8063 a_n4209_38502.t2 VSS 0.046968f
C8064 a_n4209_38502.t1 VSS 0.046968f
C8065 a_n4209_38502.n6 VSS 0.119534f
C8066 a_n4209_38502.n7 VSS 0.421353f
C8067 a_n4209_38502.n8 VSS 0.096618f
C8068 a_n4209_38502.t3 VSS 0.046968f
C8069 a_10341_43396.t1 VSS 0.033148f
C8070 a_10341_43396.t3 VSS 0.020588f
C8071 a_10341_43396.t2 VSS 0.013138f
C8072 a_10341_43396.n0 VSS 0.515287f
C8073 a_10341_43396.n1 VSS 3.74385f
C8074 a_10341_43396.t0 VSS 0.073987f
C8075 w_1575_34786.t3 VSS 0.024713f
C8076 w_1575_34786.n0 VSS 0.073491f
C8077 w_1575_34786.t1 VSS 0.08531f
C8078 w_1575_34786.n1 VSS 0.087589f
C8079 w_1575_34786.n2 VSS 0.156337f
C8080 w_1575_34786.n3 VSS 0.037194f
C8081 w_1575_34786.n4 VSS 0.026879f
C8082 w_1575_34786.n5 VSS 0.037646f
C8083 w_1575_34786.n6 VSS 0.055814f
C8084 w_1575_34786.n7 VSS 0.087338f
C8085 w_1575_34786.n8 VSS 0.028141f
C8086 w_1575_34786.t10 VSS 6.64883f
C8087 w_1575_34786.n9 VSS 0.035169f
C8088 w_1575_34786.n10 VSS 0.283024f
C8089 w_1575_34786.n11 VSS 0.035169f
C8090 w_1575_34786.n12 VSS 0.200676f
C8091 w_1575_34786.n13 VSS 0.657254f
C8092 w_1575_34786.n14 VSS 0.193395f
C8093 w_1575_34786.n15 VSS 0.032088f
C8094 w_1575_34786.n16 VSS 0.019274f
C8095 w_1575_34786.t9 VSS 0.019948f
C8096 w_1575_34786.n17 VSS 0.021382f
C8097 w_1575_34786.n18 VSS 0.024177f
C8098 w_1575_34786.n19 VSS 0.034106f
C8099 w_1575_34786.n20 VSS 0.063213f
C8100 w_1575_34786.t17 VSS 0.067657f
C8101 w_1575_34786.n21 VSS 1.42949f
C8102 w_1575_34786.n22 VSS 2.73452f
C8103 w_1575_34786.t16 VSS 0.01846f
C8104 w_1575_34786.n23 VSS 0.03768f
C8105 w_1575_34786.t14 VSS 0.086116f
C8106 w_1575_34786.n24 VSS 1.43029f
C8107 w_1575_34786.n25 VSS 0.185108f
C8108 w_1575_34786.n26 VSS 0.030618f
C8109 w_1575_34786.n27 VSS 0.111141f
C8110 w_1575_34786.n28 VSS 0.073425f
C8111 w_1575_34786.n29 VSS 0.102689f
C8112 w_1575_34786.n30 VSS 0.026102f
C8113 w_1575_34786.n31 VSS 0.011171f
C8114 w_1575_34786.n32 VSS 0.026801f
C8115 w_1575_34786.n33 VSS 0.022502f
C8116 w_1575_34786.n34 VSS 0.010057f
C8117 w_1575_34786.n35 VSS 0.010057f
C8118 w_1575_34786.n36 VSS 0.022502f
C8119 w_1575_34786.n37 VSS 0.030618f
C8120 w_1575_34786.n38 VSS 0.010057f
C8121 w_1575_34786.t8 VSS 0.165947f
C8122 w_1575_34786.n39 VSS 0.107287f
C8123 w_1575_34786.n40 VSS 0.132019f
C8124 w_1575_34786.n41 VSS 0.252653f
C8125 w_1575_34786.n42 VSS 6.43177f
C8126 w_1575_34786.t13 VSS 6.67928f
C8127 w_1575_34786.n43 VSS 3.88858f
C8128 w_1575_34786.n44 VSS 0.156921f
C8129 w_1575_34786.n45 VSS 0.143611f
C8130 w_1575_34786.n46 VSS 0.046985f
C8131 w_1575_34786.n47 VSS 0.608887f
C8132 w_1575_34786.n48 VSS 0.644966f
C8133 w_1575_34786.n49 VSS 1.4319f
C8134 w_1575_34786.t15 VSS 0.086116f
C8135 w_1575_34786.t11 VSS 0.01846f
C8136 w_1575_34786.n50 VSS 0.03768f
C8137 w_1575_34786.n51 VSS 2.73452f
C8138 w_1575_34786.t12 VSS 0.067657f
C8139 w_1575_34786.n52 VSS 1.43072f
C8140 w_1575_34786.n53 VSS 0.275517f
C8141 w_1575_34786.n54 VSS 0.663641f
C8142 w_1575_34786.n55 VSS 0.146189f
C8143 w_1575_34786.n56 VSS 0.097053f
C8144 w_1575_34786.n57 VSS 0.155341f
C8145 w_1575_34786.n58 VSS 3.60692f
C8146 w_1575_34786.n59 VSS 0.573236f
C8147 w_1575_34786.t0 VSS 0.224824f
C8148 w_1575_34786.t2 VSS 0.16688f
C8149 w_1575_34786.n60 VSS 0.111253f
C8150 w_1575_34786.t6 VSS 0.16688f
C8151 w_1575_34786.t4 VSS 0.328835f
C8152 w_1575_34786.n61 VSS 0.335938f
C8153 w_1575_34786.n62 VSS 0.027497f
C8154 w_1575_34786.n63 VSS 0.037403f
C8155 w_1575_34786.n64 VSS 0.080959f
C8156 w_1575_34786.n65 VSS 0.125932f
C8157 w_1575_34786.n66 VSS 0.163439f
C8158 w_1575_34786.n67 VSS 0.039349f
C8159 w_1575_34786.t5 VSS 0.090587f
C8160 w_1575_34786.n68 VSS 0.290963f
C8161 w_1575_34786.n69 VSS 0.055466f
C8162 w_1575_34786.t7 VSS 0.024713f
C8163 EN_VIN_BSTR_P.t6 VSS 0.030933f
C8164 EN_VIN_BSTR_P.t5 VSS 0.030933f
C8165 EN_VIN_BSTR_P.n0 VSS 0.063662f
C8166 EN_VIN_BSTR_P.t3 VSS 0.030933f
C8167 EN_VIN_BSTR_P.t4 VSS 0.030933f
C8168 EN_VIN_BSTR_P.n1 VSS 0.063662f
C8169 EN_VIN_BSTR_P.t10 VSS 0.016326f
C8170 EN_VIN_BSTR_P.t7 VSS 0.041127f
C8171 EN_VIN_BSTR_P.t16 VSS 0.04343f
C8172 EN_VIN_BSTR_P.n2 VSS 0.058307f
C8173 EN_VIN_BSTR_P.n3 VSS 0.312119f
C8174 EN_VIN_BSTR_P.n4 VSS 0.06955f
C8175 EN_VIN_BSTR_P.n5 VSS 0.074759f
C8176 EN_VIN_BSTR_P.t2 VSS 0.107508f
C8177 EN_VIN_BSTR_P.t0 VSS 0.111067f
C8178 EN_VIN_BSTR_P.t1 VSS 0.107639f
C8179 EN_VIN_BSTR_P.n6 VSS 0.285815f
C8180 EN_VIN_BSTR_P.n7 VSS 0.17615f
C8181 EN_VIN_BSTR_P.n8 VSS 0.083622f
C8182 EN_VIN_BSTR_P.t21 VSS 0.016204f
C8183 EN_VIN_BSTR_P.t17 VSS 0.01635f
C8184 EN_VIN_BSTR_P.n9 VSS 0.11489f
C8185 EN_VIN_BSTR_P.t20 VSS 0.016204f
C8186 EN_VIN_BSTR_P.t23 VSS 0.016207f
C8187 EN_VIN_BSTR_P.t15 VSS 0.020036f
C8188 EN_VIN_BSTR_P.t8 VSS 0.023039f
C8189 EN_VIN_BSTR_P.n10 VSS 0.033139f
C8190 EN_VIN_BSTR_P.t12 VSS 0.02977f
C8191 EN_VIN_BSTR_P.n11 VSS 0.061739f
C8192 EN_VIN_BSTR_P.t19 VSS 0.016182f
C8193 EN_VIN_BSTR_P.n12 VSS 0.032604f
C8194 EN_VIN_BSTR_P.t13 VSS 0.016182f
C8195 EN_VIN_BSTR_P.n13 VSS 0.038345f
C8196 EN_VIN_BSTR_P.t22 VSS 0.016182f
C8197 EN_VIN_BSTR_P.n14 VSS 0.038345f
C8198 EN_VIN_BSTR_P.t14 VSS 0.016182f
C8199 EN_VIN_BSTR_P.n15 VSS 0.02944f
C8200 EN_VIN_BSTR_P.n16 VSS 0.058941f
C8201 EN_VIN_BSTR_P.n17 VSS 0.0656f
C8202 EN_VIN_BSTR_P.n18 VSS 0.352047f
C8203 EN_VIN_BSTR_P.t11 VSS 0.08989f
C8204 EN_VIN_BSTR_P.t9 VSS 0.083309f
C8205 EN_VIN_BSTR_P.t18 VSS 0.085697f
C8206 EN_VIN_BSTR_P.n19 VSS 0.075473f
C8207 EN_VIN_BSTR_P.n20 VSS 0.086725f
C8208 EN_VIN_BSTR_P.n21 VSS 0.517007f
C8209 C10_P_btm.t20 VSS 0.122926f
C8210 C10_P_btm.t21 VSS 0.122926f
C8211 C10_P_btm.n0 VSS 0.39276f
C8212 C10_P_btm.t22 VSS 0.122926f
C8213 C10_P_btm.t17 VSS 0.122926f
C8214 C10_P_btm.n1 VSS 0.379868f
C8215 C10_P_btm.n2 VSS 1.19496f
C8216 C10_P_btm.t30 VSS 0.122926f
C8217 C10_P_btm.t19 VSS 0.122926f
C8218 C10_P_btm.n3 VSS 0.379868f
C8219 C10_P_btm.n4 VSS 0.613462f
C8220 C10_P_btm.t31 VSS 0.122926f
C8221 C10_P_btm.t27 VSS 0.122926f
C8222 C10_P_btm.n5 VSS 0.379868f
C8223 C10_P_btm.n6 VSS 0.613462f
C8224 C10_P_btm.t23 VSS 0.122926f
C8225 C10_P_btm.t29 VSS 0.122926f
C8226 C10_P_btm.n7 VSS 0.379868f
C8227 C10_P_btm.n8 VSS 0.613462f
C8228 C10_P_btm.t25 VSS 0.122926f
C8229 C10_P_btm.t18 VSS 0.122926f
C8230 C10_P_btm.n9 VSS 0.379868f
C8231 C10_P_btm.n10 VSS 0.613462f
C8232 C10_P_btm.t24 VSS 0.122926f
C8233 C10_P_btm.t28 VSS 0.122926f
C8234 C10_P_btm.n11 VSS 0.379868f
C8235 C10_P_btm.n12 VSS 0.612599f
C8236 C10_P_btm.t26 VSS 0.122926f
C8237 C10_P_btm.t16 VSS 0.122926f
C8238 C10_P_btm.n13 VSS 0.379868f
C8239 C10_P_btm.n14 VSS 1.05453f
C8240 C10_P_btm.t11 VSS 0.139882f
C8241 C10_P_btm.t13 VSS 0.139882f
C8242 C10_P_btm.n15 VSS 0.57718f
C8243 C10_P_btm.t12 VSS 0.139882f
C8244 C10_P_btm.t14 VSS 0.139882f
C8245 C10_P_btm.n16 VSS 0.563454f
C8246 C10_P_btm.n17 VSS 0.845221f
C8247 C10_P_btm.t9 VSS 0.139882f
C8248 C10_P_btm.t8 VSS 0.139882f
C8249 C10_P_btm.n18 VSS 0.563454f
C8250 C10_P_btm.n19 VSS 0.434279f
C8251 C10_P_btm.t10 VSS 0.139882f
C8252 C10_P_btm.t15 VSS 0.139882f
C8253 C10_P_btm.n20 VSS 0.563454f
C8254 C10_P_btm.n21 VSS 0.493206f
C8255 C10_P_btm.n22 VSS 0.690049f
C8256 C10_P_btm.t32 VSS 0.139882f
C8257 C10_P_btm.t33 VSS 0.139882f
C8258 C10_P_btm.n23 VSS 0.69103f
C8259 C10_P_btm.n24 VSS 0.588284f
C8260 C10_P_btm.t5 VSS 0.139882f
C8261 C10_P_btm.t2 VSS 0.139882f
C8262 C10_P_btm.n25 VSS 0.583821f
C8263 C10_P_btm.t0 VSS 0.139882f
C8264 C10_P_btm.t3 VSS 0.139882f
C8265 C10_P_btm.n26 VSS 0.569903f
C8266 C10_P_btm.n27 VSS 0.861377f
C8267 C10_P_btm.t1 VSS 0.139882f
C8268 C10_P_btm.t4 VSS 0.139882f
C8269 C10_P_btm.n28 VSS 0.569903f
C8270 C10_P_btm.n29 VSS 0.443544f
C8271 C10_P_btm.t7 VSS 0.139882f
C8272 C10_P_btm.t6 VSS 0.139882f
C8273 C10_P_btm.n30 VSS 0.569903f
C8274 C10_P_btm.n31 VSS 0.497297f
C8275 C10_P_btm.n32 VSS 2.46108f
C8276 C10_P_btm.n33 VSS 2.05058f
C8277 C10_P_btm.n34 VSS 0.908087f
C8278 C10_P_btm.n35 VSS 0.911266f
C8279 C10_P_btm.n36 VSS 0.911266f
C8280 C10_P_btm.n37 VSS 0.908087f
C8281 C10_P_btm.n38 VSS 0.911266f
C8282 C10_P_btm.n39 VSS 0.911266f
C8283 C10_P_btm.n40 VSS 0.911266f
C8284 C10_P_btm.n41 VSS 0.911266f
C8285 C10_P_btm.n42 VSS 0.908087f
C8286 C10_P_btm.n43 VSS 0.911266f
C8287 C10_P_btm.n44 VSS 0.911266f
C8288 C10_P_btm.n45 VSS 0.908087f
C8289 C10_P_btm.n46 VSS 0.911266f
C8290 C10_P_btm.n47 VSS 0.911266f
C8291 C10_P_btm.n48 VSS 0.911266f
C8292 C10_P_btm.n49 VSS 0.911266f
C8293 C10_P_btm.n50 VSS 0.908087f
C8294 C10_P_btm.n51 VSS 0.911266f
C8295 C10_P_btm.n52 VSS 0.911266f
C8296 C10_P_btm.n53 VSS 0.908087f
C8297 C10_P_btm.n54 VSS 0.911266f
C8298 C10_P_btm.n55 VSS 0.911266f
C8299 C10_P_btm.n56 VSS 0.911266f
C8300 C10_P_btm.n57 VSS 0.911266f
C8301 C10_P_btm.n58 VSS 0.908087f
C8302 C10_P_btm.n59 VSS 0.911266f
C8303 C10_P_btm.n60 VSS 0.911266f
C8304 C10_P_btm.n61 VSS 0.908087f
C8305 C10_P_btm.n62 VSS 0.911266f
C8306 C10_P_btm.n63 VSS 0.911266f
C8307 C10_P_btm.n64 VSS 0.911266f
C8308 C10_P_btm.n65 VSS 1.14567f
C8309 C10_P_btm.n66 VSS 0.911266f
C8310 C10_P_btm.n67 VSS 0.911266f
C8311 C10_P_btm.n68 VSS 0.911266f
C8312 C10_P_btm.n69 VSS 0.911266f
C8313 C10_P_btm.n70 VSS 0.911266f
C8314 C10_P_btm.n71 VSS 0.911266f
C8315 C10_P_btm.n72 VSS 0.911266f
C8316 C10_P_btm.n73 VSS 0.911266f
C8317 C10_P_btm.n74 VSS 0.911266f
C8318 C10_P_btm.n75 VSS 0.911266f
C8319 C10_P_btm.n76 VSS 0.911266f
C8320 C10_P_btm.n77 VSS 0.911266f
C8321 C10_P_btm.n78 VSS 0.670504f
C8322 C10_P_btm.n79 VSS 0.911266f
C8323 C10_P_btm.n80 VSS 0.911266f
C8324 C10_P_btm.n81 VSS 0.911266f
C8325 C10_P_btm.n82 VSS 0.911266f
C8326 C10_P_btm.n83 VSS 0.911266f
C8327 C10_P_btm.n84 VSS 0.911266f
C8328 C10_P_btm.n85 VSS 0.911266f
C8329 C10_P_btm.n86 VSS 0.911266f
C8330 C10_P_btm.n87 VSS 0.911266f
C8331 C10_P_btm.n88 VSS 0.911266f
C8332 C10_P_btm.n89 VSS 0.911266f
C8333 C10_P_btm.n90 VSS 0.911266f
C8334 C10_P_btm.n91 VSS 0.911266f
C8335 C10_P_btm.n92 VSS 0.911266f
C8336 C10_P_btm.n93 VSS 0.911266f
C8337 C10_P_btm.n94 VSS 0.911266f
C8338 C10_P_btm.n95 VSS 0.911266f
C8339 C10_P_btm.n96 VSS 0.911266f
C8340 C10_P_btm.n97 VSS 0.911266f
C8341 C10_P_btm.n98 VSS 0.911266f
C8342 C10_P_btm.n99 VSS 0.911266f
C8343 C10_P_btm.n100 VSS 0.911266f
C8344 C10_P_btm.n101 VSS 0.911266f
C8345 C10_P_btm.n102 VSS 0.911266f
C8346 C10_P_btm.n103 VSS 0.911266f
C8347 C10_P_btm.n104 VSS 0.911266f
C8348 C10_P_btm.n105 VSS 0.911266f
C8349 C10_P_btm.n106 VSS 0.911266f
C8350 C10_P_btm.n107 VSS 0.911266f
C8351 C10_P_btm.n108 VSS 0.911266f
C8352 C10_P_btm.n109 VSS 0.911266f
C8353 C10_P_btm.n110 VSS 0.911266f
C8354 C10_P_btm.n111 VSS 0.911266f
C8355 C10_P_btm.n112 VSS 2.05058f
C8356 C10_P_btm.n113 VSS 0.911266f
C8357 C10_P_btm.n114 VSS 0.911266f
C8358 C10_P_btm.n115 VSS 0.911266f
C8359 C10_P_btm.n116 VSS 0.911266f
C8360 C10_P_btm.n117 VSS 0.911266f
C8361 C10_P_btm.n118 VSS 0.911266f
C8362 C10_P_btm.n119 VSS 0.911266f
C8363 C10_P_btm.n120 VSS 0.911266f
C8364 C10_P_btm.n121 VSS 0.911266f
C8365 C10_P_btm.n122 VSS 0.911266f
C8366 C10_P_btm.n123 VSS 0.911266f
C8367 C10_P_btm.n124 VSS 0.911266f
C8368 C10_P_btm.n125 VSS 0.911266f
C8369 C10_P_btm.n126 VSS 1.16658f
C8370 C10_P_btm.n127 VSS 0.911266f
C8371 C10_P_btm.n128 VSS 0.911266f
C8372 C10_P_btm.n129 VSS 3.97703f
C8373 C10_P_btm.n130 VSS 2.82095f
C8374 C10_P_btm.n131 VSS 0.911266f
C8375 C10_P_btm.n132 VSS 0.911266f
C8376 C10_P_btm.n133 VSS 0.911266f
C8377 C10_P_btm.n134 VSS 0.908087f
C8378 C10_P_btm.n135 VSS 0.908087f
C8379 C10_P_btm.n136 VSS 0.908087f
C8380 C10_P_btm.n137 VSS 0.908087f
C8381 C10_P_btm.n138 VSS 0.908087f
C8382 C10_P_btm.n139 VSS 0.911266f
C8383 C10_P_btm.n140 VSS 0.911266f
C8384 C10_P_btm.n141 VSS 0.911266f
C8385 C10_P_btm.n142 VSS 0.908087f
C8386 C10_P_btm.n143 VSS 0.911266f
C8387 C10_P_btm.n144 VSS 0.911266f
C8388 C10_P_btm.n145 VSS 0.908087f
C8389 C10_P_btm.n146 VSS 0.911266f
C8390 C10_P_btm.n147 VSS 0.911266f
C8391 C10_P_btm.n148 VSS 0.911266f
C8392 C10_P_btm.n149 VSS 0.911266f
C8393 C10_P_btm.n150 VSS 0.911266f
C8394 C10_P_btm.n151 VSS 0.908087f
C8395 C10_P_btm.n152 VSS 0.908087f
C8396 C10_P_btm.n153 VSS 0.908087f
C8397 C10_P_btm.n154 VSS 0.908087f
C8398 C10_P_btm.n155 VSS 0.911266f
C8399 C10_P_btm.n156 VSS 0.911266f
C8400 C10_P_btm.n157 VSS 0.911266f
C8401 C10_P_btm.n158 VSS 0.911266f
C8402 C10_P_btm.n159 VSS 0.911266f
C8403 C10_P_btm.n160 VSS 0.908087f
C8404 C10_P_btm.n161 VSS 0.908087f
C8405 C10_P_btm.n162 VSS 0.908087f
C8406 C10_P_btm.n163 VSS 0.908087f
C8407 C10_P_btm.n164 VSS 0.911266f
C8408 C10_P_btm.n165 VSS 0.911266f
C8409 C10_P_btm.n166 VSS 0.911266f
C8410 C10_P_btm.n167 VSS 0.911266f
C8411 C10_P_btm.n168 VSS 0.911266f
C8412 C10_P_btm.n169 VSS 0.908087f
C8413 C10_P_btm.n170 VSS 0.908087f
C8414 C10_P_btm.n171 VSS 0.911266f
C8415 C10_P_btm.n172 VSS 0.911266f
C8416 C10_P_btm.n173 VSS 0.911266f
C8417 C10_P_btm.n174 VSS 1.42745f
C8418 C10_P_btm.n175 VSS 0.911266f
C8419 C10_P_btm.n176 VSS 0.911266f
C8420 C10_P_btm.n177 VSS 0.911266f
C8421 C10_P_btm.n178 VSS 0.670504f
C8422 C10_P_btm.n179 VSS 0.911266f
C8423 C10_P_btm.n180 VSS 0.911266f
C8424 C10_P_btm.n181 VSS 0.911266f
C8425 C10_P_btm.n182 VSS 0.911266f
C8426 C10_P_btm.n183 VSS 0.911266f
C8427 C10_P_btm.n184 VSS 0.670504f
C8428 C10_P_btm.n185 VSS 0.670504f
C8429 C10_P_btm.n186 VSS 0.911266f
C8430 C10_P_btm.n187 VSS 0.911266f
C8431 C10_P_btm.n188 VSS 0.911266f
C8432 C10_P_btm.n189 VSS 0.911266f
C8433 C10_P_btm.n190 VSS 0.911266f
C8434 C10_P_btm.n191 VSS 0.911266f
C8435 C10_P_btm.n192 VSS 0.911266f
C8436 C10_P_btm.n193 VSS 0.911266f
C8437 C10_P_btm.n194 VSS 0.911266f
C8438 C10_P_btm.n195 VSS 0.911266f
C8439 C10_P_btm.n196 VSS 0.911266f
C8440 C10_P_btm.n197 VSS 0.911266f
C8441 C10_P_btm.n198 VSS 0.911266f
C8442 C10_P_btm.n199 VSS 0.911266f
C8443 C10_P_btm.n200 VSS 0.911266f
C8444 C10_P_btm.n201 VSS 0.911266f
C8445 C10_P_btm.n202 VSS 0.911266f
C8446 C10_P_btm.n203 VSS 0.911266f
C8447 C10_P_btm.n204 VSS 0.911266f
C8448 C10_P_btm.n205 VSS 0.911266f
C8449 C10_P_btm.n206 VSS 0.911266f
C8450 C10_P_btm.n207 VSS 0.911266f
C8451 C10_P_btm.n208 VSS 0.911266f
C8452 C10_P_btm.n209 VSS 0.911266f
C8453 C10_P_btm.n210 VSS 0.911266f
C8454 C10_P_btm.n211 VSS 0.911266f
C8455 C10_P_btm.n212 VSS 0.911266f
C8456 C10_P_btm.n213 VSS 0.911266f
C8457 C10_P_btm.n214 VSS 0.911266f
C8458 C10_P_btm.n215 VSS 0.911266f
C8459 C10_P_btm.n216 VSS 0.911266f
C8460 C10_P_btm.n217 VSS 0.911266f
C8461 C10_P_btm.n218 VSS 0.911266f
C8462 C10_P_btm.n219 VSS 0.911266f
C8463 C10_P_btm.n220 VSS 0.911266f
C8464 C10_P_btm.n221 VSS 0.911266f
C8465 C10_P_btm.n222 VSS 0.911266f
C8466 C10_P_btm.n223 VSS 0.911266f
C8467 C10_P_btm.n224 VSS 0.911266f
C8468 C10_P_btm.n225 VSS 0.911266f
C8469 C10_P_btm.n226 VSS 0.911266f
C8470 C10_P_btm.n227 VSS 0.911266f
C8471 C10_P_btm.n228 VSS 0.911266f
C8472 C10_P_btm.n229 VSS 0.911266f
C8473 C10_P_btm.n230 VSS 0.911266f
C8474 C10_P_btm.n231 VSS 0.911266f
C8475 C10_P_btm.n232 VSS 0.911266f
C8476 C10_P_btm.n233 VSS 0.911266f
C8477 C10_P_btm.n234 VSS 0.911266f
C8478 C10_P_btm.n235 VSS 0.911266f
C8479 C10_P_btm.n236 VSS 0.911266f
C8480 C10_P_btm.n237 VSS 0.911266f
C8481 C10_P_btm.n238 VSS 0.911266f
C8482 C10_P_btm.n239 VSS 0.911266f
C8483 C10_P_btm.n240 VSS 0.911266f
C8484 C10_P_btm.n241 VSS 0.911266f
C8485 C10_P_btm.n242 VSS 0.911266f
C8486 C10_P_btm.n243 VSS 0.911266f
C8487 C10_P_btm.n244 VSS 0.911266f
C8488 C10_P_btm.n245 VSS 0.911266f
C8489 C10_P_btm.n246 VSS 0.911266f
C8490 C10_P_btm.n247 VSS 0.911266f
C8491 C10_P_btm.n248 VSS 0.911266f
C8492 C10_P_btm.n249 VSS 0.911266f
C8493 C10_P_btm.n250 VSS 0.911266f
C8494 C10_P_btm.n251 VSS 0.911266f
C8495 C10_P_btm.n252 VSS 0.911266f
C8496 C10_P_btm.n253 VSS 0.911266f
C8497 C10_P_btm.n254 VSS 0.911266f
C8498 C10_P_btm.n255 VSS 0.911266f
C8499 C10_P_btm.n256 VSS 0.911266f
C8500 C10_P_btm.n257 VSS 0.911266f
C8501 C10_P_btm.n258 VSS 0.911266f
C8502 C10_P_btm.n259 VSS 0.911266f
C8503 C10_P_btm.n260 VSS 0.911266f
C8504 C10_P_btm.n261 VSS 0.670504f
C8505 C10_P_btm.n262 VSS 0.670504f
C8506 C10_P_btm.n263 VSS 0.670504f
C8507 C10_P_btm.n264 VSS 1.29967f
C8508 C10_P_btm.n265 VSS 0.911266f
C8509 C10_P_btm.n266 VSS 0.911266f
C8510 C10_P_btm.n267 VSS 0.911266f
C8511 C10_P_btm.n268 VSS 1.09755f
C8512 C10_P_btm.n269 VSS 0.908087f
C8513 C10_P_btm.n270 VSS 0.908087f
C8514 C10_P_btm.n271 VSS 0.908087f
C8515 C10_P_btm.n272 VSS 0.908087f
C8516 C10_P_btm.n273 VSS 0.911266f
C8517 C10_P_btm.n274 VSS 0.911266f
C8518 C10_P_btm.n275 VSS 0.911266f
C8519 C10_P_btm.n276 VSS 0.911266f
C8520 C10_P_btm.n277 VSS 0.911266f
C8521 C10_P_btm.n278 VSS 0.911266f
C8522 C10_P_btm.n279 VSS 0.911266f
C8523 C10_P_btm.n280 VSS 0.911266f
C8524 C10_P_btm.n281 VSS 0.911266f
C8525 C10_P_btm.n282 VSS 0.911266f
C8526 C10_P_btm.n283 VSS 0.911266f
C8527 C10_P_btm.n284 VSS 0.911266f
C8528 C10_P_btm.n285 VSS 0.911266f
C8529 C10_P_btm.n286 VSS 0.911266f
C8530 C10_P_btm.n287 VSS 0.911266f
C8531 C10_P_btm.n288 VSS 0.911266f
C8532 C10_P_btm.n289 VSS 0.911266f
C8533 C10_P_btm.n290 VSS 0.911266f
C8534 C10_P_btm.n291 VSS 0.911266f
C8535 C10_P_btm.n292 VSS 0.911266f
C8536 C10_P_btm.n293 VSS 0.908087f
C8537 C10_P_btm.n294 VSS 0.908087f
C8538 C10_P_btm.n295 VSS 0.908087f
C8539 C10_P_btm.n296 VSS 0.908087f
C8540 C10_P_btm.n297 VSS 0.908087f
C8541 C10_P_btm.n298 VSS 0.911266f
C8542 C10_P_btm.n299 VSS 0.911266f
C8543 C10_P_btm.n300 VSS 0.911266f
C8544 C10_P_btm.n301 VSS 0.911266f
C8545 C10_P_btm.n302 VSS 0.911266f
C8546 C10_P_btm.n303 VSS 0.911266f
C8547 C10_P_btm.n304 VSS 0.911266f
C8548 C10_P_btm.n305 VSS 0.911266f
C8549 C10_P_btm.n306 VSS 0.911266f
C8550 C10_P_btm.n307 VSS 0.911266f
C8551 C10_P_btm.n308 VSS 0.911266f
C8552 C10_P_btm.n309 VSS 2.05058f
C8553 C10_P_btm.n310 VSS 2.05058f
C8554 C10_P_btm.n311 VSS 2.05058f
C8555 C10_P_btm.n312 VSS 2.05058f
C8556 C10_P_btm.n313 VSS 2.05058f
C8557 C10_P_btm.n314 VSS 0.911266f
C8558 C10_P_btm.n315 VSS 0.911266f
C8559 C10_P_btm.n316 VSS 0.911266f
C8560 C10_P_btm.n317 VSS 0.911266f
C8561 C10_P_btm.n318 VSS 0.911266f
C8562 C10_P_btm.n319 VSS 0.911266f
C8563 C10_P_btm.n320 VSS 0.911266f
C8564 C10_P_btm.n321 VSS 0.911266f
C8565 C10_P_btm.n322 VSS 0.911266f
C8566 C10_P_btm.n323 VSS 0.911266f
C8567 C10_P_btm.n324 VSS 0.911266f
C8568 C10_P_btm.n325 VSS 0.911266f
C8569 C10_P_btm.n326 VSS 0.911266f
C8570 C10_P_btm.n327 VSS 0.911266f
C8571 C10_P_btm.n328 VSS 0.911266f
C8572 C10_P_btm.n329 VSS 0.911266f
C8573 C10_P_btm.n330 VSS 0.911266f
C8574 C10_P_btm.n331 VSS 0.911266f
C8575 C10_P_btm.n332 VSS 0.911266f
C8576 C10_P_btm.n333 VSS 0.911266f
C8577 C10_P_btm.n334 VSS 0.911266f
C8578 C10_P_btm.n335 VSS 0.911266f
C8579 C10_P_btm.n336 VSS 0.911266f
C8580 C10_P_btm.n337 VSS 0.911266f
C8581 C10_P_btm.n338 VSS 0.911266f
C8582 C10_P_btm.n339 VSS 0.911266f
C8583 C10_P_btm.n340 VSS 0.911266f
C8584 C10_P_btm.n341 VSS 0.911266f
C8585 C10_P_btm.n342 VSS 0.911266f
C8586 C10_P_btm.n343 VSS 0.911266f
C8587 C10_P_btm.n344 VSS 0.911266f
C8588 C10_P_btm.n345 VSS 0.911266f
C8589 C10_P_btm.n346 VSS 0.911266f
C8590 C10_P_btm.n347 VSS 0.911266f
C8591 C10_P_btm.n348 VSS 0.911266f
C8592 C10_P_btm.n349 VSS 0.911266f
C8593 C10_P_btm.n350 VSS 0.911266f
C8594 C10_P_btm.n351 VSS 0.911266f
C8595 C10_P_btm.n352 VSS 0.911266f
C8596 C10_P_btm.n353 VSS 0.911266f
C8597 C10_P_btm.n354 VSS 0.911266f
C8598 C10_P_btm.n355 VSS 0.670504f
C8599 C10_P_btm.n356 VSS 0.670504f
C8600 C10_P_btm.n357 VSS 0.670504f
C8601 C10_P_btm.n358 VSS 0.911266f
C8602 C10_P_btm.n359 VSS 0.911266f
C8603 C10_P_btm.n360 VSS 0.670504f
C8604 C10_P_btm.n361 VSS 0.911266f
C8605 C10_P_btm.n362 VSS 0.911266f
C8606 C10_P_btm.n363 VSS 0.911266f
C8607 C10_P_btm.n364 VSS 0.911266f
C8608 C10_P_btm.n365 VSS 0.911266f
C8609 C10_P_btm.n366 VSS 0.911266f
C8610 C10_P_btm.n367 VSS 0.911266f
C8611 C10_P_btm.n368 VSS 0.911266f
C8612 C10_P_btm.n369 VSS 0.911266f
C8613 C10_P_btm.n370 VSS 0.911266f
C8614 C10_P_btm.n371 VSS 0.911266f
C8615 C10_P_btm.n372 VSS 0.879752f
C8616 C10_P_btm.n373 VSS 0.911266f
C8617 C10_P_btm.n374 VSS 0.911266f
C8618 C10_P_btm.n375 VSS 0.911266f
C8619 C10_P_btm.n376 VSS 0.911266f
C8620 C10_P_btm.n377 VSS 0.911266f
C8621 C10_P_btm.n378 VSS 0.911266f
C8622 C10_P_btm.n379 VSS 0.911266f
C8623 C10_P_btm.n380 VSS 0.911266f
C8624 C10_P_btm.n381 VSS 0.911266f
C8625 C10_P_btm.n382 VSS 0.911266f
C8626 C10_P_btm.n383 VSS 0.670504f
C8627 C10_P_btm.n384 VSS 0.911266f
C8628 C10_P_btm.n385 VSS 0.670504f
C8629 C10_P_btm.n386 VSS 0.670504f
C8630 C10_P_btm.n387 VSS 0.911266f
C8631 C10_P_btm.n388 VSS 0.911266f
C8632 C10_P_btm.n389 VSS 0.911266f
C8633 C10_P_btm.n390 VSS 0.911266f
C8634 C10_P_btm.n391 VSS 0.911266f
C8635 C10_P_btm.n392 VSS 0.911266f
C8636 C10_P_btm.n393 VSS 0.911266f
C8637 C10_P_btm.n394 VSS 0.670504f
C8638 C10_P_btm.n395 VSS 0.670504f
C8639 C10_P_btm.n396 VSS 0.911266f
C8640 C10_P_btm.n397 VSS 0.911266f
C8641 C10_P_btm.n398 VSS 0.911266f
C8642 C10_P_btm.n399 VSS 0.911266f
C8643 C10_P_btm.n400 VSS 0.911266f
C8644 C10_P_btm.n401 VSS 0.911266f
C8645 C10_P_btm.n402 VSS 0.911266f
C8646 C10_P_btm.n403 VSS 0.911266f
C8647 C10_P_btm.n404 VSS 0.911266f
C8648 C10_P_btm.n405 VSS 0.670504f
C8649 C10_P_btm.n406 VSS 0.911266f
C8650 C10_P_btm.n407 VSS 0.911266f
C8651 C10_P_btm.n408 VSS 0.911266f
C8652 C10_P_btm.n409 VSS 0.911266f
C8653 C10_P_btm.n410 VSS 0.911266f
C8654 C10_P_btm.n411 VSS 0.911266f
C8655 C10_P_btm.n412 VSS 0.911266f
C8656 C10_P_btm.n413 VSS 0.911266f
C8657 C10_P_btm.n414 VSS 1.14567f
C8658 C10_P_btm.n415 VSS 0.911266f
C8659 C10_P_btm.n416 VSS 0.911266f
C8660 C10_P_btm.n417 VSS 0.911266f
C8661 C10_P_btm.n418 VSS 0.911266f
C8662 C10_P_btm.n419 VSS 0.911266f
C8663 C10_P_btm.n420 VSS 0.911266f
C8664 C10_P_btm.n421 VSS 0.911266f
C8665 C10_P_btm.n422 VSS 0.911266f
C8666 C10_P_btm.n423 VSS 0.911266f
C8667 C10_P_btm.n424 VSS 0.670504f
C8668 C10_P_btm.n425 VSS 0.670504f
C8669 C10_P_btm.n426 VSS 0.670504f
C8670 C10_P_btm.n427 VSS 0.911266f
C8671 C10_P_btm.n428 VSS 0.911266f
C8672 C10_P_btm.n429 VSS 0.670504f
C8673 C10_P_btm.n430 VSS 0.911266f
C8674 C10_P_btm.n431 VSS 0.911266f
C8675 C10_P_btm.n432 VSS 0.911266f
C8676 C10_P_btm.n433 VSS 0.911266f
C8677 C10_P_btm.n434 VSS 0.911266f
C8678 C10_P_btm.n435 VSS 0.911266f
C8679 C10_P_btm.n436 VSS 0.911266f
C8680 C10_P_btm.n437 VSS 0.911266f
C8681 C10_P_btm.n438 VSS 0.911266f
C8682 C10_P_btm.n439 VSS 0.911266f
C8683 C10_P_btm.n440 VSS 0.911266f
C8684 C10_P_btm.n441 VSS 1.14567f
C8685 C10_P_btm.n442 VSS 0.911266f
C8686 C10_P_btm.n443 VSS 0.911266f
C8687 C10_P_btm.n444 VSS 0.911266f
C8688 C10_P_btm.n445 VSS 0.911266f
C8689 C10_P_btm.n446 VSS 0.911266f
C8690 C10_P_btm.n447 VSS 0.911266f
C8691 C10_P_btm.n448 VSS 0.911266f
C8692 C10_P_btm.n449 VSS 0.911266f
C8693 C10_P_btm.n450 VSS 0.911266f
C8694 C10_P_btm.n451 VSS 0.670504f
C8695 C10_P_btm.n452 VSS 0.670504f
C8696 C10_P_btm.n453 VSS 0.911266f
C8697 C10_P_btm.n454 VSS 0.911266f
C8698 C10_P_btm.n455 VSS 0.911266f
C8699 C10_P_btm.n456 VSS 0.911266f
C8700 C10_P_btm.n457 VSS 0.911266f
C8701 C10_P_btm.n458 VSS 0.911266f
C8702 C10_P_btm.n459 VSS 0.670504f
C8703 C10_P_btm.n460 VSS 0.670504f
C8704 C10_P_btm.n461 VSS 0.670504f
C8705 C10_P_btm.n462 VSS 0.911266f
C8706 C10_P_btm.n463 VSS 0.670504f
C8707 C10_P_btm.n464 VSS 0.911266f
C8708 C10_P_btm.n465 VSS 0.911266f
C8709 C10_P_btm.n466 VSS 0.911266f
C8710 C10_P_btm.n467 VSS 0.911266f
C8711 C10_P_btm.n468 VSS 0.911266f
C8712 C10_P_btm.n469 VSS 0.911266f
C8713 C10_P_btm.n470 VSS 1.14567f
C8714 C10_P_btm.n471 VSS 0.911266f
C8715 C10_P_btm.n472 VSS 0.911266f
C8716 C10_P_btm.n473 VSS 0.911266f
C8717 C10_P_btm.n474 VSS 0.911266f
C8718 C10_P_btm.n475 VSS 0.911266f
C8719 C10_P_btm.n476 VSS 0.911266f
C8720 C10_P_btm.n477 VSS 0.911266f
C8721 C10_P_btm.n478 VSS 0.911266f
C8722 C10_P_btm.n479 VSS 0.670504f
C8723 C10_P_btm.n480 VSS 0.911266f
C8724 C10_P_btm.n481 VSS 0.911266f
C8725 C10_P_btm.n482 VSS 0.911266f
C8726 C10_P_btm.n483 VSS 0.911266f
C8727 C10_P_btm.n484 VSS 0.911266f
C8728 C10_P_btm.n485 VSS 0.911266f
C8729 C10_P_btm.n486 VSS 0.911266f
C8730 C10_P_btm.n487 VSS 0.911266f
C8731 C10_P_btm.n488 VSS 0.911266f
C8732 C10_P_btm.n489 VSS 0.911266f
C8733 C10_P_btm.n490 VSS 0.911266f
C8734 C10_P_btm.n491 VSS 0.911266f
C8735 C10_P_btm.n492 VSS 0.911266f
C8736 C10_P_btm.n493 VSS 0.911266f
C8737 C10_P_btm.n494 VSS 0.908087f
C8738 C10_P_btm.n495 VSS 0.911266f
C8739 C10_P_btm.n496 VSS 0.908087f
C8740 C10_P_btm.n497 VSS 0.911266f
C8741 C10_P_btm.n498 VSS 0.911266f
C8742 C10_P_btm.n499 VSS 0.911266f
C8743 C10_P_btm.n500 VSS 0.911266f
C8744 C10_P_btm.n501 VSS 0.670504f
C8745 C10_P_btm.n502 VSS 0.911266f
C8746 C10_P_btm.n503 VSS 0.911266f
C8747 C10_P_btm.n504 VSS 0.911266f
C8748 C10_P_btm.n505 VSS 0.670504f
C8749 C10_P_btm.n506 VSS 0.670504f
C8750 C10_P_btm.n507 VSS 0.670504f
C8751 C10_P_btm.n508 VSS 0.911266f
C8752 C10_P_btm.n509 VSS 0.911266f
C8753 C10_P_btm.n510 VSS 0.911266f
C8754 C10_P_btm.n511 VSS 0.911266f
C8755 C10_P_btm.n512 VSS 0.911266f
C8756 C10_P_btm.n513 VSS 0.911266f
C8757 C10_P_btm.n514 VSS 0.911266f
C8758 C10_P_btm.n515 VSS 0.911266f
C8759 C10_P_btm.n516 VSS 0.911266f
C8760 C10_P_btm.n517 VSS 1.29961f
C8761 C10_P_btm.n518 VSS 1.42736f
C8762 C10_P_btm.n519 VSS 1.09754f
C8763 C10_P_btm.n520 VSS 0.908087f
C8764 C10_P_btm.n521 VSS 0.911266f
C8765 C10_P_btm.n522 VSS 0.911266f
C8766 C10_P_btm.n523 VSS 0.911266f
C8767 C10_P_btm.n524 VSS 0.911266f
C8768 C10_P_btm.n525 VSS 0.908087f
C8769 C10_P_btm.n526 VSS 0.908087f
C8770 C10_P_btm.n527 VSS 0.908087f
C8771 C10_P_btm.n528 VSS 0.911266f
C8772 C10_P_btm.n529 VSS 0.911266f
C8773 C10_P_btm.n530 VSS 0.908087f
C8774 C10_P_btm.n531 VSS 0.911266f
C8775 C10_P_btm.n532 VSS 0.911266f
C8776 C10_P_btm.n533 VSS 0.908087f
C8777 C10_P_btm.n534 VSS 0.911266f
C8778 C10_P_btm.n535 VSS 0.911266f
C8779 C10_P_btm.n536 VSS 0.911266f
C8780 C10_P_btm.n537 VSS 0.908087f
C8781 C10_P_btm.n538 VSS 0.911266f
C8782 C10_P_btm.n539 VSS 0.911266f
C8783 C10_P_btm.n540 VSS 0.908087f
C8784 C10_P_btm.n541 VSS 0.911266f
C8785 C10_P_btm.n542 VSS 0.911266f
C8786 C10_P_btm.n543 VSS 0.911266f
C8787 C10_P_btm.n544 VSS 0.911266f
C8788 C10_P_btm.n545 VSS 0.908087f
C8789 C10_P_btm.n546 VSS 0.911266f
C8790 C10_P_btm.n547 VSS 0.911266f
C8791 C10_P_btm.n548 VSS 0.908087f
C8792 C10_P_btm.n549 VSS 0.911266f
C8793 C10_P_btm.n550 VSS 0.911266f
C8794 C10_P_btm.n551 VSS 0.911266f
C8795 C10_P_btm.n552 VSS 0.911266f
C8796 C10_P_btm.n553 VSS 2.82105f
C8797 C10_P_btm.n554 VSS 0.911266f
C8798 C10_P_btm.n555 VSS 0.911266f
C8799 C10_P_btm.n556 VSS 2.05058f
C8800 C10_P_btm.n557 VSS 0.911266f
C8801 C10_P_btm.n558 VSS 0.911266f
C8802 C10_P_btm.n559 VSS 0.911266f
C8803 C10_P_btm.n560 VSS 0.911266f
C8804 C10_P_btm.n561 VSS 0.911266f
C8805 C10_P_btm.n562 VSS 0.911266f
C8806 C10_P_btm.n563 VSS 0.911266f
C8807 C10_P_btm.n564 VSS 0.911266f
C8808 C10_P_btm.n565 VSS 0.911266f
C8809 C10_P_btm.n566 VSS 0.911266f
C8810 C10_P_btm.n567 VSS 0.911266f
C8811 C10_P_btm.n568 VSS 0.911266f
C8812 C10_P_btm.n569 VSS 0.911266f
C8813 C10_P_btm.n570 VSS 0.911266f
C8814 C10_P_btm.n571 VSS 0.911266f
C8815 C10_P_btm.n572 VSS 0.911266f
C8816 C10_P_btm.n573 VSS 0.911266f
C8817 C10_P_btm.n574 VSS 0.911266f
C8818 C10_P_btm.n575 VSS 0.911266f
C8819 C10_P_btm.n576 VSS 0.911266f
C8820 C10_P_btm.n577 VSS 0.911266f
C8821 C10_P_btm.n578 VSS 0.911266f
C8822 C10_P_btm.n579 VSS 0.911266f
C8823 C10_P_btm.n580 VSS 0.911266f
C8824 C10_P_btm.n581 VSS 0.911266f
C8825 C10_P_btm.n582 VSS 0.911266f
C8826 C10_P_btm.n583 VSS 0.911266f
C8827 C10_P_btm.n584 VSS 0.911266f
C8828 C10_P_btm.n585 VSS 0.911266f
C8829 C10_P_btm.n586 VSS 0.911266f
C8830 C10_P_btm.n587 VSS 0.911266f
C8831 C10_P_btm.n588 VSS 0.911266f
C8832 C10_P_btm.n589 VSS 0.911266f
C8833 C10_P_btm.n590 VSS 0.911266f
C8834 C10_P_btm.n591 VSS 0.911266f
C8835 C10_P_btm.n592 VSS 0.911266f
C8836 C10_P_btm.n593 VSS 0.911266f
C8837 C10_P_btm.n594 VSS 0.911266f
C8838 C10_P_btm.n595 VSS 0.911266f
C8839 C10_P_btm.n596 VSS 0.911266f
C8840 C10_P_btm.n597 VSS 0.911266f
C8841 C10_P_btm.n598 VSS 0.911266f
C8842 C10_P_btm.n599 VSS 0.911266f
C8843 C10_P_btm.n600 VSS 0.911266f
C8844 C10_P_btm.n601 VSS 0.911266f
C8845 C10_P_btm.n602 VSS 0.911266f
C8846 C10_P_btm.n603 VSS 0.911266f
C8847 C10_P_btm.n604 VSS 0.911266f
C8848 C10_P_btm.n605 VSS 0.908087f
C8849 C10_P_btm.n606 VSS 0.911266f
C8850 C10_P_btm.n607 VSS 0.911266f
C8851 C10_P_btm.n608 VSS 0.911266f
C8852 C10_P_btm.n609 VSS 0.911266f
C8853 C10_P_btm.n610 VSS 0.908087f
C8854 C10_P_btm.n611 VSS 0.911266f
C8855 C10_P_btm.n612 VSS 0.911266f
C8856 C10_P_btm.n613 VSS 0.911266f
C8857 C10_P_btm.n614 VSS 0.911266f
C8858 C10_P_btm.n615 VSS 0.908087f
C8859 C10_P_btm.n616 VSS 0.911266f
C8860 C10_P_btm.n617 VSS 0.911266f
C8861 C10_P_btm.n618 VSS 0.911266f
C8862 C10_P_btm.n619 VSS 0.911266f
C8863 C10_P_btm.n620 VSS 0.908087f
C8864 C10_P_btm.n621 VSS 0.911266f
C8865 C10_P_btm.n622 VSS 0.911266f
C8866 C10_P_btm.n623 VSS 0.911266f
C8867 C10_P_btm.n624 VSS 0.911266f
C8868 C10_P_btm.n625 VSS 0.911266f
C8869 C10_P_btm.n626 VSS 2.05058f
C8870 C10_P_btm.n627 VSS 0.911266f
C8871 C10_P_btm.n628 VSS 0.911266f
C8872 C10_P_btm.n629 VSS 0.911266f
C8873 C10_P_btm.n630 VSS 0.911266f
C8874 C10_P_btm.n631 VSS 0.911266f
C8875 C10_P_btm.n632 VSS 0.911266f
C8876 C10_P_btm.n633 VSS 0.911266f
C8877 C10_P_btm.n634 VSS 0.911266f
C8878 C10_P_btm.n635 VSS 0.911266f
C8879 C10_P_btm.n636 VSS 0.911266f
C8880 C10_P_btm.n637 VSS 0.911266f
C8881 C10_P_btm.n638 VSS 0.911266f
C8882 C10_P_btm.n639 VSS 0.911266f
C8883 C10_P_btm.n640 VSS 0.911266f
C8884 C10_P_btm.n641 VSS 0.911266f
C8885 C10_P_btm.n642 VSS 0.911266f
C8886 C10_P_btm.n643 VSS 0.911266f
C8887 C10_P_btm.n644 VSS 0.911266f
C8888 C10_P_btm.n645 VSS 0.911266f
C8889 C10_P_btm.n646 VSS 0.911266f
C8890 C10_P_btm.n647 VSS 0.911266f
C8891 C10_P_btm.n648 VSS 0.911266f
C8892 C10_P_btm.n649 VSS 0.911266f
C8893 C10_P_btm.n650 VSS 0.911266f
C8894 C10_P_btm.n651 VSS 2.05058f
C8895 C10_P_btm.n652 VSS 3.97703f
C8896 C10_P_btm.n653 VSS 2.82095f
C8897 C10_P_btm.n654 VSS 1.16658f
C8898 C10_P_btm.n655 VSS 0.911266f
C8899 C10_P_btm.n656 VSS 0.911266f
C8900 C10_P_btm.n657 VSS 0.911266f
C8901 C10_P_btm.n658 VSS 0.908087f
C8902 C10_P_btm.n659 VSS 0.908087f
C8903 C10_P_btm.n660 VSS 0.908087f
C8904 C10_P_btm.n661 VSS 0.911266f
C8905 C10_P_btm.n662 VSS 0.911266f
C8906 C10_P_btm.n663 VSS 0.911266f
C8907 C10_P_btm.n664 VSS 0.908087f
C8908 C10_P_btm.n665 VSS 0.908087f
C8909 C10_P_btm.n666 VSS 0.908087f
C8910 C10_P_btm.n667 VSS 0.911266f
C8911 C10_P_btm.n668 VSS 0.911266f
C8912 C10_P_btm.n669 VSS 0.911266f
C8913 C10_P_btm.n670 VSS 0.908087f
C8914 C10_P_btm.n671 VSS 0.908087f
C8915 C10_P_btm.n672 VSS 0.908087f
C8916 C10_P_btm.n673 VSS 0.911266f
C8917 C10_P_btm.n674 VSS 0.911266f
C8918 C10_P_btm.n675 VSS 0.911266f
C8919 C10_P_btm.n676 VSS 0.908087f
C8920 C10_P_btm.n677 VSS 0.908087f
C8921 C10_P_btm.n678 VSS 0.908087f
C8922 C10_P_btm.n679 VSS 0.908087f
C8923 C10_P_btm.n680 VSS 0.911266f
C8924 C10_P_btm.n681 VSS 0.908087f
C8925 C10_P_btm.n682 VSS 0.911266f
C8926 C10_P_btm.n683 VSS 0.911266f
C8927 C10_P_btm.n684 VSS 0.911435f
C8928 C10_P_btm.n685 VSS 0.911266f
C8929 C10_P_btm.n686 VSS 0.911266f
C8930 C10_P_btm.n687 VSS 0.911266f
C8931 C10_P_btm.n688 VSS 0.911266f
C8932 C10_P_btm.n689 VSS 0.911266f
C8933 C10_P_btm.n690 VSS 0.911266f
C8934 C10_P_btm.n691 VSS 0.911266f
C8935 C10_P_btm.n692 VSS 0.911266f
C8936 C10_P_btm.n693 VSS 0.911266f
C8937 C10_P_btm.n694 VSS 0.911266f
C8938 C10_P_btm.n695 VSS 0.911266f
C8939 C10_P_btm.n696 VSS 0.911266f
C8940 C10_P_btm.n697 VSS 0.911266f
C8941 C10_P_btm.n698 VSS 0.911266f
C8942 C10_P_btm.n699 VSS 0.911266f
C8943 C10_P_btm.n700 VSS 0.911266f
C8944 C10_P_btm.n701 VSS 0.911266f
C8945 C10_P_btm.n702 VSS 0.911266f
C8946 C10_P_btm.n703 VSS 0.911266f
C8947 C10_P_btm.n704 VSS 0.911266f
C8948 C10_P_btm.n705 VSS 0.911266f
C8949 C10_P_btm.n706 VSS 0.911266f
C8950 C10_P_btm.n707 VSS 0.911266f
C8951 C10_P_btm.n708 VSS 0.911266f
C8952 C10_P_btm.n709 VSS 0.911266f
C8953 C10_P_btm.n710 VSS 0.911266f
C8954 C10_P_btm.n711 VSS 0.911266f
C8955 C10_P_btm.n712 VSS 0.911266f
C8956 C10_P_btm.n713 VSS 0.911266f
C8957 C10_P_btm.n714 VSS 0.911266f
C8958 C10_P_btm.n715 VSS 0.911266f
C8959 C10_P_btm.n716 VSS 0.911266f
C8960 C10_P_btm.n717 VSS 0.911266f
C8961 C10_P_btm.n718 VSS 0.911266f
C8962 C10_P_btm.n719 VSS 0.911266f
C8963 C10_P_btm.n720 VSS 0.911266f
C8964 C10_P_btm.n721 VSS 0.911266f
C8965 C10_P_btm.n722 VSS 0.911266f
C8966 C10_P_btm.n723 VSS 0.911266f
C8967 C10_P_btm.n724 VSS 0.911266f
C8968 C10_P_btm.n725 VSS 0.911266f
C8969 C10_P_btm.n726 VSS 0.911266f
C8970 C10_P_btm.n727 VSS 0.911266f
C8971 C10_P_btm.n728 VSS 0.908087f
C8972 C10_P_btm.n729 VSS 0.908087f
C8973 C10_P_btm.n730 VSS 0.908087f
C8974 C10_P_btm.n731 VSS 0.911266f
C8975 C10_P_btm.n732 VSS 0.911266f
C8976 C10_P_btm.n733 VSS 0.911266f
C8977 C10_P_btm.n734 VSS 0.911266f
C8978 C10_P_btm.n735 VSS 0.911266f
C8979 C10_P_btm.n736 VSS 0.911266f
C8980 C10_P_btm.n737 VSS 0.911266f
C8981 C10_P_btm.n738 VSS 0.911266f
C8982 C10_P_btm.n739 VSS 0.911266f
C8983 C10_P_btm.n740 VSS 0.911266f
C8984 C10_P_btm.n741 VSS 0.911266f
C8985 C10_P_btm.n742 VSS 0.911266f
C8986 C10_P_btm.n743 VSS 0.911266f
C8987 C10_P_btm.n744 VSS 0.911266f
C8988 C10_P_btm.n745 VSS 0.911266f
C8989 C10_P_btm.n746 VSS 0.911266f
C8990 C10_P_btm.n747 VSS 0.911266f
C8991 C10_P_btm.n748 VSS 0.911266f
C8992 C10_P_btm.n749 VSS 0.911266f
C8993 C10_P_btm.n750 VSS 0.911266f
C8994 C10_P_btm.n751 VSS 0.911266f
C8995 C10_P_btm.n752 VSS 0.911266f
C8996 C10_P_btm.n753 VSS 0.911266f
C8997 C10_P_btm.n754 VSS 0.911266f
C8998 C10_P_btm.n755 VSS 0.911266f
C8999 C10_P_btm.n756 VSS 0.911266f
C9000 C10_P_btm.n757 VSS 0.911266f
C9001 C10_P_btm.n758 VSS 0.911266f
C9002 C10_P_btm.n759 VSS 0.911266f
C9003 C10_P_btm.n760 VSS 0.911266f
C9004 C10_P_btm.n761 VSS 0.911266f
C9005 C10_P_btm.n762 VSS 2.05058f
C9006 C10_P_btm.n763 VSS 2.05058f
C9007 C10_P_btm.n764 VSS 3.9771f
C9008 C10_P_btm.n765 VSS 0.911266f
C9009 C10_P_btm.n766 VSS 0.911266f
C9010 C10_P_btm.n767 VSS 0.911266f
C9011 C10_P_btm.n768 VSS 1.16658f
C9012 C10_P_btm.n769 VSS 0.908087f
C9013 C10_P_btm.n770 VSS 0.908087f
C9014 C10_P_btm.n771 VSS 0.908087f
C9015 C10_P_btm.n772 VSS 0.911266f
C9016 C10_P_btm.n773 VSS 0.911266f
C9017 C10_P_btm.n774 VSS 0.911266f
C9018 C10_P_btm.n775 VSS 0.911266f
C9019 C10_P_btm.n776 VSS 0.908087f
C9020 C10_P_btm.n777 VSS 0.908087f
C9021 C10_P_btm.n778 VSS 0.908087f
C9022 C10_P_btm.n779 VSS 0.908087f
C9023 C10_P_btm.n780 VSS 0.911266f
C9024 C10_P_btm.n781 VSS 0.911266f
C9025 C10_P_btm.n782 VSS 0.911266f
C9026 C10_P_btm.n783 VSS 0.911266f
C9027 C10_P_btm.n784 VSS 0.908087f
C9028 C10_P_btm.n785 VSS 0.908087f
C9029 C10_P_btm.n786 VSS 0.908087f
C9030 C10_P_btm.n787 VSS 0.911266f
C9031 C10_P_btm.n788 VSS 0.911266f
C9032 C10_P_btm.n789 VSS 0.911266f
C9033 C10_P_btm.n790 VSS 0.911266f
C9034 C10_P_btm.n791 VSS 0.908087f
C9035 C10_P_btm.n792 VSS 0.908087f
C9036 C10_P_btm.n793 VSS 0.908087f
C9037 C10_P_btm.n794 VSS 0.908087f
C9038 C10_P_btm.n795 VSS 0.911266f
C9039 C10_P_btm.n796 VSS 0.911266f
C9040 C10_P_btm.n797 VSS 0.911266f
C9041 C10_P_btm.n798 VSS 0.911266f
C9042 C10_P_btm.n799 VSS 0.911266f
C9043 C10_P_btm.n800 VSS 0.911266f
C9044 C10_P_btm.n801 VSS 0.911266f
C9045 C10_P_btm.n802 VSS 0.911266f
C9046 C10_P_btm.n803 VSS 0.911266f
C9047 C10_P_btm.n804 VSS 0.911266f
C9048 C10_P_btm.n805 VSS 0.911266f
C9049 C10_P_btm.n806 VSS 0.911266f
C9050 C10_P_btm.n807 VSS 0.911266f
C9051 C10_P_btm.n808 VSS 0.911266f
C9052 C10_P_btm.n809 VSS 0.911266f
C9053 C10_P_btm.n810 VSS 0.911266f
C9054 C10_P_btm.n811 VSS 0.670504f
C9055 C10_P_btm.n812 VSS 0.670504f
C9056 C10_P_btm.n813 VSS 0.670504f
C9057 C10_P_btm.n814 VSS 0.911266f
C9058 C10_P_btm.n815 VSS 0.911266f
C9059 C10_P_btm.n816 VSS 0.911266f
C9060 C10_P_btm.n817 VSS 0.911266f
C9061 C10_P_btm.n818 VSS 0.911266f
C9062 C10_P_btm.n819 VSS 0.911266f
C9063 C10_P_btm.n820 VSS 0.911266f
C9064 C10_P_btm.n821 VSS 0.911266f
C9065 C10_P_btm.n822 VSS 1.14567f
C9066 C10_P_btm.n823 VSS 1.14567f
C9067 C10_P_btm.n824 VSS 1.14567f
C9068 C10_P_btm.n825 VSS 0.911266f
C9069 C10_P_btm.n826 VSS 0.911266f
C9070 C10_P_btm.n827 VSS 0.911266f
C9071 C10_P_btm.n828 VSS 0.911266f
C9072 C10_P_btm.n829 VSS 0.911266f
C9073 C10_P_btm.n830 VSS 0.911266f
C9074 C10_P_btm.n831 VSS 0.911266f
C9075 C10_P_btm.n832 VSS 0.911266f
C9076 C10_P_btm.n833 VSS 0.670504f
C9077 C10_P_btm.n834 VSS 0.670504f
C9078 C10_P_btm.n835 VSS 0.670504f
C9079 C10_P_btm.n836 VSS 0.911266f
C9080 C10_P_btm.n837 VSS 0.911266f
C9081 C10_P_btm.n838 VSS 0.911266f
C9082 C10_P_btm.n839 VSS 0.911266f
C9083 C10_P_btm.n840 VSS 0.911266f
C9084 C10_P_btm.n841 VSS 0.911266f
C9085 C10_P_btm.n842 VSS 0.911266f
C9086 C10_P_btm.n843 VSS 0.911266f
C9087 C10_P_btm.n844 VSS 1.14567f
C9088 C10_P_btm.n845 VSS 1.14567f
C9089 C10_P_btm.n846 VSS 0.911266f
C9090 C10_P_btm.n847 VSS 0.879698f
C9091 C10_P_btm.n848 VSS 0.911266f
C9092 C10_P_btm.n849 VSS 0.911266f
C9093 C10_P_btm.n850 VSS 1.14567f
C9094 C10_P_btm.n851 VSS 1.24398f
C9095 C10_P_btm.n852 VSS 0.911266f
C9096 C10_P_btm.n853 VSS 0.911266f
C9097 C10_P_btm.n854 VSS 0.911266f
C9098 C10_P_btm.n855 VSS 0.911266f
C9099 C10_P_btm.n856 VSS 0.911266f
C9100 C10_P_btm.n857 VSS 0.911266f
C9101 C10_P_btm.n858 VSS 0.911266f
C9102 C10_P_btm.n859 VSS 0.911266f
C9103 C10_P_btm.n860 VSS 0.911266f
C9104 C10_P_btm.n861 VSS 0.911266f
C9105 C10_P_btm.n862 VSS 2.22141f
C9106 C10_P_btm.n863 VSS 1.14567f
C9107 C10_P_btm.n864 VSS 1.14567f
C9108 C10_P_btm.n865 VSS 1.14567f
C9109 C10_P_btm.n866 VSS 0.911266f
C9110 C10_P_btm.n867 VSS 0.911266f
C9111 C10_P_btm.n868 VSS 0.911266f
C9112 C10_P_btm.n869 VSS 0.911266f
C9113 C10_P_btm.n870 VSS 0.911266f
C9114 C10_P_btm.n871 VSS 0.911266f
C9115 C10_P_btm.n872 VSS 0.911266f
C9116 C10_P_btm.n873 VSS 0.911266f
C9117 C10_P_btm.n874 VSS 0.911266f
C9118 C10_P_btm.n875 VSS 0.670504f
C9119 C10_P_btm.n876 VSS 0.670504f
C9120 C10_P_btm.n877 VSS 0.670504f
C9121 C10_P_btm.n878 VSS 0.670504f
C9122 C10_P_btm.n879 VSS 0.911266f
C9123 C10_P_btm.n880 VSS 0.911266f
C9124 C10_P_btm.n881 VSS 0.911266f
C9125 C10_P_btm.n882 VSS 0.911266f
C9126 C10_P_btm.n883 VSS 0.911266f
C9127 C10_P_btm.n884 VSS 0.911266f
C9128 C10_P_btm.n885 VSS 0.911266f
C9129 C10_P_btm.n886 VSS 1.14567f
C9130 C10_P_btm.n887 VSS 1.14567f
C9131 C10_P_btm.n888 VSS 1.14567f
C9132 C10_P_btm.n889 VSS 0.911266f
C9133 C10_P_btm.n890 VSS 0.911266f
C9134 C10_P_btm.n891 VSS 1.14567f
C9135 C10_P_btm.n892 VSS 0.911266f
C9136 C10_P_btm.n893 VSS 0.911266f
C9137 C10_P_btm.n894 VSS 0.911266f
C9138 C10_P_btm.n895 VSS 0.911266f
C9139 C10_P_btm.n896 VSS 0.911266f
C9140 C10_P_btm.n897 VSS 0.911266f
C9141 C10_P_btm.n898 VSS 0.911266f
C9142 C10_P_btm.n899 VSS 0.911266f
C9143 C10_P_btm.n900 VSS 1.14567f
C9144 C10_P_btm.n901 VSS 0.911266f
C9145 C10_P_btm.n902 VSS 1.14567f
C9146 C10_P_btm.n903 VSS 0.911266f
C9147 C10_P_btm.n904 VSS 0.911266f
C9148 C10_P_btm.n905 VSS 0.911266f
C9149 C10_P_btm.n906 VSS 0.911266f
C9150 C10_P_btm.n907 VSS 0.911266f
C9151 C10_P_btm.n908 VSS 0.911266f
C9152 C10_P_btm.n909 VSS 1.24386f
C9153 C10_P_btm.n910 VSS 0.911266f
C9154 C10_P_btm.n911 VSS 0.911266f
C9155 C10_P_btm.n912 VSS 0.911266f
C9156 C10_P_btm.n913 VSS 0.911266f
C9157 C10_P_btm.n914 VSS 1.14567f
C9158 C10_P_btm.n915 VSS 1.14567f
C9159 C10_P_btm.n916 VSS 1.14567f
C9160 C10_P_btm.n917 VSS 1.14567f
C9161 C10_P_btm.n918 VSS 0.911266f
C9162 C10_P_btm.n919 VSS 0.911266f
C9163 C10_P_btm.n920 VSS 0.911266f
C9164 C10_P_btm.n921 VSS 0.911266f
C9165 C10_P_btm.n922 VSS 0.911266f
C9166 C10_P_btm.n923 VSS 0.911266f
C9167 C10_P_btm.n924 VSS 0.911266f
C9168 C10_P_btm.n925 VSS 0.911266f
C9169 C10_P_btm.n926 VSS 0.911266f
C9170 C10_P_btm.n927 VSS 0.911266f
C9171 C10_P_btm.n928 VSS 0.911266f
C9172 C10_P_btm.n929 VSS 0.911266f
C9173 C10_P_btm.n930 VSS 0.911266f
C9174 C10_P_btm.n931 VSS 0.911266f
C9175 C10_P_btm.n932 VSS 0.911266f
C9176 C10_P_btm.n933 VSS 0.911266f
C9177 C10_P_btm.n934 VSS 1.14567f
C9178 C10_P_btm.n935 VSS 1.14567f
C9179 C10_P_btm.n936 VSS 1.14567f
C9180 C10_P_btm.n937 VSS 1.14567f
C9181 C10_P_btm.n938 VSS 0.911266f
C9182 C10_P_btm.n939 VSS 0.911266f
C9183 C10_P_btm.n940 VSS 0.911266f
C9184 C10_P_btm.n941 VSS 0.911266f
C9185 C10_P_btm.n942 VSS 0.911266f
C9186 C10_P_btm.n943 VSS 0.911266f
C9187 C10_P_btm.n944 VSS 0.911266f
C9188 C10_P_btm.n945 VSS 0.670504f
C9189 C10_P_btm.n946 VSS 0.670504f
C9190 C10_P_btm.n947 VSS 0.670504f
C9191 C10_P_btm.n948 VSS 0.670504f
C9192 C10_P_btm.n949 VSS 0.670504f
C9193 C10_P_btm.n950 VSS 0.670504f
C9194 C10_P_btm.n951 VSS 0.670504f
C9195 C10_P_btm.n952 VSS 0.670504f
C9196 C10_P_btm.n953 VSS 0.670504f
C9197 C10_P_btm.n954 VSS 0.670504f
C9198 C10_P_btm.n955 VSS 0.670504f
C9199 C10_P_btm.n956 VSS 0.670504f
C9200 C10_P_btm.n957 VSS 0.911266f
C9201 C10_P_btm.n958 VSS 0.911266f
C9202 C10_P_btm.n959 VSS 0.911266f
C9203 C10_P_btm.n960 VSS 0.911266f
C9204 C10_P_btm.n961 VSS 0.911266f
C9205 C10_P_btm.n962 VSS 0.911266f
C9206 C10_P_btm.n963 VSS 0.911266f
C9207 C10_P_btm.n964 VSS 0.911266f
C9208 C10_P_btm.n965 VSS 2.22148f
C9209 C10_P_btm.n966 VSS 1.14567f
C9210 C10_P_btm.n967 VSS 0.911266f
C9211 C10_P_btm.n968 VSS 1.14567f
C9212 C10_P_btm.n969 VSS 0.911266f
C9213 C10_P_btm.n970 VSS 0.911266f
C9214 C10_P_btm.n971 VSS 1.14567f
C9215 C10_P_btm.n972 VSS 1.14567f
C9216 C10_P_btm.n973 VSS 1.14567f
C9217 C10_P_btm.n974 VSS 0.911266f
C9218 C10_P_btm.n975 VSS 0.911266f
C9219 C10_P_btm.n976 VSS 0.911266f
C9220 C10_P_btm.n977 VSS 0.911266f
C9221 C10_P_btm.n978 VSS 0.911266f
C9222 C10_P_btm.n979 VSS 0.911266f
C9223 C10_P_btm.n980 VSS 0.911266f
C9224 C10_P_btm.n981 VSS 0.911266f
C9225 C10_P_btm.n982 VSS 0.911266f
C9226 C10_P_btm.n983 VSS 0.911266f
C9227 C10_P_btm.n984 VSS 0.911266f
C9228 C10_P_btm.n985 VSS 0.911266f
C9229 C10_P_btm.n986 VSS 1.14567f
C9230 C10_P_btm.n987 VSS 1.14567f
C9231 C10_P_btm.n988 VSS 1.14567f
C9232 C10_P_btm.n989 VSS 1.14567f
C9233 C10_P_btm.n990 VSS 0.911266f
C9234 C10_P_btm.n991 VSS 0.911266f
C9235 C10_P_btm.n992 VSS 0.911266f
C9236 C10_P_btm.n993 VSS 0.911266f
C9237 C10_P_btm.n994 VSS 0.911266f
C9238 C10_P_btm.n995 VSS 0.911266f
C9239 C10_P_btm.n996 VSS 0.911266f
C9240 C10_P_btm.n997 VSS 0.911266f
C9241 C10_P_btm.n998 VSS 0.911266f
C9242 C10_P_btm.n999 VSS 0.670504f
C9243 C10_P_btm.n1000 VSS 0.670504f
C9244 C10_P_btm.n1001 VSS 0.670504f
C9245 C10_P_btm.n1002 VSS 0.670504f
C9246 C10_P_btm.n1003 VSS 0.911266f
C9247 C10_P_btm.n1004 VSS 0.911266f
C9248 C10_P_btm.n1005 VSS 0.911266f
C9249 C10_P_btm.n1006 VSS 0.911266f
C9250 C10_P_btm.n1007 VSS 0.911266f
C9251 C10_P_btm.n1008 VSS 0.911266f
C9252 C10_P_btm.n1009 VSS 0.911266f
C9253 C10_P_btm.n1010 VSS 0.911266f
C9254 C10_P_btm.n1011 VSS 0.911266f
C9255 C10_P_btm.n1012 VSS 0.911266f
C9256 C10_P_btm.n1013 VSS 0.908087f
C9257 C10_P_btm.n1014 VSS 0.908087f
C9258 C10_P_btm.n1015 VSS 0.911266f
C9259 C10_P_btm.n1016 VSS 0.911266f
C9260 C10_P_btm.n1017 VSS 0.911266f
C9261 C10_P_btm.n1018 VSS 0.911266f
C9262 C10_P_btm.n1019 VSS 0.908087f
C9263 C10_P_btm.n1020 VSS 0.908087f
C9264 C10_P_btm.n1021 VSS 0.908087f
C9265 C10_P_btm.n1022 VSS 0.908087f
C9266 C10_P_btm.n1023 VSS 0.911266f
C9267 C10_P_btm.n1024 VSS 0.911266f
C9268 C10_P_btm.n1025 VSS 0.911266f
C9269 C10_P_btm.n1026 VSS 0.911266f
C9270 C10_P_btm.n1027 VSS 0.908087f
C9271 C10_P_btm.n1028 VSS 0.908087f
C9272 C10_P_btm.n1029 VSS 0.908087f
C9273 C10_P_btm.n1030 VSS 0.908087f
C9274 C10_P_btm.n1031 VSS 0.911266f
C9275 C10_P_btm.n1032 VSS 0.911266f
C9276 C10_P_btm.n1033 VSS 0.911266f
C9277 C10_P_btm.n1034 VSS 0.911266f
C9278 C10_P_btm.n1035 VSS 0.908087f
C9279 C10_P_btm.n1036 VSS 0.908087f
C9280 C10_P_btm.n1037 VSS 0.908087f
C9281 C10_P_btm.n1038 VSS 0.908087f
C9282 C10_P_btm.n1039 VSS 0.911266f
C9283 C10_P_btm.n1040 VSS 0.911266f
C9284 C10_P_btm.n1041 VSS 0.911266f
C9285 C10_P_btm.n1042 VSS 0.911266f
C9286 C10_P_btm.n1043 VSS 0.908087f
C9287 C10_P_btm.n1044 VSS 2.01139f
C9288 a_n4064_40160.t2 VSS 0.031188f
C9289 a_n4064_40160.t0 VSS 0.031188f
C9290 a_n4064_40160.t1 VSS 0.031188f
C9291 a_n4064_40160.n0 VSS 0.065553f
C9292 a_n4064_40160.t5 VSS 0.020272f
C9293 a_n4064_40160.t7 VSS 0.020272f
C9294 a_n4064_40160.n1 VSS 0.042018f
C9295 a_n4064_40160.t4 VSS 0.020272f
C9296 a_n4064_40160.t6 VSS 0.020272f
C9297 a_n4064_40160.n2 VSS 0.049863f
C9298 a_n4064_40160.n3 VSS 0.186059f
C9299 a_n4064_40160.t14 VSS 0.031826f
C9300 a_n4064_40160.t12 VSS 0.050682f
C9301 a_n4064_40160.n4 VSS 0.088983f
C9302 a_n4064_40160.n5 VSS 0.129407f
C9303 a_n4064_40160.t10 VSS 0.39598f
C9304 a_n4064_40160.t17 VSS 0.396982f
C9305 a_n4064_40160.t9 VSS 0.39598f
C9306 a_n4064_40160.t11 VSS 0.396982f
C9307 a_n4064_40160.t15 VSS 0.39598f
C9308 a_n4064_40160.t8 VSS 0.396982f
C9309 a_n4064_40160.n6 VSS 0.190289f
C9310 a_n4064_40160.t16 VSS 0.39598f
C9311 a_n4064_40160.n7 VSS 0.196709f
C9312 a_n4064_40160.n8 VSS 0.229488f
C9313 a_n4064_40160.n9 VSS 0.205528f
C9314 a_n4064_40160.n10 VSS 0.190289f
C9315 a_n4064_40160.n11 VSS 0.205528f
C9316 a_n4064_40160.n12 VSS 0.190289f
C9317 a_n4064_40160.t13 VSS 0.407333f
C9318 a_n4064_40160.n13 VSS 0.367847f
C9319 a_n4064_40160.n14 VSS 2.8676f
C9320 a_n4064_40160.n15 VSS 3.40691f
C9321 a_n4064_40160.n16 VSS 0.120772f
C9322 a_n4064_40160.n17 VSS 0.215941f
C9323 a_n4064_40160.n18 VSS 0.080373f
C9324 a_n4064_40160.t3 VSS 0.031188f
C9325 a_13467_32519.t0 VSS 0.058665f
C9326 a_13467_32519.t4 VSS 2.27165f
C9327 a_13467_32519.t2 VSS 0.038132f
C9328 a_13467_32519.t3 VSS 0.038132f
C9329 a_13467_32519.n0 VSS 0.076264f
C9330 a_13467_32519.n1 VSS 19.2825f
C9331 a_13467_32519.n2 VSS 0.176033f
C9332 a_13467_32519.t1 VSS 0.058665f
C9333 a_n3674_38680.t0 VSS 0.038341f
C9334 a_n3674_38680.t3 VSS 0.024921f
C9335 a_n3674_38680.t2 VSS 0.024921f
C9336 a_n3674_38680.n0 VSS 0.092296f
C9337 a_n3674_38680.t4 VSS 0.064051f
C9338 a_n3674_38680.t5 VSS 0.040114f
C9339 a_n3674_38680.n1 VSS 1.07573f
C9340 a_n3674_38680.n2 VSS 4.32458f
C9341 a_n3674_38680.n3 VSS 0.076712f
C9342 a_n3674_38680.t1 VSS 0.038341f
C9343 a_n4064_37984.t1 VSS 0.05638f
C9344 a_n4064_37984.t0 VSS 0.05638f
C9345 a_n4064_37984.t2 VSS 0.05638f
C9346 a_n4064_37984.n0 VSS 0.118503f
C9347 a_n4064_37984.t7 VSS 0.036647f
C9348 a_n4064_37984.t6 VSS 0.036647f
C9349 a_n4064_37984.n1 VSS 0.075958f
C9350 a_n4064_37984.t5 VSS 0.036647f
C9351 a_n4064_37984.t4 VSS 0.036647f
C9352 a_n4064_37984.n2 VSS 0.090139f
C9353 a_n4064_37984.n3 VSS 0.336347f
C9354 a_n4064_37984.t8 VSS 0.057533f
C9355 a_n4064_37984.t10 VSS 0.091621f
C9356 a_n4064_37984.n4 VSS 0.160859f
C9357 a_n4064_37984.t9 VSS 1.10909f
C9358 a_n4064_37984.n5 VSS 12.433901f
C9359 a_n4064_37984.n6 VSS 0.218325f
C9360 a_n4064_37984.n7 VSS 0.390366f
C9361 a_n4064_37984.n8 VSS 0.145294f
C9362 a_n4064_37984.t3 VSS 0.05638f
C9363 a_22612_30879.t6 VSS 0.544485f
C9364 a_22612_30879.t10 VSS 0.544569f
C9365 a_22612_30879.t8 VSS 0.544485f
C9366 a_22612_30879.n0 VSS 0.402155f
C9367 a_22612_30879.t16 VSS 0.544485f
C9368 a_22612_30879.n1 VSS 0.204694f
C9369 a_22612_30879.t14 VSS 0.544485f
C9370 a_22612_30879.n2 VSS 0.204694f
C9371 a_22612_30879.t4 VSS 0.544485f
C9372 a_22612_30879.n3 VSS 0.204694f
C9373 a_22612_30879.t11 VSS 0.544485f
C9374 a_22612_30879.n4 VSS 0.204694f
C9375 a_22612_30879.t17 VSS 0.544485f
C9376 a_22612_30879.n5 VSS 0.204694f
C9377 a_22612_30879.t7 VSS 0.544485f
C9378 a_22612_30879.n6 VSS 0.204694f
C9379 a_22612_30879.t15 VSS 0.544485f
C9380 a_22612_30879.n7 VSS 0.204694f
C9381 a_22612_30879.t19 VSS 0.544485f
C9382 a_22612_30879.n8 VSS 0.204694f
C9383 a_22612_30879.t12 VSS 0.544485f
C9384 a_22612_30879.n9 VSS 0.204694f
C9385 a_22612_30879.t9 VSS 0.544485f
C9386 a_22612_30879.n10 VSS 0.204694f
C9387 a_22612_30879.t13 VSS 0.544485f
C9388 a_22612_30879.n11 VSS 0.204694f
C9389 a_22612_30879.t18 VSS 0.544485f
C9390 a_22612_30879.n12 VSS 0.204694f
C9391 a_22612_30879.t5 VSS 0.544485f
C9392 a_22612_30879.n13 VSS 0.204301f
C9393 a_22612_30879.n14 VSS 2.25385f
C9394 a_22612_30879.t3 VSS 0.010456f
C9395 a_22612_30879.t2 VSS 0.010456f
C9396 a_22612_30879.n15 VSS 0.020912f
C9397 a_22612_30879.n16 VSS 1.74926f
C9398 a_22612_30879.t0 VSS 0.016086f
C9399 a_22612_30879.n17 VSS 0.048268f
C9400 a_22612_30879.t1 VSS 0.016086f
C9401 C7_P_btm.t3 VSS 0.15694f
C9402 C7_P_btm.t2 VSS 0.15694f
C9403 C7_P_btm.n0 VSS 0.933237f
C9404 C7_P_btm.t0 VSS 1.12025f
C9405 C7_P_btm.n1 VSS 2.0822f
C9406 C7_P_btm.t1 VSS 1.12621f
C9407 C7_P_btm.n2 VSS 1.11461f
C9408 C7_P_btm.t4 VSS 0.21231f
C9409 C7_P_btm.n3 VSS 2.69238f
C9410 a_5534_30871.t0 VSS 0.047423f
C9411 a_5534_30871.t7 VSS 0.046008f
C9412 a_5534_30871.t6 VSS 0.07377f
C9413 a_5534_30871.n0 VSS 0.231385f
C9414 a_5534_30871.t5 VSS 0.711036f
C9415 a_5534_30871.t4 VSS 0.713785f
C9416 a_5534_30871.n1 VSS 11.2661f
C9417 a_5534_30871.n2 VSS 6.98622f
C9418 a_5534_30871.t3 VSS 0.030825f
C9419 a_5534_30871.t2 VSS 0.030825f
C9420 a_5534_30871.n3 VSS 0.06165f
C9421 a_5534_30871.n4 VSS 0.611205f
C9422 a_5534_30871.n5 VSS 0.142301f
C9423 a_5534_30871.t1 VSS 0.047423f
C9424 a_6123_31319.t7 VSS 0.406419f
C9425 a_6123_31319.t4 VSS 0.379058f
C9426 a_6123_31319.n0 VSS 17.756401f
C9427 a_6123_31319.t5 VSS 0.090211f
C9428 a_6123_31319.t6 VSS 0.056261f
C9429 a_6123_31319.n1 VSS 0.212819f
C9430 a_6123_31319.n2 VSS 10.0411f
C9431 a_6123_31319.t2 VSS 0.037695f
C9432 a_6123_31319.t3 VSS 0.037695f
C9433 a_6123_31319.n3 VSS 0.075389f
C9434 a_6123_31319.n4 VSS 0.517004f
C9435 a_6123_31319.t0 VSS 0.057992f
C9436 a_6123_31319.n5 VSS 0.174014f
C9437 a_6123_31319.t1 VSS 0.057992f
C9438 a_n237_47217.t0 VSS 0.017838f
C9439 a_n237_47217.t5 VSS 0.027749f
C9440 a_n237_47217.t14 VSS 0.016352f
C9441 a_n237_47217.t6 VSS 0.027749f
C9442 a_n237_47217.t9 VSS 0.016352f
C9443 a_n237_47217.n0 VSS 0.046558f
C9444 a_n237_47217.n1 VSS 0.073165f
C9445 a_n237_47217.t7 VSS 0.018438f
C9446 a_n237_47217.t15 VSS 0.029529f
C9447 a_n237_47217.n2 VSS 0.05796f
C9448 a_n237_47217.t4 VSS 0.013443f
C9449 a_n237_47217.t8 VSS 0.019563f
C9450 a_n237_47217.n3 VSS 0.071214f
C9451 a_n237_47217.t10 VSS 0.01313f
C9452 a_n237_47217.t13 VSS 0.036091f
C9453 a_n237_47217.n4 VSS 0.107676f
C9454 a_n237_47217.t12 VSS 0.052102f
C9455 a_n237_47217.t11 VSS 0.027429f
C9456 a_n237_47217.n5 VSS 0.143667f
C9457 a_n237_47217.n6 VSS 1.54871f
C9458 a_n237_47217.n7 VSS 0.982282f
C9459 a_n237_47217.n8 VSS 0.266953f
C9460 a_n237_47217.n9 VSS 0.253519f
C9461 a_n237_47217.t3 VSS 0.011595f
C9462 a_n237_47217.t2 VSS 0.011595f
C9463 a_n237_47217.n10 VSS 0.02319f
C9464 a_n237_47217.n11 VSS 0.119003f
C9465 a_n237_47217.n12 VSS 0.049312f
C9466 a_n237_47217.t1 VSS 0.017838f
C9467 C0_P_btm.t0 VSS 1.3641f
C9468 C0_P_btm.t2 VSS 0.406352f
C9469 C0_P_btm.t1 VSS 0.273912f
C9470 C0_P_btm.n0 VSS 2.20629f
C9471 C0_P_btm.n1 VSS 3.34443f
C9472 C0_P_btm.t3 VSS 0.195052f
C9473 C0_P_btm.n2 VSS 3.77471f
C9474 a_n784_42308.t0 VSS 0.04459f
C9475 a_n784_42308.t6 VSS 0.279993f
C9476 a_n784_42308.t4 VSS 0.282765f
C9477 a_n784_42308.n0 VSS 13.8403f
C9478 a_n784_42308.t5 VSS 0.069363f
C9479 a_n784_42308.t7 VSS 0.043259f
C9480 a_n784_42308.n1 VSS 0.268838f
C9481 a_n784_42308.n2 VSS 9.314759f
C9482 a_n784_42308.t2 VSS 0.028983f
C9483 a_n784_42308.t3 VSS 0.028983f
C9484 a_n784_42308.n3 VSS 0.057967f
C9485 a_n784_42308.n4 VSS 0.461843f
C9486 a_n784_42308.n5 VSS 0.1338f
C9487 a_n784_42308.t1 VSS 0.04459f
C9488 a_4883_46098.t2 VSS 0.023367f
C9489 a_4883_46098.t6 VSS 0.034504f
C9490 a_4883_46098.n0 VSS 0.115993f
C9491 a_4883_46098.t8 VSS 0.023443f
C9492 a_4883_46098.t4 VSS 0.036737f
C9493 a_4883_46098.n1 VSS 0.134498f
C9494 a_4883_46098.t5 VSS 0.036737f
C9495 a_4883_46098.t3 VSS 0.023443f
C9496 a_4883_46098.n2 VSS 0.186466f
C9497 a_4883_46098.n3 VSS 4.20315f
C9498 a_4883_46098.t9 VSS 0.023851f
C9499 a_4883_46098.t7 VSS 0.043515f
C9500 a_4883_46098.n4 VSS 0.089775f
C9501 a_4883_46098.n5 VSS 4.7127f
C9502 a_4883_46098.n6 VSS 2.75627f
C9503 a_4883_46098.t1 VSS 0.059556f
C9504 a_4883_46098.n7 VSS 0.191111f
C9505 a_4883_46098.t0 VSS 0.104886f
C9506 a_n3565_38502.t4 VSS 0.031286f
C9507 a_n3565_38502.t6 VSS 0.031286f
C9508 a_n3565_38502.n0 VSS 0.119451f
C9509 a_n3565_38502.t5 VSS 0.031286f
C9510 a_n3565_38502.t7 VSS 0.031286f
C9511 a_n3565_38502.n1 VSS 0.071005f
C9512 a_n3565_38502.n2 VSS 0.343553f
C9513 a_n3565_38502.t8 VSS 0.081114f
C9514 a_n3565_38502.t9 VSS 0.050935f
C9515 a_n3565_38502.n3 VSS 0.128297f
C9516 a_n3565_38502.t10 VSS 1.52407f
C9517 a_n3565_38502.n4 VSS 9.105949f
C9518 a_n3565_38502.n5 VSS 0.198998f
C9519 a_n3565_38502.t0 VSS 0.048132f
C9520 a_n3565_38502.t2 VSS 0.048132f
C9521 a_n3565_38502.n6 VSS 0.099013f
C9522 a_n3565_38502.n7 VSS 0.437439f
C9523 a_n3565_38502.t1 VSS 0.048132f
C9524 a_n3565_38502.n8 VSS 0.122497f
C9525 a_n3565_38502.t3 VSS 0.048132f
C9526 a_2063_45854.t0 VSS 0.010096f
C9527 a_2063_45854.n0 VSS 0.023681f
C9528 a_2063_45854.t15 VSS 0.011072f
C9529 a_2063_45854.n1 VSS 0.039801f
C9530 a_2063_45854.t11 VSS 0.01044f
C9531 a_2063_45854.t7 VSS 0.016719f
C9532 a_2063_45854.n2 VSS 0.033687f
C9533 a_2063_45854.t4 VSS 0.016713f
C9534 a_2063_45854.t12 VSS 0.010435f
C9535 a_2063_45854.n3 VSS 0.033995f
C9536 a_2063_45854.n4 VSS 0.197778f
C9537 a_2063_45854.t16 VSS 0.016876f
C9538 a_2063_45854.t5 VSS 0.010571f
C9539 a_2063_45854.n5 VSS 0.031948f
C9540 a_2063_45854.n6 VSS 0.165042f
C9541 a_2063_45854.t9 VSS 0.010417f
C9542 a_2063_45854.t8 VSS 0.016691f
C9543 a_2063_45854.n7 VSS 0.037359f
C9544 a_2063_45854.n8 VSS 0.2501f
C9545 a_2063_45854.t10 VSS 0.020427f
C9546 a_2063_45854.n9 VSS 0.042576f
C9547 a_2063_45854.t14 VSS 0.020427f
C9548 a_2063_45854.n10 VSS 0.040582f
C9549 a_2063_45854.n11 VSS 1.15991f
C9550 a_2063_45854.n12 VSS 1.10829f
C9551 a_2063_45854.n13 VSS 0.138935f
C9552 a_2063_45854.n14 VSS 0.059541f
C9553 a_2063_45854.n15 VSS 0.020193f
C9554 a_2063_45854.t1 VSS 0.010096f
C9555 a_n2312_40392.t4 VSS 0.053743f
C9556 a_n2312_40392.t5 VSS 0.086151f
C9557 a_n2312_40392.n0 VSS 2.02155f
C9558 a_n2312_40392.t2 VSS 0.033914f
C9559 a_n2312_40392.t3 VSS 0.033914f
C9560 a_n2312_40392.n1 VSS 0.067827f
C9561 a_n2312_40392.n2 VSS 8.242f
C9562 a_n2312_40392.t0 VSS 0.052175f
C9563 a_n2312_40392.n3 VSS 0.156559f
C9564 a_n2312_40392.t1 VSS 0.052175f
C9565 a_11823_42460.t2 VSS 0.015083f
C9566 a_11823_42460.n0 VSS 0.037703f
C9567 a_11823_42460.n1 VSS 0.022401f
C9568 a_11823_42460.n2 VSS 0.124769f
C9569 a_11823_42460.t16 VSS 0.024865f
C9570 a_11823_42460.t17 VSS 0.057618f
C9571 a_11823_42460.t10 VSS 0.025418f
C9572 a_11823_42460.t19 VSS 0.015961f
C9573 a_11823_42460.n3 VSS 0.038504f
C9574 a_11823_42460.n4 VSS 0.516785f
C9575 a_11823_42460.t22 VSS 0.020441f
C9576 a_11823_42460.t23 VSS 0.013926f
C9577 a_11823_42460.n5 VSS 0.052259f
C9578 a_11823_42460.t25 VSS 0.022896f
C9579 a_11823_42460.t8 VSS 0.010857f
C9580 a_11823_42460.n6 VSS 0.092806f
C9581 a_11823_42460.n7 VSS 0.385222f
C9582 a_11823_42460.t15 VSS 0.013826f
C9583 a_11823_42460.t14 VSS 0.023462f
C9584 a_11823_42460.t12 VSS 0.013826f
C9585 a_11823_42460.t26 VSS 0.023462f
C9586 a_11823_42460.n8 VSS 0.039366f
C9587 a_11823_42460.n9 VSS 0.059333f
C9588 a_11823_42460.n10 VSS 0.094671f
C9589 a_11823_42460.n11 VSS 0.251805f
C9590 a_11823_42460.t11 VSS 0.025418f
C9591 a_11823_42460.t29 VSS 0.015961f
C9592 a_11823_42460.n12 VSS 0.041559f
C9593 a_11823_42460.t24 VSS 0.026126f
C9594 a_11823_42460.t27 VSS 0.015707f
C9595 a_11823_42460.n13 VSS 0.047099f
C9596 a_11823_42460.n14 VSS 0.471547f
C9597 a_11823_42460.n15 VSS 0.374582f
C9598 a_11823_42460.t18 VSS 0.013687f
C9599 a_11823_42460.t21 VSS 0.010347f
C9600 a_11823_42460.n16 VSS 0.034093f
C9601 a_11823_42460.t9 VSS 0.020441f
C9602 a_11823_42460.t28 VSS 0.013926f
C9603 a_11823_42460.n17 VSS 0.046271f
C9604 a_11823_42460.n18 VSS 0.210764f
C9605 a_11823_42460.n19 VSS 0.279369f
C9606 a_11823_42460.t20 VSS 0.015562f
C9607 a_11823_42460.t13 VSS 0.025119f
C9608 a_11823_42460.n20 VSS 0.052131f
C9609 a_11823_42460.n21 VSS 0.2678f
C9610 a_11823_42460.n22 VSS 0.103168f
C9611 a_11823_42460.t0 VSS 0.015083f
C9612 a_11823_42460.t1 VSS 0.015083f
C9613 a_11823_42460.n23 VSS 0.045801f
C9614 a_11823_42460.n24 VSS 0.128106f
C9615 a_11823_42460.n25 VSS 0.033686f
C9616 a_11823_42460.t3 VSS 0.015083f
C9617 a_9290_44172.n0 VSS 0.025625f
C9618 a_9290_44172.n1 VSS 0.021095f
C9619 a_9290_44172.n2 VSS 0.012533f
C9620 a_9290_44172.n3 VSS 0.069807f
C9621 a_9290_44172.t29 VSS 0.011327f
C9622 a_9290_44172.n4 VSS 0.029626f
C9623 a_9290_44172.t28 VSS 0.014106f
C9624 a_9290_44172.n5 VSS 0.027388f
C9625 a_9290_44172.t10 VSS 0.014054f
C9626 a_9290_44172.n6 VSS 0.029189f
C9627 a_9290_44172.t19 VSS 0.014221f
C9628 a_9290_44172.n7 VSS 0.022341f
C9629 a_9290_44172.t21 VSS 0.014221f
C9630 a_9290_44172.n8 VSS 0.021543f
C9631 a_9290_44172.t17 VSS 0.014221f
C9632 a_9290_44172.n9 VSS 0.022302f
C9633 a_9290_44172.n10 VSS 0.173727f
C9634 a_9290_44172.t11 VSS 0.014617f
C9635 a_9290_44172.n11 VSS 0.025352f
C9636 a_9290_44172.n12 VSS 0.172256f
C9637 a_9290_44172.t22 VSS 0.013127f
C9638 a_9290_44172.t25 VSS 0.013127f
C9639 a_9290_44172.n13 VSS 0.022025f
C9640 a_9290_44172.n14 VSS 0.046532f
C9641 a_9290_44172.t8 VSS 0.01281f
C9642 a_9290_44172.n15 VSS 0.047931f
C9643 a_9290_44172.n16 VSS 0.383849f
C9644 a_9290_44172.n17 VSS 0.222613f
C9645 a_9290_44172.n18 VSS 0.152659f
C9646 a_9290_44172.n19 VSS 0.035672f
C9647 a_9290_44172.n20 VSS 0.286132f
C9648 a_9290_44172.n21 VSS 0.048419f
C9649 a_9290_44172.n22 VSS 0.192731f
C9650 a_9290_44172.n23 VSS 0.159155f
C9651 a_9290_44172.n24 VSS 0.071641f
C9652 a_9290_44172.n25 VSS 0.071674f
C9653 a_9290_44172.n26 VSS 0.018847f
C9654 a_3483_46348.t6 VSS 0.010046f
C9655 a_3483_46348.n0 VSS 0.022168f
C9656 a_3483_46348.t9 VSS 0.01006f
C9657 a_3483_46348.n1 VSS 0.015046f
C9658 a_3483_46348.t20 VSS 0.010091f
C9659 a_3483_46348.n2 VSS 0.019803f
C9660 a_3483_46348.t11 VSS 0.010091f
C9661 a_3483_46348.n3 VSS 0.016406f
C9662 a_3483_46348.t16 VSS 0.012523f
C9663 a_3483_46348.n4 VSS 0.020823f
C9664 a_3483_46348.t22 VSS 0.012523f
C9665 a_3483_46348.n5 VSS 0.012621f
C9666 a_3483_46348.n6 VSS 0.248134f
C9667 a_3483_46348.t18 VSS 0.012523f
C9668 a_3483_46348.n7 VSS 0.012621f
C9669 a_3483_46348.n8 VSS 0.092639f
C9670 a_3483_46348.n9 VSS 0.198183f
C9671 a_3483_46348.n10 VSS 0.019472f
C9672 a_3483_46348.n11 VSS 0.233929f
C9673 a_3483_46348.n12 VSS 0.145679f
C9674 a_3483_46348.t7 VSS 0.010091f
C9675 a_3483_46348.n13 VSS 0.01522f
C9676 a_3483_46348.n14 VSS 0.112026f
C9677 a_3483_46348.n15 VSS 0.01827f
C9678 a_3483_46348.n16 VSS 0.226019f
C9679 a_3483_46348.n17 VSS 0.388552f
C9680 a_3483_46348.n18 VSS 0.223826f
C9681 a_3483_46348.n20 VSS 0.042764f
C9682 a_3483_46348.n21 VSS 0.017967f
C9683 a_10903_43370.t0 VSS 0.010526f
C9684 a_10903_43370.n0 VSS 0.029519f
C9685 a_10903_43370.t23 VSS 0.01088f
C9686 a_10903_43370.t15 VSS 0.017425f
C9687 a_10903_43370.n1 VSS 0.035368f
C9688 a_10903_43370.t4 VSS 0.017739f
C9689 a_10903_43370.t20 VSS 0.011139f
C9690 a_10903_43370.n2 VSS 0.042828f
C9691 a_10903_43370.t17 VSS 0.011022f
C9692 a_10903_43370.t19 VSS 0.017595f
C9693 a_10903_43370.n3 VSS 0.02946f
C9694 a_10903_43370.n4 VSS 0.354745f
C9695 a_10903_43370.n5 VSS 0.02859f
C9696 a_10903_43370.t8 VSS 0.017739f
C9697 a_10903_43370.t12 VSS 0.011139f
C9698 a_10903_43370.n6 VSS 0.03744f
C9699 a_10903_43370.n7 VSS 0.286184f
C9700 a_10903_43370.n8 VSS 0.074001f
C9701 a_10903_43370.t11 VSS 0.014064f
C9702 a_10903_43370.n9 VSS 0.038931f
C9703 a_10903_43370.n10 VSS 0.181184f
C9704 a_10903_43370.t16 VSS 0.017437f
C9705 a_10903_43370.t5 VSS 0.01089f
C9706 a_10903_43370.n11 VSS 0.042635f
C9707 a_10903_43370.n12 VSS 0.231089f
C9708 a_10903_43370.n13 VSS 0.10711f
C9709 a_10903_43370.t6 VSS 0.017739f
C9710 a_10903_43370.t14 VSS 0.011139f
C9711 a_10903_43370.n14 VSS 0.032605f
C9712 a_10903_43370.t18 VSS 0.014266f
C9713 a_10903_43370.n15 VSS 0.037096f
C9714 a_10903_43370.n16 VSS 0.249549f
C9715 a_10903_43370.t13 VSS 0.014266f
C9716 a_10903_43370.n17 VSS 0.034204f
C9717 a_10903_43370.n18 VSS 0.151966f
C9718 a_10903_43370.n19 VSS 0.164325f
C9719 a_10903_43370.n20 VSS 0.102169f
C9720 a_10903_43370.n21 VSS 0.021092f
C9721 a_10903_43370.t1 VSS 0.010526f
C9722 a_18184_42460.t2 VSS 0.010407f
C9723 a_18184_42460.t1 VSS 0.057251f
C9724 a_18184_42460.t3 VSS 0.016943f
C9725 a_18184_42460.t5 VSS 0.026982f
C9726 a_18184_42460.n0 VSS 0.046225f
C9727 a_18184_42460.t7 VSS 0.026982f
C9728 a_18184_42460.t8 VSS 0.016943f
C9729 a_18184_42460.n1 VSS 0.078436f
C9730 a_18184_42460.t4 VSS 0.016519f
C9731 a_18184_42460.t6 VSS 0.026665f
C9732 a_18184_42460.n2 VSS 0.081152f
C9733 a_18184_42460.n3 VSS 0.98006f
C9734 a_18184_42460.n4 VSS 0.41829f
C9735 a_18184_42460.n5 VSS 0.232974f
C9736 a_18184_42460.n6 VSS 0.053761f
C9737 a_18184_42460.t0 VSS 0.010407f
C9738 a_5891_43370.n0 VSS 0.022129f
C9739 a_5891_43370.n1 VSS 0.013148f
C9740 a_5891_43370.n2 VSS 0.057903f
C9741 a_5891_43370.t18 VSS 0.014797f
C9742 a_5891_43370.n3 VSS 0.03246f
C9743 a_5891_43370.n4 VSS 0.027286f
C9744 a_5891_43370.t16 VSS 0.014743f
C9745 a_5891_43370.n5 VSS 0.032111f
C9746 a_5891_43370.t23 VSS 0.014635f
C9747 a_5891_43370.n6 VSS 0.032496f
C9748 a_5891_43370.t15 VSS 0.015332f
C9749 a_5891_43370.n7 VSS 0.027933f
C9750 a_5891_43370.n8 VSS 0.16771f
C9751 a_5891_43370.t11 VSS 0.014919f
C9752 a_5891_43370.n9 VSS 0.021192f
C9753 a_5891_43370.n10 VSS 0.15574f
C9754 a_5891_43370.n11 VSS 0.171802f
C9755 a_5891_43370.n12 VSS 0.179308f
C9756 a_5891_43370.n13 VSS 0.01973f
C9757 a_5891_43370.n14 VSS 0.121979f
C9758 a_5891_43370.n15 VSS 0.033492f
C9759 a_5891_43370.n16 VSS 0.150438f
C9760 a_5891_43370.n17 VSS 0.022885f
C9761 a_5891_43370.n18 VSS 0.173109f
C9762 a_5891_43370.n19 VSS 0.232398f
C9763 a_5891_43370.n20 VSS 0.037611f
C9764 a_5891_43370.n21 VSS 0.019771f
C9765 a_5891_43370.n22 VSS 0.089402f
C9766 a_5891_43370.n23 VSS 0.026882f
C9767 a_15493_43396.t1 VSS 0.106935f
C9768 a_15493_43396.t2 VSS 0.029253f
C9769 a_15493_43396.t3 VSS 0.023425f
C9770 a_15493_43396.n0 VSS 0.272145f
C9771 a_15493_43396.n1 VSS 1.75455f
C9772 a_15493_43396.t0 VSS 0.113691f
C9773 a_n2438_43548.t9 VSS 0.010683f
C9774 a_n2438_43548.t2 VSS 0.010683f
C9775 a_n2438_43548.t7 VSS 0.010683f
C9776 a_n2438_43548.n0 VSS 0.022518f
C9777 a_n2438_43548.t5 VSS 0.010683f
C9778 a_n2438_43548.t0 VSS 0.010683f
C9779 a_n2438_43548.n1 VSS 0.022225f
C9780 a_n2438_43548.n2 VSS 0.015932f
C9781 a_n2438_43548.n3 VSS 0.010243f
C9782 a_n2438_43548.n4 VSS 0.06472f
C9783 a_n2438_43548.n5 VSS 0.010243f
C9784 a_n2438_43548.n6 VSS 0.038902f
C9785 a_n2438_43548.n7 VSS 0.010249f
C9786 a_n2438_43548.n8 VSS 0.040128f
C9787 a_n2438_43548.n9 VSS 0.010243f
C9788 a_n2438_43548.n10 VSS 0.038902f
C9789 a_n2438_43548.n11 VSS 0.010243f
C9790 a_n2438_43548.n12 VSS 0.039096f
C9791 a_n2438_43548.n13 VSS 0.010243f
C9792 a_n2438_43548.n14 VSS 0.033583f
C9793 a_n2438_43548.n16 VSS 0.104217f
C9794 a_n2438_43548.n17 VSS 0.125472f
C9795 a_n2438_43548.n18 VSS 0.050772f
C9796 a_n2438_43548.t34 VSS 0.016721f
C9797 a_n2438_43548.t32 VSS 0.011188f
C9798 a_n2438_43548.n19 VSS 0.036537f
C9799 a_n2438_43548.t35 VSS 0.011188f
C9800 a_n2438_43548.t43 VSS 0.016721f
C9801 a_n2438_43548.n20 VSS 0.034959f
C9802 a_n2438_43548.t38 VSS 0.016721f
C9803 a_n2438_43548.t45 VSS 0.011188f
C9804 a_n2438_43548.n21 VSS 0.036185f
C9805 a_n2438_43548.n22 VSS 0.220257f
C9806 a_n2438_43548.t39 VSS 0.011188f
C9807 a_n2438_43548.t42 VSS 0.016721f
C9808 a_n2438_43548.n23 VSS 0.034279f
C9809 a_n2438_43548.n24 VSS 0.121158f
C9810 a_n2438_43548.t44 VSS 0.016721f
C9811 a_n2438_43548.t41 VSS 0.011188f
C9812 a_n2438_43548.n25 VSS 0.036185f
C9813 a_n2438_43548.n26 VSS 0.197022f
C9814 a_n2438_43548.t36 VSS 0.011188f
C9815 a_n2438_43548.t40 VSS 0.016721f
C9816 a_n2438_43548.n27 VSS 0.033839f
C9817 a_n2438_43548.n28 VSS 0.265675f
C9818 a_n2438_43548.t33 VSS 0.016721f
C9819 a_n2438_43548.t37 VSS 0.011188f
C9820 a_n2438_43548.n29 VSS 0.033932f
C9821 a_n2438_43548.n30 VSS 0.278153f
C9822 a_n2438_43548.n31 VSS 0.438366f
C9823 a_n2438_43548.t1 VSS 0.010683f
C9824 a_n2438_43548.t4 VSS 0.010683f
C9825 a_n2438_43548.n32 VSS 0.021365f
C9826 a_n2438_43548.n33 VSS 0.07388f
C9827 a_n2438_43548.n34 VSS 0.035618f
C9828 a_n2438_43548.t12 VSS 0.010683f
C9829 a_n2438_43548.t8 VSS 0.010683f
C9830 a_n2438_43548.n35 VSS 0.022518f
C9831 a_n2438_43548.n36 VSS 0.058839f
C9832 a_n2438_43548.t3 VSS 0.010683f
C9833 a_n2438_43548.t10 VSS 0.010683f
C9834 a_n2438_43548.n37 VSS 0.022518f
C9835 a_n2438_43548.n38 VSS 0.058839f
C9836 a_n2438_43548.t14 VSS 0.010683f
C9837 a_n2438_43548.t6 VSS 0.010683f
C9838 a_n2438_43548.n39 VSS 0.022518f
C9839 a_n2438_43548.n40 VSS 0.059113f
C9840 a_n2438_43548.t11 VSS 0.010683f
C9841 a_n2438_43548.t13 VSS 0.010683f
C9842 a_n2438_43548.n41 VSS 0.027137f
C9843 a_n2438_43548.n42 VSS 0.10262f
C9844 a_n2438_43548.n43 VSS 0.022518f
C9845 a_n2438_43548.t15 VSS 0.010683f
C9846 a_3090_45724.t0 VSS 0.016601f
C9847 a_3090_45724.t3 VSS 0.02029f
C9848 a_3090_45724.t2 VSS 0.02029f
C9849 a_3090_45724.n0 VSS 0.043668f
C9850 a_3090_45724.t4 VSS 0.01079f
C9851 a_3090_45724.t5 VSS 0.01079f
C9852 a_3090_45724.n1 VSS 0.021846f
C9853 a_3090_45724.t10 VSS 0.015328f
C9854 a_3090_45724.t17 VSS 0.012219f
C9855 a_3090_45724.n2 VSS 0.058703f
C9856 a_3090_45724.t18 VSS 0.027509f
C9857 a_3090_45724.t13 VSS 0.017182f
C9858 a_3090_45724.n3 VSS 0.060665f
C9859 a_3090_45724.t7 VSS 0.017382f
C9860 a_3090_45724.t19 VSS 0.027749f
C9861 a_3090_45724.n4 VSS 0.05631f
C9862 a_3090_45724.t16 VSS 0.017217f
C9863 a_3090_45724.t15 VSS 0.027551f
C9864 a_3090_45724.n5 VSS 0.052589f
C9865 a_3090_45724.t11 VSS 0.027509f
C9866 a_3090_45724.t9 VSS 0.017182f
C9867 a_3090_45724.n6 VSS 0.080821f
C9868 a_3090_45724.t21 VSS 0.02749f
C9869 a_3090_45724.t12 VSS 0.017166f
C9870 a_3090_45724.n7 VSS 0.055226f
C9871 a_3090_45724.n8 VSS 0.849085f
C9872 a_3090_45724.n9 VSS 0.456865f
C9873 a_3090_45724.t8 VSS 0.017182f
C9874 a_3090_45724.t14 VSS 0.027509f
C9875 a_3090_45724.n10 VSS 0.058968f
C9876 a_3090_45724.n11 VSS 1.96205f
C9877 a_3090_45724.n12 VSS 1.92093f
C9878 a_3090_45724.n13 VSS 1.74078f
C9879 a_3090_45724.t20 VSS 0.027976f
C9880 a_3090_45724.t6 VSS 0.017567f
C9881 a_3090_45724.n14 VSS 0.039369f
C9882 a_3090_45724.n15 VSS 0.550891f
C9883 a_3090_45724.n16 VSS 0.576918f
C9884 a_3090_45724.n17 VSS 0.048799f
C9885 a_3090_45724.n18 VSS 0.180842f
C9886 a_3090_45724.n19 VSS 0.047587f
C9887 a_3090_45724.t1 VSS 0.016601f
C9888 a_11206_38545.t4 VSS 0.031106f
C9889 a_11206_38545.t3 VSS 1.21993f
C9890 a_11206_38545.t2 VSS 1.02548f
C9891 a_11206_38545.n0 VSS 2.85069f
C9892 a_11206_38545.t1 VSS 1.02548f
C9893 a_11206_38545.n1 VSS 2.55854f
C9894 a_11206_38545.n2 VSS 0.157657f
C9895 a_11206_38545.t0 VSS 0.031106f
C9896 a_7754_40130.n0 VSS 0.11668f
C9897 a_7754_40130.n1 VSS 0.230022f
C9898 a_7754_40130.n2 VSS 0.230022f
C9899 a_7754_40130.n3 VSS 0.436037f
C9900 a_7754_40130.t12 VSS 0.441623f
C9901 a_7754_40130.t6 VSS 0.44132f
C9902 a_7754_40130.n4 VSS 0.436037f
C9903 a_7754_40130.n5 VSS 0.230022f
C9904 a_7754_40130.t7 VSS 0.44132f
C9905 a_7754_40130.n6 VSS 0.230022f
C9906 a_7754_40130.t5 VSS 0.44132f
C9907 a_7754_40130.n7 VSS 0.230022f
C9908 a_7754_40130.n8 VSS 0.230022f
C9909 a_7754_40130.t15 VSS 0.44132f
C9910 a_7754_40130.n9 VSS 0.230022f
C9911 a_7754_40130.t10 VSS 0.44132f
C9912 a_7754_40130.n10 VSS 0.230022f
C9913 a_7754_40130.n11 VSS 0.199574f
C9914 a_7754_40130.t0 VSS 0.44132f
C9915 a_7754_40130.n12 VSS 0.199574f
C9916 a_7754_40130.n13 VSS 0.230022f
C9917 a_7754_40130.n14 VSS 0.230022f
C9918 a_7754_40130.t11 VSS 0.441479f
C9919 a_7754_40130.t3 VSS 0.077849f
C9920 a_7754_40130.t2 VSS 0.04413f
C9921 a_7754_40130.n15 VSS 0.926275f
C9922 a_7754_40130.n16 VSS 0.361406f
C9923 a_7754_40130.n17 VSS 0.22704f
C9924 a_7754_40130.t9 VSS 0.44132f
C9925 a_7754_40130.n18 VSS 0.434782f
C9926 a_7754_40130.t13 VSS 0.44132f
C9927 a_7754_40130.n19 VSS 0.230022f
C9928 a_7754_40130.n20 VSS 0.230022f
C9929 a_7754_40130.t4 VSS 0.44132f
C9930 a_7754_40130.n21 VSS 0.230022f
C9931 a_7754_40130.t14 VSS 0.44132f
C9932 a_7754_40130.n22 VSS 0.230022f
C9933 a_7754_40130.n23 VSS 0.21778f
C9934 a_7754_40130.t8 VSS 0.44132f
C9935 a_7754_40130.n24 VSS 0.21778f
C9936 a_7754_40130.n25 VSS 0.116902f
C9937 a_7754_40130.n26 VSS 0.396147f
C9938 a_7754_40130.t1 VSS 0.33407f
C9939 a_10227_46804.n0 VSS 0.016334f
C9940 a_10227_46804.n1 VSS 0.015293f
C9941 a_10227_46804.n2 VSS 0.175875f
C9942 a_10227_46804.n3 VSS 0.014827f
C9943 a_10227_46804.n4 VSS 0.234326f
C9944 a_10227_46804.n5 VSS 0.01594f
C9945 a_10227_46804.n6 VSS 0.015476f
C9946 a_10227_46804.n7 VSS 0.163436f
C9947 a_10227_46804.n8 VSS 0.01594f
C9948 a_10227_46804.n9 VSS 0.015476f
C9949 a_10227_46804.n10 VSS 0.132924f
C9950 a_10227_46804.n11 VSS 0.326035f
C9951 a_10227_46804.n12 VSS 0.015823f
C9952 a_10227_46804.n13 VSS 0.01548f
C9953 a_10227_46804.n14 VSS 0.090662f
C9954 a_10227_46804.n15 VSS 0.015291f
C9955 a_10227_46804.n16 VSS 0.016361f
C9956 a_10227_46804.n17 VSS 0.085253f
C9957 a_10227_46804.n18 VSS 0.015913f
C9958 a_10227_46804.n19 VSS 0.015484f
C9959 a_10227_46804.n20 VSS 0.253005f
C9960 a_10227_46804.n21 VSS 0.189655f
C9961 a_10227_46804.n22 VSS 0.136777f
C9962 a_10227_46804.n23 VSS 0.01594f
C9963 a_10227_46804.n24 VSS 0.015476f
C9964 a_10227_46804.n25 VSS 0.089585f
C9965 a_10227_46804.n26 VSS 0.09486f
C9966 a_10227_46804.n27 VSS 0.225422f
C9967 a_10227_46804.n28 VSS 0.106723f
C9968 a_10227_46804.n30 VSS 0.033964f
C9969 a_10227_46804.n31 VSS 0.016099f
C9970 C6_P_btm.t2 VSS 1.67804f
C9971 C6_P_btm.t3 VSS 0.051941f
C9972 C6_P_btm.t4 VSS 0.051941f
C9973 C6_P_btm.n0 VSS 0.138138f
C9974 C6_P_btm.t1 VSS 0.051941f
C9975 C6_P_btm.t0 VSS 0.051941f
C9976 C6_P_btm.n1 VSS 0.247039f
C9977 C6_P_btm.n2 VSS 1.35068f
C9978 C6_P_btm.n3 VSS 2.10571f
C9979 C6_P_btm.t5 VSS 0.120999f
C9980 C6_P_btm.n4 VSS 2.99527f
C9981 a_n3565_39304.t1 VSS 0.043965f
C9982 a_n3565_39304.t4 VSS 0.028577f
C9983 a_n3565_39304.t7 VSS 0.028577f
C9984 a_n3565_39304.n0 VSS 0.109108f
C9985 a_n3565_39304.t5 VSS 0.028577f
C9986 a_n3565_39304.t6 VSS 0.028577f
C9987 a_n3565_39304.n1 VSS 0.064856f
C9988 a_n3565_39304.n2 VSS 0.313806f
C9989 a_n3565_39304.t9 VSS 0.046525f
C9990 a_n3565_39304.t10 VSS 0.074091f
C9991 a_n3565_39304.n3 VSS 0.118665f
C9992 a_n3565_39304.t8 VSS 1.91876f
C9993 a_n3565_39304.n4 VSS 8.88085f
C9994 a_n3565_39304.n5 VSS 0.181275f
C9995 a_n3565_39304.t2 VSS 0.043965f
C9996 a_n3565_39304.t0 VSS 0.043965f
C9997 a_n3565_39304.n6 VSS 0.09044f
C9998 a_n3565_39304.n7 VSS 0.399563f
C9999 a_n3565_39304.n8 VSS 0.111891f
C10000 a_n3565_39304.t3 VSS 0.043965f
C10001 a_n4064_39072.t1 VSS 0.042953f
C10002 a_n4064_39072.t5 VSS 0.027919f
C10003 a_n4064_39072.t4 VSS 0.027919f
C10004 a_n4064_39072.n0 VSS 0.057867f
C10005 a_n4064_39072.t7 VSS 0.027919f
C10006 a_n4064_39072.t6 VSS 0.027919f
C10007 a_n4064_39072.n1 VSS 0.068671f
C10008 a_n4064_39072.n2 VSS 0.256241f
C10009 a_n4064_39072.t10 VSS 0.04383f
C10010 a_n4064_39072.t8 VSS 0.0698f
C10011 a_n4064_39072.n3 VSS 0.122548f
C10012 a_n4064_39072.t9 VSS 0.819006f
C10013 a_n4064_39072.n4 VSS 8.813861f
C10014 a_n4064_39072.n5 VSS 0.166328f
C10015 a_n4064_39072.t2 VSS 0.042953f
C10016 a_n4064_39072.t0 VSS 0.042953f
C10017 a_n4064_39072.n6 VSS 0.11069f
C10018 a_n4064_39072.n7 VSS 0.297395f
C10019 a_n4064_39072.n8 VSS 0.09028f
C10020 a_n4064_39072.t3 VSS 0.042953f
C10021 a_n3674_37592.t4 VSS 0.023944f
C10022 a_n3674_37592.t5 VSS 0.014996f
C10023 a_n3674_37592.n0 VSS 0.464718f
C10024 a_n3674_37592.n1 VSS 0.018633f
C10025 a_n3674_37592.n2 VSS 2.4874f
C10026 a_n3674_37592.t0 VSS 0.014333f
C10027 a_n3674_37592.n3 VSS 0.043008f
C10028 a_n3674_37592.t1 VSS 0.014333f
C10029 a_n2017_45002.t0 VSS 0.03412f
C10030 a_n2017_45002.t2 VSS 0.022178f
C10031 a_n2017_45002.t3 VSS 0.022178f
C10032 a_n2017_45002.n0 VSS 0.071202f
C10033 a_n2017_45002.t5 VSS 0.033102f
C10034 a_n2017_45002.t4 VSS 0.053077f
C10035 a_n2017_45002.n1 VSS 3.40334f
C10036 a_n2017_45002.n2 VSS 14.1582f
C10037 a_n2017_45002.n3 VSS 0.068512f
C10038 a_n2017_45002.t1 VSS 0.03412f
C10039 a_6171_45002.t1 VSS 0.058026f
C10040 a_6171_45002.n0 VSS 0.093334f
C10041 a_6171_45002.t4 VSS 0.019345f
C10042 a_6171_45002.t2 VSS 0.030807f
C10043 a_6171_45002.n1 VSS 0.077327f
C10044 a_6171_45002.t3 VSS 0.030222f
C10045 a_6171_45002.t5 VSS 0.018861f
C10046 a_6171_45002.n2 VSS 0.069678f
C10047 a_6171_45002.n3 VSS 4.40008f
C10048 a_6171_45002.n4 VSS 0.238394f
C10049 a_6171_45002.t0 VSS 0.06393f
C10050 a_13258_32519.t2 VSS 0.024064f
C10051 a_13258_32519.t3 VSS 0.024064f
C10052 a_13258_32519.n0 VSS 0.089119f
C10053 a_13258_32519.t4 VSS 1.72561f
C10054 a_13258_32519.n1 VSS 12.189f
C10055 a_13258_32519.t0 VSS 0.037021f
C10056 a_13258_32519.n2 VSS 0.074072f
C10057 a_13258_32519.t1 VSS 0.037021f
C10058 a_n97_42460.t7 VSS 0.013459f
C10059 a_n97_42460.n0 VSS 0.021686f
C10060 a_n97_42460.t10 VSS 0.013459f
C10061 a_n97_42460.n1 VSS 0.021443f
C10062 a_n97_42460.t22 VSS 0.013459f
C10063 a_n97_42460.n2 VSS 0.026011f
C10064 a_n97_42460.t20 VSS 0.01328f
C10065 a_n97_42460.n3 VSS 0.0286f
C10066 a_n97_42460.n4 VSS 0.226253f
C10067 a_n97_42460.t21 VSS 0.013459f
C10068 a_n97_42460.n5 VSS 0.021658f
C10069 a_n97_42460.n6 VSS 0.349093f
C10070 a_n97_42460.t18 VSS 0.013459f
C10071 a_n97_42460.n7 VSS 0.020575f
C10072 a_n97_42460.n8 VSS 0.415646f
C10073 a_n97_42460.n9 VSS 0.235886f
C10074 a_n97_42460.t5 VSS 0.013459f
C10075 a_n97_42460.n10 VSS 0.024127f
C10076 a_n97_42460.n11 VSS 0.303952f
C10077 a_n97_42460.t8 VSS 0.013459f
C10078 a_n97_42460.n12 VSS 0.024127f
C10079 a_n97_42460.n13 VSS 0.251521f
C10080 a_n97_42460.n14 VSS 0.289149f
C10081 a_n97_42460.t23 VSS 0.013459f
C10082 a_n97_42460.n15 VSS 0.021853f
C10083 a_n97_42460.t17 VSS 0.01328f
C10084 a_n97_42460.n16 VSS 0.025154f
C10085 a_n97_42460.n17 VSS 0.126177f
C10086 a_n97_42460.n18 VSS 0.679265f
C10087 a_n97_42460.n19 VSS 0.010414f
C10088 a_n97_42460.n20 VSS 0.208562f
C10089 a_n97_42460.n21 VSS 0.024038f
C10090 a_n2956_39768.t0 VSS 0.058317f
C10091 a_n2956_39768.t3 VSS 0.037906f
C10092 a_n2956_39768.t2 VSS 0.037906f
C10093 a_n2956_39768.n0 VSS 0.140383f
C10094 a_n2956_39768.t5 VSS 0.096293f
C10095 a_n2956_39768.t4 VSS 0.060069f
C10096 a_n2956_39768.n1 VSS 2.65786f
C10097 a_n2956_39768.n2 VSS 9.13627f
C10098 a_n2956_39768.n3 VSS 0.11668f
C10099 a_n2956_39768.t1 VSS 0.058317f
C10100 a_13747_46662.t2 VSS 0.018356f
C10101 a_13747_46662.t1 VSS 0.060727f
C10102 a_13747_46662.t8 VSS 0.018981f
C10103 a_13747_46662.t10 VSS 0.030397f
C10104 a_13747_46662.n0 VSS 0.060283f
C10105 a_13747_46662.t5 VSS 0.016826f
C10106 a_13747_46662.t4 VSS 0.028554f
C10107 a_13747_46662.t11 VSS 0.016826f
C10108 a_13747_46662.t3 VSS 0.028554f
C10109 a_13747_46662.n1 VSS 0.04791f
C10110 a_13747_46662.n2 VSS 0.110701f
C10111 a_13747_46662.n3 VSS 0.822651f
C10112 a_13747_46662.t6 VSS 0.030628f
C10113 a_13747_46662.t12 VSS 0.016788f
C10114 a_13747_46662.n4 VSS 0.059578f
C10115 a_13747_46662.t9 VSS 0.020426f
C10116 a_13747_46662.t7 VSS 0.014064f
C10117 a_13747_46662.n5 VSS 0.072355f
C10118 a_13747_46662.n6 VSS 0.950898f
C10119 a_13747_46662.n7 VSS 0.832316f
C10120 a_13747_46662.n8 VSS 0.378621f
C10121 a_13747_46662.n9 VSS 0.045204f
C10122 a_13747_46662.t0 VSS 0.018356f
C10123 a_n4209_38216.t2 VSS 0.047234f
C10124 a_n4209_38216.t6 VSS 0.030702f
C10125 a_n4209_38216.t4 VSS 0.030702f
C10126 a_n4209_38216.n0 VSS 0.117223f
C10127 a_n4209_38216.t5 VSS 0.030702f
C10128 a_n4209_38216.t7 VSS 0.030702f
C10129 a_n4209_38216.n1 VSS 0.06968f
C10130 a_n4209_38216.n2 VSS 0.377154f
C10131 a_n4209_38216.t9 VSS 0.049985f
C10132 a_n4209_38216.t8 VSS 0.079601f
C10133 a_n4209_38216.n3 VSS 0.169374f
C10134 a_n4209_38216.t10 VSS 1.43719f
C10135 a_n4209_38216.n4 VSS 9.1866f
C10136 a_n4209_38216.n5 VSS 0.192045f
C10137 a_n4209_38216.t1 VSS 0.047234f
C10138 a_n4209_38216.t0 VSS 0.047234f
C10139 a_n4209_38216.n6 VSS 0.097166f
C10140 a_n4209_38216.n7 VSS 0.392021f
C10141 a_n4209_38216.n8 VSS 0.120212f
C10142 a_n4209_38216.t3 VSS 0.047234f
C10143 VREF_GND.t21 VSS 0.279548f
C10144 VREF_GND.t44 VSS 0.275287f
C10145 VREF_GND.n0 VSS 0.753594f
C10146 VREF_GND.t18 VSS 0.275287f
C10147 VREF_GND.n1 VSS 0.396367f
C10148 VREF_GND.t33 VSS 0.275287f
C10149 VREF_GND.n2 VSS 0.396367f
C10150 VREF_GND.t32 VSS 0.275287f
C10151 VREF_GND.n3 VSS 0.396367f
C10152 VREF_GND.t19 VSS 0.076737f
C10153 VREF_GND.t23 VSS 0.076737f
C10154 VREF_GND.n4 VSS 0.193169f
C10155 VREF_GND.n5 VSS 0.339262f
C10156 VREF_GND.t20 VSS 0.275287f
C10157 VREF_GND.n6 VSS 1.66922f
C10158 VREF_GND.t31 VSS 0.306946f
C10159 VREF_GND.t22 VSS 0.306946f
C10160 VREF_GND.n7 VSS 1.02045f
C10161 VREF_GND.n8 VSS 1.82943f
C10162 VREF_GND.t8 VSS 0.306946f
C10163 VREF_GND.t30 VSS 0.306946f
C10164 VREF_GND.n9 VSS 1.02045f
C10165 VREF_GND.n10 VSS 0.702822f
C10166 VREF_GND.t9 VSS 0.306946f
C10167 VREF_GND.t7 VSS 0.306946f
C10168 VREF_GND.n11 VSS 1.02045f
C10169 VREF_GND.n12 VSS 0.702822f
C10170 VREF_GND.t12 VSS 0.306946f
C10171 VREF_GND.t6 VSS 0.306946f
C10172 VREF_GND.n13 VSS 1.02045f
C10173 VREF_GND.n14 VSS 0.702822f
C10174 VREF_GND.t16 VSS 0.306946f
C10175 VREF_GND.t13 VSS 0.306946f
C10176 VREF_GND.n15 VSS 1.02045f
C10177 VREF_GND.n16 VSS 0.705147f
C10178 VREF_GND.t15 VSS 0.306946f
C10179 VREF_GND.t14 VSS 0.306946f
C10180 VREF_GND.n17 VSS 1.02045f
C10181 VREF_GND.n18 VSS 0.705147f
C10182 VREF_GND.t11 VSS 0.306946f
C10183 VREF_GND.t10 VSS 0.306946f
C10184 VREF_GND.n19 VSS 1.02045f
C10185 VREF_GND.n20 VSS 0.702822f
C10186 VREF_GND.t17 VSS 1.36818f
C10187 VREF_GND.n21 VSS 11.8345f
C10188 VREF_GND.t45 VSS 0.279548f
C10189 VREF_GND.t25 VSS 0.275287f
C10190 VREF_GND.n22 VSS 0.753594f
C10191 VREF_GND.t27 VSS 0.275287f
C10192 VREF_GND.n23 VSS 0.396367f
C10193 VREF_GND.t43 VSS 0.275287f
C10194 VREF_GND.n24 VSS 0.396367f
C10195 VREF_GND.t24 VSS 0.275287f
C10196 VREF_GND.n25 VSS 0.396367f
C10197 VREF_GND.t26 VSS 0.076737f
C10198 VREF_GND.t5 VSS 0.076737f
C10199 VREF_GND.n26 VSS 0.193169f
C10200 VREF_GND.n27 VSS 0.339262f
C10201 VREF_GND.t4 VSS 0.275287f
C10202 VREF_GND.n28 VSS 1.66922f
C10203 VREF_GND.t42 VSS 0.306946f
C10204 VREF_GND.t28 VSS 0.306946f
C10205 VREF_GND.n29 VSS 1.02045f
C10206 VREF_GND.n30 VSS 1.82943f
C10207 VREF_GND.t29 VSS 0.306946f
C10208 VREF_GND.t3 VSS 0.306946f
C10209 VREF_GND.n31 VSS 1.02045f
C10210 VREF_GND.n32 VSS 0.702822f
C10211 VREF_GND.t0 VSS 0.306946f
C10212 VREF_GND.t2 VSS 0.306946f
C10213 VREF_GND.n33 VSS 1.02045f
C10214 VREF_GND.n34 VSS 0.702822f
C10215 VREF_GND.t1 VSS 0.306946f
C10216 VREF_GND.t40 VSS 0.306946f
C10217 VREF_GND.n35 VSS 1.02045f
C10218 VREF_GND.n36 VSS 0.702822f
C10219 VREF_GND.t34 VSS 0.306946f
C10220 VREF_GND.t39 VSS 0.306946f
C10221 VREF_GND.n37 VSS 1.02045f
C10222 VREF_GND.n38 VSS 0.705147f
C10223 VREF_GND.t37 VSS 0.306946f
C10224 VREF_GND.t35 VSS 0.306946f
C10225 VREF_GND.n39 VSS 1.02045f
C10226 VREF_GND.n40 VSS 0.705147f
C10227 VREF_GND.t41 VSS 0.306946f
C10228 VREF_GND.t36 VSS 0.306946f
C10229 VREF_GND.n41 VSS 1.02045f
C10230 VREF_GND.n42 VSS 0.702822f
C10231 VREF_GND.t38 VSS 1.36818f
C10232 VREF_GND.n43 VSS 11.8959f
C10233 a_18114_32519.t0 VSS 0.038616f
C10234 a_18114_32519.t2 VSS 0.0251f
C10235 a_18114_32519.t3 VSS 0.0251f
C10236 a_18114_32519.n0 VSS 0.092957f
C10237 a_18114_32519.n1 VSS 0.166159f
C10238 a_18114_32519.t8 VSS 0.508439f
C10239 a_18114_32519.t11 VSS 0.523017f
C10240 a_18114_32519.t5 VSS 0.509726f
C10241 a_18114_32519.t6 VSS 0.508439f
C10242 a_18114_32519.t9 VSS 0.509726f
C10243 a_18114_32519.t4 VSS 0.508439f
C10244 a_18114_32519.t7 VSS 0.509726f
C10245 a_18114_32519.n2 VSS 0.244332f
C10246 a_18114_32519.t10 VSS 0.508439f
C10247 a_18114_32519.n3 VSS 0.252575f
C10248 a_18114_32519.n4 VSS 0.294663f
C10249 a_18114_32519.n5 VSS 0.263898f
C10250 a_18114_32519.n6 VSS 0.244332f
C10251 a_18114_32519.n7 VSS 0.263898f
C10252 a_18114_32519.n8 VSS 0.244332f
C10253 a_18114_32519.n9 VSS 0.472316f
C10254 a_18114_32519.n10 VSS 6.10861f
C10255 a_18114_32519.n11 VSS 5.16128f
C10256 a_18114_32519.n12 VSS 0.077262f
C10257 a_18114_32519.t1 VSS 0.038616f
C10258 a_4646_46812.n0 VSS 0.02296f
C10259 a_4646_46812.n1 VSS 0.019052f
C10260 a_4646_46812.n2 VSS 0.086824f
C10261 a_4646_46812.n3 VSS 0.019052f
C10262 a_4646_46812.n4 VSS 0.050014f
C10263 a_4646_46812.n5 VSS 0.019052f
C10264 a_4646_46812.n6 VSS 0.049782f
C10265 a_4646_46812.n7 VSS 0.019052f
C10266 a_4646_46812.n8 VSS 0.049782f
C10267 a_4646_46812.t34 VSS 0.014148f
C10268 a_4646_46812.n9 VSS 0.027596f
C10269 a_4646_46812.t41 VSS 0.014148f
C10270 a_4646_46812.n10 VSS 0.039253f
C10271 a_4646_46812.n11 VSS 0.339789f
C10272 a_4646_46812.t40 VSS 0.014148f
C10273 a_4646_46812.n12 VSS 0.030615f
C10274 a_4646_46812.n13 VSS 0.184686f
C10275 a_4646_46812.t32 VSS 0.014148f
C10276 a_4646_46812.n14 VSS 0.032038f
C10277 a_4646_46812.t39 VSS 0.014148f
C10278 a_4646_46812.n15 VSS 0.035435f
C10279 a_4646_46812.n16 VSS 0.366686f
C10280 a_4646_46812.n17 VSS 0.155423f
C10281 a_4646_46812.n18 VSS 0.018077f
C10282 a_4646_46812.n19 VSS 0.016189f
C10283 a_4646_46812.n20 VSS 0.030136f
C10284 a_4646_46812.n21 VSS 0.018804f
C10285 a_4646_46812.n22 VSS 0.01348f
C10286 a_4646_46812.n24 VSS 0.054758f
C10287 a_4646_46812.n26 VSS 0.032914f
C10288 a_4646_46812.n28 VSS 0.033951f
C10289 a_4646_46812.n30 VSS 0.032914f
C10290 a_4646_46812.n32 VSS 0.033078f
C10291 a_4646_46812.n34 VSS 0.028414f
C10292 a_4646_46812.n36 VSS 0.088175f
C10293 a_4646_46812.n37 VSS 0.106159f
C10294 a_4646_46812.n38 VSS 0.042957f
C10295 a_4646_46812.n39 VSS 0.019052f
C10296 SMPL_ON_N.t7 VSS 0.022613f
C10297 SMPL_ON_N.t5 VSS 0.022613f
C10298 SMPL_ON_N.n0 VSS 0.069791f
C10299 SMPL_ON_N.t4 VSS 0.022613f
C10300 SMPL_ON_N.t6 VSS 0.022613f
C10301 SMPL_ON_N.n1 VSS 0.049941f
C10302 SMPL_ON_N.n2 VSS 0.270239f
C10303 SMPL_ON_N.t1 VSS 0.034789f
C10304 SMPL_ON_N.t3 VSS 0.034789f
C10305 SMPL_ON_N.n3 VSS 0.10593f
C10306 SMPL_ON_N.t0 VSS 0.034789f
C10307 SMPL_ON_N.t2 VSS 0.034789f
C10308 SMPL_ON_N.n4 VSS 0.077065f
C10309 SMPL_ON_N.n5 VSS 0.367794f
C10310 SMPL_ON_N.n6 VSS 3.58136f
C10311 SMPL_ON_N.t9 VSS 0.033751f
C10312 SMPL_ON_N.t8 VSS 0.054116f
C10313 SMPL_ON_N.n7 VSS 0.16577f
C10314 a_3422_30871.t0 VSS 0.024908f
C10315 a_3422_30871.t2 VSS 0.01619f
C10316 a_3422_30871.t3 VSS 0.01619f
C10317 a_3422_30871.n0 VSS 0.0563f
C10318 a_3422_30871.n1 VSS 0.125783f
C10319 a_3422_30871.t11 VSS 0.327959f
C10320 a_3422_30871.t16 VSS 0.337737f
C10321 a_3422_30871.t12 VSS 0.328512f
C10322 a_3422_30871.t20 VSS 0.327959f
C10323 a_3422_30871.t6 VSS 0.328512f
C10324 a_3422_30871.t7 VSS 0.327959f
C10325 a_3422_30871.t13 VSS 0.328512f
C10326 a_3422_30871.n2 VSS 0.150752f
C10327 a_3422_30871.t8 VSS 0.327959f
C10328 a_3422_30871.n3 VSS 0.162119f
C10329 a_3422_30871.n4 VSS 0.220887f
C10330 a_3422_30871.n5 VSS 0.16864f
C10331 a_3422_30871.n6 VSS 0.150752f
C10332 a_3422_30871.n7 VSS 0.16864f
C10333 a_3422_30871.n8 VSS 0.150752f
C10334 a_3422_30871.n9 VSS 0.297892f
C10335 a_3422_30871.n10 VSS 1.13984f
C10336 a_3422_30871.n11 VSS 0.125783f
C10337 a_3422_30871.t9 VSS 0.327959f
C10338 a_3422_30871.t10 VSS 0.328512f
C10339 a_3422_30871.t18 VSS 0.327959f
C10340 a_3422_30871.t5 VSS 0.328512f
C10341 a_3422_30871.t19 VSS 0.327959f
C10342 a_3422_30871.t17 VSS 0.328512f
C10343 a_3422_30871.n12 VSS 0.150752f
C10344 a_3422_30871.t21 VSS 0.327959f
C10345 a_3422_30871.n13 VSS 0.162119f
C10346 a_3422_30871.n14 VSS 0.220887f
C10347 a_3422_30871.n15 VSS 0.16864f
C10348 a_3422_30871.n16 VSS 0.150752f
C10349 a_3422_30871.n17 VSS 0.16864f
C10350 a_3422_30871.n18 VSS 0.150752f
C10351 a_3422_30871.t15 VSS 0.337737f
C10352 a_3422_30871.n19 VSS 0.297892f
C10353 a_3422_30871.n20 VSS 1.27603f
C10354 a_3422_30871.n21 VSS 5.13817f
C10355 a_3422_30871.t14 VSS 0.038747f
C10356 a_3422_30871.t4 VSS 0.024165f
C10357 a_3422_30871.n22 VSS 0.150662f
C10358 a_3422_30871.n23 VSS 4.04291f
C10359 a_3422_30871.n24 VSS 0.33736f
C10360 a_3422_30871.n25 VSS 0.050969f
C10361 a_3422_30871.t1 VSS 0.024908f
C10362 a_4223_44672.t0 VSS 0.028881f
C10363 a_4223_44672.t3 VSS 0.018773f
C10364 a_4223_44672.t2 VSS 0.018773f
C10365 a_4223_44672.n0 VSS 0.090458f
C10366 a_4223_44672.t8 VSS 0.047612f
C10367 a_4223_44672.t4 VSS 0.117982f
C10368 a_4223_44672.t7 VSS 0.048671f
C10369 a_4223_44672.t6 VSS 0.030563f
C10370 a_4223_44672.n1 VSS 0.065425f
C10371 a_4223_44672.t5 VSS 0.048098f
C10372 a_4223_44672.t9 VSS 0.029798f
C10373 a_4223_44672.n2 VSS 0.105228f
C10374 a_4223_44672.n3 VSS 0.491756f
C10375 a_4223_44672.n4 VSS 1.52867f
C10376 a_4223_44672.n5 VSS 0.24244f
C10377 a_4223_44672.n6 VSS 0.057992f
C10378 a_4223_44672.t1 VSS 0.028881f
C10379 VIN_N.t3 VSS 0.265616f
C10380 VIN_N.t2 VSS 0.268837f
C10381 VIN_N.n0 VSS 1.60996f
C10382 VIN_N.t5 VSS 0.144996f
C10383 VIN_N.t7 VSS 0.144996f
C10384 VIN_N.n1 VSS 0.513004f
C10385 VIN_N.t6 VSS 0.062178f
C10386 VIN_N.t13 VSS 0.060662f
C10387 VIN_N.n2 VSS 0.20897f
C10388 VIN_N.t10 VSS 0.06066f
C10389 VIN_N.n3 VSS 0.113566f
C10390 VIN_N.t8 VSS 0.064106f
C10391 VIN_N.n4 VSS 0.172747f
C10392 VIN_N.t11 VSS 0.063671f
C10393 VIN_N.n5 VSS 0.140791f
C10394 VIN_N.t15 VSS 0.063671f
C10395 VIN_N.n6 VSS 0.152702f
C10396 VIN_N.t9 VSS 0.063671f
C10397 VIN_N.n7 VSS 0.152702f
C10398 VIN_N.t14 VSS 0.063671f
C10399 VIN_N.n8 VSS 0.163687f
C10400 VIN_N.t1 VSS 0.036249f
C10401 VIN_N.t12 VSS 0.036249f
C10402 VIN_N.n9 VSS 0.098859f
C10403 VIN_N.n10 VSS 0.216413f
C10404 VIN_N.t0 VSS 0.136218f
C10405 VIN_N.n11 VSS 0.814626f
C10406 VIN_N.n12 VSS 0.960503f
C10407 VIN_N.t4 VSS 0.674566f
C10408 VIN_N.n13 VSS 1.45115f
C10409 VIN_N.n14 VSS 6.8455f
C10410 a_10890_34112.t1 VSS 0.036613f
C10411 a_10890_34112.n0 VSS 1.87509f
C10412 a_10890_34112.n1 VSS 1.90362f
C10413 a_10890_34112.t6 VSS 5.31306f
C10414 a_10890_34112.n2 VSS 0.577033f
C10415 a_10890_34112.n3 VSS 0.483993f
C10416 a_10890_34112.n4 VSS 0.445202f
C10417 a_10890_34112.n5 VSS 1.81073f
C10418 a_10890_34112.t7 VSS 5.31306f
C10419 a_10890_34112.n6 VSS 4.34368f
C10420 a_10890_34112.t4 VSS 5.31306f
C10421 a_10890_34112.n7 VSS 1.73865f
C10422 a_10890_34112.n8 VSS 0.21528f
C10423 a_10890_34112.n9 VSS 0.174568f
C10424 a_10890_34112.n10 VSS 0.420325f
C10425 a_10890_34112.n11 VSS 0.446058f
C10426 a_10890_34112.t5 VSS 5.31306f
C10427 a_10890_34112.n12 VSS 4.14877f
C10428 a_10890_34112.n13 VSS 0.47303f
C10429 a_10890_34112.n14 VSS 0.49298f
C10430 a_10890_34112.t2 VSS 0.036613f
C10431 a_10890_34112.t3 VSS 0.036613f
C10432 a_10890_34112.n15 VSS 0.099794f
C10433 a_10890_34112.n16 VSS 0.559191f
C10434 a_10890_34112.n17 VSS 0.093314f
C10435 a_10890_34112.t0 VSS 0.036613f
C10436 EN_VIN_BSTR_N.t2 VSS 0.111063f
C10437 EN_VIN_BSTR_N.t1 VSS 0.107644f
C10438 EN_VIN_BSTR_N.n0 VSS 0.285814f
C10439 EN_VIN_BSTR_N.t0 VSS 0.107508f
C10440 EN_VIN_BSTR_N.n1 VSS 0.17615f
C10441 EN_VIN_BSTR_N.t4 VSS 0.030933f
C10442 EN_VIN_BSTR_N.t5 VSS 0.030933f
C10443 EN_VIN_BSTR_N.n2 VSS 0.063662f
C10444 EN_VIN_BSTR_N.t6 VSS 0.030933f
C10445 EN_VIN_BSTR_N.t3 VSS 0.030933f
C10446 EN_VIN_BSTR_N.n3 VSS 0.063662f
C10447 EN_VIN_BSTR_N.t22 VSS 0.041127f
C10448 EN_VIN_BSTR_N.t16 VSS 0.04343f
C10449 EN_VIN_BSTR_N.n4 VSS 0.058307f
C10450 EN_VIN_BSTR_N.t13 VSS 0.016326f
C10451 EN_VIN_BSTR_N.n5 VSS 0.312119f
C10452 EN_VIN_BSTR_N.n6 VSS 0.06955f
C10453 EN_VIN_BSTR_N.n7 VSS 0.074759f
C10454 EN_VIN_BSTR_N.n8 VSS 0.0838f
C10455 EN_VIN_BSTR_N.t21 VSS 0.016204f
C10456 EN_VIN_BSTR_N.t17 VSS 0.01635f
C10457 EN_VIN_BSTR_N.n9 VSS 0.11489f
C10458 EN_VIN_BSTR_N.t19 VSS 0.016204f
C10459 EN_VIN_BSTR_N.t7 VSS 0.020036f
C10460 EN_VIN_BSTR_N.t8 VSS 0.023039f
C10461 EN_VIN_BSTR_N.n10 VSS 0.033139f
C10462 EN_VIN_BSTR_N.t12 VSS 0.02977f
C10463 EN_VIN_BSTR_N.n11 VSS 0.061739f
C10464 EN_VIN_BSTR_N.t14 VSS 0.016182f
C10465 EN_VIN_BSTR_N.n12 VSS 0.032604f
C10466 EN_VIN_BSTR_N.t9 VSS 0.016182f
C10467 EN_VIN_BSTR_N.n13 VSS 0.038345f
C10468 EN_VIN_BSTR_N.t20 VSS 0.016182f
C10469 EN_VIN_BSTR_N.n14 VSS 0.038345f
C10470 EN_VIN_BSTR_N.t10 VSS 0.016182f
C10471 EN_VIN_BSTR_N.n15 VSS 0.02944f
C10472 EN_VIN_BSTR_N.t23 VSS 0.016207f
C10473 EN_VIN_BSTR_N.n16 VSS 0.058941f
C10474 EN_VIN_BSTR_N.n17 VSS 0.0656f
C10475 EN_VIN_BSTR_N.n18 VSS 0.352047f
C10476 EN_VIN_BSTR_N.t18 VSS 0.08989f
C10477 EN_VIN_BSTR_N.t15 VSS 0.083309f
C10478 EN_VIN_BSTR_N.t11 VSS 0.085697f
C10479 EN_VIN_BSTR_N.n19 VSS 0.075473f
C10480 EN_VIN_BSTR_N.n20 VSS 0.086725f
C10481 EN_VIN_BSTR_N.n21 VSS 0.516963f
C10482 a_17730_32519.t0 VSS 0.049614f
C10483 a_17730_32519.t5 VSS 0.653249f
C10484 a_17730_32519.n0 VSS 0.32448f
C10485 a_17730_32519.t7 VSS 0.653249f
C10486 a_17730_32519.t4 VSS 0.671978f
C10487 a_17730_32519.t6 VSS 0.654902f
C10488 a_17730_32519.n1 VSS 0.31392f
C10489 a_17730_32519.n2 VSS 0.606838f
C10490 a_17730_32519.n3 VSS 7.49599f
C10491 a_17730_32519.t3 VSS 0.032249f
C10492 a_17730_32519.t2 VSS 0.032249f
C10493 a_17730_32519.n4 VSS 0.064498f
C10494 a_17730_32519.n5 VSS 6.84829f
C10495 a_17730_32519.n6 VSS 0.148875f
C10496 a_17730_32519.t1 VSS 0.049614f
C10497 a_n1151_42308.t0 VSS 0.011346f
C10498 a_n1151_42308.n0 VSS 0.012184f
C10499 a_n1151_42308.t11 VSS 0.033139f
C10500 a_n1151_42308.t9 VSS 0.017446f
C10501 a_n1151_42308.n1 VSS 0.085275f
C10502 a_n1151_42308.t6 VSS 0.022955f
C10503 a_n1151_42308.n2 VSS 0.094921f
C10504 a_n1151_42308.t10 VSS 0.033139f
C10505 a_n1151_42308.t18 VSS 0.017446f
C10506 a_n1151_42308.n3 VSS 0.079676f
C10507 a_n1151_42308.n4 VSS 1.10806f
C10508 a_n1151_42308.t16 VSS 0.022955f
C10509 a_n1151_42308.n5 VSS 0.040583f
C10510 a_n1151_42308.n6 VSS 0.290815f
C10511 a_n1151_42308.t7 VSS 0.022955f
C10512 a_n1151_42308.n7 VSS 0.049003f
C10513 a_n1151_42308.n8 VSS 0.375682f
C10514 a_n1151_42308.t4 VSS 0.022955f
C10515 a_n1151_42308.n9 VSS 0.040583f
C10516 a_n1151_42308.n10 VSS 0.32164f
C10517 a_n1151_42308.t12 VSS 0.022955f
C10518 a_n1151_42308.n11 VSS 0.042881f
C10519 a_n1151_42308.n12 VSS 1.51515f
C10520 a_n1151_42308.t17 VSS 0.012443f
C10521 a_n1151_42308.n13 VSS 0.034491f
C10522 a_n1151_42308.n14 VSS 0.476542f
C10523 a_n1151_42308.n15 VSS 0.447102f
C10524 a_n1151_42308.n16 VSS 0.247501f
C10525 a_n1151_42308.n17 VSS 0.026998f
C10526 a_n1151_42308.t1 VSS 0.011346f
C10527 a_3537_45260.t0 VSS 0.013646f
C10528 a_3537_45260.t1 VSS 0.013646f
C10529 a_3537_45260.t2 VSS 0.013646f
C10530 a_3537_45260.n0 VSS 0.041439f
C10531 a_3537_45260.n1 VSS 0.034113f
C10532 a_3537_45260.n2 VSS 0.020268f
C10533 a_3537_45260.n3 VSS 0.112886f
C10534 a_3537_45260.t16 VSS 0.022497f
C10535 a_3537_45260.t26 VSS 0.049316f
C10536 a_3537_45260.t17 VSS 0.021794f
C10537 a_3537_45260.t22 VSS 0.0422f
C10538 a_3537_45260.t13 VSS 0.022727f
C10539 a_3537_45260.t24 VSS 0.01408f
C10540 a_3537_45260.n4 VSS 0.048983f
C10541 a_3537_45260.t28 VSS 0.014441f
C10542 a_3537_45260.t12 VSS 0.022997f
C10543 a_3537_45260.n5 VSS 0.033493f
C10544 a_3537_45260.t23 VSS 0.014288f
C10545 a_3537_45260.t9 VSS 0.022811f
C10546 a_3537_45260.n6 VSS 0.040615f
C10547 a_3537_45260.n7 VSS 0.331626f
C10548 a_3537_45260.t21 VSS 0.014288f
C10549 a_3537_45260.t14 VSS 0.022811f
C10550 a_3537_45260.n8 VSS 0.037426f
C10551 a_3537_45260.n9 VSS 0.075868f
C10552 a_3537_45260.t11 VSS 0.012509f
C10553 a_3537_45260.t18 VSS 0.021228f
C10554 a_3537_45260.t8 VSS 0.012509f
C10555 a_3537_45260.t29 VSS 0.021228f
C10556 a_3537_45260.n10 VSS 0.035617f
C10557 a_3537_45260.n11 VSS 0.053714f
C10558 a_3537_45260.t20 VSS 0.014441f
C10559 a_3537_45260.t27 VSS 0.022997f
C10560 a_3537_45260.n12 VSS 0.035021f
C10561 a_3537_45260.n13 VSS 0.214882f
C10562 a_3537_45260.n14 VSS 0.222535f
C10563 a_3537_45260.t25 VSS 0.014441f
C10564 a_3537_45260.t15 VSS 0.022997f
C10565 a_3537_45260.n15 VSS 0.034728f
C10566 a_3537_45260.n16 VSS 0.279908f
C10567 a_3537_45260.t10 VSS 0.014441f
C10568 a_3537_45260.t19 VSS 0.022997f
C10569 a_3537_45260.n17 VSS 0.032668f
C10570 a_3537_45260.n18 VSS 0.30792f
C10571 a_3537_45260.n19 VSS 0.394117f
C10572 a_3537_45260.n20 VSS 0.351525f
C10573 a_3537_45260.n21 VSS 0.381509f
C10574 a_3537_45260.n22 VSS 0.078654f
C10575 a_3537_45260.n23 VSS 0.115906f
C10576 a_3537_45260.n24 VSS 0.030478f
C10577 a_3537_45260.t3 VSS 0.013646f
C10578 a_4185_45028.t2 VSS 0.034622f
C10579 a_4185_45028.t1 VSS 0.16497f
C10580 a_4185_45028.t5 VSS 0.031121f
C10581 a_4185_45028.t3 VSS 0.04877f
C10582 a_4185_45028.n0 VSS 2.23592f
C10583 a_4185_45028.t6 VSS 0.035785f
C10584 a_4185_45028.t4 VSS 0.057313f
C10585 a_4185_45028.n1 VSS 0.144088f
C10586 a_4185_45028.n2 VSS 8.02056f
C10587 a_4185_45028.n3 VSS 0.322709f
C10588 a_4185_45028.n4 VSS 0.069519f
C10589 a_4185_45028.t0 VSS 0.034622f
C10590 a_n2442_46660.t2 VSS 0.036264f
C10591 a_n2442_46660.t3 VSS 0.036264f
C10592 a_n2442_46660.n0 VSS 0.134301f
C10593 a_n2442_46660.t4 VSS 0.092121f
C10594 a_n2442_46660.t5 VSS 0.057467f
C10595 a_n2442_46660.n1 VSS 2.53127f
C10596 a_n2442_46660.n2 VSS 9.28911f
C10597 a_n2442_46660.t0 VSS 0.05579f
C10598 a_n2442_46660.n3 VSS 0.111626f
C10599 a_n2442_46660.t1 VSS 0.05579f
C10600 a_11691_44458.t0 VSS 0.019529f
C10601 a_11691_44458.t3 VSS 0.012694f
C10602 a_11691_44458.t2 VSS 0.012694f
C10603 a_11691_44458.n0 VSS 0.061167f
C10604 a_11691_44458.t9 VSS 0.032557f
C10605 a_11691_44458.t6 VSS 0.020376f
C10606 a_11691_44458.n1 VSS 0.118058f
C10607 a_11691_44458.t4 VSS 0.05704f
C10608 a_11691_44458.t7 VSS 0.030029f
C10609 a_11691_44458.n2 VSS 0.14527f
C10610 a_11691_44458.n3 VSS 1.42138f
C10611 a_11691_44458.t8 VSS 0.032911f
C10612 a_11691_44458.t5 VSS 0.020667f
C10613 a_11691_44458.n4 VSS 0.046752f
C10614 a_11691_44458.n5 VSS 0.868404f
C10615 a_11691_44458.n6 VSS 0.341727f
C10616 a_11691_44458.n7 VSS 0.039214f
C10617 a_11691_44458.t1 VSS 0.019529f
C10618 a_8049_45260.t2 VSS 0.011355f
C10619 a_8049_45260.t1 VSS 0.054106f
C10620 a_8049_45260.t3 VSS 0.015995f
C10621 a_8049_45260.t4 VSS 0.010207f
C10622 a_8049_45260.n0 VSS 0.149081f
C10623 a_8049_45260.t6 VSS 0.011737f
C10624 a_8049_45260.t5 VSS 0.018797f
C10625 a_8049_45260.n1 VSS 0.043326f
C10626 a_8049_45260.n2 VSS 3.93103f
C10627 a_8049_45260.n3 VSS 0.120211f
C10628 a_8049_45260.n4 VSS 0.0228f
C10629 a_8049_45260.t0 VSS 0.011355f
C10630 a_n4318_39768.t0 VSS 0.041093f
C10631 a_n4318_39768.t2 VSS 0.026711f
C10632 a_n4318_39768.t3 VSS 0.026711f
C10633 a_n4318_39768.n0 VSS 0.092883f
C10634 a_n4318_39768.t4 VSS 0.06865f
C10635 a_n4318_39768.t5 VSS 0.042994f
C10636 a_n4318_39768.n1 VSS 0.865599f
C10637 a_n4318_39768.n2 VSS 4.51018f
C10638 a_n4318_39768.n3 VSS 0.084088f
C10639 a_n4318_39768.t1 VSS 0.041093f
C10640 a_13661_43548.t0 VSS 0.014155f
C10641 a_13661_43548.n0 VSS 0.034074f
C10642 a_13661_43548.t23 VSS 0.010114f
C10643 a_13661_43548.n1 VSS 0.039828f
C10644 a_13661_43548.t15 VSS 0.022018f
C10645 a_13661_43548.t22 VSS 0.012975f
C10646 a_13661_43548.t21 VSS 0.022018f
C10647 a_13661_43548.t16 VSS 0.012975f
C10648 a_13661_43548.n2 VSS 0.03729f
C10649 a_13661_43548.n3 VSS 0.060219f
C10650 a_13661_43548.t7 VSS 0.023854f
C10651 a_13661_43548.t18 VSS 0.014979f
C10652 a_13661_43548.n4 VSS 0.041199f
C10653 a_13661_43548.n5 VSS 0.355964f
C10654 a_13661_43548.t5 VSS 0.023854f
C10655 a_13661_43548.t25 VSS 0.014979f
C10656 a_13661_43548.n6 VSS 0.036082f
C10657 a_13661_43548.t14 VSS 0.021487f
C10658 a_13661_43548.t24 VSS 0.010189f
C10659 a_13661_43548.n7 VSS 0.080015f
C10660 a_13661_43548.t13 VSS 0.014821f
C10661 a_13661_43548.t9 VSS 0.02366f
C10662 a_13661_43548.n8 VSS 0.038076f
C10663 a_13661_43548.t12 VSS 0.023854f
C10664 a_13661_43548.t11 VSS 0.014979f
C10665 a_13661_43548.n9 VSS 0.037562f
C10666 a_13661_43548.t6 VSS 0.018718f
C10667 a_13661_43548.t19 VSS 0.012675f
C10668 a_13661_43548.n10 VSS 0.064891f
C10669 a_13661_43548.n11 VSS 0.548106f
C10670 a_13661_43548.n12 VSS 0.264285f
C10671 a_13661_43548.n13 VSS 0.181588f
C10672 a_13661_43548.n14 VSS 0.426773f
C10673 a_13661_43548.n15 VSS 0.354892f
C10674 a_13661_43548.t20 VSS 0.01474f
C10675 a_13661_43548.t17 VSS 0.024515f
C10676 a_13661_43548.n16 VSS 0.041415f
C10677 a_13661_43548.n17 VSS 0.117101f
C10678 a_13661_43548.n18 VSS 0.258123f
C10679 a_13661_43548.t4 VSS 0.010114f
C10680 a_13661_43548.n19 VSS 0.041229f
C10681 a_13661_43548.n20 VSS 0.311461f
C10682 a_13661_43548.n21 VSS 0.088391f
C10683 a_13661_43548.n22 VSS 0.028321f
C10684 a_13661_43548.t1 VSS 0.014155f
C10685 a_n3565_39590.t0 VSS 0.027653f
C10686 a_n3565_39590.t5 VSS 0.017974f
C10687 a_n3565_39590.t6 VSS 0.017974f
C10688 a_n3565_39590.n0 VSS 0.068626f
C10689 a_n3565_39590.t4 VSS 0.017974f
C10690 a_n3565_39590.t7 VSS 0.017974f
C10691 a_n3565_39590.n1 VSS 0.040793f
C10692 a_n3565_39590.n2 VSS 0.197375f
C10693 a_n3565_39590.t11 VSS 0.046601f
C10694 a_n3565_39590.t8 VSS 0.029263f
C10695 a_n3565_39590.n3 VSS 0.073708f
C10696 a_n3565_39590.t9 VSS 0.936152f
C10697 a_n3565_39590.t12 VSS 0.936008f
C10698 a_n3565_39590.n4 VSS 0.69338f
C10699 a_n3565_39590.t10 VSS 0.936008f
C10700 a_n3565_39590.n5 VSS 0.35119f
C10701 a_n3565_39590.t13 VSS 0.936008f
C10702 a_n3565_39590.n6 VSS 2.93853f
C10703 a_n3565_39590.n7 VSS 2.84095f
C10704 a_n3565_39590.n8 VSS 0.114326f
C10705 a_n3565_39590.t2 VSS 0.027653f
C10706 a_n3565_39590.t1 VSS 0.027653f
C10707 a_n3565_39590.n9 VSS 0.056884f
C10708 a_n3565_39590.n10 VSS 0.251313f
C10709 a_n3565_39590.n11 VSS 0.070376f
C10710 a_n3565_39590.t3 VSS 0.027653f
C10711 C9_P_btm.t12 VSS 0.137574f
C10712 C9_P_btm.t11 VSS 0.137574f
C10713 C9_P_btm.n0 VSS 0.439559f
C10714 C9_P_btm.t14 VSS 0.137574f
C10715 C9_P_btm.t9 VSS 0.137574f
C10716 C9_P_btm.n1 VSS 0.425131f
C10717 C9_P_btm.n2 VSS 1.33616f
C10718 C9_P_btm.t13 VSS 0.137574f
C10719 C9_P_btm.t15 VSS 0.137574f
C10720 C9_P_btm.n3 VSS 0.425131f
C10721 C9_P_btm.n4 VSS 0.684408f
C10722 C9_P_btm.t10 VSS 0.137574f
C10723 C9_P_btm.t8 VSS 0.137574f
C10724 C9_P_btm.n5 VSS 0.425131f
C10725 C9_P_btm.n6 VSS 1.08525f
C10726 C9_P_btm.t2 VSS 0.156549f
C10727 C9_P_btm.t1 VSS 0.156549f
C10728 C9_P_btm.n7 VSS 0.630592f
C10729 C9_P_btm.t3 VSS 0.156549f
C10730 C9_P_btm.t0 VSS 0.156549f
C10731 C9_P_btm.n8 VSS 0.645454f
C10732 C9_P_btm.n9 VSS 1.02683f
C10733 C9_P_btm.n10 VSS 0.61298f
C10734 C9_P_btm.t16 VSS 0.961787f
C10735 C9_P_btm.n11 VSS 0.767348f
C10736 C9_P_btm.t6 VSS 0.156549f
C10737 C9_P_btm.t4 VSS 0.156549f
C10738 C9_P_btm.n12 VSS 0.651901f
C10739 C9_P_btm.t7 VSS 0.156549f
C10740 C9_P_btm.t5 VSS 0.156549f
C10741 C9_P_btm.n13 VSS 0.63781f
C10742 C9_P_btm.n14 VSS 1.03801f
C10743 C9_P_btm.n15 VSS 2.51243f
C10744 C9_P_btm.n16 VSS 2.29491f
C10745 C9_P_btm.n17 VSS 1.01629f
C10746 C9_P_btm.n18 VSS 1.01985f
C10747 C9_P_btm.n19 VSS 1.01985f
C10748 C9_P_btm.n20 VSS 1.01629f
C10749 C9_P_btm.n21 VSS 1.01985f
C10750 C9_P_btm.n22 VSS 1.01985f
C10751 C9_P_btm.n23 VSS 1.01985f
C10752 C9_P_btm.n24 VSS 1.01985f
C10753 C9_P_btm.n25 VSS 1.01629f
C10754 C9_P_btm.n26 VSS 1.01985f
C10755 C9_P_btm.n27 VSS 1.01985f
C10756 C9_P_btm.n28 VSS 1.01629f
C10757 C9_P_btm.n29 VSS 1.01985f
C10758 C9_P_btm.n30 VSS 1.01985f
C10759 C9_P_btm.n31 VSS 1.01985f
C10760 C9_P_btm.n32 VSS 1.01985f
C10761 C9_P_btm.n33 VSS 1.01629f
C10762 C9_P_btm.n34 VSS 1.01985f
C10763 C9_P_btm.n35 VSS 1.01985f
C10764 C9_P_btm.n36 VSS 1.01629f
C10765 C9_P_btm.n37 VSS 1.01985f
C10766 C9_P_btm.n38 VSS 1.01985f
C10767 C9_P_btm.n39 VSS 1.01985f
C10768 C9_P_btm.n40 VSS 1.28218f
C10769 C9_P_btm.n41 VSS 1.01985f
C10770 C9_P_btm.n42 VSS 1.01985f
C10771 C9_P_btm.n43 VSS 1.01985f
C10772 C9_P_btm.n44 VSS 1.01985f
C10773 C9_P_btm.n45 VSS 1.01985f
C10774 C9_P_btm.n46 VSS 1.01985f
C10775 C9_P_btm.n47 VSS 1.01985f
C10776 C9_P_btm.n48 VSS 1.01985f
C10777 C9_P_btm.n49 VSS 1.01985f
C10778 C9_P_btm.n50 VSS 1.01985f
C10779 C9_P_btm.n51 VSS 0.750398f
C10780 C9_P_btm.n52 VSS 1.01985f
C10781 C9_P_btm.n53 VSS 1.01985f
C10782 C9_P_btm.n54 VSS 1.01985f
C10783 C9_P_btm.n55 VSS 1.01985f
C10784 C9_P_btm.n56 VSS 1.01985f
C10785 C9_P_btm.n57 VSS 1.01985f
C10786 C9_P_btm.n58 VSS 1.01985f
C10787 C9_P_btm.n59 VSS 1.01985f
C10788 C9_P_btm.n60 VSS 1.01985f
C10789 C9_P_btm.n61 VSS 1.01985f
C10790 C9_P_btm.n62 VSS 1.01985f
C10791 C9_P_btm.n63 VSS 1.01985f
C10792 C9_P_btm.n64 VSS 1.01985f
C10793 C9_P_btm.n65 VSS 1.01985f
C10794 C9_P_btm.n66 VSS 1.01985f
C10795 C9_P_btm.n67 VSS 1.01985f
C10796 C9_P_btm.n68 VSS 1.01985f
C10797 C9_P_btm.n69 VSS 1.01985f
C10798 C9_P_btm.n70 VSS 1.01985f
C10799 C9_P_btm.n71 VSS 1.01985f
C10800 C9_P_btm.n72 VSS 1.01985f
C10801 C9_P_btm.n73 VSS 1.01985f
C10802 C9_P_btm.n74 VSS 1.01629f
C10803 C9_P_btm.n75 VSS 1.01629f
C10804 C9_P_btm.n76 VSS 1.01985f
C10805 C9_P_btm.n77 VSS 1.01985f
C10806 C9_P_btm.n78 VSS 1.01985f
C10807 C9_P_btm.n79 VSS 1.01985f
C10808 C9_P_btm.n80 VSS 0.750398f
C10809 C9_P_btm.n81 VSS 1.45454f
C10810 C9_P_btm.n82 VSS 1.59754f
C10811 C9_P_btm.n83 VSS 1.22832f
C10812 C9_P_btm.n84 VSS 1.01985f
C10813 C9_P_btm.n85 VSS 1.01985f
C10814 C9_P_btm.n86 VSS 1.01985f
C10815 C9_P_btm.n87 VSS 1.01985f
C10816 C9_P_btm.n88 VSS 1.01629f
C10817 C9_P_btm.n89 VSS 1.01629f
C10818 C9_P_btm.n90 VSS 1.01629f
C10819 C9_P_btm.n91 VSS 1.01629f
C10820 C9_P_btm.n92 VSS 1.01629f
C10821 C9_P_btm.n93 VSS 1.01629f
C10822 C9_P_btm.n94 VSS 1.01629f
C10823 C9_P_btm.n95 VSS 1.01629f
C10824 C9_P_btm.n96 VSS 1.01629f
C10825 C9_P_btm.n97 VSS 1.01629f
C10826 C9_P_btm.n98 VSS 1.01629f
C10827 C9_P_btm.n99 VSS 1.01629f
C10828 C9_P_btm.n100 VSS 1.01629f
C10829 C9_P_btm.n101 VSS 1.01629f
C10830 C9_P_btm.n102 VSS 1.01629f
C10831 C9_P_btm.n103 VSS 1.01629f
C10832 C9_P_btm.n104 VSS 1.30558f
C10833 C9_P_btm.n105 VSS 3.15708f
C10834 C9_P_btm.n106 VSS 2.29491f
C10835 C9_P_btm.n107 VSS 4.45091f
C10836 C9_P_btm.n108 VSS 1.01985f
C10837 C9_P_btm.n109 VSS 1.01985f
C10838 C9_P_btm.n110 VSS 1.01985f
C10839 C9_P_btm.n111 VSS 1.01985f
C10840 C9_P_btm.n112 VSS 1.01985f
C10841 C9_P_btm.n113 VSS 1.01985f
C10842 C9_P_btm.n114 VSS 1.01985f
C10843 C9_P_btm.n115 VSS 1.01985f
C10844 C9_P_btm.n116 VSS 1.01985f
C10845 C9_P_btm.n117 VSS 1.01985f
C10846 C9_P_btm.n118 VSS 1.01985f
C10847 C9_P_btm.n119 VSS 1.01985f
C10848 C9_P_btm.n120 VSS 1.01985f
C10849 C9_P_btm.n121 VSS 1.01985f
C10850 C9_P_btm.n122 VSS 1.01985f
C10851 C9_P_btm.n123 VSS 1.01985f
C10852 C9_P_btm.n124 VSS 1.01985f
C10853 C9_P_btm.n125 VSS 1.01985f
C10854 C9_P_btm.n126 VSS 1.01985f
C10855 C9_P_btm.n127 VSS 1.01985f
C10856 C9_P_btm.n128 VSS 1.01985f
C10857 C9_P_btm.n129 VSS 1.01985f
C10858 C9_P_btm.n130 VSS 1.01985f
C10859 C9_P_btm.n131 VSS 1.01985f
C10860 C9_P_btm.n132 VSS 1.01985f
C10861 C9_P_btm.n133 VSS 1.01985f
C10862 C9_P_btm.n134 VSS 1.01985f
C10863 C9_P_btm.n135 VSS 1.01985f
C10864 C9_P_btm.n136 VSS 1.01985f
C10865 C9_P_btm.n137 VSS 0.750398f
C10866 C9_P_btm.n138 VSS 0.750398f
C10867 C9_P_btm.n139 VSS 1.01985f
C10868 C9_P_btm.n140 VSS 1.01985f
C10869 C9_P_btm.n141 VSS 1.01985f
C10870 C9_P_btm.n142 VSS 1.01985f
C10871 C9_P_btm.n143 VSS 1.01985f
C10872 C9_P_btm.n144 VSS 1.45454f
C10873 C9_P_btm.n145 VSS 1.01985f
C10874 C9_P_btm.n146 VSS 1.01985f
C10875 C9_P_btm.n147 VSS 1.01985f
C10876 C9_P_btm.n148 VSS 1.01985f
C10877 C9_P_btm.n149 VSS 1.01985f
C10878 C9_P_btm.n150 VSS 1.01985f
C10879 C9_P_btm.n151 VSS 1.01985f
C10880 C9_P_btm.n152 VSS 1.01985f
C10881 C9_P_btm.n153 VSS 1.01985f
C10882 C9_P_btm.n154 VSS 1.01985f
C10883 C9_P_btm.n155 VSS 1.39208f
C10884 C9_P_btm.n156 VSS 1.01985f
C10885 C9_P_btm.n157 VSS 1.01985f
C10886 C9_P_btm.n158 VSS 1.01985f
C10887 C9_P_btm.n159 VSS 1.01985f
C10888 C9_P_btm.n160 VSS 1.01985f
C10889 C9_P_btm.n161 VSS 1.01985f
C10890 C9_P_btm.n162 VSS 1.01985f
C10891 C9_P_btm.n163 VSS 1.01985f
C10892 C9_P_btm.n164 VSS 1.01985f
C10893 C9_P_btm.n165 VSS 1.01985f
C10894 C9_P_btm.n166 VSS 0.750398f
C10895 C9_P_btm.n167 VSS 1.01985f
C10896 C9_P_btm.n168 VSS 0.750398f
C10897 C9_P_btm.n169 VSS 1.01985f
C10898 C9_P_btm.n170 VSS 1.01985f
C10899 C9_P_btm.n171 VSS 1.01985f
C10900 C9_P_btm.n172 VSS 1.01985f
C10901 C9_P_btm.n173 VSS 1.01985f
C10902 C9_P_btm.n174 VSS 1.01985f
C10903 C9_P_btm.n175 VSS 1.01985f
C10904 C9_P_btm.n176 VSS 0.750398f
C10905 C9_P_btm.n177 VSS 0.750398f
C10906 C9_P_btm.n178 VSS 0.750398f
C10907 C9_P_btm.n179 VSS 1.01985f
C10908 C9_P_btm.n180 VSS 1.01985f
C10909 C9_P_btm.n181 VSS 0.750398f
C10910 C9_P_btm.n182 VSS 1.01985f
C10911 C9_P_btm.n183 VSS 1.01985f
C10912 C9_P_btm.n184 VSS 1.01985f
C10913 C9_P_btm.n185 VSS 1.01985f
C10914 C9_P_btm.n186 VSS 1.01985f
C10915 C9_P_btm.n187 VSS 1.01985f
C10916 C9_P_btm.n188 VSS 1.01985f
C10917 C9_P_btm.n189 VSS 1.01985f
C10918 C9_P_btm.n190 VSS 1.01985f
C10919 C9_P_btm.n191 VSS 1.01985f
C10920 C9_P_btm.n192 VSS 1.01985f
C10921 C9_P_btm.n193 VSS 1.28218f
C10922 C9_P_btm.n194 VSS 1.01985f
C10923 C9_P_btm.n195 VSS 1.01985f
C10924 C9_P_btm.n196 VSS 1.01985f
C10925 C9_P_btm.n197 VSS 1.01985f
C10926 C9_P_btm.n198 VSS 1.01985f
C10927 C9_P_btm.n199 VSS 1.01985f
C10928 C9_P_btm.n200 VSS 1.01985f
C10929 C9_P_btm.n201 VSS 1.01985f
C10930 C9_P_btm.n202 VSS 1.45446f
C10931 C9_P_btm.n203 VSS 0.575755f
C10932 C9_P_btm.n204 VSS 1.01985f
C10933 C9_P_btm.n205 VSS 1.01985f
C10934 C9_P_btm.n206 VSS 1.01985f
C10935 C9_P_btm.n207 VSS 1.01985f
C10936 C9_P_btm.n208 VSS 1.01985f
C10937 C9_P_btm.n209 VSS 1.23727f
C10938 C9_P_btm.n210 VSS 0.750398f
C10939 C9_P_btm.n211 VSS 0.750398f
C10940 C9_P_btm.n212 VSS 1.01985f
C10941 C9_P_btm.n213 VSS 1.01985f
C10942 C9_P_btm.n214 VSS 1.01985f
C10943 C9_P_btm.n215 VSS 1.01985f
C10944 C9_P_btm.n216 VSS 1.01985f
C10945 C9_P_btm.n217 VSS 1.01985f
C10946 C9_P_btm.n218 VSS 1.01985f
C10947 C9_P_btm.n219 VSS 1.01985f
C10948 C9_P_btm.n220 VSS 1.01985f
C10949 C9_P_btm.n221 VSS 1.01629f
C10950 C9_P_btm.n222 VSS 1.01985f
C10951 C9_P_btm.n223 VSS 1.01985f
C10952 C9_P_btm.n224 VSS 1.01985f
C10953 C9_P_btm.n225 VSS 1.01985f
C10954 C9_P_btm.n226 VSS 1.01985f
C10955 C9_P_btm.n227 VSS 1.01985f
C10956 C9_P_btm.n228 VSS 1.01985f
C10957 C9_P_btm.n229 VSS 1.01629f
C10958 C9_P_btm.n230 VSS 1.01985f
C10959 C9_P_btm.n231 VSS 1.01985f
C10960 C9_P_btm.n232 VSS 1.01629f
C10961 C9_P_btm.n233 VSS 1.01985f
C10962 C9_P_btm.n234 VSS 1.01985f
C10963 C9_P_btm.n235 VSS 1.01985f
C10964 C9_P_btm.n236 VSS 1.01985f
C10965 C9_P_btm.n237 VSS 1.01985f
C10966 C9_P_btm.n238 VSS 0.750398f
C10967 C9_P_btm.n239 VSS 1.01985f
C10968 C9_P_btm.n240 VSS 1.01985f
C10969 C9_P_btm.n241 VSS 1.01985f
C10970 C9_P_btm.n242 VSS 1.01985f
C10971 C9_P_btm.n243 VSS 1.01985f
C10972 C9_P_btm.n244 VSS 1.01985f
C10973 C9_P_btm.n245 VSS 1.01985f
C10974 C9_P_btm.n246 VSS 0.750398f
C10975 C9_P_btm.n247 VSS 0.750398f
C10976 C9_P_btm.n248 VSS 0.750398f
C10977 C9_P_btm.n249 VSS 0.750398f
C10978 C9_P_btm.n250 VSS 1.01985f
C10979 C9_P_btm.n251 VSS 1.01985f
C10980 C9_P_btm.n252 VSS 1.01985f
C10981 C9_P_btm.n253 VSS 1.01985f
C10982 C9_P_btm.n254 VSS 1.01985f
C10983 C9_P_btm.n255 VSS 1.01985f
C10984 C9_P_btm.n256 VSS 1.01985f
C10985 C9_P_btm.n257 VSS 1.01985f
C10986 C9_P_btm.n258 VSS 1.01985f
C10987 C9_P_btm.n259 VSS 1.01985f
C10988 C9_P_btm.n260 VSS 1.01985f
C10989 C9_P_btm.n261 VSS 1.01985f
C10990 C9_P_btm.n262 VSS 1.01985f
C10991 C9_P_btm.n263 VSS 1.45446f
C10992 C9_P_btm.n264 VSS 1.59744f
C10993 C9_P_btm.n265 VSS 1.22832f
C10994 C9_P_btm.n266 VSS 1.01629f
C10995 C9_P_btm.n267 VSS 1.01629f
C10996 C9_P_btm.n268 VSS 1.01985f
C10997 C9_P_btm.n269 VSS 1.01985f
C10998 C9_P_btm.n270 VSS 1.01985f
C10999 C9_P_btm.n271 VSS 1.01985f
C11000 C9_P_btm.n272 VSS 1.01629f
C11001 C9_P_btm.n273 VSS 1.01629f
C11002 C9_P_btm.n274 VSS 1.01629f
C11003 C9_P_btm.n275 VSS 1.01629f
C11004 C9_P_btm.n276 VSS 1.01985f
C11005 C9_P_btm.n277 VSS 1.01985f
C11006 C9_P_btm.n278 VSS 1.01629f
C11007 C9_P_btm.n279 VSS 1.01985f
C11008 C9_P_btm.n280 VSS 1.01985f
C11009 C9_P_btm.n281 VSS 1.01629f
C11010 C9_P_btm.n282 VSS 1.01985f
C11011 C9_P_btm.n283 VSS 1.01985f
C11012 C9_P_btm.n284 VSS 1.01985f
C11013 C9_P_btm.n285 VSS 1.01985f
C11014 C9_P_btm.n286 VSS 1.30559f
C11015 C9_P_btm.n287 VSS 1.01985f
C11016 C9_P_btm.n288 VSS 1.01985f
C11017 C9_P_btm.n289 VSS 3.15719f
C11018 C9_P_btm.n290 VSS 1.01985f
C11019 C9_P_btm.n291 VSS 1.30558f
C11020 C9_P_btm.n292 VSS 1.01985f
C11021 C9_P_btm.n293 VSS 1.01985f
C11022 C9_P_btm.n294 VSS 1.01629f
C11023 C9_P_btm.n295 VSS 1.01629f
C11024 C9_P_btm.n296 VSS 1.01985f
C11025 C9_P_btm.n297 VSS 1.01985f
C11026 C9_P_btm.n298 VSS 1.01985f
C11027 C9_P_btm.n299 VSS 1.01985f
C11028 C9_P_btm.n300 VSS 1.01985f
C11029 C9_P_btm.n301 VSS 1.01985f
C11030 C9_P_btm.n302 VSS 1.01629f
C11031 C9_P_btm.n303 VSS 1.01629f
C11032 C9_P_btm.n304 VSS 1.01629f
C11033 C9_P_btm.n305 VSS 1.01629f
C11034 C9_P_btm.n306 VSS 1.01629f
C11035 C9_P_btm.n307 VSS 1.01985f
C11036 C9_P_btm.n308 VSS 1.01629f
C11037 C9_P_btm.n309 VSS 1.01985f
C11038 C9_P_btm.n310 VSS 1.01985f
C11039 C9_P_btm.n311 VSS 1.01985f
C11040 C9_P_btm.n312 VSS 1.01985f
C11041 C9_P_btm.n313 VSS 1.01985f
C11042 C9_P_btm.n314 VSS 1.01985f
C11043 C9_P_btm.n315 VSS 1.01629f
C11044 C9_P_btm.n316 VSS 1.01629f
C11045 C9_P_btm.n317 VSS 1.01629f
C11046 C9_P_btm.n318 VSS 1.01629f
C11047 C9_P_btm.n319 VSS 1.01985f
C11048 C9_P_btm.n320 VSS 1.01985f
C11049 C9_P_btm.n321 VSS 1.01985f
C11050 C9_P_btm.n322 VSS 1.01985f
C11051 C9_P_btm.n323 VSS 1.01985f
C11052 C9_P_btm.n324 VSS 1.01985f
C11053 C9_P_btm.n325 VSS 1.01985f
C11054 C9_P_btm.n326 VSS 1.01985f
C11055 C9_P_btm.n327 VSS 1.01985f
C11056 C9_P_btm.n328 VSS 1.01985f
C11057 C9_P_btm.n329 VSS 1.01985f
C11058 C9_P_btm.n330 VSS 1.01985f
C11059 C9_P_btm.n331 VSS 1.01985f
C11060 C9_P_btm.n332 VSS 3.15708f
C11061 C9_P_btm.n333 VSS 4.45092f
C11062 C9_P_btm.n334 VSS 4.45099f
C11063 C9_P_btm.n335 VSS 1.01985f
C11064 C9_P_btm.n336 VSS 1.01985f
C11065 C9_P_btm.n337 VSS 1.01985f
C11066 C9_P_btm.n338 VSS 1.01985f
C11067 C9_P_btm.n339 VSS 1.01629f
C11068 C9_P_btm.n340 VSS 1.01629f
C11069 C9_P_btm.n341 VSS 1.01629f
C11070 C9_P_btm.n342 VSS 1.01629f
C11071 C9_P_btm.n343 VSS 1.01985f
C11072 C9_P_btm.n344 VSS 1.01985f
C11073 C9_P_btm.n345 VSS 1.01985f
C11074 C9_P_btm.n346 VSS 1.01985f
C11075 C9_P_btm.n347 VSS 1.01629f
C11076 C9_P_btm.n348 VSS 1.01629f
C11077 C9_P_btm.n349 VSS 1.01629f
C11078 C9_P_btm.n350 VSS 1.01629f
C11079 C9_P_btm.n351 VSS 1.01985f
C11080 C9_P_btm.n352 VSS 1.01985f
C11081 C9_P_btm.n353 VSS 1.01985f
C11082 C9_P_btm.n354 VSS 1.01985f
C11083 C9_P_btm.n355 VSS 1.01985f
C11084 C9_P_btm.n356 VSS 1.01985f
C11085 C9_P_btm.n357 VSS 1.01985f
C11086 C9_P_btm.n358 VSS 1.01985f
C11087 C9_P_btm.n359 VSS 1.01629f
C11088 C9_P_btm.n360 VSS 1.02004f
C11089 C9_P_btm.n361 VSS 1.01985f
C11090 C9_P_btm.n362 VSS 1.28218f
C11091 C9_P_btm.n363 VSS 1.01985f
C11092 C9_P_btm.n364 VSS 1.01985f
C11093 C9_P_btm.n365 VSS 1.01985f
C11094 C9_P_btm.n366 VSS 1.01985f
C11095 C9_P_btm.n367 VSS 1.28218f
C11096 C9_P_btm.n368 VSS 1.28218f
C11097 C9_P_btm.n369 VSS 1.28218f
C11098 C9_P_btm.n370 VSS 1.28218f
C11099 C9_P_btm.n371 VSS 1.01985f
C11100 C9_P_btm.n372 VSS 1.01985f
C11101 C9_P_btm.n373 VSS 1.01985f
C11102 C9_P_btm.n374 VSS 1.01985f
C11103 C9_P_btm.n375 VSS 1.01985f
C11104 C9_P_btm.n376 VSS 1.01985f
C11105 C9_P_btm.n377 VSS 1.01985f
C11106 C9_P_btm.n378 VSS 1.01985f
C11107 C9_P_btm.n379 VSS 0.750398f
C11108 C9_P_btm.n380 VSS 0.750398f
C11109 C9_P_btm.n381 VSS 0.750398f
C11110 C9_P_btm.n382 VSS 1.01985f
C11111 C9_P_btm.n383 VSS 1.01985f
C11112 C9_P_btm.n384 VSS 1.01985f
C11113 C9_P_btm.n385 VSS 1.01985f
C11114 C9_P_btm.n386 VSS 1.01985f
C11115 C9_P_btm.n387 VSS 1.01985f
C11116 C9_P_btm.n388 VSS 1.28218f
C11117 C9_P_btm.n389 VSS 1.28218f
C11118 C9_P_btm.n390 VSS 1.01985f
C11119 C9_P_btm.n391 VSS 0.984518f
C11120 C9_P_btm.n392 VSS 1.01985f
C11121 C9_P_btm.n393 VSS 1.01985f
C11122 C9_P_btm.n394 VSS 1.28218f
C11123 C9_P_btm.n395 VSS 1.28218f
C11124 C9_P_btm.n396 VSS 1.39221f
C11125 C9_P_btm.n397 VSS 1.01985f
C11126 C9_P_btm.n398 VSS 1.01985f
C11127 C9_P_btm.n399 VSS 1.01985f
C11128 C9_P_btm.n400 VSS 1.01985f
C11129 C9_P_btm.n401 VSS 1.01985f
C11130 C9_P_btm.n402 VSS 1.01985f
C11131 C9_P_btm.n403 VSS 1.01985f
C11132 C9_P_btm.n404 VSS 1.01985f
C11133 C9_P_btm.n405 VSS 1.01985f
C11134 C9_P_btm.n406 VSS 1.01985f
C11135 C9_P_btm.n407 VSS 2.48611f
C11136 C9_P_btm.n408 VSS 1.28218f
C11137 C9_P_btm.n409 VSS 1.28218f
C11138 C9_P_btm.n410 VSS 1.28218f
C11139 C9_P_btm.n411 VSS 1.01985f
C11140 C9_P_btm.n412 VSS 1.01985f
C11141 C9_P_btm.n413 VSS 1.01985f
C11142 C9_P_btm.n414 VSS 1.01985f
C11143 C9_P_btm.n415 VSS 1.01985f
C11144 C9_P_btm.n416 VSS 1.01985f
C11145 C9_P_btm.n417 VSS 1.01985f
C11146 C9_P_btm.n418 VSS 1.01985f
C11147 C9_P_btm.n419 VSS 1.01985f
C11148 C9_P_btm.n420 VSS 0.750398f
C11149 C9_P_btm.n421 VSS 0.750398f
C11150 C9_P_btm.n422 VSS 0.750398f
C11151 C9_P_btm.n423 VSS 0.750398f
C11152 C9_P_btm.n424 VSS 1.01985f
C11153 C9_P_btm.n425 VSS 1.01985f
C11154 C9_P_btm.n426 VSS 1.01985f
C11155 C9_P_btm.n427 VSS 1.01985f
C11156 C9_P_btm.n428 VSS 1.01985f
C11157 C9_P_btm.n429 VSS 1.01985f
C11158 C9_P_btm.n430 VSS 1.01985f
C11159 C9_P_btm.n431 VSS 1.01985f
C11160 C9_P_btm.n432 VSS 1.01985f
C11161 C9_P_btm.n433 VSS 0.984579f
C11162 C9_P_btm.n434 VSS 2.48618f
C11163 C9_P_btm.n435 VSS 1.28218f
C11164 C9_P_btm.n436 VSS 1.01985f
C11165 C9_P_btm.n437 VSS 1.01985f
C11166 C9_P_btm.n438 VSS 1.01985f
C11167 C9_P_btm.n439 VSS 1.01985f
C11168 C9_P_btm.n440 VSS 1.01985f
C11169 C9_P_btm.n441 VSS 1.01985f
C11170 C9_P_btm.n442 VSS 1.01985f
C11171 C9_P_btm.n443 VSS 1.28218f
C11172 C9_P_btm.n444 VSS 1.28218f
C11173 C9_P_btm.n445 VSS 1.28218f
C11174 C9_P_btm.n446 VSS 1.01985f
C11175 C9_P_btm.n447 VSS 1.01985f
C11176 C9_P_btm.n448 VSS 1.01985f
C11177 C9_P_btm.n449 VSS 1.28218f
C11178 C9_P_btm.n450 VSS 1.28218f
C11179 C9_P_btm.n451 VSS 1.28218f
C11180 C9_P_btm.n452 VSS 1.01985f
C11181 C9_P_btm.n453 VSS 1.01985f
C11182 C9_P_btm.n454 VSS 1.01985f
C11183 C9_P_btm.n455 VSS 1.01985f
C11184 C9_P_btm.n456 VSS 1.01985f
C11185 C9_P_btm.n457 VSS 1.01985f
C11186 C9_P_btm.n458 VSS 1.01985f
C11187 C9_P_btm.n459 VSS 1.01985f
C11188 C9_P_btm.n460 VSS 1.01985f
C11189 C9_P_btm.n461 VSS 1.01985f
C11190 C9_P_btm.n462 VSS 1.01985f
C11191 C9_P_btm.n463 VSS 1.01985f
C11192 C9_P_btm.n464 VSS 1.28218f
C11193 C9_P_btm.n465 VSS 1.28218f
C11194 C9_P_btm.n466 VSS 1.28218f
C11195 C9_P_btm.n467 VSS 1.01985f
C11196 C9_P_btm.n468 VSS 1.01985f
C11197 C9_P_btm.n469 VSS 1.01985f
C11198 C9_P_btm.n470 VSS 1.01985f
C11199 C9_P_btm.n471 VSS 1.01985f
C11200 C9_P_btm.n472 VSS 1.01985f
C11201 C9_P_btm.n473 VSS 1.01985f
C11202 C9_P_btm.n474 VSS 1.01985f
C11203 C9_P_btm.n475 VSS 0.575815f
C11204 C9_P_btm.n476 VSS 1.23713f
C11205 C9_P_btm.n477 VSS 0.750398f
C11206 C9_P_btm.n478 VSS 0.750398f
C11207 C9_P_btm.n479 VSS 0.750398f
C11208 C9_P_btm.n480 VSS 0.750398f
C11209 C9_P_btm.n481 VSS 0.750398f
C11210 C9_P_btm.n482 VSS 0.750398f
C11211 C9_P_btm.n483 VSS 1.01985f
C11212 C9_P_btm.n484 VSS 1.01985f
C11213 C9_P_btm.n485 VSS 1.01985f
C11214 C9_P_btm.n486 VSS 1.01985f
C11215 C9_P_btm.n487 VSS 1.01985f
C11216 C9_P_btm.n488 VSS 1.01985f
C11217 C9_P_btm.n489 VSS 1.01985f
C11218 C9_P_btm.n490 VSS 1.01985f
C11219 C9_P_btm.n491 VSS 1.01629f
C11220 C9_P_btm.n492 VSS 1.01985f
C11221 C9_P_btm.n493 VSS 1.01985f
C11222 C9_P_btm.n494 VSS 1.01985f
C11223 C9_P_btm.n495 VSS 1.01985f
C11224 C9_P_btm.n496 VSS 1.01629f
C11225 C9_P_btm.n497 VSS 1.01629f
C11226 C9_P_btm.n498 VSS 1.01629f
C11227 C9_P_btm.n499 VSS 1.01629f
C11228 C9_P_btm.n500 VSS 1.01985f
C11229 C9_P_btm.n501 VSS 1.01985f
C11230 C9_P_btm.n502 VSS 1.01985f
C11231 C9_P_btm.n503 VSS 1.01985f
C11232 C9_P_btm.n504 VSS 1.01629f
C11233 C9_P_btm.n505 VSS 1.01629f
C11234 C9_P_btm.n506 VSS 1.01629f
C11235 C9_P_btm.n507 VSS 1.01629f
C11236 C9_P_btm.n508 VSS 1.01985f
C11237 C9_P_btm.n509 VSS 1.01985f
C11238 C9_P_btm.n510 VSS 1.01985f
C11239 C9_P_btm.n511 VSS 1.01985f
C11240 C9_P_btm.n512 VSS 1.01629f
C11241 C9_P_btm.n513 VSS 2.28426f
C11242 a_4958_30871.t3 VSS 0.02704f
C11243 a_4958_30871.t2 VSS 0.02704f
C11244 a_4958_30871.n0 VSS 0.10014f
C11245 a_4958_30871.t4 VSS 0.547724f
C11246 a_4958_30871.t12 VSS 0.564055f
C11247 a_4958_30871.n1 VSS 0.497511f
C11248 a_4958_30871.t6 VSS 0.547724f
C11249 a_4958_30871.t13 VSS 0.548649f
C11250 a_4958_30871.n2 VSS 0.251771f
C11251 a_4958_30871.n3 VSS 0.270725f
C11252 a_4958_30871.n4 VSS 1.67307f
C11253 a_4958_30871.t10 VSS 0.547724f
C11254 a_4958_30871.n5 VSS 0.270725f
C11255 a_4958_30871.t7 VSS 0.547724f
C11256 a_4958_30871.t11 VSS 0.548649f
C11257 a_4958_30871.n6 VSS 0.251771f
C11258 a_4958_30871.t8 VSS 0.564055f
C11259 a_4958_30871.n7 VSS 0.497511f
C11260 a_4958_30871.n8 VSS 1.81725f
C11261 a_4958_30871.n9 VSS 6.81446f
C11262 a_4958_30871.t9 VSS 0.064711f
C11263 a_4958_30871.t5 VSS 0.040358f
C11264 a_4958_30871.n10 VSS 0.167042f
C11265 a_4958_30871.n11 VSS 4.61925f
C11266 a_4958_30871.n12 VSS 0.42689f
C11267 a_4958_30871.t0 VSS 0.041599f
C11268 a_4958_30871.n13 VSS 0.083232f
C11269 a_4958_30871.t1 VSS 0.041599f
C11270 a_n971_45724.t0 VSS 0.016532f
C11271 a_n971_45724.t24 VSS 0.022191f
C11272 a_n971_45724.t18 VSS 0.015085f
C11273 a_n971_45724.n0 VSS 0.128881f
C11274 a_n971_45724.t28 VSS 0.0189f
C11275 a_n971_45724.t15 VSS 0.015265f
C11276 a_n971_45724.n1 VSS 0.107761f
C11277 a_n971_45724.t7 VSS 0.012169f
C11278 a_n971_45724.t26 VSS 0.022135f
C11279 a_n971_45724.n2 VSS 0.041341f
C11280 a_n971_45724.n3 VSS 0.134941f
C11281 a_n971_45724.n4 VSS 1.2489f
C11282 a_n971_45724.t4 VSS 0.017495f
C11283 a_n971_45724.t27 VSS 0.027861f
C11284 a_n971_45724.n5 VSS 0.04447f
C11285 a_n971_45724.t17 VSS 0.0112f
C11286 a_n971_45724.t9 VSS 0.012005f
C11287 a_n971_45724.n6 VSS 0.036846f
C11288 a_n971_45724.n7 VSS 0.332438f
C11289 a_n971_45724.t12 VSS 0.011813f
C11290 a_n971_45724.t5 VSS 0.011031f
C11291 a_n971_45724.n8 VSS 0.046519f
C11292 a_n971_45724.n9 VSS 0.397644f
C11293 a_n971_45724.n10 VSS 0.774569f
C11294 a_n971_45724.t19 VSS 0.015265f
C11295 a_n971_45724.t22 VSS 0.0189f
C11296 a_n971_45724.n11 VSS 0.107761f
C11297 a_n971_45724.t13 VSS 0.022135f
C11298 a_n971_45724.t14 VSS 0.012169f
C11299 a_n971_45724.n12 VSS 0.041341f
C11300 a_n971_45724.n13 VSS 0.140388f
C11301 a_n971_45724.n14 VSS 0.377129f
C11302 a_n971_45724.t29 VSS 0.015265f
C11303 a_n971_45724.t8 VSS 0.0189f
C11304 a_n971_45724.n15 VSS 0.107761f
C11305 a_n971_45724.t23 VSS 0.022135f
C11306 a_n971_45724.t20 VSS 0.012169f
C11307 a_n971_45724.n16 VSS 0.041341f
C11308 a_n971_45724.n17 VSS 0.134941f
C11309 a_n971_45724.n18 VSS 0.557982f
C11310 a_n971_45724.t25 VSS 0.027635f
C11311 a_n971_45724.t6 VSS 0.01731f
C11312 a_n971_45724.n19 VSS 0.044345f
C11313 a_n971_45724.n20 VSS 0.688064f
C11314 a_n971_45724.t16 VSS 0.028637f
C11315 a_n971_45724.t21 VSS 0.017216f
C11316 a_n971_45724.n21 VSS 0.057296f
C11317 a_n971_45724.n22 VSS 0.611138f
C11318 a_n971_45724.t10 VSS 0.027861f
C11319 a_n971_45724.t11 VSS 0.017495f
C11320 a_n971_45724.n23 VSS 0.049713f
C11321 a_n971_45724.n24 VSS 0.142308f
C11322 a_n971_45724.t3 VSS 0.010746f
C11323 a_n971_45724.t2 VSS 0.010746f
C11324 a_n971_45724.n25 VSS 0.021492f
C11325 a_n971_45724.n26 VSS 0.108285f
C11326 a_n971_45724.n27 VSS 0.049609f
C11327 a_n971_45724.t1 VSS 0.016532f
C11328 a_11599_46634.t4 VSS 0.015208f
C11329 a_11599_46634.t2 VSS 0.015208f
C11330 a_11599_46634.t9 VSS 0.015208f
C11331 a_11599_46634.n0 VSS 0.038632f
C11332 a_11599_46634.t7 VSS 0.015208f
C11333 a_11599_46634.t12 VSS 0.015208f
C11334 a_11599_46634.n1 VSS 0.032056f
C11335 a_11599_46634.n2 VSS 0.146088f
C11336 a_11599_46634.n3 VSS 0.022681f
C11337 a_11599_46634.n4 VSS 0.014581f
C11338 a_11599_46634.n5 VSS 0.092134f
C11339 a_11599_46634.n6 VSS 0.014581f
C11340 a_11599_46634.n7 VSS 0.05538f
C11341 a_11599_46634.n8 VSS 0.01459f
C11342 a_11599_46634.n9 VSS 0.057125f
C11343 a_11599_46634.n10 VSS 0.014581f
C11344 a_11599_46634.n11 VSS 0.05538f
C11345 a_11599_46634.n12 VSS 0.014581f
C11346 a_11599_46634.n13 VSS 0.055657f
C11347 a_11599_46634.n14 VSS 0.014581f
C11348 a_11599_46634.n15 VSS 0.047808f
C11349 a_11599_46634.n16 VSS 0.014029f
C11350 a_11599_46634.t32 VSS 0.015926f
C11351 a_11599_46634.t35 VSS 0.023804f
C11352 a_11599_46634.n17 VSS 0.04837f
C11353 a_11599_46634.t34 VSS 0.023804f
C11354 a_11599_46634.t49 VSS 0.015926f
C11355 a_11599_46634.n18 VSS 0.050358f
C11356 a_11599_46634.t47 VSS 0.023804f
C11357 a_11599_46634.t43 VSS 0.015926f
C11358 a_11599_46634.n19 VSS 0.048306f
C11359 a_11599_46634.t36 VSS 0.023804f
C11360 a_11599_46634.t41 VSS 0.015926f
C11361 a_11599_46634.n20 VSS 0.05765f
C11362 a_11599_46634.n21 VSS 0.406193f
C11363 a_11599_46634.n22 VSS 0.306573f
C11364 a_11599_46634.n23 VSS 0.329864f
C11365 a_11599_46634.t39 VSS 0.015926f
C11366 a_11599_46634.t37 VSS 0.023804f
C11367 a_11599_46634.n24 VSS 0.04861f
C11368 a_11599_46634.t40 VSS 0.023804f
C11369 a_11599_46634.t46 VSS 0.015926f
C11370 a_11599_46634.n25 VSS 0.046432f
C11371 a_11599_46634.t45 VSS 0.023804f
C11372 a_11599_46634.t44 VSS 0.015926f
C11373 a_11599_46634.n26 VSS 0.046547f
C11374 a_11599_46634.n27 VSS 0.272214f
C11375 a_11599_46634.n28 VSS 0.508784f
C11376 a_11599_46634.t38 VSS 0.015926f
C11377 a_11599_46634.t42 VSS 0.023804f
C11378 a_11599_46634.n29 VSS 0.054859f
C11379 a_11599_46634.t48 VSS 0.023804f
C11380 a_11599_46634.t33 VSS 0.015926f
C11381 a_11599_46634.n30 VSS 0.049498f
C11382 a_11599_46634.n31 VSS 0.415496f
C11383 a_11599_46634.n32 VSS 0.313667f
C11384 a_11599_46634.n33 VSS 0.29198f
C11385 a_11599_46634.t3 VSS 0.015208f
C11386 a_11599_46634.t10 VSS 0.015208f
C11387 a_11599_46634.n34 VSS 0.031412f
C11388 a_11599_46634.n35 VSS 0.14228f
C11389 a_11599_46634.n36 VSS 0.086499f
C11390 a_11599_46634.n37 VSS 0.06822f
C11391 a_11599_46634.t5 VSS 0.015208f
C11392 a_11599_46634.t1 VSS 0.015208f
C11393 a_11599_46634.n38 VSS 0.032056f
C11394 a_11599_46634.n39 VSS 0.072522f
C11395 a_11599_46634.t6 VSS 0.015208f
C11396 a_11599_46634.t13 VSS 0.015208f
C11397 a_11599_46634.n40 VSS 0.032056f
C11398 a_11599_46634.n41 VSS 0.084153f
C11399 a_11599_46634.t11 VSS 0.015208f
C11400 a_11599_46634.t0 VSS 0.015208f
C11401 a_11599_46634.n42 VSS 0.032056f
C11402 a_11599_46634.n43 VSS 0.083762f
C11403 a_11599_46634.t8 VSS 0.015208f
C11404 a_11599_46634.t14 VSS 0.015208f
C11405 a_11599_46634.n44 VSS 0.032056f
C11406 a_11599_46634.n45 VSS 0.083762f
C11407 a_11599_46634.n46 VSS 0.084153f
C11408 a_11599_46634.n47 VSS 0.032056f
C11409 a_11599_46634.t15 VSS 0.015208f
C11410 a_n4209_39590.t1 VSS 0.020737f
C11411 a_n4209_39590.t7 VSS 0.013479f
C11412 a_n4209_39590.t6 VSS 0.013479f
C11413 a_n4209_39590.n0 VSS 0.051465f
C11414 a_n4209_39590.t5 VSS 0.013479f
C11415 a_n4209_39590.t4 VSS 0.013479f
C11416 a_n4209_39590.n1 VSS 0.030592f
C11417 a_n4209_39590.n2 VSS 0.15047f
C11418 a_n4209_39590.t14 VSS 0.034947f
C11419 a_n4209_39590.t10 VSS 0.021945f
C11420 a_n4209_39590.n3 VSS 0.073397f
C11421 a_n4209_39590.t8 VSS 0.702048f
C11422 a_n4209_39590.t16 VSS 0.701939f
C11423 a_n4209_39590.n4 VSS 0.520753f
C11424 a_n4209_39590.t9 VSS 0.701939f
C11425 a_n4209_39590.n5 VSS 0.263887f
C11426 a_n4209_39590.t17 VSS 0.701939f
C11427 a_n4209_39590.n6 VSS 0.263887f
C11428 a_n4209_39590.t12 VSS 0.701939f
C11429 a_n4209_39590.n7 VSS 0.263887f
C11430 a_n4209_39590.t13 VSS 0.701939f
C11431 a_n4209_39590.n8 VSS 0.263887f
C11432 a_n4209_39590.t15 VSS 0.701939f
C11433 a_n4209_39590.n9 VSS 0.26301f
C11434 a_n4209_39590.t11 VSS 0.701941f
C11435 a_n4209_39590.n10 VSS 2.04036f
C11436 a_n4209_39590.n11 VSS 2.23805f
C11437 a_n4209_39590.n12 VSS 0.0855f
C11438 a_n4209_39590.t2 VSS 0.020737f
C11439 a_n4209_39590.t0 VSS 0.020737f
C11440 a_n4209_39590.n13 VSS 0.042659f
C11441 a_n4209_39590.n14 VSS 0.186037f
C11442 a_n4209_39590.n15 VSS 0.052777f
C11443 a_n4209_39590.t3 VSS 0.020737f
C11444 a_11967_42832.n0 VSS 0.011068f
C11445 a_11967_42832.n2 VSS 0.044961f
C11446 a_11967_42832.n4 VSS 0.027025f
C11447 a_11967_42832.n6 VSS 0.027877f
C11448 a_11967_42832.n8 VSS 0.027025f
C11449 a_11967_42832.n10 VSS 0.02716f
C11450 a_11967_42832.n12 VSS 0.02333f
C11451 a_11967_42832.n14 VSS 0.025775f
C11452 a_11967_42832.t47 VSS 0.011132f
C11453 a_11967_42832.t33 VSS 0.011132f
C11454 a_11967_42832.n15 VSS 0.018678f
C11455 a_11967_42832.n16 VSS 0.02818f
C11456 a_11967_42832.t40 VSS 0.011616f
C11457 a_11967_42832.n17 VSS 0.022659f
C11458 a_11967_42832.n18 VSS 0.139616f
C11459 a_11967_42832.t41 VSS 0.011616f
C11460 a_11967_42832.n19 VSS 0.023573f
C11461 a_11967_42832.n20 VSS 0.181535f
C11462 a_11967_42832.t32 VSS 0.011616f
C11463 a_11967_42832.n21 VSS 0.022693f
C11464 a_11967_42832.t44 VSS 0.011616f
C11465 a_11967_42832.n22 VSS 0.025698f
C11466 a_11967_42832.t38 VSS 0.011616f
C11467 a_11967_42832.n23 VSS 0.022659f
C11468 a_11967_42832.t43 VSS 0.011616f
C11469 a_11967_42832.n24 VSS 0.023047f
C11470 a_11967_42832.n25 VSS 0.229661f
C11471 a_11967_42832.n26 VSS 0.263153f
C11472 a_11967_42832.t45 VSS 0.011616f
C11473 a_11967_42832.n27 VSS 0.029549f
C11474 a_11967_42832.n28 VSS 0.187675f
C11475 a_11967_42832.n29 VSS 0.112002f
C11476 a_11967_42832.n30 VSS 0.194593f
C11477 a_11967_42832.n31 VSS 0.087866f
C11478 a_11967_42832.n32 VSS 0.015433f
C11479 a_11967_42832.n33 VSS 0.084896f
C11480 a_11967_42832.n34 VSS 0.015643f
C11481 a_11967_42832.n35 VSS 0.03539f
C11482 a_11967_42832.n36 VSS 0.015643f
C11483 a_11967_42832.n37 VSS 0.041066f
C11484 a_11967_42832.n38 VSS 0.015643f
C11485 a_11967_42832.n39 VSS 0.040875f
C11486 a_11967_42832.n40 VSS 0.015643f
C11487 a_11967_42832.n41 VSS 0.040875f
C11488 a_11967_42832.n42 VSS 0.015643f
C11489 a_11967_42832.n43 VSS 0.041066f
C11490 a_11967_42832.n44 VSS 0.015643f
C11491 a_11967_42832.n45 VSS 0.07129f
C11492 a_11967_42832.n46 VSS 0.018852f
C11493 VCM.t22 VSS 0.212736f
C11494 VCM.t61 VSS 0.209711f
C11495 VCM.n0 VSS 0.697234f
C11496 VCM.t19 VSS 0.209711f
C11497 VCM.n1 VSS 0.369146f
C11498 VCM.t0 VSS 0.209711f
C11499 VCM.n2 VSS 0.369146f
C11500 VCM.t20 VSS 0.209711f
C11501 VCM.n3 VSS 0.369146f
C11502 VCM.t43 VSS 0.209711f
C11503 VCM.n4 VSS 0.369146f
C11504 VCM.t25 VSS 0.055783f
C11505 VCM.t62 VSS 0.055783f
C11506 VCM.n5 VSS 0.15224f
C11507 VCM.n6 VSS 0.323503f
C11508 VCM.t27 VSS 0.209711f
C11509 VCM.n7 VSS 0.893101f
C11510 VCM.t28 VSS 0.223132f
C11511 VCM.t41 VSS 0.223132f
C11512 VCM.n8 VSS 0.926112f
C11513 VCM.t33 VSS 0.223132f
C11514 VCM.t29 VSS 0.223132f
C11515 VCM.n9 VSS 0.904283f
C11516 VCM.n10 VSS 1.8485f
C11517 VCM.t32 VSS 0.223132f
C11518 VCM.t39 VSS 0.223132f
C11519 VCM.n11 VSS 0.904283f
C11520 VCM.n12 VSS 0.702776f
C11521 VCM.t9 VSS 0.223132f
C11522 VCM.t38 VSS 0.223132f
C11523 VCM.n13 VSS 0.904283f
C11524 VCM.n14 VSS 0.704698f
C11525 VCM.t6 VSS 0.223132f
C11526 VCM.t3 VSS 0.223132f
C11527 VCM.n15 VSS 0.904283f
C11528 VCM.n16 VSS 0.704698f
C11529 VCM.t7 VSS 0.223132f
C11530 VCM.t2 VSS 0.223132f
C11531 VCM.n17 VSS 0.904283f
C11532 VCM.n18 VSS 0.703008f
C11533 VCM.t5 VSS 0.223132f
C11534 VCM.t4 VSS 0.223132f
C11535 VCM.n19 VSS 0.904283f
C11536 VCM.n20 VSS 0.703008f
C11537 VCM.t47 VSS 0.223132f
C11538 VCM.t8 VSS 0.223132f
C11539 VCM.n21 VSS 0.904283f
C11540 VCM.n22 VSS 0.704698f
C11541 VCM.t46 VSS 0.223132f
C11542 VCM.t52 VSS 0.223132f
C11543 VCM.n23 VSS 0.904283f
C11544 VCM.n24 VSS 0.704698f
C11545 VCM.t59 VSS 0.223132f
C11546 VCM.t45 VSS 0.223132f
C11547 VCM.n25 VSS 0.904283f
C11548 VCM.n26 VSS 0.703008f
C11549 VCM.t50 VSS 0.223132f
C11550 VCM.t51 VSS 0.223132f
C11551 VCM.n27 VSS 0.904283f
C11552 VCM.n28 VSS 0.703008f
C11553 VCM.t54 VSS 1.14389f
C11554 VCM.n29 VSS 8.814361f
C11555 VCM.t40 VSS 0.223132f
C11556 VCM.t31 VSS 0.223132f
C11557 VCM.n30 VSS 0.926112f
C11558 VCM.t23 VSS 0.212736f
C11559 VCM.t60 VSS 0.209711f
C11560 VCM.n31 VSS 0.697234f
C11561 VCM.t18 VSS 0.209711f
C11562 VCM.n32 VSS 0.369146f
C11563 VCM.t1 VSS 0.209711f
C11564 VCM.n33 VSS 0.369146f
C11565 VCM.t21 VSS 0.209711f
C11566 VCM.n34 VSS 0.369146f
C11567 VCM.t42 VSS 0.209711f
C11568 VCM.n35 VSS 0.369146f
C11569 VCM.t63 VSS 0.055783f
C11570 VCM.t24 VSS 0.055783f
C11571 VCM.n36 VSS 0.15224f
C11572 VCM.n37 VSS 0.323503f
C11573 VCM.t26 VSS 0.209711f
C11574 VCM.n38 VSS 0.893101f
C11575 VCM.t30 VSS 0.223132f
C11576 VCM.t36 VSS 0.223132f
C11577 VCM.n39 VSS 0.904283f
C11578 VCM.n40 VSS 1.8485f
C11579 VCM.t37 VSS 0.223132f
C11580 VCM.t34 VSS 0.223132f
C11581 VCM.n41 VSS 0.904283f
C11582 VCM.n42 VSS 0.702776f
C11583 VCM.t35 VSS 0.223132f
C11584 VCM.t15 VSS 0.223132f
C11585 VCM.n43 VSS 0.904283f
C11586 VCM.n44 VSS 0.704698f
C11587 VCM.t12 VSS 0.223132f
C11588 VCM.t10 VSS 0.223132f
C11589 VCM.n45 VSS 0.904283f
C11590 VCM.n46 VSS 0.704698f
C11591 VCM.t13 VSS 0.223132f
C11592 VCM.t11 VSS 0.223132f
C11593 VCM.n47 VSS 0.904283f
C11594 VCM.n48 VSS 0.703008f
C11595 VCM.t14 VSS 0.223132f
C11596 VCM.t17 VSS 0.223132f
C11597 VCM.n49 VSS 0.904283f
C11598 VCM.n50 VSS 0.703008f
C11599 VCM.t16 VSS 0.223132f
C11600 VCM.t58 VSS 0.223132f
C11601 VCM.n51 VSS 0.904283f
C11602 VCM.n52 VSS 0.704698f
C11603 VCM.t55 VSS 0.223132f
C11604 VCM.t57 VSS 0.223132f
C11605 VCM.n53 VSS 0.904283f
C11606 VCM.n54 VSS 0.704698f
C11607 VCM.t44 VSS 0.223132f
C11608 VCM.t56 VSS 0.223132f
C11609 VCM.n55 VSS 0.904283f
C11610 VCM.n56 VSS 0.703008f
C11611 VCM.t49 VSS 0.223132f
C11612 VCM.t48 VSS 0.223132f
C11613 VCM.n57 VSS 0.904283f
C11614 VCM.n58 VSS 0.703008f
C11615 VCM.t53 VSS 1.14389f
C11616 VCM.n59 VSS 8.85736f
C11617 C10_N_btm.t12 VSS 0.122926f
C11618 C10_N_btm.t14 VSS 0.122926f
C11619 C10_N_btm.n0 VSS 0.39276f
C11620 C10_N_btm.t18 VSS 0.122926f
C11621 C10_N_btm.t20 VSS 0.122926f
C11622 C10_N_btm.n1 VSS 0.379868f
C11623 C10_N_btm.n2 VSS 1.19496f
C11624 C10_N_btm.t15 VSS 0.122926f
C11625 C10_N_btm.t8 VSS 0.122926f
C11626 C10_N_btm.n3 VSS 0.379868f
C11627 C10_N_btm.n4 VSS 0.613462f
C11628 C10_N_btm.t11 VSS 0.122926f
C11629 C10_N_btm.t21 VSS 0.122926f
C11630 C10_N_btm.n5 VSS 0.379868f
C11631 C10_N_btm.n6 VSS 0.613462f
C11632 C10_N_btm.t23 VSS 0.122926f
C11633 C10_N_btm.t19 VSS 0.122926f
C11634 C10_N_btm.n7 VSS 0.379868f
C11635 C10_N_btm.n8 VSS 0.613462f
C11636 C10_N_btm.t13 VSS 0.122926f
C11637 C10_N_btm.t16 VSS 0.122926f
C11638 C10_N_btm.n9 VSS 0.379868f
C11639 C10_N_btm.n10 VSS 0.613462f
C11640 C10_N_btm.t22 VSS 0.122926f
C11641 C10_N_btm.t17 VSS 0.122926f
C11642 C10_N_btm.n11 VSS 0.379868f
C11643 C10_N_btm.n12 VSS 0.612599f
C11644 C10_N_btm.t10 VSS 0.122926f
C11645 C10_N_btm.t9 VSS 0.122926f
C11646 C10_N_btm.n13 VSS 0.379868f
C11647 C10_N_btm.n14 VSS 1.05453f
C11648 C10_N_btm.t27 VSS 0.139882f
C11649 C10_N_btm.t30 VSS 0.139882f
C11650 C10_N_btm.n15 VSS 0.57718f
C11651 C10_N_btm.t29 VSS 0.139882f
C11652 C10_N_btm.t24 VSS 0.139882f
C11653 C10_N_btm.n16 VSS 0.563454f
C11654 C10_N_btm.n17 VSS 0.84522f
C11655 C10_N_btm.t25 VSS 0.139882f
C11656 C10_N_btm.t26 VSS 0.139882f
C11657 C10_N_btm.n18 VSS 0.563454f
C11658 C10_N_btm.n19 VSS 0.434278f
C11659 C10_N_btm.t31 VSS 0.139882f
C11660 C10_N_btm.t28 VSS 0.139882f
C11661 C10_N_btm.n20 VSS 0.563454f
C11662 C10_N_btm.n21 VSS 0.493206f
C11663 C10_N_btm.n22 VSS 0.690049f
C11664 C10_N_btm.t32 VSS 0.139882f
C11665 C10_N_btm.t33 VSS 0.139882f
C11666 C10_N_btm.n23 VSS 0.69103f
C11667 C10_N_btm.n24 VSS 0.588284f
C11668 C10_N_btm.t6 VSS 0.139882f
C11669 C10_N_btm.t3 VSS 0.139882f
C11670 C10_N_btm.n25 VSS 0.569903f
C11671 C10_N_btm.t1 VSS 0.139882f
C11672 C10_N_btm.t7 VSS 0.139882f
C11673 C10_N_btm.n26 VSS 0.583821f
C11674 C10_N_btm.t0 VSS 0.139882f
C11675 C10_N_btm.t4 VSS 0.139882f
C11676 C10_N_btm.n27 VSS 0.569903f
C11677 C10_N_btm.n28 VSS 0.861377f
C11678 C10_N_btm.t2 VSS 0.139882f
C11679 C10_N_btm.t5 VSS 0.139882f
C11680 C10_N_btm.n29 VSS 0.569903f
C11681 C10_N_btm.n30 VSS 0.443544f
C11682 C10_N_btm.n31 VSS 0.497297f
C11683 C10_N_btm.n32 VSS 2.46311f
C11684 C10_N_btm.n33 VSS 2.05041f
C11685 C10_N_btm.n34 VSS 0.908086f
C11686 C10_N_btm.n35 VSS 0.911266f
C11687 C10_N_btm.n36 VSS 0.911266f
C11688 C10_N_btm.n37 VSS 0.908086f
C11689 C10_N_btm.n38 VSS 0.911266f
C11690 C10_N_btm.n39 VSS 0.911266f
C11691 C10_N_btm.n40 VSS 0.911266f
C11692 C10_N_btm.n41 VSS 0.911266f
C11693 C10_N_btm.n42 VSS 0.908086f
C11694 C10_N_btm.n43 VSS 0.911266f
C11695 C10_N_btm.n44 VSS 0.911266f
C11696 C10_N_btm.n45 VSS 0.908086f
C11697 C10_N_btm.n46 VSS 0.911266f
C11698 C10_N_btm.n47 VSS 0.911266f
C11699 C10_N_btm.n48 VSS 0.911266f
C11700 C10_N_btm.n49 VSS 0.911266f
C11701 C10_N_btm.n50 VSS 0.908086f
C11702 C10_N_btm.n51 VSS 0.911266f
C11703 C10_N_btm.n52 VSS 0.911266f
C11704 C10_N_btm.n53 VSS 0.908086f
C11705 C10_N_btm.n54 VSS 0.911266f
C11706 C10_N_btm.n55 VSS 0.911266f
C11707 C10_N_btm.n56 VSS 0.911266f
C11708 C10_N_btm.n57 VSS 0.911266f
C11709 C10_N_btm.n58 VSS 0.908086f
C11710 C10_N_btm.n59 VSS 0.911266f
C11711 C10_N_btm.n60 VSS 0.911266f
C11712 C10_N_btm.n61 VSS 0.908086f
C11713 C10_N_btm.n62 VSS 0.911266f
C11714 C10_N_btm.n63 VSS 0.911266f
C11715 C10_N_btm.n64 VSS 0.911266f
C11716 C10_N_btm.n65 VSS 1.1455f
C11717 C10_N_btm.n66 VSS 0.911266f
C11718 C10_N_btm.n67 VSS 0.911266f
C11719 C10_N_btm.n68 VSS 0.911266f
C11720 C10_N_btm.n69 VSS 0.911266f
C11721 C10_N_btm.n70 VSS 0.911266f
C11722 C10_N_btm.n71 VSS 0.911266f
C11723 C10_N_btm.n72 VSS 0.911266f
C11724 C10_N_btm.n73 VSS 0.911266f
C11725 C10_N_btm.n74 VSS 0.911266f
C11726 C10_N_btm.n75 VSS 0.911266f
C11727 C10_N_btm.n76 VSS 0.911266f
C11728 C10_N_btm.n77 VSS 0.911266f
C11729 C10_N_btm.n78 VSS 0.911266f
C11730 C10_N_btm.n79 VSS 0.911266f
C11731 C10_N_btm.n80 VSS 0.911266f
C11732 C10_N_btm.n81 VSS 0.911266f
C11733 C10_N_btm.n82 VSS 0.911266f
C11734 C10_N_btm.n83 VSS 0.911266f
C11735 C10_N_btm.n84 VSS 0.911266f
C11736 C10_N_btm.n85 VSS 0.911266f
C11737 C10_N_btm.n86 VSS 0.911266f
C11738 C10_N_btm.n87 VSS 0.911266f
C11739 C10_N_btm.n88 VSS 0.911266f
C11740 C10_N_btm.n89 VSS 0.911266f
C11741 C10_N_btm.n90 VSS 0.911266f
C11742 C10_N_btm.n91 VSS 0.911266f
C11743 C10_N_btm.n92 VSS 0.911266f
C11744 C10_N_btm.n93 VSS 0.911266f
C11745 C10_N_btm.n94 VSS 0.911266f
C11746 C10_N_btm.n95 VSS 0.911266f
C11747 C10_N_btm.n96 VSS 0.911266f
C11748 C10_N_btm.n97 VSS 0.911266f
C11749 C10_N_btm.n98 VSS 0.911266f
C11750 C10_N_btm.n99 VSS 0.911266f
C11751 C10_N_btm.n100 VSS 0.911266f
C11752 C10_N_btm.n101 VSS 0.911266f
C11753 C10_N_btm.n102 VSS 0.911266f
C11754 C10_N_btm.n103 VSS 0.911266f
C11755 C10_N_btm.n104 VSS 0.911266f
C11756 C10_N_btm.n105 VSS 0.911266f
C11757 C10_N_btm.n106 VSS 0.911266f
C11758 C10_N_btm.n107 VSS 0.911266f
C11759 C10_N_btm.n108 VSS 0.911266f
C11760 C10_N_btm.n109 VSS 0.911266f
C11761 C10_N_btm.n110 VSS 0.911266f
C11762 C10_N_btm.n111 VSS 0.911266f
C11763 C10_N_btm.n112 VSS 0.911266f
C11764 C10_N_btm.n113 VSS 0.911266f
C11765 C10_N_btm.n114 VSS 0.911266f
C11766 C10_N_btm.n115 VSS 0.911266f
C11767 C10_N_btm.n116 VSS 0.911266f
C11768 C10_N_btm.n117 VSS 0.911266f
C11769 C10_N_btm.n118 VSS 0.911266f
C11770 C10_N_btm.n119 VSS 0.911266f
C11771 C10_N_btm.n120 VSS 0.911266f
C11772 C10_N_btm.n121 VSS 0.911266f
C11773 C10_N_btm.n122 VSS 0.911266f
C11774 C10_N_btm.n123 VSS 0.911266f
C11775 C10_N_btm.n124 VSS 0.911266f
C11776 C10_N_btm.n125 VSS 0.911266f
C11777 C10_N_btm.n126 VSS 0.911266f
C11778 C10_N_btm.n127 VSS 0.911266f
C11779 C10_N_btm.n128 VSS 2.05041f
C11780 C10_N_btm.n129 VSS 2.05041f
C11781 C10_N_btm.n130 VSS 0.911266f
C11782 C10_N_btm.n131 VSS 3.97683f
C11783 C10_N_btm.n132 VSS 0.911266f
C11784 C10_N_btm.n133 VSS 0.911266f
C11785 C10_N_btm.n134 VSS 0.911266f
C11786 C10_N_btm.n135 VSS 0.911266f
C11787 C10_N_btm.n136 VSS 0.911266f
C11788 C10_N_btm.n137 VSS 0.911266f
C11789 C10_N_btm.n138 VSS 0.911266f
C11790 C10_N_btm.n139 VSS 0.911266f
C11791 C10_N_btm.n140 VSS 0.911266f
C11792 C10_N_btm.n141 VSS 0.911266f
C11793 C10_N_btm.n142 VSS 0.911266f
C11794 C10_N_btm.n143 VSS 0.911266f
C11795 C10_N_btm.n144 VSS 0.911266f
C11796 C10_N_btm.n145 VSS 0.911266f
C11797 C10_N_btm.n146 VSS 0.911266f
C11798 C10_N_btm.n147 VSS 0.911266f
C11799 C10_N_btm.n148 VSS 0.911266f
C11800 C10_N_btm.n149 VSS 0.911266f
C11801 C10_N_btm.n150 VSS 0.911266f
C11802 C10_N_btm.n151 VSS 0.911266f
C11803 C10_N_btm.n152 VSS 0.911266f
C11804 C10_N_btm.n153 VSS 0.911266f
C11805 C10_N_btm.n154 VSS 0.911266f
C11806 C10_N_btm.n155 VSS 0.911266f
C11807 C10_N_btm.n156 VSS 0.911266f
C11808 C10_N_btm.n157 VSS 0.911266f
C11809 C10_N_btm.n158 VSS 0.911266f
C11810 C10_N_btm.n159 VSS 0.911266f
C11811 C10_N_btm.n160 VSS 0.911266f
C11812 C10_N_btm.n161 VSS 0.911266f
C11813 C10_N_btm.n162 VSS 0.911266f
C11814 C10_N_btm.n163 VSS 0.911266f
C11815 C10_N_btm.n164 VSS 0.911266f
C11816 C10_N_btm.n165 VSS 0.911266f
C11817 C10_N_btm.n166 VSS 0.911266f
C11818 C10_N_btm.n167 VSS 0.911266f
C11819 C10_N_btm.n168 VSS 0.911266f
C11820 C10_N_btm.n169 VSS 0.911266f
C11821 C10_N_btm.n170 VSS 0.911266f
C11822 C10_N_btm.n171 VSS 0.911266f
C11823 C10_N_btm.n172 VSS 0.911266f
C11824 C10_N_btm.n173 VSS 0.911266f
C11825 C10_N_btm.n174 VSS 0.911266f
C11826 C10_N_btm.n175 VSS 0.911266f
C11827 C10_N_btm.n176 VSS 0.911266f
C11828 C10_N_btm.n177 VSS 0.911266f
C11829 C10_N_btm.n178 VSS 0.911435f
C11830 C10_N_btm.n179 VSS 0.911266f
C11831 C10_N_btm.n180 VSS 0.911435f
C11832 C10_N_btm.n181 VSS 2.82097f
C11833 C10_N_btm.n182 VSS 1.16658f
C11834 C10_N_btm.n183 VSS 0.908086f
C11835 C10_N_btm.n184 VSS 0.911266f
C11836 C10_N_btm.n185 VSS 0.908086f
C11837 C10_N_btm.n186 VSS 0.908086f
C11838 C10_N_btm.n187 VSS 0.908086f
C11839 C10_N_btm.n188 VSS 0.908086f
C11840 C10_N_btm.n189 VSS 0.911266f
C11841 C10_N_btm.n190 VSS 0.908086f
C11842 C10_N_btm.n191 VSS 0.908086f
C11843 C10_N_btm.n192 VSS 0.908086f
C11844 C10_N_btm.n193 VSS 0.908086f
C11845 C10_N_btm.n194 VSS 0.911266f
C11846 C10_N_btm.n195 VSS 0.908086f
C11847 C10_N_btm.n196 VSS 0.908086f
C11848 C10_N_btm.n197 VSS 0.908086f
C11849 C10_N_btm.n198 VSS 0.908086f
C11850 C10_N_btm.n199 VSS 0.911266f
C11851 C10_N_btm.n200 VSS 0.908086f
C11852 C10_N_btm.n201 VSS 0.908086f
C11853 C10_N_btm.n202 VSS 0.908086f
C11854 C10_N_btm.n203 VSS 0.908086f
C11855 C10_N_btm.n204 VSS 0.911266f
C11856 C10_N_btm.n205 VSS 0.908086f
C11857 C10_N_btm.n206 VSS 0.908086f
C11858 C10_N_btm.n207 VSS 0.908086f
C11859 C10_N_btm.n208 VSS 0.908086f
C11860 C10_N_btm.n209 VSS 0.911266f
C11861 C10_N_btm.n210 VSS 0.908086f
C11862 C10_N_btm.n211 VSS 0.908086f
C11863 C10_N_btm.n212 VSS 0.908086f
C11864 C10_N_btm.n213 VSS 0.908086f
C11865 C10_N_btm.n214 VSS 0.911266f
C11866 C10_N_btm.n215 VSS 0.908086f
C11867 C10_N_btm.n216 VSS 1.09754f
C11868 C10_N_btm.n217 VSS 1.42736f
C11869 C10_N_btm.n218 VSS 0.911435f
C11870 C10_N_btm.n219 VSS 0.670503f
C11871 C10_N_btm.n220 VSS 0.911266f
C11872 C10_N_btm.n221 VSS 0.911435f
C11873 C10_N_btm.n222 VSS 0.911266f
C11874 C10_N_btm.n223 VSS 0.911266f
C11875 C10_N_btm.n224 VSS 0.911266f
C11876 C10_N_btm.n225 VSS 0.911266f
C11877 C10_N_btm.n226 VSS 0.911266f
C11878 C10_N_btm.n227 VSS 0.911266f
C11879 C10_N_btm.n228 VSS 0.911266f
C11880 C10_N_btm.n229 VSS 0.911266f
C11881 C10_N_btm.n230 VSS 0.911266f
C11882 C10_N_btm.n231 VSS 0.911266f
C11883 C10_N_btm.n232 VSS 0.911266f
C11884 C10_N_btm.n233 VSS 0.911266f
C11885 C10_N_btm.n234 VSS 0.911266f
C11886 C10_N_btm.n235 VSS 0.911435f
C11887 C10_N_btm.n236 VSS 0.670503f
C11888 C10_N_btm.n237 VSS 0.911435f
C11889 C10_N_btm.n238 VSS 0.670503f
C11890 C10_N_btm.n239 VSS 0.911266f
C11891 C10_N_btm.n240 VSS 0.911435f
C11892 C10_N_btm.n241 VSS 0.911266f
C11893 C10_N_btm.n242 VSS 0.911266f
C11894 C10_N_btm.n243 VSS 0.911266f
C11895 C10_N_btm.n244 VSS 0.911266f
C11896 C10_N_btm.n245 VSS 0.911266f
C11897 C10_N_btm.n246 VSS 1.1455f
C11898 C10_N_btm.n247 VSS 0.911266f
C11899 C10_N_btm.n248 VSS 0.911266f
C11900 C10_N_btm.n249 VSS 0.911266f
C11901 C10_N_btm.n250 VSS 0.911266f
C11902 C10_N_btm.n251 VSS 0.911266f
C11903 C10_N_btm.n252 VSS 0.911266f
C11904 C10_N_btm.n253 VSS 0.911266f
C11905 C10_N_btm.n254 VSS 0.911435f
C11906 C10_N_btm.n255 VSS 0.670503f
C11907 C10_N_btm.n256 VSS 0.911435f
C11908 C10_N_btm.n257 VSS 0.670503f
C11909 C10_N_btm.n258 VSS 0.911435f
C11910 C10_N_btm.n259 VSS 0.911266f
C11911 C10_N_btm.n260 VSS 0.911266f
C11912 C10_N_btm.n261 VSS 0.911266f
C11913 C10_N_btm.n262 VSS 0.911266f
C11914 C10_N_btm.n263 VSS 0.911266f
C11915 C10_N_btm.n264 VSS 0.911266f
C11916 C10_N_btm.n265 VSS 0.911266f
C11917 C10_N_btm.n266 VSS 0.911266f
C11918 C10_N_btm.n267 VSS 0.911266f
C11919 C10_N_btm.n268 VSS 0.911266f
C11920 C10_N_btm.n269 VSS 1.1455f
C11921 C10_N_btm.n270 VSS 1.1455f
C11922 C10_N_btm.n271 VSS 0.911266f
C11923 C10_N_btm.n272 VSS 0.879621f
C11924 C10_N_btm.n273 VSS 0.911266f
C11925 C10_N_btm.n274 VSS 0.911266f
C11926 C10_N_btm.n275 VSS 0.911266f
C11927 C10_N_btm.n276 VSS 0.911266f
C11928 C10_N_btm.n277 VSS 0.911266f
C11929 C10_N_btm.n278 VSS 0.911266f
C11930 C10_N_btm.n279 VSS 0.911266f
C11931 C10_N_btm.n280 VSS 0.911266f
C11932 C10_N_btm.n281 VSS 0.911266f
C11933 C10_N_btm.n282 VSS 0.911435f
C11934 C10_N_btm.n283 VSS 0.670503f
C11935 C10_N_btm.n284 VSS 0.911435f
C11936 C10_N_btm.n285 VSS 0.911266f
C11937 C10_N_btm.n286 VSS 0.911266f
C11938 C10_N_btm.n287 VSS 0.911266f
C11939 C10_N_btm.n288 VSS 0.911266f
C11940 C10_N_btm.n289 VSS 1.24381f
C11941 C10_N_btm.n290 VSS 0.911266f
C11942 C10_N_btm.n291 VSS 0.911266f
C11943 C10_N_btm.n292 VSS 0.911266f
C11944 C10_N_btm.n293 VSS 0.911266f
C11945 C10_N_btm.n294 VSS 0.911266f
C11946 C10_N_btm.n295 VSS 0.911266f
C11947 C10_N_btm.n296 VSS 0.911266f
C11948 C10_N_btm.n297 VSS 0.911266f
C11949 C10_N_btm.n298 VSS 0.911266f
C11950 C10_N_btm.n299 VSS 0.911266f
C11951 C10_N_btm.n300 VSS 0.911266f
C11952 C10_N_btm.n301 VSS 0.911266f
C11953 C10_N_btm.n302 VSS 0.911266f
C11954 C10_N_btm.n303 VSS 0.911266f
C11955 C10_N_btm.n304 VSS 0.911266f
C11956 C10_N_btm.n305 VSS 2.22115f
C11957 C10_N_btm.n306 VSS 0.911266f
C11958 C10_N_btm.n307 VSS 0.911266f
C11959 C10_N_btm.n308 VSS 0.911266f
C11960 C10_N_btm.n309 VSS 0.911266f
C11961 C10_N_btm.n310 VSS 0.911266f
C11962 C10_N_btm.n311 VSS 0.911266f
C11963 C10_N_btm.n312 VSS 0.911266f
C11964 C10_N_btm.n313 VSS 0.911435f
C11965 C10_N_btm.n314 VSS 0.911266f
C11966 C10_N_btm.n315 VSS 0.911435f
C11967 C10_N_btm.n316 VSS 0.670503f
C11968 C10_N_btm.n317 VSS 0.911435f
C11969 C10_N_btm.n318 VSS 0.911266f
C11970 C10_N_btm.n319 VSS 0.911266f
C11971 C10_N_btm.n320 VSS 0.911266f
C11972 C10_N_btm.n321 VSS 0.911266f
C11973 C10_N_btm.n322 VSS 0.911266f
C11974 C10_N_btm.n323 VSS 0.911266f
C11975 C10_N_btm.n324 VSS 0.911266f
C11976 C10_N_btm.n325 VSS 0.911266f
C11977 C10_N_btm.n326 VSS 1.1455f
C11978 C10_N_btm.n327 VSS 0.911266f
C11979 C10_N_btm.n328 VSS 0.911266f
C11980 C10_N_btm.n329 VSS 0.911266f
C11981 C10_N_btm.n330 VSS 0.911266f
C11982 C10_N_btm.n331 VSS 0.911266f
C11983 C10_N_btm.n332 VSS 0.911266f
C11984 C10_N_btm.n333 VSS 1.1455f
C11985 C10_N_btm.n334 VSS 1.1455f
C11986 C10_N_btm.n335 VSS 1.1455f
C11987 C10_N_btm.n336 VSS 0.911266f
C11988 C10_N_btm.n337 VSS 0.911266f
C11989 C10_N_btm.n338 VSS 1.1455f
C11990 C10_N_btm.n339 VSS 0.911266f
C11991 C10_N_btm.n340 VSS 0.911266f
C11992 C10_N_btm.n341 VSS 0.911266f
C11993 C10_N_btm.n342 VSS 0.911266f
C11994 C10_N_btm.n343 VSS 0.911266f
C11995 C10_N_btm.n344 VSS 0.911266f
C11996 C10_N_btm.n345 VSS 0.911266f
C11997 C10_N_btm.n346 VSS 0.911266f
C11998 C10_N_btm.n347 VSS 0.911435f
C11999 C10_N_btm.n348 VSS 0.911266f
C12000 C10_N_btm.n349 VSS 0.911435f
C12001 C10_N_btm.n350 VSS 0.670503f
C12002 C10_N_btm.n351 VSS 0.911435f
C12003 C10_N_btm.n352 VSS 0.911266f
C12004 C10_N_btm.n353 VSS 0.911266f
C12005 C10_N_btm.n354 VSS 0.911266f
C12006 C10_N_btm.n355 VSS 0.911266f
C12007 C10_N_btm.n356 VSS 0.911266f
C12008 C10_N_btm.n357 VSS 0.911266f
C12009 C10_N_btm.n358 VSS 0.911266f
C12010 C10_N_btm.n359 VSS 0.911266f
C12011 C10_N_btm.n360 VSS 0.911266f
C12012 C10_N_btm.n361 VSS 0.911266f
C12013 C10_N_btm.n362 VSS 0.911266f
C12014 C10_N_btm.n363 VSS 0.911266f
C12015 C10_N_btm.n364 VSS 0.911266f
C12016 C10_N_btm.n365 VSS 0.911266f
C12017 C10_N_btm.n366 VSS 0.911266f
C12018 C10_N_btm.n367 VSS 1.1455f
C12019 C10_N_btm.n368 VSS 0.911266f
C12020 C10_N_btm.n369 VSS 0.911266f
C12021 C10_N_btm.n370 VSS 0.911266f
C12022 C10_N_btm.n371 VSS 0.911266f
C12023 C10_N_btm.n372 VSS 0.911266f
C12024 C10_N_btm.n373 VSS 0.911266f
C12025 C10_N_btm.n374 VSS 0.907917f
C12026 C10_N_btm.n375 VSS 0.908086f
C12027 C10_N_btm.n376 VSS 0.911266f
C12028 C10_N_btm.n377 VSS 0.911266f
C12029 C10_N_btm.n378 VSS 0.911266f
C12030 C10_N_btm.n379 VSS 0.908086f
C12031 C10_N_btm.n380 VSS 0.911266f
C12032 C10_N_btm.n381 VSS 0.911266f
C12033 C10_N_btm.n382 VSS 0.908086f
C12034 C10_N_btm.n383 VSS 0.911266f
C12035 C10_N_btm.n384 VSS 0.911266f
C12036 C10_N_btm.n385 VSS 0.911266f
C12037 C10_N_btm.n386 VSS 0.911266f
C12038 C10_N_btm.n387 VSS 0.911266f
C12039 C10_N_btm.n388 VSS 0.908086f
C12040 C10_N_btm.n389 VSS 0.908086f
C12041 C10_N_btm.n390 VSS 0.908086f
C12042 C10_N_btm.n391 VSS 0.908086f
C12043 C10_N_btm.n392 VSS 0.911266f
C12044 C10_N_btm.n393 VSS 0.911266f
C12045 C10_N_btm.n394 VSS 0.911266f
C12046 C10_N_btm.n395 VSS 0.911266f
C12047 C10_N_btm.n396 VSS 0.911266f
C12048 C10_N_btm.n397 VSS 0.908086f
C12049 C10_N_btm.n398 VSS 0.908086f
C12050 C10_N_btm.n399 VSS 0.908086f
C12051 C10_N_btm.n400 VSS 0.908086f
C12052 C10_N_btm.n401 VSS 0.911266f
C12053 C10_N_btm.n402 VSS 0.911266f
C12054 C10_N_btm.n403 VSS 0.911266f
C12055 C10_N_btm.n404 VSS 0.911266f
C12056 C10_N_btm.n405 VSS 0.911266f
C12057 C10_N_btm.n406 VSS 0.908086f
C12058 C10_N_btm.n407 VSS 0.908086f
C12059 C10_N_btm.n408 VSS 0.908086f
C12060 C10_N_btm.n409 VSS 0.908086f
C12061 C10_N_btm.n410 VSS 0.911266f
C12062 C10_N_btm.n411 VSS 0.911266f
C12063 C10_N_btm.n412 VSS 0.911266f
C12064 C10_N_btm.n413 VSS 0.911266f
C12065 C10_N_btm.n414 VSS 0.911266f
C12066 C10_N_btm.n415 VSS 0.911266f
C12067 C10_N_btm.n416 VSS 2.05041f
C12068 C10_N_btm.n417 VSS 0.911266f
C12069 C10_N_btm.n418 VSS 0.911266f
C12070 C10_N_btm.n419 VSS 0.911266f
C12071 C10_N_btm.n420 VSS 0.911266f
C12072 C10_N_btm.n421 VSS 0.911266f
C12073 C10_N_btm.n422 VSS 0.911266f
C12074 C10_N_btm.n423 VSS 0.911266f
C12075 C10_N_btm.n424 VSS 2.82087f
C12076 C10_N_btm.n425 VSS 3.97677f
C12077 C10_N_btm.n426 VSS 0.911266f
C12078 C10_N_btm.n427 VSS 0.911266f
C12079 C10_N_btm.n428 VSS 0.911266f
C12080 C10_N_btm.n429 VSS 1.16658f
C12081 C10_N_btm.n430 VSS 0.908086f
C12082 C10_N_btm.n431 VSS 0.908086f
C12083 C10_N_btm.n432 VSS 0.911266f
C12084 C10_N_btm.n433 VSS 0.911266f
C12085 C10_N_btm.n434 VSS 0.908086f
C12086 C10_N_btm.n435 VSS 0.911266f
C12087 C10_N_btm.n436 VSS 0.911266f
C12088 C10_N_btm.n437 VSS 0.908086f
C12089 C10_N_btm.n438 VSS 0.911266f
C12090 C10_N_btm.n439 VSS 0.911266f
C12091 C10_N_btm.n440 VSS 0.911266f
C12092 C10_N_btm.n441 VSS 0.911266f
C12093 C10_N_btm.n442 VSS 0.908086f
C12094 C10_N_btm.n443 VSS 0.911266f
C12095 C10_N_btm.n444 VSS 0.911266f
C12096 C10_N_btm.n445 VSS 0.908086f
C12097 C10_N_btm.n446 VSS 0.911266f
C12098 C10_N_btm.n447 VSS 0.911266f
C12099 C10_N_btm.n448 VSS 0.911266f
C12100 C10_N_btm.n449 VSS 0.911266f
C12101 C10_N_btm.n450 VSS 0.908086f
C12102 C10_N_btm.n451 VSS 0.911266f
C12103 C10_N_btm.n452 VSS 0.911266f
C12104 C10_N_btm.n453 VSS 0.908086f
C12105 C10_N_btm.n454 VSS 0.911266f
C12106 C10_N_btm.n455 VSS 0.911266f
C12107 C10_N_btm.n456 VSS 0.911266f
C12108 C10_N_btm.n457 VSS 0.911266f
C12109 C10_N_btm.n458 VSS 0.908086f
C12110 C10_N_btm.n459 VSS 0.911266f
C12111 C10_N_btm.n460 VSS 0.911266f
C12112 C10_N_btm.n461 VSS 0.908086f
C12113 C10_N_btm.n462 VSS 0.911266f
C12114 C10_N_btm.n463 VSS 0.911266f
C12115 C10_N_btm.n464 VSS 0.911435f
C12116 C10_N_btm.n465 VSS 0.670503f
C12117 C10_N_btm.n466 VSS 0.911435f
C12118 C10_N_btm.n467 VSS 0.911266f
C12119 C10_N_btm.n468 VSS 0.911266f
C12120 C10_N_btm.n469 VSS 0.911266f
C12121 C10_N_btm.n470 VSS 0.911266f
C12122 C10_N_btm.n471 VSS 0.911266f
C12123 C10_N_btm.n472 VSS 0.911266f
C12124 C10_N_btm.n473 VSS 0.911266f
C12125 C10_N_btm.n474 VSS 0.911266f
C12126 C10_N_btm.n475 VSS 0.911266f
C12127 C10_N_btm.n476 VSS 0.911266f
C12128 C10_N_btm.n477 VSS 0.911266f
C12129 C10_N_btm.n478 VSS 0.911266f
C12130 C10_N_btm.n479 VSS 0.911266f
C12131 C10_N_btm.n480 VSS 0.911266f
C12132 C10_N_btm.n481 VSS 0.911266f
C12133 C10_N_btm.n482 VSS 0.911266f
C12134 C10_N_btm.n483 VSS 0.911266f
C12135 C10_N_btm.n484 VSS 0.911266f
C12136 C10_N_btm.n485 VSS 0.911266f
C12137 C10_N_btm.n486 VSS 0.911266f
C12138 C10_N_btm.n487 VSS 0.911266f
C12139 C10_N_btm.n488 VSS 0.911266f
C12140 C10_N_btm.n489 VSS 0.911266f
C12141 C10_N_btm.n490 VSS 0.911266f
C12142 C10_N_btm.n491 VSS 0.911266f
C12143 C10_N_btm.n492 VSS 0.911266f
C12144 C10_N_btm.n493 VSS 0.911266f
C12145 C10_N_btm.n494 VSS 0.911266f
C12146 C10_N_btm.n495 VSS 0.911266f
C12147 C10_N_btm.n496 VSS 0.911266f
C12148 C10_N_btm.n497 VSS 0.911266f
C12149 C10_N_btm.n498 VSS 0.911266f
C12150 C10_N_btm.n499 VSS 0.911266f
C12151 C10_N_btm.n500 VSS 0.911266f
C12152 C10_N_btm.n501 VSS 0.911266f
C12153 C10_N_btm.n502 VSS 0.911266f
C12154 C10_N_btm.n503 VSS 0.911266f
C12155 C10_N_btm.n504 VSS 0.911266f
C12156 C10_N_btm.n505 VSS 0.911266f
C12157 C10_N_btm.n506 VSS 0.911266f
C12158 C10_N_btm.n507 VSS 0.911266f
C12159 C10_N_btm.n508 VSS 0.911266f
C12160 C10_N_btm.n509 VSS 0.911266f
C12161 C10_N_btm.n510 VSS 0.911266f
C12162 C10_N_btm.n511 VSS 0.911266f
C12163 C10_N_btm.n512 VSS 0.911266f
C12164 C10_N_btm.n513 VSS 0.911266f
C12165 C10_N_btm.n514 VSS 0.911266f
C12166 C10_N_btm.n515 VSS 0.911435f
C12167 C10_N_btm.n516 VSS 0.670503f
C12168 C10_N_btm.n517 VSS 0.670503f
C12169 C10_N_btm.n518 VSS 0.670503f
C12170 C10_N_btm.n519 VSS 0.911435f
C12171 C10_N_btm.n520 VSS 0.911266f
C12172 C10_N_btm.n521 VSS 0.911266f
C12173 C10_N_btm.n522 VSS 0.911266f
C12174 C10_N_btm.n523 VSS 0.911266f
C12175 C10_N_btm.n524 VSS 0.911266f
C12176 C10_N_btm.n525 VSS 0.911266f
C12177 C10_N_btm.n526 VSS 0.911266f
C12178 C10_N_btm.n527 VSS 0.911266f
C12179 C10_N_btm.n528 VSS 0.911266f
C12180 C10_N_btm.n529 VSS 0.911266f
C12181 C10_N_btm.n530 VSS 0.911266f
C12182 C10_N_btm.n531 VSS 0.911266f
C12183 C10_N_btm.n532 VSS 0.911266f
C12184 C10_N_btm.n533 VSS 0.911266f
C12185 C10_N_btm.n534 VSS 0.911266f
C12186 C10_N_btm.n535 VSS 0.911266f
C12187 C10_N_btm.n536 VSS 0.911266f
C12188 C10_N_btm.n537 VSS 0.911266f
C12189 C10_N_btm.n538 VSS 0.911266f
C12190 C10_N_btm.n539 VSS 0.911266f
C12191 C10_N_btm.n540 VSS 0.911266f
C12192 C10_N_btm.n541 VSS 0.911266f
C12193 C10_N_btm.n542 VSS 0.911266f
C12194 C10_N_btm.n543 VSS 0.911266f
C12195 C10_N_btm.n544 VSS 0.911266f
C12196 C10_N_btm.n545 VSS 0.911266f
C12197 C10_N_btm.n546 VSS 0.911266f
C12198 C10_N_btm.n547 VSS 0.911266f
C12199 C10_N_btm.n548 VSS 0.911266f
C12200 C10_N_btm.n549 VSS 0.911266f
C12201 C10_N_btm.n550 VSS 0.911266f
C12202 C10_N_btm.n551 VSS 0.911266f
C12203 C10_N_btm.n552 VSS 0.911266f
C12204 C10_N_btm.n553 VSS 0.911266f
C12205 C10_N_btm.n554 VSS 0.911266f
C12206 C10_N_btm.n555 VSS 0.911266f
C12207 C10_N_btm.n556 VSS 0.911266f
C12208 C10_N_btm.n557 VSS 0.911266f
C12209 C10_N_btm.n558 VSS 0.911266f
C12210 C10_N_btm.n559 VSS 0.911266f
C12211 C10_N_btm.n560 VSS 0.911266f
C12212 C10_N_btm.n561 VSS 0.911266f
C12213 C10_N_btm.n562 VSS 0.911266f
C12214 C10_N_btm.n563 VSS 0.911266f
C12215 C10_N_btm.n564 VSS 0.911266f
C12216 C10_N_btm.n565 VSS 0.911266f
C12217 C10_N_btm.n566 VSS 0.911266f
C12218 C10_N_btm.n567 VSS 0.911266f
C12219 C10_N_btm.n568 VSS 0.911266f
C12220 C10_N_btm.n569 VSS 0.911266f
C12221 C10_N_btm.n570 VSS 0.911266f
C12222 C10_N_btm.n571 VSS 0.911266f
C12223 C10_N_btm.n572 VSS 0.911266f
C12224 C10_N_btm.n573 VSS 0.911266f
C12225 C10_N_btm.n574 VSS 0.911266f
C12226 C10_N_btm.n575 VSS 0.911266f
C12227 C10_N_btm.n576 VSS 0.911266f
C12228 C10_N_btm.n577 VSS 0.911266f
C12229 C10_N_btm.n578 VSS 0.911266f
C12230 C10_N_btm.n579 VSS 0.911266f
C12231 C10_N_btm.n580 VSS 0.911266f
C12232 C10_N_btm.n581 VSS 0.911266f
C12233 C10_N_btm.n582 VSS 0.911266f
C12234 C10_N_btm.n583 VSS 0.911266f
C12235 C10_N_btm.n584 VSS 0.911266f
C12236 C10_N_btm.n585 VSS 0.911266f
C12237 C10_N_btm.n586 VSS 0.911266f
C12238 C10_N_btm.n587 VSS 0.911266f
C12239 C10_N_btm.n588 VSS 0.911266f
C12240 C10_N_btm.n589 VSS 0.911266f
C12241 C10_N_btm.n590 VSS 0.911266f
C12242 C10_N_btm.n591 VSS 0.911266f
C12243 C10_N_btm.n592 VSS 0.911266f
C12244 C10_N_btm.n593 VSS 0.911266f
C12245 C10_N_btm.n594 VSS 0.911435f
C12246 C10_N_btm.n595 VSS 0.911435f
C12247 C10_N_btm.n596 VSS 1.29961f
C12248 C10_N_btm.n597 VSS 1.4275f
C12249 C10_N_btm.n598 VSS 1.09757f
C12250 C10_N_btm.n599 VSS 0.911266f
C12251 C10_N_btm.n600 VSS 0.911266f
C12252 C10_N_btm.n601 VSS 0.911266f
C12253 C10_N_btm.n602 VSS 0.911266f
C12254 C10_N_btm.n603 VSS 0.908086f
C12255 C10_N_btm.n604 VSS 0.908086f
C12256 C10_N_btm.n605 VSS 0.908086f
C12257 C10_N_btm.n606 VSS 0.908086f
C12258 C10_N_btm.n607 VSS 0.911266f
C12259 C10_N_btm.n608 VSS 0.911266f
C12260 C10_N_btm.n609 VSS 0.911266f
C12261 C10_N_btm.n610 VSS 0.911266f
C12262 C10_N_btm.n611 VSS 0.908086f
C12263 C10_N_btm.n612 VSS 0.908086f
C12264 C10_N_btm.n613 VSS 0.908086f
C12265 C10_N_btm.n614 VSS 0.908086f
C12266 C10_N_btm.n615 VSS 0.911266f
C12267 C10_N_btm.n616 VSS 0.911266f
C12268 C10_N_btm.n617 VSS 0.911266f
C12269 C10_N_btm.n618 VSS 0.911266f
C12270 C10_N_btm.n619 VSS 0.908086f
C12271 C10_N_btm.n620 VSS 0.908086f
C12272 C10_N_btm.n621 VSS 0.908086f
C12273 C10_N_btm.n622 VSS 0.908086f
C12274 C10_N_btm.n623 VSS 0.911266f
C12275 C10_N_btm.n624 VSS 0.911266f
C12276 C10_N_btm.n625 VSS 0.911266f
C12277 C10_N_btm.n626 VSS 0.911266f
C12278 C10_N_btm.n627 VSS 0.908086f
C12279 C10_N_btm.n628 VSS 0.908086f
C12280 C10_N_btm.n629 VSS 0.908086f
C12281 C10_N_btm.n630 VSS 0.908086f
C12282 C10_N_btm.n631 VSS 0.911266f
C12283 C10_N_btm.n632 VSS 0.911266f
C12284 C10_N_btm.n633 VSS 0.911266f
C12285 C10_N_btm.n634 VSS 0.911266f
C12286 C10_N_btm.n635 VSS 0.911266f
C12287 C10_N_btm.n636 VSS 0.911266f
C12288 C10_N_btm.n637 VSS 0.911266f
C12289 C10_N_btm.n638 VSS 0.911266f
C12290 C10_N_btm.n639 VSS 2.05041f
C12291 C10_N_btm.n640 VSS 2.05041f
C12292 C10_N_btm.n641 VSS 2.05041f
C12293 C10_N_btm.n642 VSS 2.05041f
C12294 C10_N_btm.n643 VSS 3.97683f
C12295 C10_N_btm.n644 VSS 1.16658f
C12296 C10_N_btm.n645 VSS 2.82097f
C12297 C10_N_btm.n646 VSS 0.911266f
C12298 C10_N_btm.n647 VSS 0.911266f
C12299 C10_N_btm.n648 VSS 0.911266f
C12300 C10_N_btm.n649 VSS 0.911266f
C12301 C10_N_btm.n650 VSS 0.911266f
C12302 C10_N_btm.n651 VSS 0.911266f
C12303 C10_N_btm.n652 VSS 0.911266f
C12304 C10_N_btm.n653 VSS 0.911266f
C12305 C10_N_btm.n654 VSS 0.911266f
C12306 C10_N_btm.n655 VSS 0.911266f
C12307 C10_N_btm.n656 VSS 0.911266f
C12308 C10_N_btm.n657 VSS 0.911266f
C12309 C10_N_btm.n658 VSS 0.911266f
C12310 C10_N_btm.n659 VSS 0.911266f
C12311 C10_N_btm.n660 VSS 0.911266f
C12312 C10_N_btm.n661 VSS 0.911266f
C12313 C10_N_btm.n662 VSS 0.911266f
C12314 C10_N_btm.n663 VSS 0.911266f
C12315 C10_N_btm.n664 VSS 0.911266f
C12316 C10_N_btm.n665 VSS 0.911266f
C12317 C10_N_btm.n666 VSS 0.911266f
C12318 C10_N_btm.n667 VSS 0.911266f
C12319 C10_N_btm.n668 VSS 0.911266f
C12320 C10_N_btm.n669 VSS 0.911266f
C12321 C10_N_btm.n670 VSS 0.911266f
C12322 C10_N_btm.n671 VSS 0.908086f
C12323 C10_N_btm.n672 VSS 0.908086f
C12324 C10_N_btm.n673 VSS 0.908086f
C12325 C10_N_btm.n674 VSS 0.908086f
C12326 C10_N_btm.n675 VSS 0.908086f
C12327 C10_N_btm.n676 VSS 0.911266f
C12328 C10_N_btm.n677 VSS 0.911266f
C12329 C10_N_btm.n678 VSS 0.911266f
C12330 C10_N_btm.n679 VSS 0.911266f
C12331 C10_N_btm.n680 VSS 0.911266f
C12332 C10_N_btm.n681 VSS 0.911266f
C12333 C10_N_btm.n682 VSS 0.911266f
C12334 C10_N_btm.n683 VSS 0.911266f
C12335 C10_N_btm.n684 VSS 0.911266f
C12336 C10_N_btm.n685 VSS 0.911266f
C12337 C10_N_btm.n686 VSS 0.911266f
C12338 C10_N_btm.n687 VSS 0.911266f
C12339 C10_N_btm.n688 VSS 0.911435f
C12340 C10_N_btm.n689 VSS 0.670503f
C12341 C10_N_btm.n690 VSS 0.670503f
C12342 C10_N_btm.n691 VSS 0.670503f
C12343 C10_N_btm.n692 VSS 0.911435f
C12344 C10_N_btm.n693 VSS 0.911266f
C12345 C10_N_btm.n694 VSS 0.911435f
C12346 C10_N_btm.n695 VSS 0.670503f
C12347 C10_N_btm.n696 VSS 0.670503f
C12348 C10_N_btm.n697 VSS 0.670503f
C12349 C10_N_btm.n698 VSS 0.911435f
C12350 C10_N_btm.n699 VSS 0.911266f
C12351 C10_N_btm.n700 VSS 0.911266f
C12352 C10_N_btm.n701 VSS 0.911266f
C12353 C10_N_btm.n702 VSS 0.911266f
C12354 C10_N_btm.n703 VSS 0.911266f
C12355 C10_N_btm.n704 VSS 0.911266f
C12356 C10_N_btm.n705 VSS 0.911266f
C12357 C10_N_btm.n706 VSS 0.911266f
C12358 C10_N_btm.n707 VSS 0.911266f
C12359 C10_N_btm.n708 VSS 0.911435f
C12360 C10_N_btm.n709 VSS 0.911435f
C12361 C10_N_btm.n710 VSS 0.670503f
C12362 C10_N_btm.n711 VSS 0.670503f
C12363 C10_N_btm.n712 VSS 0.670503f
C12364 C10_N_btm.n713 VSS 0.911435f
C12365 C10_N_btm.n714 VSS 0.911266f
C12366 C10_N_btm.n715 VSS 0.911266f
C12367 C10_N_btm.n716 VSS 0.911266f
C12368 C10_N_btm.n717 VSS 0.911266f
C12369 C10_N_btm.n718 VSS 0.911266f
C12370 C10_N_btm.n719 VSS 0.911266f
C12371 C10_N_btm.n720 VSS 0.911266f
C12372 C10_N_btm.n721 VSS 0.911266f
C12373 C10_N_btm.n722 VSS 1.1455f
C12374 C10_N_btm.n723 VSS 1.1455f
C12375 C10_N_btm.n724 VSS 1.1455f
C12376 C10_N_btm.n725 VSS 1.1455f
C12377 C10_N_btm.n726 VSS 0.911266f
C12378 C10_N_btm.n727 VSS 0.911266f
C12379 C10_N_btm.n728 VSS 0.911266f
C12380 C10_N_btm.n729 VSS 0.911266f
C12381 C10_N_btm.n730 VSS 0.911266f
C12382 C10_N_btm.n731 VSS 0.911266f
C12383 C10_N_btm.n732 VSS 0.911266f
C12384 C10_N_btm.n733 VSS 0.911435f
C12385 C10_N_btm.n734 VSS 0.670503f
C12386 C10_N_btm.n735 VSS 0.670503f
C12387 C10_N_btm.n736 VSS 0.670503f
C12388 C10_N_btm.n737 VSS 0.911435f
C12389 C10_N_btm.n738 VSS 0.911266f
C12390 C10_N_btm.n739 VSS 0.911266f
C12391 C10_N_btm.n740 VSS 0.911266f
C12392 C10_N_btm.n741 VSS 0.911266f
C12393 C10_N_btm.n742 VSS 0.911266f
C12394 C10_N_btm.n743 VSS 0.911435f
C12395 C10_N_btm.n744 VSS 0.670503f
C12396 C10_N_btm.n745 VSS 0.670503f
C12397 C10_N_btm.n746 VSS 0.670503f
C12398 C10_N_btm.n747 VSS 0.911435f
C12399 C10_N_btm.n748 VSS 0.911435f
C12400 C10_N_btm.n749 VSS 0.670503f
C12401 C10_N_btm.n750 VSS 0.911266f
C12402 C10_N_btm.n751 VSS 0.911435f
C12403 C10_N_btm.n752 VSS 0.911266f
C12404 C10_N_btm.n753 VSS 0.911266f
C12405 C10_N_btm.n754 VSS 0.911266f
C12406 C10_N_btm.n755 VSS 0.911266f
C12407 C10_N_btm.n756 VSS 0.911266f
C12408 C10_N_btm.n757 VSS 0.911266f
C12409 C10_N_btm.n758 VSS 0.911266f
C12410 C10_N_btm.n759 VSS 0.911266f
C12411 C10_N_btm.n760 VSS 0.911266f
C12412 C10_N_btm.n761 VSS 0.911266f
C12413 C10_N_btm.n762 VSS 0.911266f
C12414 C10_N_btm.n763 VSS 0.911266f
C12415 C10_N_btm.n764 VSS 0.911266f
C12416 C10_N_btm.n765 VSS 0.911266f
C12417 C10_N_btm.n766 VSS 0.911266f
C12418 C10_N_btm.n767 VSS 0.911435f
C12419 C10_N_btm.n768 VSS 0.670503f
C12420 C10_N_btm.n769 VSS 0.670503f
C12421 C10_N_btm.n770 VSS 0.670503f
C12422 C10_N_btm.n771 VSS 0.911435f
C12423 C10_N_btm.n772 VSS 0.911435f
C12424 C10_N_btm.n773 VSS 0.911266f
C12425 C10_N_btm.n774 VSS 0.911266f
C12426 C10_N_btm.n775 VSS 0.911266f
C12427 C10_N_btm.n776 VSS 0.911266f
C12428 C10_N_btm.n777 VSS 0.911266f
C12429 C10_N_btm.n778 VSS 0.911266f
C12430 C10_N_btm.n779 VSS 0.911266f
C12431 C10_N_btm.n780 VSS 0.911435f
C12432 C10_N_btm.n781 VSS 0.670503f
C12433 C10_N_btm.n782 VSS 0.670503f
C12434 C10_N_btm.n783 VSS 0.670503f
C12435 C10_N_btm.n784 VSS 0.670503f
C12436 C10_N_btm.n785 VSS 0.911435f
C12437 C10_N_btm.n786 VSS 0.911435f
C12438 C10_N_btm.n787 VSS 0.911266f
C12439 C10_N_btm.n788 VSS 0.911266f
C12440 C10_N_btm.n789 VSS 0.911266f
C12441 C10_N_btm.n790 VSS 0.911266f
C12442 C10_N_btm.n791 VSS 0.911266f
C12443 C10_N_btm.n792 VSS 0.911266f
C12444 C10_N_btm.n793 VSS 0.911266f
C12445 C10_N_btm.n794 VSS 0.911266f
C12446 C10_N_btm.n795 VSS 0.911435f
C12447 C10_N_btm.n796 VSS 0.911435f
C12448 C10_N_btm.n797 VSS 0.670503f
C12449 C10_N_btm.n798 VSS 0.670503f
C12450 C10_N_btm.n799 VSS 0.670503f
C12451 C10_N_btm.n800 VSS 0.670503f
C12452 C10_N_btm.n801 VSS 0.911435f
C12453 C10_N_btm.n802 VSS 0.911435f
C12454 C10_N_btm.n803 VSS 0.911266f
C12455 C10_N_btm.n804 VSS 0.911266f
C12456 C10_N_btm.n805 VSS 0.911266f
C12457 C10_N_btm.n806 VSS 0.911266f
C12458 C10_N_btm.n807 VSS 0.911266f
C12459 C10_N_btm.n808 VSS 0.911266f
C12460 C10_N_btm.n809 VSS 0.911266f
C12461 C10_N_btm.n810 VSS 0.911266f
C12462 C10_N_btm.n811 VSS 0.911435f
C12463 C10_N_btm.n812 VSS 0.911435f
C12464 C10_N_btm.n813 VSS 0.670503f
C12465 C10_N_btm.n814 VSS 0.670503f
C12466 C10_N_btm.n815 VSS 0.670503f
C12467 C10_N_btm.n816 VSS 0.911435f
C12468 C10_N_btm.n817 VSS 0.911266f
C12469 C10_N_btm.n818 VSS 0.911266f
C12470 C10_N_btm.n819 VSS 0.911266f
C12471 C10_N_btm.n820 VSS 0.911266f
C12472 C10_N_btm.n821 VSS 0.911266f
C12473 C10_N_btm.n822 VSS 0.911266f
C12474 C10_N_btm.n823 VSS 0.911266f
C12475 C10_N_btm.n824 VSS 0.879621f
C12476 C10_N_btm.n825 VSS 1.24381f
C12477 C10_N_btm.n826 VSS 1.1455f
C12478 C10_N_btm.n827 VSS 1.1455f
C12479 C10_N_btm.n828 VSS 1.1455f
C12480 C10_N_btm.n829 VSS 1.1455f
C12481 C10_N_btm.n830 VSS 1.1455f
C12482 C10_N_btm.n831 VSS 1.1455f
C12483 C10_N_btm.n832 VSS 1.1455f
C12484 C10_N_btm.n833 VSS 1.1455f
C12485 C10_N_btm.n834 VSS 1.1455f
C12486 C10_N_btm.n835 VSS 1.1455f
C12487 C10_N_btm.n836 VSS 1.1455f
C12488 C10_N_btm.n837 VSS 1.1455f
C12489 C10_N_btm.n838 VSS 1.1455f
C12490 C10_N_btm.n839 VSS 1.1455f
C12491 C10_N_btm.n840 VSS 1.1455f
C12492 C10_N_btm.n841 VSS 1.1455f
C12493 C10_N_btm.n842 VSS 0.911266f
C12494 C10_N_btm.n843 VSS 0.911266f
C12495 C10_N_btm.n844 VSS 0.911266f
C12496 C10_N_btm.n845 VSS 0.911266f
C12497 C10_N_btm.n846 VSS 0.911266f
C12498 C10_N_btm.n847 VSS 0.911435f
C12499 C10_N_btm.n848 VSS 0.670503f
C12500 C10_N_btm.n849 VSS 0.670503f
C12501 C10_N_btm.n850 VSS 0.670503f
C12502 C10_N_btm.n851 VSS 0.911266f
C12503 C10_N_btm.n852 VSS 0.911435f
C12504 C10_N_btm.n853 VSS 0.670503f
C12505 C10_N_btm.n854 VSS 0.670503f
C12506 C10_N_btm.n855 VSS 0.911435f
C12507 C10_N_btm.n856 VSS 0.911435f
C12508 C10_N_btm.n857 VSS 0.911266f
C12509 C10_N_btm.n858 VSS 0.911266f
C12510 C10_N_btm.n859 VSS 0.911266f
C12511 C10_N_btm.n860 VSS 0.911266f
C12512 C10_N_btm.n861 VSS 0.911266f
C12513 C10_N_btm.n862 VSS 0.911266f
C12514 C10_N_btm.n863 VSS 0.911266f
C12515 C10_N_btm.n864 VSS 2.22115f
C12516 C10_N_btm.n865 VSS 1.1455f
C12517 C10_N_btm.n866 VSS 1.1455f
C12518 C10_N_btm.n867 VSS 1.1455f
C12519 C10_N_btm.n868 VSS 0.911266f
C12520 C10_N_btm.n869 VSS 0.911266f
C12521 C10_N_btm.n870 VSS 0.911266f
C12522 C10_N_btm.n871 VSS 0.911266f
C12523 C10_N_btm.n872 VSS 0.911266f
C12524 C10_N_btm.n873 VSS 0.911266f
C12525 C10_N_btm.n874 VSS 0.911435f
C12526 C10_N_btm.n875 VSS 0.670503f
C12527 C10_N_btm.n876 VSS 0.670504f
C12528 C10_N_btm.n877 VSS 0.670503f
C12529 C10_N_btm.n878 VSS 0.670503f
C12530 C10_N_btm.n879 VSS 0.911435f
C12531 C10_N_btm.n880 VSS 0.911266f
C12532 C10_N_btm.n881 VSS 0.911266f
C12533 C10_N_btm.n882 VSS 0.911266f
C12534 C10_N_btm.n883 VSS 0.911266f
C12535 C10_N_btm.n884 VSS 0.911266f
C12536 C10_N_btm.n885 VSS 0.911266f
C12537 C10_N_btm.n886 VSS 0.911266f
C12538 C10_N_btm.n887 VSS 1.1455f
C12539 C10_N_btm.n888 VSS 1.1455f
C12540 C10_N_btm.n889 VSS 1.1455f
C12541 C10_N_btm.n890 VSS 0.911266f
C12542 C10_N_btm.n891 VSS 0.911266f
C12543 C10_N_btm.n892 VSS 0.911266f
C12544 C10_N_btm.n893 VSS 0.911266f
C12545 C10_N_btm.n894 VSS 0.911266f
C12546 C10_N_btm.n895 VSS 0.911266f
C12547 C10_N_btm.n896 VSS 0.911266f
C12548 C10_N_btm.n897 VSS 0.911435f
C12549 C10_N_btm.n898 VSS 0.911435f
C12550 C10_N_btm.n899 VSS 0.670503f
C12551 C10_N_btm.n900 VSS 0.670503f
C12552 C10_N_btm.n901 VSS 0.670503f
C12553 C10_N_btm.n902 VSS 0.670503f
C12554 C10_N_btm.n903 VSS 0.911435f
C12555 C10_N_btm.n904 VSS 0.911266f
C12556 C10_N_btm.n905 VSS 0.911266f
C12557 C10_N_btm.n906 VSS 0.911266f
C12558 C10_N_btm.n907 VSS 0.911266f
C12559 C10_N_btm.n908 VSS 0.911266f
C12560 C10_N_btm.n909 VSS 0.911266f
C12561 C10_N_btm.n910 VSS 0.911266f
C12562 C10_N_btm.n911 VSS 0.911266f
C12563 C10_N_btm.n912 VSS 0.911266f
C12564 C10_N_btm.n913 VSS 0.911266f
C12565 C10_N_btm.n914 VSS 0.911266f
C12566 C10_N_btm.n915 VSS 0.911266f
C12567 C10_N_btm.n916 VSS 0.911266f
C12568 C10_N_btm.n917 VSS 0.911266f
C12569 C10_N_btm.n918 VSS 0.911435f
C12570 C10_N_btm.n919 VSS 0.911435f
C12571 C10_N_btm.n920 VSS 0.670503f
C12572 C10_N_btm.n921 VSS 0.670503f
C12573 C10_N_btm.n922 VSS 0.670503f
C12574 C10_N_btm.n923 VSS 1.29961f
C12575 C10_N_btm.n924 VSS 0.911435f
C12576 C10_N_btm.n925 VSS 0.911266f
C12577 C10_N_btm.n926 VSS 0.911266f
C12578 C10_N_btm.n927 VSS 0.911266f
C12579 C10_N_btm.n928 VSS 0.911266f
C12580 C10_N_btm.n929 VSS 0.911266f
C12581 C10_N_btm.n930 VSS 0.911266f
C12582 C10_N_btm.n931 VSS 0.911266f
C12583 C10_N_btm.n932 VSS 0.911266f
C12584 C10_N_btm.n933 VSS 0.911266f
C12585 C10_N_btm.n934 VSS 0.911266f
C12586 C10_N_btm.n935 VSS 0.911266f
C12587 C10_N_btm.n936 VSS 0.911266f
C12588 C10_N_btm.n937 VSS 0.911266f
C12589 C10_N_btm.n938 VSS 0.911266f
C12590 C10_N_btm.n939 VSS 0.911266f
C12591 C10_N_btm.n940 VSS 0.911266f
C12592 C10_N_btm.n941 VSS 0.911266f
C12593 C10_N_btm.n942 VSS 0.911266f
C12594 C10_N_btm.n943 VSS 0.911266f
C12595 C10_N_btm.n944 VSS 0.911266f
C12596 C10_N_btm.n945 VSS 0.911266f
C12597 C10_N_btm.n946 VSS 0.911266f
C12598 C10_N_btm.n947 VSS 0.911266f
C12599 C10_N_btm.n948 VSS 0.911266f
C12600 C10_N_btm.n949 VSS 0.911266f
C12601 C10_N_btm.n950 VSS 0.911266f
C12602 C10_N_btm.n951 VSS 0.911266f
C12603 C10_N_btm.n952 VSS 0.911266f
C12604 C10_N_btm.n953 VSS 0.911266f
C12605 C10_N_btm.n954 VSS 0.911266f
C12606 C10_N_btm.n955 VSS 0.911266f
C12607 C10_N_btm.n956 VSS 0.911266f
C12608 C10_N_btm.n957 VSS 0.911266f
C12609 C10_N_btm.n958 VSS 0.911266f
C12610 C10_N_btm.n959 VSS 0.911266f
C12611 C10_N_btm.n960 VSS 0.911266f
C12612 C10_N_btm.n961 VSS 0.911266f
C12613 C10_N_btm.n962 VSS 0.911266f
C12614 C10_N_btm.n963 VSS 0.911266f
C12615 C10_N_btm.n964 VSS 0.911266f
C12616 C10_N_btm.n965 VSS 0.911266f
C12617 C10_N_btm.n966 VSS 0.911266f
C12618 C10_N_btm.n967 VSS 0.911266f
C12619 C10_N_btm.n968 VSS 0.911266f
C12620 C10_N_btm.n969 VSS 2.05041f
C12621 C10_N_btm.n970 VSS 2.05041f
C12622 C10_N_btm.n971 VSS 2.05041f
C12623 C10_N_btm.n972 VSS 2.05041f
C12624 C10_N_btm.n973 VSS 0.911266f
C12625 C10_N_btm.n974 VSS 0.911266f
C12626 C10_N_btm.n975 VSS 0.911266f
C12627 C10_N_btm.n976 VSS 0.911266f
C12628 C10_N_btm.n977 VSS 0.911266f
C12629 C10_N_btm.n978 VSS 0.911266f
C12630 C10_N_btm.n979 VSS 0.911266f
C12631 C10_N_btm.n980 VSS 0.911266f
C12632 C10_N_btm.n981 VSS 0.911266f
C12633 C10_N_btm.n982 VSS 0.911266f
C12634 C10_N_btm.n983 VSS 0.911266f
C12635 C10_N_btm.n984 VSS 0.911266f
C12636 C10_N_btm.n985 VSS 0.911266f
C12637 C10_N_btm.n986 VSS 0.911266f
C12638 C10_N_btm.n987 VSS 0.911266f
C12639 C10_N_btm.n988 VSS 0.911266f
C12640 C10_N_btm.n989 VSS 0.911266f
C12641 C10_N_btm.n990 VSS 0.911266f
C12642 C10_N_btm.n991 VSS 0.911266f
C12643 C10_N_btm.n992 VSS 0.911266f
C12644 C10_N_btm.n993 VSS 0.911266f
C12645 C10_N_btm.n994 VSS 0.911266f
C12646 C10_N_btm.n995 VSS 0.911266f
C12647 C10_N_btm.n996 VSS 0.911266f
C12648 C10_N_btm.n997 VSS 0.911266f
C12649 C10_N_btm.n998 VSS 0.911266f
C12650 C10_N_btm.n999 VSS 0.911266f
C12651 C10_N_btm.n1000 VSS 0.911266f
C12652 C10_N_btm.n1001 VSS 0.911266f
C12653 C10_N_btm.n1002 VSS 0.911266f
C12654 C10_N_btm.n1003 VSS 0.911266f
C12655 C10_N_btm.n1004 VSS 0.911266f
C12656 C10_N_btm.n1005 VSS 0.911266f
C12657 C10_N_btm.n1006 VSS 0.911266f
C12658 C10_N_btm.n1007 VSS 0.911266f
C12659 C10_N_btm.n1008 VSS 0.911266f
C12660 C10_N_btm.n1009 VSS 0.911266f
C12661 C10_N_btm.n1010 VSS 0.911266f
C12662 C10_N_btm.n1011 VSS 0.911266f
C12663 C10_N_btm.n1012 VSS 0.911266f
C12664 C10_N_btm.n1013 VSS 0.908086f
C12665 C10_N_btm.n1014 VSS 0.908086f
C12666 C10_N_btm.n1015 VSS 0.911266f
C12667 C10_N_btm.n1016 VSS 0.911266f
C12668 C10_N_btm.n1017 VSS 0.911266f
C12669 C10_N_btm.n1018 VSS 0.911266f
C12670 C10_N_btm.n1019 VSS 0.908086f
C12671 C10_N_btm.n1020 VSS 0.908086f
C12672 C10_N_btm.n1021 VSS 0.908086f
C12673 C10_N_btm.n1022 VSS 0.908086f
C12674 C10_N_btm.n1023 VSS 0.911266f
C12675 C10_N_btm.n1024 VSS 0.911266f
C12676 C10_N_btm.n1025 VSS 0.911266f
C12677 C10_N_btm.n1026 VSS 0.911266f
C12678 C10_N_btm.n1027 VSS 0.908086f
C12679 C10_N_btm.n1028 VSS 0.908086f
C12680 C10_N_btm.n1029 VSS 0.908086f
C12681 C10_N_btm.n1030 VSS 0.908086f
C12682 C10_N_btm.n1031 VSS 0.911266f
C12683 C10_N_btm.n1032 VSS 0.911266f
C12684 C10_N_btm.n1033 VSS 0.911266f
C12685 C10_N_btm.n1034 VSS 0.911266f
C12686 C10_N_btm.n1035 VSS 0.908086f
C12687 C10_N_btm.n1036 VSS 0.908086f
C12688 C10_N_btm.n1037 VSS 0.908086f
C12689 C10_N_btm.n1038 VSS 0.908086f
C12690 C10_N_btm.n1039 VSS 0.911266f
C12691 C10_N_btm.n1040 VSS 0.911266f
C12692 C10_N_btm.n1041 VSS 0.911266f
C12693 C10_N_btm.n1042 VSS 0.911266f
C12694 C10_N_btm.n1043 VSS 0.908086f
C12695 C10_N_btm.n1044 VSS 2.01002f
C12696 a_4190_30871.t0 VSS 0.030815f
C12697 a_4190_30871.t3 VSS 0.02003f
C12698 a_4190_30871.t2 VSS 0.02003f
C12699 a_4190_30871.n0 VSS 0.074179f
C12700 a_4190_30871.n1 VSS 0.15561f
C12701 a_4190_30871.t18 VSS 0.405728f
C12702 a_4190_30871.t16 VSS 0.417826f
C12703 a_4190_30871.t4 VSS 0.406413f
C12704 a_4190_30871.t7 VSS 0.405728f
C12705 a_4190_30871.t15 VSS 0.406413f
C12706 a_4190_30871.t11 VSS 0.405728f
C12707 a_4190_30871.t5 VSS 0.406413f
C12708 a_4190_30871.n2 VSS 0.1865f
C12709 a_4190_30871.t14 VSS 0.405728f
C12710 a_4190_30871.n3 VSS 0.200549f
C12711 a_4190_30871.n4 VSS 0.267802f
C12712 a_4190_30871.n5 VSS 0.20863f
C12713 a_4190_30871.n6 VSS 0.1865f
C12714 a_4190_30871.n7 VSS 0.20863f
C12715 a_4190_30871.n8 VSS 0.1865f
C12716 a_4190_30871.n9 VSS 0.368532f
C12717 a_4190_30871.n10 VSS 1.26949f
C12718 a_4190_30871.n11 VSS 0.15561f
C12719 a_4190_30871.t10 VSS 0.405728f
C12720 a_4190_30871.t20 VSS 0.406413f
C12721 a_4190_30871.t12 VSS 0.405728f
C12722 a_4190_30871.t19 VSS 0.406413f
C12723 a_4190_30871.t13 VSS 0.405728f
C12724 a_4190_30871.t8 VSS 0.406413f
C12725 a_4190_30871.n12 VSS 0.1865f
C12726 a_4190_30871.t6 VSS 0.405728f
C12727 a_4190_30871.n13 VSS 0.200549f
C12728 a_4190_30871.n14 VSS 0.267802f
C12729 a_4190_30871.n15 VSS 0.20863f
C12730 a_4190_30871.n16 VSS 0.1865f
C12731 a_4190_30871.n17 VSS 0.20863f
C12732 a_4190_30871.n18 VSS 0.1865f
C12733 a_4190_30871.t21 VSS 0.417826f
C12734 a_4190_30871.n19 VSS 0.368532f
C12735 a_4190_30871.n20 VSS 1.40705f
C12736 a_4190_30871.n21 VSS 5.61859f
C12737 a_4190_30871.t17 VSS 0.047935f
C12738 a_4190_30871.t9 VSS 0.029895f
C12739 a_4190_30871.n22 VSS 0.22738f
C12740 a_4190_30871.n23 VSS 4.7428f
C12741 a_4190_30871.n24 VSS 0.360882f
C12742 a_4190_30871.n25 VSS 0.061654f
C12743 a_4190_30871.t1 VSS 0.030815f
C12744 a_6151_47436.t1 VSS 0.054923f
C12745 a_6151_47436.t4 VSS 0.018223f
C12746 a_6151_47436.t3 VSS 0.028557f
C12747 a_6151_47436.n0 VSS 0.071023f
C12748 a_6151_47436.t6 VSS 0.018579f
C12749 a_6151_47436.t8 VSS 0.034014f
C12750 a_6151_47436.n1 VSS 0.074158f
C12751 a_6151_47436.t9 VSS 0.032583f
C12752 a_6151_47436.t5 VSS 0.013907f
C12753 a_6151_47436.n2 VSS 0.057844f
C12754 a_6151_47436.t7 VSS 0.028361f
C12755 a_6151_47436.t10 VSS 0.017862f
C12756 a_6151_47436.n3 VSS 0.061452f
C12757 a_6151_47436.n4 VSS 0.527464f
C12758 a_6151_47436.n5 VSS 0.77723f
C12759 a_6151_47436.t12 VSS 0.032583f
C12760 a_6151_47436.t11 VSS 0.013907f
C12761 a_6151_47436.n6 VSS 0.060137f
C12762 a_6151_47436.t2 VSS 0.028361f
C12763 a_6151_47436.t13 VSS 0.017862f
C12764 a_6151_47436.n7 VSS 0.058509f
C12765 a_6151_47436.n8 VSS 0.332287f
C12766 a_6151_47436.n9 VSS 0.877859f
C12767 a_6151_47436.n10 VSS 0.958869f
C12768 a_6151_47436.n11 VSS 0.150234f
C12769 a_6151_47436.t0 VSS 0.053212f
C12770 a_10193_42453.t0 VSS 0.01942f
C12771 a_10193_42453.t16 VSS 0.020072f
C12772 a_10193_42453.t13 VSS 0.032147f
C12773 a_10193_42453.n0 VSS 0.062643f
C12774 a_10193_42453.t11 VSS 0.020551f
C12775 a_10193_42453.t20 VSS 0.032727f
C12776 a_10193_42453.n1 VSS 0.046023f
C12777 a_10193_42453.n2 VSS 0.135819f
C12778 a_10193_42453.t10 VSS 0.020572f
C12779 a_10193_42453.t5 VSS 0.040617f
C12780 a_10193_42453.n3 VSS 0.048039f
C12781 a_10193_42453.t9 VSS 0.020551f
C12782 a_10193_42453.t18 VSS 0.032727f
C12783 a_10193_42453.n4 VSS 0.099524f
C12784 a_10193_42453.n5 VSS 1.03f
C12785 a_10193_42453.t23 VSS 0.032727f
C12786 a_10193_42453.t6 VSS 0.020551f
C12787 a_10193_42453.n6 VSS 0.088861f
C12788 a_10193_42453.t14 VSS 0.032727f
C12789 a_10193_42453.t17 VSS 0.020551f
C12790 a_10193_42453.n7 VSS 0.049351f
C12791 a_10193_42453.n8 VSS 1.08476f
C12792 a_10193_42453.t4 VSS 0.040617f
C12793 a_10193_42453.t15 VSS 0.020572f
C12794 a_10193_42453.n9 VSS 0.042422f
C12795 a_10193_42453.n10 VSS 0.436748f
C12796 a_10193_42453.t12 VSS 0.040617f
C12797 a_10193_42453.t19 VSS 0.020572f
C12798 a_10193_42453.n11 VSS 0.062712f
C12799 a_10193_42453.n12 VSS 0.67121f
C12800 a_10193_42453.t8 VSS 0.040617f
C12801 a_10193_42453.t22 VSS 0.020572f
C12802 a_10193_42453.n13 VSS 0.049081f
C12803 a_10193_42453.n14 VSS 1.06069f
C12804 a_10193_42453.t7 VSS 0.032727f
C12805 a_10193_42453.t21 VSS 0.020551f
C12806 a_10193_42453.n15 VSS 0.050516f
C12807 a_10193_42453.n16 VSS 0.556624f
C12808 a_10193_42453.n17 VSS 0.719928f
C12809 a_10193_42453.n18 VSS 0.747127f
C12810 a_10193_42453.t3 VSS 0.012623f
C12811 a_10193_42453.t2 VSS 0.012623f
C12812 a_10193_42453.n19 VSS 0.025246f
C12813 a_10193_42453.n20 VSS 0.146968f
C12814 a_10193_42453.n21 VSS 0.058272f
C12815 a_10193_42453.t1 VSS 0.01942f
C12816 a_n2312_39304.t0 VSS 0.053828f
C12817 a_n2312_39304.t3 VSS 0.034988f
C12818 a_n2312_39304.t2 VSS 0.034988f
C12819 a_n2312_39304.n0 VSS 0.129578f
C12820 a_n2312_39304.t5 VSS 0.055446f
C12821 a_n2312_39304.t4 VSS 0.088882f
C12822 a_n2312_39304.n1 VSS 2.43072f
C12823 a_n2312_39304.n2 VSS 9.31004f
C12824 a_n2312_39304.n3 VSS 0.1077f
C12825 a_n2312_39304.t1 VSS 0.053828f
C12826 a_19237_31679.t3 VSS 0.038924f
C12827 a_19237_31679.t2 VSS 0.038924f
C12828 a_19237_31679.n0 VSS 0.144154f
C12829 a_19237_31679.t4 VSS 2.9556f
C12830 a_19237_31679.n1 VSS 14.4828f
C12831 a_19237_31679.t0 VSS 0.059883f
C12832 a_19237_31679.n2 VSS 0.119815f
C12833 a_19237_31679.t1 VSS 0.059883f
C12834 a_n3420_39072.t0 VSS 0.045098f
C12835 a_n3420_39072.t5 VSS 0.029314f
C12836 a_n3420_39072.t7 VSS 0.029314f
C12837 a_n3420_39072.n0 VSS 0.060758f
C12838 a_n3420_39072.t6 VSS 0.029314f
C12839 a_n3420_39072.t4 VSS 0.029314f
C12840 a_n3420_39072.n1 VSS 0.072102f
C12841 a_n3420_39072.n2 VSS 0.269042f
C12842 a_n3420_39072.t9 VSS 0.137711f
C12843 a_n3420_39072.t10 VSS 0.158352f
C12844 a_n3420_39072.n3 VSS 2.11232f
C12845 a_n3420_39072.t11 VSS 0.04602f
C12846 a_n3420_39072.t8 VSS 0.073287f
C12847 a_n3420_39072.n4 VSS 0.10638f
C12848 a_n3420_39072.n5 VSS 8.36947f
C12849 a_n3420_39072.n6 VSS 0.173645f
C12850 a_n3420_39072.t2 VSS 0.045098f
C12851 a_n3420_39072.t1 VSS 0.045098f
C12852 a_n3420_39072.n7 VSS 0.11622f
C12853 a_n3420_39072.n8 VSS 0.312252f
C12854 a_n3420_39072.n9 VSS 0.09479f
C12855 a_n3420_39072.t3 VSS 0.045098f
C12856 a_1666_39043.t2 VSS 0.09052f
C12857 a_1666_39043.t1 VSS 0.314741f
C12858 a_1666_39043.n0 VSS 0.583025f
C12859 a_1666_39043.t3 VSS 0.020581f
C12860 a_1666_39043.t6 VSS 0.032955f
C12861 a_1666_39043.n1 VSS 0.067673f
C12862 a_1666_39043.t5 VSS 0.12908f
C12863 a_1666_39043.t4 VSS 0.07125f
C12864 a_1666_39043.n2 VSS 0.789511f
C12865 a_1666_39043.n3 VSS 0.369162f
C12866 a_1666_39043.n4 VSS 0.352324f
C12867 a_1666_39043.t0 VSS 0.079176f
C12868 a_3232_43370.t0 VSS 0.011595f
C12869 a_3232_43370.n0 VSS 0.017194f
C12870 a_3232_43370.t7 VSS 0.020162f
C12871 a_3232_43370.t23 VSS 0.020098f
C12872 a_3232_43370.t22 VSS 0.010178f
C12873 a_3232_43370.n1 VSS 0.024607f
C12874 a_3232_43370.t21 VSS 0.011466f
C12875 a_3232_43370.n2 VSS 0.013978f
C12876 a_3232_43370.n3 VSS 0.029899f
C12877 a_3232_43370.t6 VSS 0.019194f
C12878 a_3232_43370.t20 VSS 0.020098f
C12879 a_3232_43370.t18 VSS 0.010178f
C12880 a_3232_43370.n4 VSS 0.024607f
C12881 a_3232_43370.t16 VSS 0.010371f
C12882 a_3232_43370.n5 VSS 0.021558f
C12883 a_3232_43370.n6 VSS 0.026301f
C12884 a_3232_43370.n7 VSS 0.208755f
C12885 a_3232_43370.t13 VSS 0.012222f
C12886 a_3232_43370.t11 VSS 0.019481f
C12887 a_3232_43370.n8 VSS 0.034256f
C12888 a_3232_43370.t8 VSS 0.018037f
C12889 a_3232_43370.t9 VSS 0.012919f
C12890 a_3232_43370.n9 VSS 0.049104f
C12891 a_3232_43370.t10 VSS 0.019194f
C12892 a_3232_43370.t17 VSS 0.011984f
C12893 a_3232_43370.n10 VSS 0.038414f
C12894 a_3232_43370.n11 VSS 0.202144f
C12895 a_3232_43370.t19 VSS 0.019509f
C12896 a_3232_43370.t12 VSS 0.012245f
C12897 a_3232_43370.n12 VSS 0.038953f
C12898 a_3232_43370.n13 VSS 0.200182f
C12899 a_3232_43370.t14 VSS 0.013511f
C12900 a_3232_43370.t15 VSS 0.01561f
C12901 a_3232_43370.n14 VSS 0.039634f
C12902 a_3232_43370.n15 VSS 0.465358f
C12903 a_3232_43370.n16 VSS 0.629802f
C12904 a_3232_43370.n17 VSS 0.340125f
C12905 a_3232_43370.n18 VSS 0.066153f
C12906 a_3232_43370.t2 VSS 0.011595f
C12907 a_3232_43370.t3 VSS 0.011595f
C12908 a_3232_43370.n19 VSS 0.025775f
C12909 a_3232_43370.n20 VSS 0.130085f
C12910 a_3232_43370.n21 VSS 0.035206f
C12911 a_3232_43370.t1 VSS 0.011595f
C12912 a_n2293_43922.t3 VSS 0.012f
C12913 a_n2293_43922.n0 VSS 0.471053f
C12914 a_n2293_43922.t2 VSS 0.016814f
C12915 a_n2293_43922.n1 VSS 1.54681f
C12916 a_n2293_43922.n2 VSS 0.028626f
C12917 a_n4064_39616.t0 VSS 0.039069f
C12918 a_n4064_39616.t4 VSS 0.025395f
C12919 a_n4064_39616.t5 VSS 0.025395f
C12920 a_n4064_39616.n0 VSS 0.052635f
C12921 a_n4064_39616.t7 VSS 0.025395f
C12922 a_n4064_39616.t6 VSS 0.025395f
C12923 a_n4064_39616.n1 VSS 0.062462f
C12924 a_n4064_39616.n2 VSS 0.235466f
C12925 a_n4064_39616.t12 VSS 0.063489f
C12926 a_n4064_39616.t10 VSS 0.039867f
C12927 a_n4064_39616.n3 VSS 0.114063f
C12928 a_n4064_39616.t8 VSS 0.496037f
C12929 a_n4064_39616.n4 VSS 0.24639f
C12930 a_n4064_39616.t13 VSS 0.496037f
C12931 a_n4064_39616.t11 VSS 0.497293f
C12932 a_n4064_39616.n5 VSS 0.238372f
C12933 a_n4064_39616.t9 VSS 0.510259f
C12934 a_n4064_39616.n6 VSS 0.460795f
C12935 a_n4064_39616.n7 VSS 3.78678f
C12936 a_n4064_39616.n8 VSS 4.34086f
C12937 a_n4064_39616.n9 VSS 0.150761f
C12938 a_n4064_39616.t2 VSS 0.039069f
C12939 a_n4064_39616.t1 VSS 0.039069f
C12940 a_n4064_39616.n10 VSS 0.100682f
C12941 a_n4064_39616.n11 VSS 0.267779f
C12942 a_n4064_39616.n12 VSS 0.082117f
C12943 a_n4064_39616.t3 VSS 0.039069f
C12944 a_743_42282.t0 VSS 0.021324f
C12945 a_743_42282.t3 VSS 0.021324f
C12946 a_743_42282.t2 VSS 0.021324f
C12947 a_743_42282.n0 VSS 0.043524f
C12948 a_743_42282.t6 VSS 0.032807f
C12949 a_743_42282.t4 VSS 0.032807f
C12950 a_743_42282.n1 VSS 0.081713f
C12951 a_743_42282.n2 VSS 0.168227f
C12952 a_743_42282.t5 VSS 0.021324f
C12953 a_743_42282.t7 VSS 0.021324f
C12954 a_743_42282.n3 VSS 0.043247f
C12955 a_743_42282.t9 VSS 0.044562f
C12956 a_743_42282.t8 VSS 0.028436f
C12957 a_743_42282.n4 VSS 2.08561f
C12958 a_743_42282.n5 VSS 12.505501f
C12959 a_743_42282.n6 VSS 0.05119f
C12960 a_743_42282.n7 VSS 0.185908f
C12961 a_743_42282.n8 VSS 0.068546f
C12962 a_743_42282.t1 VSS 0.021324f
C12963 a_12549_44172.t0 VSS 0.013562f
C12964 a_12549_44172.n0 VSS 0.032647f
C12965 a_12549_44172.t26 VSS 0.014352f
C12966 a_12549_44172.t14 VSS 0.022855f
C12967 a_12549_44172.n1 VSS 0.033718f
C12968 a_12549_44172.t29 VSS 0.016524f
C12969 a_12549_44172.t25 VSS 0.013875f
C12970 a_12549_44172.n2 VSS 0.056865f
C12971 a_12549_44172.t31 VSS 0.018146f
C12972 a_12549_44172.n3 VSS 0.051035f
C12973 a_12549_44172.t24 VSS 0.021096f
C12974 a_12549_44172.t17 VSS 0.012432f
C12975 a_12549_44172.n4 VSS 0.026943f
C12976 a_12549_44172.t15 VSS 0.021096f
C12977 a_12549_44172.t23 VSS 0.012432f
C12978 a_12549_44172.n5 VSS 0.029927f
C12979 a_12549_44172.n6 VSS 0.045707f
C12980 a_12549_44172.t11 VSS 0.021096f
C12981 a_12549_44172.t7 VSS 0.012432f
C12982 a_12549_44172.n7 VSS 0.027772f
C12983 a_12549_44172.t20 VSS 0.021096f
C12984 a_12549_44172.t16 VSS 0.012432f
C12985 a_12549_44172.n8 VSS 0.030258f
C12986 a_12549_44172.n9 VSS 0.023313f
C12987 a_12549_44172.n10 VSS 0.424319f
C12988 a_12549_44172.n11 VSS 1.37361f
C12989 a_12549_44172.t19 VSS 0.016524f
C12990 a_12549_44172.t22 VSS 0.013875f
C12991 a_12549_44172.n12 VSS 0.051141f
C12992 a_12549_44172.n13 VSS 0.353699f
C12993 a_12549_44172.n14 VSS 0.337416f
C12994 a_12549_44172.n15 VSS 0.397216f
C12995 a_12549_44172.t4 VSS 0.022521f
C12996 a_12549_44172.t9 VSS 0.04491f
C12997 a_12549_44172.n16 VSS 1.50627f
C12998 a_12549_44172.t8 VSS 0.015092f
C12999 a_12549_44172.t27 VSS 0.010391f
C13000 a_12549_44172.n17 VSS 0.040996f
C13001 a_12549_44172.n18 VSS 0.786103f
C13002 a_12549_44172.t5 VSS 0.021096f
C13003 a_12549_44172.t30 VSS 0.012432f
C13004 a_12549_44172.n19 VSS 0.034076f
C13005 a_12549_44172.t18 VSS 0.021096f
C13006 a_12549_44172.t10 VSS 0.012432f
C13007 a_12549_44172.n20 VSS 0.041013f
C13008 a_12549_44172.n21 VSS 0.025555f
C13009 a_12549_44172.t13 VSS 0.014024f
C13010 a_12549_44172.t28 VSS 0.022458f
C13011 a_12549_44172.n22 VSS 0.050636f
C13012 a_12549_44172.t21 VSS 0.020587f
C13013 a_12549_44172.n23 VSS 0.076564f
C13014 a_12549_44172.n24 VSS 0.360511f
C13015 a_12549_44172.n25 VSS 0.25078f
C13016 a_12549_44172.n26 VSS 0.345566f
C13017 a_12549_44172.n27 VSS 0.128213f
C13018 a_12549_44172.n28 VSS 0.027135f
C13019 a_12549_44172.t1 VSS 0.013562f
C13020 a_n1925_42282.t2 VSS 0.028923f
C13021 a_n1925_42282.t1 VSS 0.137814f
C13022 a_n1925_42282.t4 VSS 0.040742f
C13023 a_n1925_42282.t3 VSS 0.025998f
C13024 a_n1925_42282.n0 VSS 0.868647f
C13025 a_n1925_42282.n1 VSS 3.21088f
C13026 a_n1925_42282.n2 VSS 0.058075f
C13027 a_n1925_42282.t0 VSS 0.028923f
C13028 a_n1696_34930.n0 VSS 0.021712f
C13029 a_n1696_34930.n1 VSS 0.015537f
C13030 a_n1696_34930.n2 VSS 0.084871f
C13031 a_n1696_34930.t8 VSS 0.070589f
C13032 a_n1696_34930.t14 VSS 0.074374f
C13033 a_n1696_34930.n3 VSS 0.093245f
C13034 a_n1696_34930.t9 VSS 0.070589f
C13035 a_n1696_34930.t10 VSS 0.070589f
C13036 a_n1696_34930.n4 VSS 0.052936f
C13037 a_n1696_34930.n5 VSS 0.049222f
C13038 a_n1696_34930.n6 VSS 0.230592f
C13039 a_n1696_34930.t12 VSS 0.070348f
C13040 a_n1696_34930.t11 VSS 0.074288f
C13041 a_n1696_34930.n7 VSS 0.08614f
C13042 a_n1696_34930.n8 VSS 0.361783f
C13043 a_n1696_34930.t13 VSS 0.070348f
C13044 a_n1696_34930.t15 VSS 0.074288f
C13045 a_n1696_34930.n9 VSS 0.08614f
C13046 a_n1696_34930.n10 VSS 0.232589f
C13047 a_n1696_34930.n11 VSS 0.067856f
C13048 a_n1696_34930.t0 VSS 0.010823f
C13049 a_n1696_34930.t2 VSS 0.010823f
C13050 a_n1696_34930.n12 VSS 0.023975f
C13051 a_n1696_34930.n13 VSS 0.113606f
C13052 a_n1696_34930.t1 VSS 0.010823f
C13053 a_n1696_34930.n14 VSS 0.032955f
C13054 a_n1696_34930.t3 VSS 0.010823f
C13055 a_n1794_35082.t2 VSS 0.015848f
C13056 a_n1794_35082.t3 VSS 0.015848f
C13057 a_n1794_35082.n0 VSS 0.05511f
C13058 a_n1794_35082.t10 VSS 0.037927f
C13059 a_n1794_35082.t11 VSS 0.02235f
C13060 a_n1794_35082.n1 VSS 0.086077f
C13061 a_n1794_35082.n2 VSS 0.067594f
C13062 a_n1794_35082.t17 VSS 0.037927f
C13063 a_n1794_35082.t7 VSS 0.02235f
C13064 a_n1794_35082.t13 VSS 0.037927f
C13065 a_n1794_35082.t14 VSS 0.02235f
C13066 a_n1794_35082.t18 VSS 0.037927f
C13067 a_n1794_35082.t15 VSS 0.02235f
C13068 a_n1794_35082.n3 VSS 0.051121f
C13069 a_n1794_35082.n4 VSS 0.029229f
C13070 a_n1794_35082.n5 VSS 0.054697f
C13071 a_n1794_35082.n6 VSS 0.025032f
C13072 a_n1794_35082.n7 VSS 0.054697f
C13073 a_n1794_35082.n8 VSS 0.025032f
C13074 a_n1794_35082.n9 VSS 0.035252f
C13075 a_n1794_35082.n10 VSS 3.78969f
C13076 a_n1794_35082.t6 VSS 0.037927f
C13077 a_n1794_35082.t9 VSS 0.02235f
C13078 a_n1794_35082.n11 VSS 0.086077f
C13079 a_n1794_35082.n12 VSS 0.067594f
C13080 a_n1794_35082.t5 VSS 0.037927f
C13081 a_n1794_35082.t19 VSS 0.02235f
C13082 a_n1794_35082.t16 VSS 0.037927f
C13083 a_n1794_35082.t4 VSS 0.02235f
C13084 a_n1794_35082.t8 VSS 0.037927f
C13085 a_n1794_35082.t12 VSS 0.02235f
C13086 a_n1794_35082.n13 VSS 0.051121f
C13087 a_n1794_35082.n14 VSS 0.029229f
C13088 a_n1794_35082.n15 VSS 0.054697f
C13089 a_n1794_35082.n16 VSS 0.025032f
C13090 a_n1794_35082.n17 VSS 0.054697f
C13091 a_n1794_35082.n18 VSS 0.025032f
C13092 a_n1794_35082.n19 VSS 0.035233f
C13093 a_n1794_35082.n20 VSS 1.27199f
C13094 a_n1794_35082.n21 VSS 6.43814f
C13095 a_n1794_35082.n22 VSS 1.47506f
C13096 a_n1794_35082.t0 VSS 0.024382f
C13097 a_n1794_35082.n23 VSS 0.049892f
C13098 a_n1794_35082.t1 VSS 0.024382f
C13099 a_n1059_45260.t0 VSS 0.033396f
C13100 a_n1059_45260.t6 VSS 0.021707f
C13101 a_n1059_45260.t5 VSS 0.021707f
C13102 a_n1059_45260.n0 VSS 0.083481f
C13103 a_n1059_45260.t4 VSS 0.021707f
C13104 a_n1059_45260.t7 VSS 0.021707f
C13105 a_n1059_45260.n1 VSS 0.0496f
C13106 a_n1059_45260.n2 VSS 0.218438f
C13107 a_n1059_45260.t8 VSS 0.056279f
C13108 a_n1059_45260.t13 VSS 0.03534f
C13109 a_n1059_45260.n3 VSS 0.081865f
C13110 a_n1059_45260.t16 VSS 0.04462f
C13111 a_n1059_45260.t17 VSS 0.030298f
C13112 a_n1059_45260.n4 VSS 0.121503f
C13113 a_n1059_45260.n5 VSS 0.549435f
C13114 a_n1059_45260.t23 VSS 0.034777f
C13115 a_n1059_45260.t22 VSS 0.05784f
C13116 a_n1059_45260.n6 VSS 0.096815f
C13117 a_n1059_45260.t15 VSS 0.03534f
C13118 a_n1059_45260.t9 VSS 0.056279f
C13119 a_n1059_45260.n7 VSS 0.084597f
C13120 a_n1059_45260.t12 VSS 0.055054f
C13121 a_n1059_45260.t21 VSS 0.103996f
C13122 a_n1059_45260.t11 VSS 0.034456f
C13123 a_n1059_45260.t20 VSS 0.055617f
C13124 a_n1059_45260.n8 VSS 0.236991f
C13125 a_n1059_45260.n9 VSS 1.85405f
C13126 a_n1059_45260.t18 VSS 0.023862f
C13127 a_n1059_45260.t10 VSS 0.022283f
C13128 a_n1059_45260.n10 VSS 0.097822f
C13129 a_n1059_45260.n11 VSS 2.36231f
C13130 a_n1059_45260.t19 VSS 0.030134f
C13131 a_n1059_45260.t14 VSS 0.026116f
C13132 a_n1059_45260.n12 VSS 0.10888f
C13133 a_n1059_45260.n13 VSS 8.52017f
C13134 a_n1059_45260.n14 VSS 1.33814f
C13135 a_n1059_45260.n15 VSS 0.459107f
C13136 a_n1059_45260.n16 VSS 0.588582f
C13137 a_n1059_45260.n17 VSS 0.212257f
C13138 a_n1059_45260.t1 VSS 0.033396f
C13139 a_n1059_45260.t2 VSS 0.033396f
C13140 a_n1059_45260.n18 VSS 0.074585f
C13141 a_n1059_45260.n19 VSS 0.337267f
C13142 a_n1059_45260.n20 VSS 0.10141f
C13143 a_n1059_45260.t3 VSS 0.033396f
C13144 a_2107_46812.t1 VSS 0.042099f
C13145 a_2107_46812.t3 VSS 0.022383f
C13146 a_2107_46812.t2 VSS 0.014021f
C13147 a_2107_46812.n0 VSS 0.420918f
C13148 a_2107_46812.n1 VSS 2.44944f
C13149 a_2107_46812.t0 VSS 0.05114f
C13150 a_584_46384.n0 VSS 0.026356f
C13151 a_584_46384.n1 VSS 0.021696f
C13152 a_584_46384.n2 VSS 0.012891f
C13153 a_584_46384.n3 VSS 0.056771f
C13154 a_584_46384.t17 VSS 0.02535f
C13155 a_584_46384.t10 VSS 0.013346f
C13156 a_584_46384.n4 VSS 0.111514f
C13157 a_584_46384.t15 VSS 0.02535f
C13158 a_584_46384.t21 VSS 0.013346f
C13159 a_584_46384.n5 VSS 0.077665f
C13160 a_584_46384.t20 VSS 0.014627f
C13161 a_584_46384.n6 VSS 0.021967f
C13162 a_584_46384.t19 VSS 0.013501f
C13163 a_584_46384.t22 VSS 0.013501f
C13164 a_584_46384.n7 VSS 0.022653f
C13165 a_584_46384.n8 VSS 0.042234f
C13166 a_584_46384.t16 VSS 0.014416f
C13167 a_584_46384.n9 VSS 0.042051f
C13168 a_584_46384.t13 VSS 0.014508f
C13169 a_584_46384.n10 VSS 0.022424f
C13170 a_584_46384.n11 VSS 0.06835f
C13171 a_584_46384.n12 VSS 0.456232f
C13172 a_584_46384.n13 VSS 0.380237f
C13173 a_584_46384.t9 VSS 0.014627f
C13174 a_584_46384.n14 VSS 0.020583f
C13175 a_584_46384.n15 VSS 0.21734f
C13176 a_584_46384.n16 VSS 0.274116f
C13177 a_584_46384.n17 VSS 0.199244f
C13178 a_584_46384.n18 VSS 0.04641f
C13179 a_584_46384.n19 VSS 0.087654f
C13180 a_584_46384.n20 VSS 0.019384f
C13181 a_n2661_43370.t1 VSS 0.013862f
C13182 a_n2661_43370.t4 VSS 0.019527f
C13183 a_n2661_43370.t3 VSS 0.012461f
C13184 a_n2661_43370.n0 VSS 0.635036f
C13185 a_n2661_43370.t2 VSS 0.062521f
C13186 a_n2661_43370.n1 VSS 4.21397f
C13187 a_n2661_43370.n2 VSS 0.02876f
C13188 a_n2661_43370.t0 VSS 0.013862f
C13189 a_n913_45002.t1 VSS 0.019423f
C13190 a_n913_45002.t8 VSS 0.012625f
C13191 a_n913_45002.t10 VSS 0.012625f
C13192 a_n913_45002.n0 VSS 0.031488f
C13193 a_n913_45002.t9 VSS 0.012625f
C13194 a_n913_45002.t11 VSS 0.012625f
C13195 a_n913_45002.n1 VSS 0.02525f
C13196 a_n913_45002.n2 VSS 0.073705f
C13197 a_n913_45002.t7 VSS 0.019423f
C13198 a_n913_45002.t4 VSS 0.019423f
C13199 a_n913_45002.n3 VSS 0.041965f
C13200 a_n913_45002.t6 VSS 0.019423f
C13201 a_n913_45002.t5 VSS 0.019423f
C13202 a_n913_45002.n4 VSS 0.063872f
C13203 a_n913_45002.n5 VSS 0.177472f
C13204 a_n913_45002.n6 VSS 0.07788f
C13205 a_n913_45002.t0 VSS 0.019423f
C13206 a_n913_45002.t2 VSS 0.019423f
C13207 a_n913_45002.n7 VSS 0.043176f
C13208 a_n913_45002.n8 VSS 0.124427f
C13209 a_n913_45002.t28 VSS 0.032163f
C13210 a_n913_45002.t19 VSS 0.020084f
C13211 a_n913_45002.n9 VSS 0.062344f
C13212 a_n913_45002.t31 VSS 0.032163f
C13213 a_n913_45002.t18 VSS 0.020084f
C13214 a_n913_45002.n10 VSS 0.062344f
C13215 a_n913_45002.t13 VSS 0.032163f
C13216 a_n913_45002.t32 VSS 0.020084f
C13217 a_n913_45002.n11 VSS 0.062344f
C13218 a_n913_45002.t30 VSS 0.032163f
C13219 a_n913_45002.t29 VSS 0.020084f
C13220 a_n913_45002.n12 VSS 0.062294f
C13221 a_n913_45002.t17 VSS 0.032163f
C13222 a_n913_45002.t16 VSS 0.020084f
C13223 a_n913_45002.n13 VSS 0.068192f
C13224 a_n913_45002.n14 VSS 1.20379f
C13225 a_n913_45002.t26 VSS 0.020084f
C13226 a_n913_45002.t23 VSS 0.032163f
C13227 a_n913_45002.n15 VSS 0.062294f
C13228 a_n913_45002.n16 VSS 1.17355f
C13229 a_n913_45002.t14 VSS 0.032163f
C13230 a_n913_45002.t20 VSS 0.020084f
C13231 a_n913_45002.n17 VSS 0.071362f
C13232 a_n913_45002.n18 VSS 0.654182f
C13233 a_n913_45002.t22 VSS 0.032163f
C13234 a_n913_45002.t33 VSS 0.020084f
C13235 a_n913_45002.n19 VSS 0.068811f
C13236 a_n913_45002.n20 VSS 0.720409f
C13237 a_n913_45002.t21 VSS 0.032163f
C13238 a_n913_45002.t24 VSS 0.020084f
C13239 a_n913_45002.n21 VSS 0.062294f
C13240 a_n913_45002.n22 VSS 0.428991f
C13241 a_n913_45002.n23 VSS 0.270174f
C13242 a_n913_45002.n24 VSS 0.262968f
C13243 a_n913_45002.n25 VSS 0.456875f
C13244 a_n913_45002.t27 VSS 0.032163f
C13245 a_n913_45002.t25 VSS 0.020084f
C13246 a_n913_45002.n26 VSS 0.062448f
C13247 a_n913_45002.n27 VSS 0.469632f
C13248 a_n913_45002.t12 VSS 0.020084f
C13249 a_n913_45002.t15 VSS 0.032163f
C13250 a_n913_45002.n28 VSS 0.152273f
C13251 a_n913_45002.n29 VSS 1.21462f
C13252 a_n913_45002.n30 VSS 0.068959f
C13253 a_n913_45002.n31 VSS 0.039f
C13254 a_n913_45002.t3 VSS 0.019423f
C13255 a_1307_43914.t0 VSS 0.024861f
C13256 a_1307_43914.t7 VSS 0.010441f
C13257 a_1307_43914.t4 VSS 0.010441f
C13258 a_1307_43914.n0 VSS 0.036972f
C13259 a_1307_43914.t22 VSS 0.025119f
C13260 a_1307_43914.t33 VSS 0.040094f
C13261 a_1307_43914.n1 VSS 0.080102f
C13262 a_1307_43914.t12 VSS 0.025119f
C13263 a_1307_43914.t29 VSS 0.040094f
C13264 a_1307_43914.n2 VSS 0.067674f
C13265 a_1307_43914.t13 VSS 0.017645f
C13266 a_1307_43914.t18 VSS 0.021374f
C13267 a_1307_43914.n3 VSS 0.072289f
C13268 a_1307_43914.t10 VSS 0.021975f
C13269 a_1307_43914.t26 VSS 0.037291f
C13270 a_1307_43914.n4 VSS 0.050263f
C13271 a_1307_43914.n5 VSS 0.030243f
C13272 a_1307_43914.t19 VSS 0.021975f
C13273 a_1307_43914.t24 VSS 0.037291f
C13274 a_1307_43914.n6 VSS 0.053779f
C13275 a_1307_43914.t21 VSS 0.021975f
C13276 a_1307_43914.t14 VSS 0.037291f
C13277 a_1307_43914.t8 VSS 0.021975f
C13278 a_1307_43914.t20 VSS 0.037291f
C13279 a_1307_43914.n7 VSS 0.062569f
C13280 a_1307_43914.n8 VSS 0.066085f
C13281 a_1307_43914.n9 VSS 0.026196f
C13282 a_1307_43914.n10 VSS 0.187593f
C13283 a_1307_43914.n11 VSS 0.490765f
C13284 a_1307_43914.n12 VSS 0.217581f
C13285 a_1307_43914.n13 VSS 0.511509f
C13286 a_1307_43914.t16 VSS 0.024734f
C13287 a_1307_43914.t32 VSS 0.039924f
C13288 a_1307_43914.n14 VSS 0.083049f
C13289 a_1307_43914.t30 VSS 0.024826f
C13290 a_1307_43914.t23 VSS 0.039741f
C13291 a_1307_43914.n15 VSS 0.075374f
C13292 a_1307_43914.t11 VSS 0.024734f
C13293 a_1307_43914.t34 VSS 0.039924f
C13294 a_1307_43914.n16 VSS 0.083049f
C13295 a_1307_43914.t17 VSS 0.025369f
C13296 a_1307_43914.t9 VSS 0.0404f
C13297 a_1307_43914.n17 VSS 0.207022f
C13298 a_1307_43914.t35 VSS 0.025119f
C13299 a_1307_43914.t15 VSS 0.040094f
C13300 a_1307_43914.n18 VSS 0.070396f
C13301 a_1307_43914.n19 VSS 6.28264f
C13302 a_1307_43914.n20 VSS 0.307297f
C13303 a_1307_43914.n21 VSS 0.27065f
C13304 a_1307_43914.t25 VSS 0.022135f
C13305 a_1307_43914.t27 VSS 0.027406f
C13306 a_1307_43914.n22 VSS 0.156259f
C13307 a_1307_43914.t28 VSS 0.032097f
C13308 a_1307_43914.t31 VSS 0.017645f
C13309 a_1307_43914.n23 VSS 0.059947f
C13310 a_1307_43914.n24 VSS 0.293486f
C13311 a_1307_43914.n25 VSS 0.365001f
C13312 a_1307_43914.n26 VSS 0.188307f
C13313 a_1307_43914.n27 VSS 0.296943f
C13314 a_1307_43914.t6 VSS 0.010441f
C13315 a_1307_43914.t5 VSS 0.010441f
C13316 a_1307_43914.n28 VSS 0.020883f
C13317 a_1307_43914.n29 VSS 0.089306f
C13318 a_1307_43914.n30 VSS 0.195769f
C13319 a_1307_43914.t2 VSS 0.024861f
C13320 a_1307_43914.t1 VSS 0.024861f
C13321 a_1307_43914.n31 VSS 0.050896f
C13322 a_1307_43914.n32 VSS 0.221265f
C13323 a_1307_43914.n33 VSS 0.056968f
C13324 a_1307_43914.t3 VSS 0.024861f
C13325 a_n3565_37414.t7 VSS 0.028251f
C13326 a_n3565_37414.t5 VSS 0.028251f
C13327 a_n3565_37414.n0 VSS 0.107864f
C13328 a_n3565_37414.t4 VSS 0.028251f
C13329 a_n3565_37414.t6 VSS 0.028251f
C13330 a_n3565_37414.n1 VSS 0.064117f
C13331 a_n3565_37414.n2 VSS 0.310226f
C13332 a_n3565_37414.t9 VSS 0.073246f
C13333 a_n3565_37414.t10 VSS 0.045994f
C13334 a_n3565_37414.n3 VSS 0.115851f
C13335 a_n3565_37414.t8 VSS 1.35413f
C13336 a_n3565_37414.n4 VSS 8.067f
C13337 a_n3565_37414.n5 VSS 0.179694f
C13338 a_n3565_37414.t1 VSS 0.043463f
C13339 a_n3565_37414.t0 VSS 0.043463f
C13340 a_n3565_37414.n6 VSS 0.089408f
C13341 a_n3565_37414.n7 VSS 0.395005f
C13342 a_n3565_37414.t2 VSS 0.043463f
C13343 a_n3565_37414.n8 VSS 0.110614f
C13344 a_n3565_37414.t3 VSS 0.043463f
C13345 VREF.t64 VSS 0.575652f
C13346 VREF.t70 VSS 0.568008f
C13347 VREF.n0 VSS 1.59734f
C13348 VREF.t71 VSS 0.568008f
C13349 VREF.n1 VSS 0.826404f
C13350 VREF.t33 VSS 0.568008f
C13351 VREF.n2 VSS 0.826404f
C13352 VREF.t51 VSS 0.568008f
C13353 VREF.n3 VSS 0.824013f
C13354 VREF.t50 VSS 0.568008f
C13355 VREF.n4 VSS 0.824013f
C13356 VREF.t28 VSS 0.277371f
C13357 VREF.t32 VSS 0.277371f
C13358 VREF.n5 VSS 0.698227f
C13359 VREF.n6 VSS 0.847783f
C13360 VREF.t0 VSS 0.277371f
C13361 VREF.t29 VSS 0.277371f
C13362 VREF.n7 VSS 0.698227f
C13363 VREF.n8 VSS 0.852565f
C13364 VREF.t2 VSS 0.277371f
C13365 VREF.t1 VSS 0.277371f
C13366 VREF.n9 VSS 0.698227f
C13367 VREF.n10 VSS 0.850174f
C13368 VREF.t8 VSS 0.277371f
C13369 VREF.t3 VSS 0.277371f
C13370 VREF.n11 VSS 0.698227f
C13371 VREF.n12 VSS 0.850174f
C13372 VREF.t11 VSS 0.277371f
C13373 VREF.t4 VSS 0.277371f
C13374 VREF.n13 VSS 0.698227f
C13375 VREF.n14 VSS 0.852565f
C13376 VREF.t9 VSS 0.277371f
C13377 VREF.t7 VSS 0.277371f
C13378 VREF.n15 VSS 0.698227f
C13379 VREF.n16 VSS 0.850174f
C13380 VREF.t5 VSS 0.277371f
C13381 VREF.t10 VSS 0.277371f
C13382 VREF.n17 VSS 0.698227f
C13383 VREF.n18 VSS 0.850174f
C13384 VREF.t18 VSS 0.277371f
C13385 VREF.t6 VSS 0.277371f
C13386 VREF.n19 VSS 0.698227f
C13387 VREF.n20 VSS 0.850174f
C13388 VREF.t24 VSS 0.277371f
C13389 VREF.t16 VSS 0.277371f
C13390 VREF.n21 VSS 0.698227f
C13391 VREF.n22 VSS 0.850174f
C13392 VREF.t12 VSS 0.277371f
C13393 VREF.t22 VSS 0.277371f
C13394 VREF.n23 VSS 0.698227f
C13395 VREF.n24 VSS 0.852565f
C13396 VREF.t25 VSS 0.277371f
C13397 VREF.t19 VSS 0.277371f
C13398 VREF.n25 VSS 0.698227f
C13399 VREF.n26 VSS 0.850174f
C13400 VREF.t23 VSS 0.277371f
C13401 VREF.t15 VSS 0.277371f
C13402 VREF.n27 VSS 0.698227f
C13403 VREF.n28 VSS 0.850174f
C13404 VREF.t20 VSS 0.277371f
C13405 VREF.t27 VSS 0.277371f
C13406 VREF.n29 VSS 0.698227f
C13407 VREF.n30 VSS 0.850174f
C13408 VREF.t21 VSS 0.277371f
C13409 VREF.t17 VSS 0.277371f
C13410 VREF.n31 VSS 0.698227f
C13411 VREF.n32 VSS 0.850174f
C13412 VREF.t13 VSS 0.277371f
C13413 VREF.t26 VSS 0.277371f
C13414 VREF.n33 VSS 0.698227f
C13415 VREF.n34 VSS 0.852565f
C13416 VREF.t14 VSS 1.15117f
C13417 VREF.n35 VSS 14.191099f
C13418 VREF.t53 VSS 0.575652f
C13419 VREF.t72 VSS 0.568008f
C13420 VREF.n36 VSS 1.59734f
C13421 VREF.t73 VSS 0.568008f
C13422 VREF.n37 VSS 0.826404f
C13423 VREF.t62 VSS 0.568008f
C13424 VREF.n38 VSS 0.826404f
C13425 VREF.t63 VSS 0.568008f
C13426 VREF.n39 VSS 0.824013f
C13427 VREF.t52 VSS 0.568008f
C13428 VREF.n40 VSS 0.824013f
C13429 VREF.t65 VSS 0.277371f
C13430 VREF.t31 VSS 0.277371f
C13431 VREF.n41 VSS 0.698227f
C13432 VREF.n42 VSS 0.847783f
C13433 VREF.t30 VSS 0.277371f
C13434 VREF.t66 VSS 0.277371f
C13435 VREF.n43 VSS 0.698227f
C13436 VREF.n44 VSS 0.852565f
C13437 VREF.t68 VSS 0.277371f
C13438 VREF.t67 VSS 0.277371f
C13439 VREF.n45 VSS 0.698227f
C13440 VREF.n46 VSS 0.850174f
C13441 VREF.t69 VSS 0.277371f
C13442 VREF.t54 VSS 0.277371f
C13443 VREF.n47 VSS 0.698227f
C13444 VREF.n48 VSS 0.850174f
C13445 VREF.t60 VSS 0.277371f
C13446 VREF.t55 VSS 0.277371f
C13447 VREF.n49 VSS 0.698227f
C13448 VREF.n50 VSS 0.852565f
C13449 VREF.t61 VSS 0.277371f
C13450 VREF.t57 VSS 0.277371f
C13451 VREF.n51 VSS 0.698227f
C13452 VREF.n52 VSS 0.850174f
C13453 VREF.t58 VSS 0.277371f
C13454 VREF.t59 VSS 0.277371f
C13455 VREF.n53 VSS 0.698227f
C13456 VREF.n54 VSS 0.850174f
C13457 VREF.t56 VSS 0.277371f
C13458 VREF.t38 VSS 0.277371f
C13459 VREF.n55 VSS 0.698227f
C13460 VREF.n56 VSS 0.850174f
C13461 VREF.t39 VSS 0.277371f
C13462 VREF.t40 VSS 0.277371f
C13463 VREF.n57 VSS 0.698227f
C13464 VREF.n58 VSS 0.850174f
C13465 VREF.t35 VSS 0.277371f
C13466 VREF.t48 VSS 0.277371f
C13467 VREF.n59 VSS 0.698227f
C13468 VREF.n60 VSS 0.852565f
C13469 VREF.t37 VSS 0.277371f
C13470 VREF.t49 VSS 0.277371f
C13471 VREF.n61 VSS 0.698227f
C13472 VREF.n62 VSS 0.850174f
C13473 VREF.t45 VSS 0.277371f
C13474 VREF.t41 VSS 0.277371f
C13475 VREF.n63 VSS 0.698227f
C13476 VREF.n64 VSS 0.850174f
C13477 VREF.t47 VSS 0.277371f
C13478 VREF.t43 VSS 0.277371f
C13479 VREF.n65 VSS 0.698227f
C13480 VREF.n66 VSS 0.850174f
C13481 VREF.t36 VSS 0.277371f
C13482 VREF.t42 VSS 0.277371f
C13483 VREF.n67 VSS 0.698227f
C13484 VREF.n68 VSS 0.850174f
C13485 VREF.t46 VSS 0.277371f
C13486 VREF.t44 VSS 0.277371f
C13487 VREF.n69 VSS 0.698227f
C13488 VREF.n70 VSS 0.852565f
C13489 VREF.t34 VSS 1.15117f
C13490 VREF.n71 VSS 14.264299f
C13491 C8_N_btm.t3 VSS 0.1469f
C13492 C8_N_btm.t2 VSS 0.1469f
C13493 C8_N_btm.n0 VSS 0.453952f
C13494 C8_N_btm.t1 VSS 0.1469f
C13495 C8_N_btm.t0 VSS 0.1469f
C13496 C8_N_btm.n1 VSS 0.468327f
C13497 C8_N_btm.n2 VSS 1.81139f
C13498 C8_N_btm.t6 VSS 0.167162f
C13499 C8_N_btm.t7 VSS 0.167162f
C13500 C8_N_btm.n3 VSS 0.847137f
C13501 C8_N_btm.n4 VSS 1.20098f
C13502 C8_N_btm.t5 VSS 0.167162f
C13503 C8_N_btm.t4 VSS 0.167162f
C13504 C8_N_btm.n5 VSS 0.853379f
C13505 C8_N_btm.n6 VSS 0.927507f
C13506 C8_N_btm.t9 VSS 0.041791f
C13507 C8_N_btm.t8 VSS 0.041791f
C13508 C8_N_btm.n7 VSS 0.156641f
C13509 C8_N_btm.n8 VSS 2.6195f
C13510 C8_N_btm.n9 VSS 2.45029f
C13511 C8_N_btm.n10 VSS 1.08519f
C13512 C8_N_btm.n11 VSS 1.08899f
C13513 C8_N_btm.n12 VSS 1.08899f
C13514 C8_N_btm.n13 VSS 1.08519f
C13515 C8_N_btm.n14 VSS 1.08899f
C13516 C8_N_btm.n15 VSS 1.08899f
C13517 C8_N_btm.n16 VSS 1.08899f
C13518 C8_N_btm.n17 VSS 1.08899f
C13519 C8_N_btm.n18 VSS 1.08519f
C13520 C8_N_btm.n19 VSS 1.08899f
C13521 C8_N_btm.n20 VSS 1.08899f
C13522 C8_N_btm.n21 VSS 1.08519f
C13523 C8_N_btm.n22 VSS 1.08899f
C13524 C8_N_btm.n23 VSS 1.08899f
C13525 C8_N_btm.n24 VSS 1.08899f
C13526 C8_N_btm.n25 VSS 1.05117f
C13527 C8_N_btm.n26 VSS 1.08899f
C13528 C8_N_btm.n27 VSS 1.08899f
C13529 C8_N_btm.n28 VSS 1.08899f
C13530 C8_N_btm.n29 VSS 1.08899f
C13531 C8_N_btm.n30 VSS 1.08919f
C13532 C8_N_btm.n31 VSS 1.08899f
C13533 C8_N_btm.n32 VSS 1.08919f
C13534 C8_N_btm.n33 VSS 0.801269f
C13535 C8_N_btm.n34 VSS 1.08919f
C13536 C8_N_btm.n35 VSS 1.08899f
C13537 C8_N_btm.n36 VSS 1.3689f
C13538 C8_N_btm.n37 VSS 1.08919f
C13539 C8_N_btm.n38 VSS 1.08899f
C13540 C8_N_btm.n39 VSS 1.08919f
C13541 C8_N_btm.n40 VSS 0.801269f
C13542 C8_N_btm.n41 VSS 1.08919f
C13543 C8_N_btm.n42 VSS 1.08899f
C13544 C8_N_btm.n43 VSS 1.3689f
C13545 C8_N_btm.n44 VSS 1.08899f
C13546 C8_N_btm.n45 VSS 1.3689f
C13547 C8_N_btm.n46 VSS 1.08919f
C13548 C8_N_btm.n47 VSS 1.08899f
C13549 C8_N_btm.n48 VSS 1.08919f
C13550 C8_N_btm.n49 VSS 0.801269f
C13551 C8_N_btm.n50 VSS 1.08919f
C13552 C8_N_btm.n51 VSS 1.08899f
C13553 C8_N_btm.n52 VSS 1.3689f
C13554 C8_N_btm.n53 VSS 1.08899f
C13555 C8_N_btm.n54 VSS 1.3689f
C13556 C8_N_btm.n55 VSS 1.08919f
C13557 C8_N_btm.n56 VSS 1.08899f
C13558 C8_N_btm.n57 VSS 1.08919f
C13559 C8_N_btm.n58 VSS 0.801269f
C13560 C8_N_btm.n59 VSS 1.08919f
C13561 C8_N_btm.n60 VSS 1.08899f
C13562 C8_N_btm.n61 VSS 1.3689f
C13563 C8_N_btm.n62 VSS 2.37442f
C13564 C8_N_btm.n63 VSS 1.08899f
C13565 C8_N_btm.n64 VSS 1.08899f
C13566 C8_N_btm.n65 VSS 1.08899f
C13567 C8_N_btm.n66 VSS 1.08899f
C13568 C8_N_btm.n67 VSS 1.08899f
C13569 C8_N_btm.n68 VSS 1.08899f
C13570 C8_N_btm.n69 VSS 1.08899f
C13571 C8_N_btm.n70 VSS 1.08899f
C13572 C8_N_btm.n71 VSS 1.08899f
C13573 C8_N_btm.n72 VSS 1.08899f
C13574 C8_N_btm.n73 VSS 1.08498f
C13575 C8_N_btm.n74 VSS 1.08519f
C13576 C8_N_btm.n75 VSS 1.08519f
C13577 C8_N_btm.n76 VSS 1.08519f
C13578 C8_N_btm.n77 VSS 1.08899f
C13579 C8_N_btm.n78 VSS 1.08519f
C13580 C8_N_btm.n79 VSS 1.08519f
C13581 C8_N_btm.n80 VSS 1.08899f
C13582 C8_N_btm.n81 VSS 1.08899f
C13583 C8_N_btm.n82 VSS 1.08899f
C13584 C8_N_btm.n83 VSS 1.08899f
C13585 C8_N_btm.n84 VSS 1.08899f
C13586 C8_N_btm.n85 VSS 1.08899f
C13587 C8_N_btm.n86 VSS 1.08899f
C13588 C8_N_btm.n87 VSS 1.08519f
C13589 C8_N_btm.n88 VSS 1.08519f
C13590 C8_N_btm.n89 VSS 1.08519f
C13591 C8_N_btm.n90 VSS 1.3941f
C13592 C8_N_btm.n91 VSS 1.08899f
C13593 C8_N_btm.n92 VSS 1.31162f
C13594 C8_N_btm.n93 VSS 1.08899f
C13595 C8_N_btm.n94 VSS 1.7059f
C13596 C8_N_btm.n95 VSS 1.08919f
C13597 C8_N_btm.n96 VSS 1.08919f
C13598 C8_N_btm.n97 VSS 0.801269f
C13599 C8_N_btm.n98 VSS 0.801269f
C13600 C8_N_btm.n99 VSS 1.55307f
C13601 C8_N_btm.n100 VSS 1.08919f
C13602 C8_N_btm.n101 VSS 1.08919f
C13603 C8_N_btm.n102 VSS 1.08899f
C13604 C8_N_btm.n103 VSS 1.08899f
C13605 C8_N_btm.n104 VSS 1.08519f
C13606 C8_N_btm.n105 VSS 1.08519f
C13607 C8_N_btm.n106 VSS 1.08519f
C13608 C8_N_btm.n107 VSS 1.08519f
C13609 C8_N_btm.n108 VSS 1.08519f
C13610 C8_N_btm.n109 VSS 1.08519f
C13611 C8_N_btm.n110 VSS 1.08899f
C13612 C8_N_btm.n111 VSS 1.08899f
C13613 C8_N_btm.n112 VSS 1.08519f
C13614 C8_N_btm.n113 VSS 1.08519f
C13615 C8_N_btm.n114 VSS 1.08519f
C13616 C8_N_btm.n115 VSS 1.08519f
C13617 C8_N_btm.n116 VSS 1.08519f
C13618 C8_N_btm.n117 VSS 1.39409f
C13619 C8_N_btm.n118 VSS 1.08899f
C13620 C8_N_btm.n119 VSS 1.08899f
C13621 C8_N_btm.n120 VSS 3.37102f
C13622 C8_N_btm.n121 VSS 7.05447f
C13623 C8_N_btm.n122 VSS 3.37113f
C13624 C8_N_btm.n123 VSS 1.08899f
C13625 C8_N_btm.n124 VSS 1.08899f
C13626 C8_N_btm.n125 VSS 1.08899f
C13627 C8_N_btm.n126 VSS 1.08899f
C13628 C8_N_btm.n127 VSS 1.08899f
C13629 C8_N_btm.n128 VSS 1.08899f
C13630 C8_N_btm.n129 VSS 1.08899f
C13631 C8_N_btm.n130 VSS 1.08899f
C13632 C8_N_btm.n131 VSS 1.08899f
C13633 C8_N_btm.n132 VSS 1.08899f
C13634 C8_N_btm.n133 VSS 1.08899f
C13635 C8_N_btm.n134 VSS 1.08899f
C13636 C8_N_btm.n135 VSS 1.08899f
C13637 C8_N_btm.n136 VSS 1.08899f
C13638 C8_N_btm.n137 VSS 1.08899f
C13639 C8_N_btm.n138 VSS 1.08899f
C13640 C8_N_btm.n139 VSS 1.08899f
C13641 C8_N_btm.n140 VSS 1.08899f
C13642 C8_N_btm.n141 VSS 1.08899f
C13643 C8_N_btm.n142 VSS 1.05117f
C13644 C8_N_btm.n143 VSS 1.48639f
C13645 C8_N_btm.n144 VSS 1.08899f
C13646 C8_N_btm.n145 VSS 1.08919f
C13647 C8_N_btm.n146 VSS 0.801269f
C13648 C8_N_btm.n147 VSS 0.801269f
C13649 C8_N_btm.n148 VSS 1.08919f
C13650 C8_N_btm.n149 VSS 0.801269f
C13651 C8_N_btm.n150 VSS 0.801269f
C13652 C8_N_btm.n151 VSS 0.801269f
C13653 C8_N_btm.n152 VSS 1.08919f
C13654 C8_N_btm.n153 VSS 1.08899f
C13655 C8_N_btm.n154 VSS 1.08899f
C13656 C8_N_btm.n155 VSS 1.3689f
C13657 C8_N_btm.n156 VSS 1.3689f
C13658 C8_N_btm.n157 VSS 1.3689f
C13659 C8_N_btm.n158 VSS 1.3689f
C13660 C8_N_btm.n159 VSS 1.08899f
C13661 C8_N_btm.n160 VSS 1.08919f
C13662 C8_N_btm.n161 VSS 0.801269f
C13663 C8_N_btm.n162 VSS 0.801269f
C13664 C8_N_btm.n163 VSS 1.08919f
C13665 C8_N_btm.n164 VSS 0.801269f
C13666 C8_N_btm.n165 VSS 1.87973f
C13667 C8_N_btm.n166 VSS 1.89339f
C13668 C8_N_btm.n167 VSS 1.08899f
C13669 C8_N_btm.n168 VSS 1.08899f
C13670 C8_N_btm.n169 VSS 1.08899f
C13671 C8_N_btm.n170 VSS 1.3689f
C13672 C8_N_btm.n171 VSS 1.3689f
C13673 C8_N_btm.n172 VSS 1.3689f
C13674 C8_N_btm.n173 VSS 1.3689f
C13675 C8_N_btm.n174 VSS 1.08899f
C13676 C8_N_btm.n175 VSS 1.08919f
C13677 C8_N_btm.n176 VSS 0.801269f
C13678 C8_N_btm.n177 VSS 0.801269f
C13679 C8_N_btm.n178 VSS 0.801269f
C13680 C8_N_btm.n179 VSS 1.08919f
C13681 C8_N_btm.n180 VSS 0.801269f
C13682 C8_N_btm.n181 VSS 0.801269f
C13683 C8_N_btm.n182 VSS 0.801269f
C13684 C8_N_btm.n183 VSS 1.08919f
C13685 C8_N_btm.n184 VSS 1.08899f
C13686 C8_N_btm.n185 VSS 1.08899f
C13687 C8_N_btm.n186 VSS 1.3689f
C13688 C8_N_btm.n187 VSS 1.3689f
C13689 C8_N_btm.n188 VSS 1.48639f
C13690 C8_N_btm.n189 VSS 1.08899f
C13691 C8_N_btm.n190 VSS 1.08899f
C13692 C8_N_btm.n191 VSS 1.08919f
C13693 C8_N_btm.n192 VSS 1.08919f
C13694 C8_N_btm.n193 VSS 0.801269f
C13695 C8_N_btm.n194 VSS 0.801269f
C13696 C8_N_btm.n195 VSS 1.08519f
C13697 C8_N_btm.n196 VSS 1.08519f
C13698 C8_N_btm.n197 VSS 1.08519f
C13699 C8_N_btm.n198 VSS 1.08519f
C13700 C8_N_btm.n199 VSS 1.08519f
C13701 C8_N_btm.n200 VSS 1.08519f
C13702 C8_N_btm.n201 VSS 1.08519f
C13703 C8_N_btm.n202 VSS 1.08519f
C13704 C8_N_btm.n203 VSS 1.08519f
C13705 C8_N_btm.n204 VSS 1.08519f
C13706 C8_N_btm.n205 VSS 1.3941f
C13707 C8_N_btm.n206 VSS 4.75242f
C13708 C8_N_btm.n207 VSS 3.37113f
C13709 C8_N_btm.n208 VSS 1.08899f
C13710 C8_N_btm.n209 VSS 1.08899f
C13711 C8_N_btm.n210 VSS 1.08899f
C13712 C8_N_btm.n211 VSS 1.08899f
C13713 C8_N_btm.n212 VSS 1.08899f
C13714 C8_N_btm.n213 VSS 1.08899f
C13715 C8_N_btm.n214 VSS 1.08899f
C13716 C8_N_btm.n215 VSS 1.08899f
C13717 C8_N_btm.n216 VSS 1.08899f
C13718 C8_N_btm.n217 VSS 1.08899f
C13719 C8_N_btm.n218 VSS 1.08899f
C13720 C8_N_btm.n219 VSS 1.08899f
C13721 C8_N_btm.n220 VSS 1.08899f
C13722 C8_N_btm.n221 VSS 1.08899f
C13723 C8_N_btm.n222 VSS 1.08899f
C13724 C8_N_btm.n223 VSS 1.08899f
C13725 C8_N_btm.n224 VSS 1.08899f
C13726 C8_N_btm.n225 VSS 1.08519f
C13727 C8_N_btm.n226 VSS 1.31159f
C13728 C8_N_btm.n227 VSS 1.70573f
C13729 C8_N_btm.n228 VSS 1.55307f
C13730 C8_N_btm.n229 VSS 1.08919f
C13731 C8_N_btm.n230 VSS 1.08899f
C13732 C8_N_btm.n231 VSS 1.08899f
C13733 C8_N_btm.n232 VSS 1.08899f
C13734 C8_N_btm.n233 VSS 1.08899f
C13735 C8_N_btm.n234 VSS 2.37442f
C13736 C8_N_btm.n235 VSS 1.08519f
C13737 C8_N_btm.n236 VSS 1.08519f
C13738 C8_N_btm.n237 VSS 1.08899f
C13739 C8_N_btm.n238 VSS 1.08899f
C13740 C8_N_btm.n239 VSS 1.08899f
C13741 C8_N_btm.n240 VSS 1.08899f
C13742 C8_N_btm.n241 VSS 1.08519f
C13743 C8_N_btm.n242 VSS 1.08519f
C13744 C8_N_btm.n243 VSS 1.08519f
C13745 C8_N_btm.n244 VSS 1.08519f
C13746 C8_N_btm.n245 VSS 1.08899f
C13747 C8_N_btm.n246 VSS 1.08899f
C13748 C8_N_btm.n247 VSS 1.08899f
C13749 C8_N_btm.n248 VSS 1.08899f
C13750 C8_N_btm.n249 VSS 1.08519f
C13751 C8_N_btm.n250 VSS 2.45819f
C13752 a_21076_30879.t5 VSS 1.26097f
C13753 a_21076_30879.t4 VSS 1.26078f
C13754 a_21076_30879.n0 VSS 0.933964f
C13755 a_21076_30879.t6 VSS 1.26078f
C13756 a_21076_30879.n1 VSS 0.473043f
C13757 a_21076_30879.t7 VSS 1.26078f
C13758 a_21076_30879.n2 VSS 5.6323f
C13759 a_21076_30879.t3 VSS 0.024211f
C13760 a_21076_30879.t2 VSS 0.024211f
C13761 a_21076_30879.n3 VSS 0.048421f
C13762 a_21076_30879.n4 VSS 4.53429f
C13763 a_21076_30879.t0 VSS 0.037247f
C13764 a_21076_30879.n5 VSS 0.111767f
C13765 a_21076_30879.t1 VSS 0.037247f
C13766 a_14021_43940.t1 VSS 0.050229f
C13767 a_14021_43940.t3 VSS 0.02181f
C13768 a_14021_43940.t2 VSS 0.013917f
C13769 a_14021_43940.n0 VSS 0.447484f
C13770 a_14021_43940.n1 VSS 2.51054f
C13771 a_14021_43940.t0 VSS 0.056022f
C13772 a_3626_43646.t0 VSS 0.030173f
C13773 a_3626_43646.t2 VSS 0.030173f
C13774 a_3626_43646.t5 VSS 0.030173f
C13775 a_3626_43646.n0 VSS 0.061305f
C13776 a_3626_43646.t3 VSS 0.019612f
C13777 a_3626_43646.t4 VSS 0.019612f
C13778 a_3626_43646.n1 VSS 0.039772f
C13779 a_3626_43646.t6 VSS 0.040985f
C13780 a_3626_43646.t7 VSS 0.026154f
C13781 a_3626_43646.n2 VSS 1.63441f
C13782 a_3626_43646.n3 VSS 9.535339f
C13783 a_3626_43646.n4 VSS 0.229142f
C13784 a_3626_43646.n5 VSS 0.072972f
C13785 a_3626_43646.t1 VSS 0.030173f
C13786 a_n2810_45028.t5 VSS 0.095357f
C13787 a_n2810_45028.t4 VSS 0.059485f
C13788 a_n2810_45028.n0 VSS 2.16904f
C13789 a_n2810_45028.t2 VSS 0.037537f
C13790 a_n2810_45028.t3 VSS 0.037537f
C13791 a_n2810_45028.n1 VSS 0.075075f
C13792 a_n2810_45028.n2 VSS 9.03718f
C13793 a_n2810_45028.t0 VSS 0.05775f
C13794 a_n2810_45028.n3 VSS 0.173288f
C13795 a_n2810_45028.t1 VSS 0.05775f
C13796 VDAC_Ni.t9 VSS 0.031209f
C13797 VDAC_Ni.t10 VSS 0.089861f
C13798 VDAC_Ni.t4 VSS 0.106007f
C13799 VDAC_Ni.n0 VSS 1.2327f
C13800 VDAC_Ni.t1 VSS 0.02843f
C13801 VDAC_Ni.t2 VSS 0.02843f
C13802 VDAC_Ni.n1 VSS 0.062743f
C13803 VDAC_Ni.t0 VSS 0.02843f
C13804 VDAC_Ni.t3 VSS 0.02843f
C13805 VDAC_Ni.n2 VSS 0.062352f
C13806 VDAC_Ni.n3 VSS 0.429559f
C13807 VDAC_Ni.n4 VSS 0.242952f
C13808 VDAC_Ni.t5 VSS 0.02843f
C13809 VDAC_Ni.t6 VSS 0.02843f
C13810 VDAC_Ni.n5 VSS 0.072657f
C13811 VDAC_Ni.n6 VSS 0.158267f
C13812 VDAC_Ni.t7 VSS 0.02843f
C13813 VDAC_Ni.t8 VSS 0.02843f
C13814 VDAC_Ni.n7 VSS 0.072657f
C13815 VDAC_Ni.n8 VSS 0.163297f
C13816 VDAC_Ni.n9 VSS 0.038628f
C13817 a_2437_43646.t1 VSS 0.013323f
C13818 a_2437_43646.t2 VSS 0.013323f
C13819 a_2437_43646.n0 VSS 0.026753f
C13820 a_2437_43646.t3 VSS 0.018768f
C13821 a_2437_43646.t4 VSS 0.011976f
C13822 a_2437_43646.n1 VSS 1.52651f
C13823 a_2437_43646.n2 VSS 5.52586f
C13824 a_2437_43646.t0 VSS 0.063485f
C13825 a_n443_46116.t0 VSS 0.012987f
C13826 a_n443_46116.t2 VSS 0.012987f
C13827 a_n443_46116.t1 VSS 0.012987f
C13828 a_n443_46116.n0 VSS 0.039437f
C13829 a_n443_46116.n1 VSS 0.032464f
C13830 a_n443_46116.n2 VSS 0.019289f
C13831 a_n443_46116.n3 VSS 0.107432f
C13832 a_n443_46116.t20 VSS 0.037932f
C13833 a_n443_46116.t23 VSS 0.01997f
C13834 a_n443_46116.n4 VSS 0.104594f
C13835 a_n443_46116.t24 VSS 0.021708f
C13836 a_n443_46116.t15 VSS 0.013598f
C13837 a_n443_46116.n5 VSS 0.052648f
C13838 a_n443_46116.n6 VSS 0.658435f
C13839 a_n443_46116.t14 VSS 0.021886f
C13840 a_n443_46116.t17 VSS 0.013743f
C13841 a_n443_46116.n7 VSS 0.047404f
C13842 a_n443_46116.t21 VSS 0.021708f
C13843 a_n443_46116.t10 VSS 0.013598f
C13844 a_n443_46116.n8 VSS 0.063076f
C13845 a_n443_46116.t18 VSS 0.021572f
C13846 a_n443_46116.t13 VSS 0.013473f
C13847 a_n443_46116.n9 VSS 0.041694f
C13848 a_n443_46116.n10 VSS 0.09651f
C13849 a_n443_46116.t9 VSS 0.021498f
C13850 a_n443_46116.t19 VSS 0.013423f
C13851 a_n443_46116.n11 VSS 0.04202f
C13852 a_n443_46116.n12 VSS 0.075939f
C13853 a_n443_46116.n13 VSS 0.29872f
C13854 a_n443_46116.t8 VSS 0.013743f
C13855 a_n443_46116.t11 VSS 0.021886f
C13856 a_n443_46116.n14 VSS 0.03206f
C13857 a_n443_46116.n15 VSS 0.302639f
C13858 a_n443_46116.n16 VSS 0.468214f
C13859 a_n443_46116.t25 VSS 0.02147f
C13860 a_n443_46116.t22 VSS 0.013399f
C13861 a_n443_46116.n17 VSS 0.044202f
C13862 a_n443_46116.n18 VSS 0.18702f
C13863 a_n443_46116.t12 VSS 0.037932f
C13864 a_n443_46116.t16 VSS 0.01997f
C13865 a_n443_46116.n19 VSS 0.097609f
C13866 a_n443_46116.n20 VSS 0.359625f
C13867 a_n443_46116.n21 VSS 0.141433f
C13868 a_n443_46116.n22 VSS 0.110305f
C13869 a_n443_46116.n23 VSS 0.029005f
C13870 a_n443_46116.t3 VSS 0.012987f
C13871 a_16327_47482.n0 VSS 0.012337f
C13872 a_16327_47482.n3 VSS 0.042856f
C13873 a_16327_47482.n4 VSS 0.015425f
C13874 a_16327_47482.n5 VSS 0.014976f
C13875 a_16327_47482.n6 VSS 0.091623f
C13876 a_16327_47482.n7 VSS 0.01543f
C13877 a_16327_47482.n8 VSS 0.014951f
C13878 a_16327_47482.n9 VSS 0.104834f
C13879 a_16327_47482.n10 VSS 0.021633f
C13880 a_16327_47482.n11 VSS 0.014797f
C13881 a_16327_47482.n12 VSS 0.015832f
C13882 a_16327_47482.n13 VSS 0.15431f
C13883 a_16327_47482.n14 VSS 0.015425f
C13884 a_16327_47482.n15 VSS 0.014976f
C13885 a_16327_47482.n16 VSS 0.086605f
C13886 a_16327_47482.n17 VSS 0.069143f
C13887 a_16327_47482.n18 VSS 0.015425f
C13888 a_16327_47482.n19 VSS 0.014976f
C13889 a_16327_47482.n20 VSS 0.17056f
C13890 a_16327_47482.n21 VSS 0.129153f
C13891 a_16327_47482.n22 VSS 0.157797f
C13892 a_16327_47482.n23 VSS 0.014951f
C13893 a_16327_47482.n24 VSS 0.015429f
C13894 a_16327_47482.n25 VSS 0.095238f
C13895 a_16327_47482.n26 VSS 0.085419f
C13896 a_16327_47482.n27 VSS 0.020983f
C13897 a_16327_47482.n28 VSS 0.014312f
C13898 a_16327_47482.n29 VSS 0.015787f
C13899 a_16327_47482.n30 VSS 0.071652f
C13900 a_16327_47482.n31 VSS 0.011591f
C13901 a_16327_47482.n32 VSS 0.032013f
C13902 a_16327_47482.n33 VSS 0.015398f
C13903 a_16327_47482.n34 VSS 0.014984f
C13904 a_16327_47482.n35 VSS 0.095142f
C13905 a_16327_47482.n36 VSS 0.036674f
C13906 a_16327_47482.n37 VSS 0.096742f
C13907 a_16327_47482.n38 VSS 0.015398f
C13908 a_16327_47482.n39 VSS 0.014984f
C13909 a_16327_47482.n40 VSS 0.102981f
C13910 a_16327_47482.n41 VSS 0.392319f
C13911 a_16327_47482.n42 VSS 0.107563f
C13912 a_16327_47482.n43 VSS 0.025729f
C13913 a_16327_47482.n44 VSS 0.033747f
C13914 a_16327_47482.n45 VSS 0.011022f
C13915 a_n1613_43370.t25 VSS 0.012263f
C13916 a_n1613_43370.n0 VSS 0.026692f
C13917 a_n1613_43370.t40 VSS 0.014088f
C13918 a_n1613_43370.n1 VSS 0.024986f
C13919 a_n1613_43370.n2 VSS 0.249079f
C13920 a_n1613_43370.t27 VSS 0.014088f
C13921 a_n1613_43370.n3 VSS 0.026044f
C13922 a_n1613_43370.t43 VSS 0.012263f
C13923 a_n1613_43370.n4 VSS 0.025286f
C13924 a_n1613_43370.n5 VSS 0.146136f
C13925 a_n1613_43370.n6 VSS 0.292344f
C13926 a_n1613_43370.n7 VSS 0.277067f
C13927 a_n1613_43370.t32 VSS 0.012263f
C13928 a_n1613_43370.n8 VSS 0.025286f
C13929 a_n1613_43370.n9 VSS 0.092573f
C13930 a_n1613_43370.n10 VSS 0.034616f
C13931 a_n1613_43370.t8 VSS 0.014088f
C13932 a_n1613_43370.n11 VSS 0.026045f
C13933 a_n1613_43370.t23 VSS 0.012263f
C13934 a_n1613_43370.n12 VSS 0.025286f
C13935 a_n1613_43370.n13 VSS 0.172491f
C13936 a_n1613_43370.t13 VSS 0.014088f
C13937 a_n1613_43370.n14 VSS 0.026044f
C13938 a_n1613_43370.t30 VSS 0.012263f
C13939 a_n1613_43370.n15 VSS 0.025286f
C13940 a_n1613_43370.n16 VSS 0.192441f
C13941 a_n1613_43370.n17 VSS 0.116568f
C13942 a_n1613_43370.t38 VSS 0.014088f
C13943 a_n1613_43370.n18 VSS 0.026045f
C13944 a_n1613_43370.t45 VSS 0.012263f
C13945 a_n1613_43370.n19 VSS 0.025286f
C13946 a_n1613_43370.n20 VSS 0.159451f
C13947 a_n1613_43370.n21 VSS 0.051079f
C13948 a_n1613_43370.t9 VSS 0.014088f
C13949 a_n1613_43370.n22 VSS 0.025998f
C13950 a_n1613_43370.t41 VSS 0.012263f
C13951 a_n1613_43370.n23 VSS 0.025299f
C13952 a_n1613_43370.n24 VSS 0.182978f
C13953 a_n1613_43370.n25 VSS 0.145875f
C13954 a_n1613_43370.t14 VSS 0.014088f
C13955 a_n1613_43370.n26 VSS 0.026f
C13956 a_n1613_43370.t42 VSS 0.012263f
C13957 a_n1613_43370.n27 VSS 0.025299f
C13958 a_n1613_43370.n28 VSS 0.165759f
C13959 a_n1613_43370.n29 VSS 0.216549f
C13960 a_n1613_43370.t46 VSS 0.014088f
C13961 a_n1613_43370.n30 VSS 0.025853f
C13962 a_n1613_43370.t37 VSS 0.012263f
C13963 a_n1613_43370.n31 VSS 0.025293f
C13964 a_n1613_43370.n32 VSS 0.165832f
C13965 a_n1613_43370.n33 VSS 0.297949f
C13966 a_n1613_43370.t36 VSS 0.014088f
C13967 a_n1613_43370.n34 VSS 0.026002f
C13968 a_n1613_43370.t28 VSS 0.012263f
C13969 a_n1613_43370.n35 VSS 0.025299f
C13970 a_n1613_43370.n36 VSS 0.143676f
C13971 a_n1613_43370.n37 VSS 0.190996f
C13972 a_n1613_43370.t12 VSS 0.014088f
C13973 a_n1613_43370.n38 VSS 0.024165f
C13974 a_n1613_43370.n39 VSS 0.01957f
C13975 a_n1613_43370.n40 VSS 0.075455f
C13976 a_n1613_43370.n41 VSS 0.066842f
C13977 a_n1613_43370.n42 VSS 0.147376f
C13978 a_n1613_43370.n43 VSS 0.018181f
C13979 a_n1613_43370.n44 VSS 0.036992f
C13980 a_n1613_43370.n45 VSS 0.013519f
C13981 a_n1613_43370.n47 VSS 0.081565f
C13982 a_n1613_43370.n48 VSS 0.055964f
C13983 a_n1613_43370.n49 VSS 0.01861f
C13984 a_5937_45572.t0 VSS 0.011931f
C13985 a_5937_45572.t14 VSS 0.013084f
C13986 a_5937_45572.n0 VSS 0.043652f
C13987 a_5937_45572.t13 VSS 0.01989f
C13988 a_5937_45572.t7 VSS 0.012448f
C13989 a_5937_45572.n1 VSS 0.034945f
C13990 a_5937_45572.t6 VSS 0.020075f
C13991 a_5937_45572.t19 VSS 0.0126f
C13992 a_5937_45572.n2 VSS 0.036311f
C13993 a_5937_45572.t16 VSS 0.01231f
C13994 a_5937_45572.t8 VSS 0.019725f
C13995 a_5937_45572.n3 VSS 0.045426f
C13996 a_5937_45572.n4 VSS 0.248331f
C13997 a_5937_45572.n5 VSS 0.207625f
C13998 a_5937_45572.t12 VSS 0.012493f
C13999 a_5937_45572.t10 VSS 0.019943f
C14000 a_5937_45572.n6 VSS 0.043141f
C14001 a_5937_45572.n7 VSS 0.224045f
C14002 a_5937_45572.t15 VSS 0.012332f
C14003 a_5937_45572.t4 VSS 0.019751f
C14004 a_5937_45572.n8 VSS 0.038554f
C14005 a_5937_45572.n9 VSS 0.140166f
C14006 a_5937_45572.t5 VSS 0.012626f
C14007 a_5937_45572.t17 VSS 0.020107f
C14008 a_5937_45572.n10 VSS 0.029197f
C14009 a_5937_45572.t18 VSS 0.012626f
C14010 a_5937_45572.t11 VSS 0.020107f
C14011 a_5937_45572.n11 VSS 0.035877f
C14012 a_5937_45572.n12 VSS 0.225037f
C14013 a_5937_45572.n13 VSS 0.143874f
C14014 a_5937_45572.n14 VSS 0.26234f
C14015 a_5937_45572.n15 VSS 0.015511f
C14016 a_5937_45572.n16 VSS 0.104507f
C14017 a_5937_45572.n17 VSS 0.032982f
C14018 a_5937_45572.t1 VSS 0.011931f
C14019 a_n755_45592.t1 VSS 0.013731f
C14020 a_n755_45592.t2 VSS 0.013731f
C14021 a_n755_45592.t0 VSS 0.013731f
C14022 a_n755_45592.n0 VSS 0.041696f
C14023 a_n755_45592.n1 VSS 0.034324f
C14024 a_n755_45592.n2 VSS 0.020393f
C14025 a_n755_45592.n3 VSS 0.113586f
C14026 a_n755_45592.n4 VSS 0.035828f
C14027 a_n755_45592.t25 VSS 0.014167f
C14028 a_n755_45592.t11 VSS 0.0227f
C14029 a_n755_45592.n5 VSS 0.046011f
C14030 a_n755_45592.t20 VSS 0.022636f
C14031 a_n755_45592.t14 VSS 0.05417f
C14032 a_n755_45592.t8 VSS 0.022952f
C14033 a_n755_45592.t18 VSS 0.014377f
C14034 a_n755_45592.n6 VSS 0.037017f
C14035 a_n755_45592.n7 VSS 0.581893f
C14036 a_n755_45592.n8 VSS 0.229005f
C14037 a_n755_45592.n9 VSS 0.037214f
C14038 a_n755_45592.n10 VSS 0.163441f
C14039 a_n755_45592.n11 VSS 0.275218f
C14040 a_n755_45592.t10 VSS 0.022867f
C14041 a_n755_45592.t27 VSS 0.014167f
C14042 a_n755_45592.n12 VSS 0.047568f
C14043 a_n755_45592.t26 VSS 0.01246f
C14044 a_n755_45592.n13 VSS 0.02997f
C14045 a_n755_45592.t21 VSS 0.018609f
C14046 a_n755_45592.t9 VSS 0.012678f
C14047 a_n755_45592.n14 VSS 0.166044f
C14048 a_n755_45592.n15 VSS 1.10975f
C14049 a_n755_45592.n16 VSS 0.322955f
C14050 a_n755_45592.t23 VSS 0.02314f
C14051 a_n755_45592.t16 VSS 0.01453f
C14052 a_n755_45592.n17 VSS 0.035164f
C14053 a_n755_45592.n18 VSS 0.284269f
C14054 a_n755_45592.t24 VSS 0.014299f
C14055 a_n755_45592.t13 VSS 0.023782f
C14056 a_n755_45592.n19 VSS 0.040175f
C14057 a_n755_45592.n20 VSS 0.225564f
C14058 a_n755_45592.n21 VSS 0.252591f
C14059 a_n755_45592.n22 VSS 0.077209f
C14060 a_n755_45592.n23 VSS 0.116624f
C14061 a_n755_45592.n24 VSS 0.030667f
C14062 a_n755_45592.t3 VSS 0.013731f
C14063 a_526_44458.t1 VSS 0.01078f
C14064 a_526_44458.n0 VSS 0.016031f
C14065 a_526_44458.n1 VSS 0.010031f
C14066 a_526_44458.n2 VSS 0.096721f
C14067 a_526_44458.t0 VSS 0.01078f
C14068 a_526_44458.t2 VSS 0.01078f
C14069 a_526_44458.n3 VSS 0.022069f
C14070 a_526_44458.n4 VSS 0.066363f
C14071 a_526_44458.t11 VSS 0.016169f
C14072 a_526_44458.n5 VSS 0.021794f
C14073 a_526_44458.t16 VSS 0.016169f
C14074 a_526_44458.n6 VSS 0.021794f
C14075 a_526_44458.n7 VSS 0.014024f
C14076 a_526_44458.t23 VSS 0.011f
C14077 a_526_44458.t20 VSS 0.017517f
C14078 a_526_44458.n8 VSS 0.033303f
C14079 a_526_44458.n9 VSS 0.226931f
C14080 a_526_44458.t26 VSS 0.011011f
C14081 a_526_44458.t28 VSS 0.02174f
C14082 a_526_44458.n10 VSS 0.021942f
C14083 a_526_44458.t15 VSS 0.02174f
C14084 a_526_44458.t14 VSS 0.011011f
C14085 a_526_44458.n11 VSS 0.088498f
C14086 a_526_44458.n12 VSS 0.713793f
C14087 a_526_44458.t29 VSS 0.011f
C14088 a_526_44458.t22 VSS 0.017517f
C14089 a_526_44458.n13 VSS 0.023875f
C14090 a_526_44458.t34 VSS 0.02174f
C14091 a_526_44458.t12 VSS 0.011011f
C14092 a_526_44458.n14 VSS 0.029605f
C14093 a_526_44458.n15 VSS 0.231774f
C14094 a_526_44458.n16 VSS 0.129067f
C14095 a_526_44458.t17 VSS 0.017331f
C14096 a_526_44458.t9 VSS 0.010884f
C14097 a_526_44458.n17 VSS 0.045055f
C14098 a_526_44458.t13 VSS 0.017464f
C14099 a_526_44458.t30 VSS 0.010957f
C14100 a_526_44458.n18 VSS 0.032458f
C14101 a_526_44458.n19 VSS 0.509129f
C14102 a_526_44458.n20 VSS 0.030142f
C14103 a_526_44458.t10 VSS 0.016169f
C14104 a_526_44458.t21 VSS 0.016169f
C14105 a_526_44458.t18 VSS 0.016169f
C14106 a_526_44458.n21 VSS 0.021794f
C14107 a_526_44458.n22 VSS 0.012676f
C14108 a_526_44458.n23 VSS 0.023319f
C14109 a_526_44458.n24 VSS 0.010672f
C14110 a_526_44458.n25 VSS 0.026346f
C14111 a_526_44458.t8 VSS 0.016169f
C14112 a_526_44458.n26 VSS 0.035847f
C14113 a_526_44458.n28 VSS 0.044853f
C14114 a_526_44458.n29 VSS 0.298278f
C14115 a_526_44458.n30 VSS 0.533208f
C14116 a_526_44458.n31 VSS 0.175291f
C14117 a_526_44458.t32 VSS 0.017331f
C14118 a_526_44458.t24 VSS 0.010884f
C14119 a_526_44458.n32 VSS 0.041036f
C14120 a_526_44458.n33 VSS 0.357664f
C14121 a_526_44458.n34 VSS 0.049714f
C14122 a_526_44458.n35 VSS 0.021559f
C14123 a_526_44458.t3 VSS 0.01078f
C14124 a_12861_44030.t26 VSS 0.014867f
C14125 a_12861_44030.n0 VSS 0.043853f
C14126 a_12861_44030.n1 VSS 0.032523f
C14127 a_12861_44030.n2 VSS 0.336865f
C14128 a_12861_44030.n3 VSS 0.021252f
C14129 a_12861_44030.n4 VSS 0.445109f
C14130 a_12861_44030.t29 VSS 0.013887f
C14131 a_12861_44030.n5 VSS 0.016208f
C14132 a_12861_44030.t13 VSS 0.013887f
C14133 a_12861_44030.t25 VSS 0.013887f
C14134 a_12861_44030.n7 VSS 0.0233f
C14135 a_12861_44030.n8 VSS 0.03769f
C14136 a_12861_44030.t21 VSS 0.013887f
C14137 a_12861_44030.n9 VSS 0.029835f
C14138 a_12861_44030.n10 VSS 0.022945f
C14139 a_12861_44030.n11 VSS 0.028125f
C14140 a_12861_44030.t32 VSS 0.011805f
C14141 a_12861_44030.n12 VSS 0.035913f
C14142 a_12861_44030.t31 VSS 0.011805f
C14143 a_12861_44030.n13 VSS 0.035402f
C14144 a_12861_44030.n14 VSS 0.025916f
C14145 a_12861_44030.n15 VSS 0.305785f
C14146 a_12861_44030.n16 VSS 0.222375f
C14147 a_12861_44030.t33 VSS 0.015044f
C14148 a_12861_44030.n17 VSS 0.02274f
C14149 a_12861_44030.n18 VSS 0.192093f
C14150 a_12861_44030.t11 VSS 0.010229f
C14151 a_12861_44030.n19 VSS 0.097331f
C14152 a_12861_44030.n20 VSS 0.542661f
C14153 a_12861_44030.t35 VSS 0.013887f
C14154 a_12861_44030.t14 VSS 0.013887f
C14155 a_12861_44030.n21 VSS 0.0233f
C14156 a_12861_44030.n22 VSS 0.035117f
C14157 a_12861_44030.n23 VSS 0.134726f
C14158 a_12861_44030.n24 VSS 0.089838f
C14159 a_12861_44030.n25 VSS 0.210602f
C14160 a_12861_44030.n26 VSS 0.018515f
C14161 a_12861_44030.n27 VSS 0.044715f
C14162 a_12861_44030.n28 VSS 0.013768f
C14163 a_12861_44030.n30 VSS 0.083066f
C14164 a_12861_44030.n31 VSS 0.056994f
C14165 a_12861_44030.n32 VSS 0.018953f
C14166 a_3080_42308.t0 VSS 0.047281f
C14167 a_3080_42308.t5 VSS 0.073549f
C14168 a_3080_42308.t4 VSS 0.04587f
C14169 a_3080_42308.n0 VSS 0.212734f
C14170 a_3080_42308.t6 VSS 0.315812f
C14171 a_3080_42308.t7 VSS 0.308951f
C14172 a_3080_42308.n1 VSS 13.4591f
C14173 a_3080_42308.n2 VSS 8.08834f
C14174 a_3080_42308.t3 VSS 0.030732f
C14175 a_3080_42308.t2 VSS 0.030732f
C14176 a_3080_42308.n3 VSS 0.061465f
C14177 a_3080_42308.n4 VSS 0.436325f
C14178 a_3080_42308.n5 VSS 0.141874f
C14179 a_3080_42308.t1 VSS 0.047281f
C14180 CAL_N.n0 VSS 2.19473f
C14181 CAL_N.t5 VSS 6.07059f
C14182 CAL_N.n1 VSS 4.24689f
C14183 CAL_N.t3 VSS 5.40859f
C14184 CAL_N.n2 VSS 4.24598f
C14185 CAL_N.t6 VSS 6.05896f
C14186 CAL_N.n3 VSS 2.12538f
C14187 CAL_N.n4 VSS 0.2083f
C14188 CAL_N.t1 VSS 0.01784f
C14189 CAL_N.n6 VSS 0.409935f
C14190 CAL_N.n7 VSS 0.414784f
C14191 CAL_N.t4 VSS 0.120027f
C14192 a_2324_44458.t1 VSS 0.011277f
C14193 a_2324_44458.n0 VSS 0.016818f
C14194 a_2324_44458.n1 VSS 0.010812f
C14195 a_2324_44458.n2 VSS 0.068318f
C14196 a_2324_44458.n3 VSS 0.010812f
C14197 a_2324_44458.n4 VSS 0.041064f
C14198 a_2324_44458.n5 VSS 0.010818f
C14199 a_2324_44458.n6 VSS 0.042359f
C14200 a_2324_44458.n7 VSS 0.010812f
C14201 a_2324_44458.n8 VSS 0.041064f
C14202 a_2324_44458.t61 VSS 0.015888f
C14203 a_2324_44458.t45 VSS 0.015888f
C14204 a_2324_44458.t41 VSS 0.015888f
C14205 a_2324_44458.t59 VSS 0.015888f
C14206 a_2324_44458.n10 VSS 0.03627f
C14207 a_2324_44458.n11 VSS 0.047773f
C14208 a_2324_44458.n12 VSS 0.047773f
C14209 a_2324_44458.n13 VSS 0.063696f
C14210 a_2324_44458.t50 VSS 0.015888f
C14211 a_2324_44458.t40 VSS 0.015888f
C14212 a_2324_44458.t63 VSS 0.015888f
C14213 a_2324_44458.t35 VSS 0.015888f
C14214 a_2324_44458.n14 VSS 0.03627f
C14215 a_2324_44458.n15 VSS 0.047773f
C14216 a_2324_44458.n16 VSS 0.047773f
C14217 a_2324_44458.n17 VSS 0.06491f
C14218 a_2324_44458.n18 VSS 0.921909f
C14219 a_2324_44458.t55 VSS 0.015888f
C14220 a_2324_44458.t57 VSS 0.015888f
C14221 a_2324_44458.t62 VSS 0.015888f
C14222 a_2324_44458.t43 VSS 0.015888f
C14223 a_2324_44458.n19 VSS 0.03627f
C14224 a_2324_44458.n20 VSS 0.047773f
C14225 a_2324_44458.n21 VSS 0.047773f
C14226 a_2324_44458.n22 VSS 0.08003f
C14227 a_2324_44458.t34 VSS 0.015888f
C14228 a_2324_44458.t48 VSS 0.015888f
C14229 a_2324_44458.t39 VSS 0.015888f
C14230 a_2324_44458.t49 VSS 0.015888f
C14231 a_2324_44458.n23 VSS 0.03627f
C14232 a_2324_44458.n24 VSS 0.047773f
C14233 a_2324_44458.n25 VSS 0.047773f
C14234 a_2324_44458.n26 VSS 0.059667f
C14235 a_2324_44458.n27 VSS 0.651008f
C14236 a_2324_44458.n28 VSS 1.19234f
C14237 a_2324_44458.n29 VSS 0.015985f
C14238 a_2324_44458.n30 VSS 0.026484f
C14239 a_2324_44458.n31 VSS 0.010812f
C14240 a_2324_44458.n32 VSS 0.03545f
C14241 a_2324_44458.n33 VSS 0.010524f
C14242 a_2324_44458.n34 VSS 0.110482f
C14243 a_2324_44458.t10 VSS 0.011277f
C14244 a_2324_44458.t3 VSS 0.011277f
C14245 a_2324_44458.n35 VSS 0.023451f
C14246 a_2324_44458.n36 VSS 0.131814f
C14247 a_2324_44458.t2 VSS 0.011277f
C14248 a_2324_44458.t9 VSS 0.011277f
C14249 a_2324_44458.n37 VSS 0.02377f
C14250 a_2324_44458.n38 VSS 0.053776f
C14251 a_2324_44458.t5 VSS 0.011277f
C14252 a_2324_44458.t0 VSS 0.011277f
C14253 a_2324_44458.n39 VSS 0.02377f
C14254 a_2324_44458.n40 VSS 0.0624f
C14255 a_2324_44458.t4 VSS 0.011277f
C14256 a_2324_44458.t13 VSS 0.011277f
C14257 a_2324_44458.n41 VSS 0.028646f
C14258 a_2324_44458.t14 VSS 0.011277f
C14259 a_2324_44458.t12 VSS 0.011277f
C14260 a_2324_44458.n42 VSS 0.02377f
C14261 a_2324_44458.n43 VSS 0.108325f
C14262 a_2324_44458.t7 VSS 0.011277f
C14263 a_2324_44458.t6 VSS 0.011277f
C14264 a_2324_44458.n44 VSS 0.02377f
C14265 a_2324_44458.n45 VSS 0.0624f
C14266 a_2324_44458.t8 VSS 0.011277f
C14267 a_2324_44458.t11 VSS 0.011277f
C14268 a_2324_44458.n46 VSS 0.02377f
C14269 a_2324_44458.n47 VSS 0.06211f
C14270 a_2324_44458.n48 VSS 0.06211f
C14271 a_2324_44458.n49 VSS 0.02377f
C14272 a_2324_44458.t15 VSS 0.011277f
C14273 VDD.t3645 VSS 0.016552f
C14274 VDD.n5 VSS 0.428084f
C14275 VDD.t3824 VSS 0.196177f
C14276 VDD.n6 VSS 0.074208f
C14277 VDD.t3805 VSS 0.196175f
C14278 VDD.n7 VSS 0.073454f
C14279 VDD.n8 VSS 0.082501f
C14280 VDD.t3783 VSS 0.197136f
C14281 VDD.n9 VSS 0.192011f
C14282 VDD.n10 VSS 0.21833f
C14283 VDD.n11 VSS 0.50592f
C14284 VDD.n12 VSS 0.19641f
C14285 VDD.n13 VSS 0.180192f
C14286 VDD.n14 VSS 0.171526f
C14287 VDD.n15 VSS 0.171526f
C14288 VDD.n16 VSS 0.20197f
C14289 VDD.n17 VSS 0.225568f
C14290 VDD.n18 VSS 0.525294f
C14291 VDD.t2955 VSS 0.592128f
C14292 VDD.t3761 VSS 0.640657f
C14293 VDD.t3766 VSS 0.640657f
C14294 VDD.t3096 VSS 0.640657f
C14295 VDD.t3231 VSS 0.640657f
C14296 VDD.t2921 VSS 0.644628f
C14297 VDD.t3604 VSS 0.493729f
C14298 VDD.t1972 VSS 0.33886f
C14299 VDD.t1969 VSS 0.33886f
C14300 VDD.t3609 VSS 0.33886f
C14301 VDD.t3613 VSS 0.33886f
C14302 VDD.t3610 VSS 0.33886f
C14303 VDD.t3614 VSS 0.33886f
C14304 VDD.t3072 VSS 0.33886f
C14305 VDD.t3079 VSS 0.33886f
C14306 VDD.t3073 VSS 0.199874f
C14307 VDD.n19 VSS 0.070155f
C14308 VDD.n20 VSS 0.138985f
C14309 VDD.t3080 VSS 0.268705f
C14310 VDD.t3075 VSS 0.33886f
C14311 VDD.t3076 VSS 0.33886f
C14312 VDD.t3078 VSS 0.33886f
C14313 VDD.t3074 VSS 0.33886f
C14314 VDD.t2072 VSS 0.33886f
C14315 VDD.t2073 VSS 0.33886f
C14316 VDD.t2074 VSS 0.33886f
C14317 VDD.t2069 VSS 0.33886f
C14318 VDD.t2084 VSS 0.33886f
C14319 VDD.t2071 VSS 0.33886f
C14320 VDD.t2085 VSS 0.33886f
C14321 VDD.t2081 VSS 0.33886f
C14322 VDD.t2075 VSS 0.33886f
C14323 VDD.t2083 VSS 0.33886f
C14324 VDD.t2077 VSS 0.33886f
C14325 VDD.t2070 VSS 0.33886f
C14326 VDD.t2076 VSS 0.33886f
C14327 VDD.t2082 VSS 0.33886f
C14328 VDD.t2080 VSS 0.33886f
C14329 VDD.t2068 VSS 0.434851f
C14330 VDD.n21 VSS 0.518436f
C14331 VDD.n22 VSS 0.196597f
C14332 VDD.n23 VSS 0.193559f
C14333 VDD.n24 VSS 0.175072f
C14334 VDD.n25 VSS 0.486357f
C14335 VDD.n26 VSS 0.391578f
C14336 VDD.t2195 VSS 0.10507f
C14337 VDD.t3059 VSS 0.031978f
C14338 VDD.t2193 VSS 0.031978f
C14339 VDD.t3066 VSS 0.035023f
C14340 VDD.t3055 VSS 0.063956f
C14341 VDD.t3057 VSS 0.041114f
C14342 VDD.t2409 VSS 0.041114f
C14343 VDD.t2405 VSS 0.063956f
C14344 VDD.t2403 VSS 0.04987f
C14345 VDD.t2407 VSS 0.173303f
C14346 VDD.n28 VSS 0.017977f
C14347 VDD.t2408 VSS 0.01271f
C14348 VDD.n29 VSS 0.037969f
C14349 VDD.t2194 VSS 0.01447f
C14350 VDD.t2196 VSS 0.014207f
C14351 VDD.t3060 VSS 0.012671f
C14352 VDD.n33 VSS 0.014179f
C14353 VDD.n34 VSS 0.023611f
C14354 VDD.n35 VSS 0.011881f
C14355 VDD.n37 VSS 0.023783f
C14356 VDD.t2410 VSS 0.014487f
C14357 VDD.n38 VSS 0.020035f
C14358 VDD.t3058 VSS 0.014487f
C14359 VDD.n41 VSS 0.020424f
C14360 VDD.n42 VSS 0.043128f
C14361 VDD.n43 VSS 0.058405f
C14362 VDD.n44 VSS 1.09625f
C14363 VDD.n45 VSS 1.44135f
C14364 VDD.n46 VSS 0.486367f
C14365 VDD.n47 VSS 0.50592f
C14366 VDD.n48 VSS 0.175072f
C14367 VDD.n49 VSS 0.180192f
C14368 VDD.n50 VSS 0.171526f
C14369 VDD.n51 VSS 0.171526f
C14370 VDD.n52 VSS 0.196417f
C14371 VDD.n53 VSS 0.201985f
C14372 VDD.n54 VSS 0.225547f
C14373 VDD.n55 VSS 0.525294f
C14374 VDD.t3547 VSS 0.592128f
C14375 VDD.t3663 VSS 0.640657f
C14376 VDD.t3702 VSS 0.640657f
C14377 VDD.t2033 VSS 0.640657f
C14378 VDD.t2893 VSS 0.640657f
C14379 VDD.t2102 VSS 0.644628f
C14380 VDD.t2001 VSS 0.493729f
C14381 VDD.t1963 VSS 0.33886f
C14382 VDD.t1964 VSS 0.33886f
C14383 VDD.t3555 VSS 0.33886f
C14384 VDD.t3554 VSS 0.33886f
C14385 VDD.t3556 VSS 0.33886f
C14386 VDD.t3557 VSS 0.33886f
C14387 VDD.t1777 VSS 0.33886f
C14388 VDD.t1773 VSS 0.33886f
C14389 VDD.t1780 VSS 0.199874f
C14390 VDD.n56 VSS 0.070155f
C14391 VDD.n57 VSS 0.138985f
C14392 VDD.t1776 VSS 0.268705f
C14393 VDD.t1778 VSS 0.33886f
C14394 VDD.t1779 VSS 0.33886f
C14395 VDD.t1774 VSS 0.33886f
C14396 VDD.t1775 VSS 0.33886f
C14397 VDD.t1945 VSS 0.33886f
C14398 VDD.t1943 VSS 0.33886f
C14399 VDD.t1951 VSS 0.33886f
C14400 VDD.t1949 VSS 0.33886f
C14401 VDD.t1939 VSS 0.33886f
C14402 VDD.t1946 VSS 0.33886f
C14403 VDD.t1952 VSS 0.33886f
C14404 VDD.t1942 VSS 0.33886f
C14405 VDD.t1950 VSS 0.33886f
C14406 VDD.t1954 VSS 0.33886f
C14407 VDD.t1947 VSS 0.33886f
C14408 VDD.t1944 VSS 0.33886f
C14409 VDD.t1948 VSS 0.33886f
C14410 VDD.t1953 VSS 0.33886f
C14411 VDD.t1940 VSS 0.33886f
C14412 VDD.t1941 VSS 0.434851f
C14413 VDD.n58 VSS 0.518436f
C14414 VDD.n59 VSS 0.196597f
C14415 VDD.n60 VSS 0.193559f
C14416 VDD.n61 VSS 0.218326f
C14417 VDD.n62 VSS 0.391572f
C14418 VDD.n63 VSS 0.043193f
C14419 VDD.n64 VSS 0.011881f
C14420 VDD.t1658 VSS 0.173303f
C14421 VDD.t1656 VSS 0.10507f
C14422 VDD.t3070 VSS 0.031978f
C14423 VDD.t1654 VSS 0.031978f
C14424 VDD.t3064 VSS 0.035023f
C14425 VDD.t3068 VSS 0.063956f
C14426 VDD.t3061 VSS 0.041114f
C14427 VDD.t1660 VSS 0.041114f
C14428 VDD.t1662 VSS 0.063956f
C14429 VDD.t1664 VSS 0.04987f
C14430 VDD.n66 VSS 0.017977f
C14431 VDD.t1659 VSS 0.01271f
C14432 VDD.n67 VSS 0.037968f
C14433 VDD.t3062 VSS 0.014487f
C14434 VDD.n70 VSS 0.020424f
C14435 VDD.t1661 VSS 0.014487f
C14436 VDD.t1655 VSS 0.01447f
C14437 VDD.t3071 VSS 0.012671f
C14438 VDD.t1657 VSS 0.014207f
C14439 VDD.n73 VSS 0.014179f
C14440 VDD.n74 VSS 0.023611f
C14441 VDD.n76 VSS 0.023783f
C14442 VDD.n77 VSS 0.020035f
C14443 VDD.n79 VSS 0.058374f
C14444 VDD.n80 VSS 1.13691f
C14445 VDD.t3785 VSS 0.197137f
C14446 VDD.n81 VSS 0.431813f
C14447 VDD.t3133 VSS 0.01655f
C14448 VDD.n82 VSS 0.427848f
C14449 VDD.t3825 VSS 0.196175f
C14450 VDD.t3786 VSS 0.196177f
C14451 VDD.n83 VSS 0.074082f
C14452 VDD.n84 VSS 0.07358f
C14453 VDD.n85 VSS 0.054535f
C14454 VDD.n86 VSS 2.42454f
C14455 VDD.n87 VSS 0.354856f
C14456 VDD.t3434 VSS 0.143093f
C14457 VDD.n88 VSS 0.499455f
C14458 VDD.n89 VSS 0.372351f
C14459 VDD.n90 VSS 0.375148f
C14460 VDD.n91 VSS 0.342447f
C14461 VDD.n92 VSS 0.08955f
C14462 VDD.n93 VSS 0.103727f
C14463 VDD.n94 VSS 0.12653f
C14464 VDD.t1755 VSS 10.2697f
C14465 VDD.t1758 VSS 10.2697f
C14466 VDD.n95 VSS 0.199365f
C14467 VDD.n96 VSS 0.126325f
C14468 VDD.n97 VSS 0.126325f
C14469 VDD.n98 VSS 4.00715f
C14470 VDD.n99 VSS 0.126325f
C14471 VDD.n100 VSS 0.050115f
C14472 VDD.n101 VSS 0.018273f
C14473 VDD.n102 VSS 0.013607f
C14474 VDD.n103 VSS 0.014158f
C14475 VDD.n104 VSS 0.197231f
C14476 VDD.n105 VSS 0.677889f
C14477 VDD.n106 VSS 0.129852f
C14478 VDD.n107 VSS 0.0141f
C14479 VDD.n108 VSS 0.025952f
C14480 VDD.t660 VSS 0.081848f
C14481 VDD.t935 VSS 0.090849f
C14482 VDD.n109 VSS 0.013607f
C14483 VDD.n110 VSS 0.018273f
C14484 VDD.n111 VSS 0.016511f
C14485 VDD.n112 VSS 0.016212f
C14486 VDD.n113 VSS 0.016511f
C14487 VDD.n114 VSS 0.018273f
C14488 VDD.n115 VSS 0.016212f
C14489 VDD.n116 VSS 0.016212f
C14490 VDD.t2391 VSS 0.162771f
C14491 VDD.n117 VSS 0.16908f
C14492 VDD.n118 VSS 0.016212f
C14493 VDD.n119 VSS 0.036827f
C14494 VDD.n120 VSS 0.025883f
C14495 VDD.n121 VSS 0.018273f
C14496 VDD.n122 VSS 0.060566f
C14497 VDD.t3480 VSS 0.090849f
C14498 VDD.t1242 VSS 0.141952f
C14499 VDD.t1612 VSS 0.01449f
C14500 VDD.t1611 VSS 0.01449f
C14501 VDD.n123 VSS 0.038176f
C14502 VDD.n124 VSS 0.011881f
C14503 VDD.t1938 VSS 0.014485f
C14504 VDD.t2638 VSS 0.014485f
C14505 VDD.t2390 VSS 0.01447f
C14506 VDD.t937 VSS 0.01447f
C14507 VDD.n125 VSS 0.029398f
C14508 VDD.n126 VSS 0.928837f
C14509 VDD.t3433 VSS 0.039011f
C14510 VDD.n127 VSS 0.928837f
C14511 VDD.n128 VSS 0.079563f
C14512 VDD.t3430 VSS 0.078021f
C14513 VDD.n129 VSS 0.079563f
C14514 VDD.t3432 VSS 0.182104f
C14515 VDD.n130 VSS 0.497625f
C14516 VDD.n131 VSS 0.011881f
C14517 VDD.t2283 VSS 0.014453f
C14518 VDD.t3481 VSS 0.089462f
C14519 VDD.t1245 VSS 0.102786f
C14520 VDD.t1608 VSS 0.036546f
C14521 VDD.t662 VSS 0.052916f
C14522 VDD.t2282 VSS 0.114684f
C14523 VDD.n133 VSS 0.063478f
C14524 VDD.t1609 VSS 0.01447f
C14525 VDD.n135 VSS 0.015032f
C14526 VDD.n136 VSS 0.013517f
C14527 VDD.n138 VSS 0.039405f
C14528 VDD.n139 VSS 0.011881f
C14529 VDD.t3482 VSS 0.01447f
C14530 VDD.n141 VSS 0.015466f
C14531 VDD.t661 VSS 0.01447f
C14532 VDD.n143 VSS 0.016845f
C14533 VDD.n144 VSS 0.0184f
C14534 VDD.n145 VSS 0.928837f
C14535 VDD.t1759 VSS 0.039011f
C14536 VDD.t1760 VSS 0.143093f
C14537 VDD.n146 VSS 0.499455f
C14538 VDD.n147 VSS 0.928837f
C14539 VDD.n148 VSS 0.079563f
C14540 VDD.t1754 VSS 0.078021f
C14541 VDD.n149 VSS 0.079563f
C14542 VDD.t1756 VSS 0.182104f
C14543 VDD.n150 VSS 0.542117f
C14544 VDD.n151 VSS 0.044737f
C14545 VDD.n152 VSS 0.069654f
C14546 VDD.n153 VSS 0.036362f
C14547 VDD.n154 VSS 0.065816f
C14548 VDD.n155 VSS 0.057906f
C14549 VDD.n156 VSS 0.059902f
C14550 VDD.n157 VSS 0.214683f
C14551 VDD.n158 VSS 0.026743f
C14552 VDD.n159 VSS 0.01368f
C14553 VDD.n161 VSS 0.036303f
C14554 VDD.n163 VSS 0.034516f
C14555 VDD.n164 VSS 0.13311f
C14556 VDD.t1610 VSS 0.128608f
C14557 VDD.t1937 VSS 0.119156f
C14558 VDD.t936 VSS 0.169026f
C14559 VDD.n165 VSS 0.412837f
C14560 VDD.n166 VSS 3.83711f
C14561 VDD.n167 VSS 0.10359f
C14562 VDD.n168 VSS 0.021792f
C14563 VDD.n169 VSS 0.054857f
C14564 VDD.n170 VSS 0.014951f
C14565 VDD.n171 VSS 0.016177f
C14566 VDD.n172 VSS 0.023992f
C14567 VDD.n173 VSS 0.237196f
C14568 VDD.n174 VSS 0.228732f
C14569 VDD.n175 VSS 0.295297f
C14570 VDD.n176 VSS 0.199365f
C14571 VDD.t1753 VSS 13.205299f
C14572 VDD.n177 VSS 0.146403f
C14573 VDD.n178 VSS 0.144756f
C14574 VDD.n179 VSS 0.15156f
C14575 VDD.n180 VSS 0.078425f
C14576 VDD.n181 VSS 0.141245f
C14577 VDD.n182 VSS 0.273443f
C14578 VDD.n183 VSS 0.365097f
C14579 VDD.n184 VSS 5.69147f
C14580 VDD.t3594 VSS 0.121419f
C14581 VDD.t3593 VSS 0.123336f
C14582 VDD.n185 VSS 0.314863f
C14583 VDD.t3596 VSS 0.1217f
C14584 VDD.t3597 VSS 0.123641f
C14585 VDD.n186 VSS 0.307912f
C14586 VDD.n187 VSS 0.363667f
C14587 VDD.n188 VSS 0.480693f
C14588 VDD.n189 VSS 0.118319f
C14589 VDD.n190 VSS 0.094333f
C14590 VDD.n191 VSS 0.076651f
C14591 VDD.n192 VSS 0.094333f
C14592 VDD.t3592 VSS 0.634898f
C14593 VDD.t1766 VSS 0.158444f
C14594 VDD.n193 VSS 0.094913f
C14595 VDD.t3590 VSS 0.742762f
C14596 VDD.n194 VSS 0.017014f
C14597 VDD.n195 VSS 0.068655f
C14598 VDD.n196 VSS 0.106529f
C14599 VDD.n197 VSS 0.053888f
C14600 VDD.n198 VSS 0.016867f
C14601 VDD.n199 VSS 0.027369f
C14602 VDD.n200 VSS 0.046194f
C14603 VDD.t1757 VSS 0.124783f
C14604 VDD.n201 VSS 0.118049f
C14605 VDD.n202 VSS 0.027369f
C14606 VDD.t3431 VSS 0.124783f
C14607 VDD.n203 VSS 0.118049f
C14608 VDD.n204 VSS 0.018788f
C14609 VDD.n205 VSS 0.046194f
C14610 VDD.n206 VSS 0.01675f
C14611 VDD.n207 VSS 0.048937f
C14612 VDD.t1767 VSS 0.014204f
C14613 VDD.n208 VSS 0.042946f
C14614 VDD.n209 VSS 0.29422f
C14615 VDD.n210 VSS 0.127167f
C14616 VDD.n211 VSS 0.038914f
C14617 VDD.n212 VSS 0.048266f
C14618 VDD.n213 VSS 0.082908f
C14619 VDD.n214 VSS 0.036993f
C14620 VDD.n215 VSS 0.037918f
C14621 VDD.n216 VSS 0.038242f
C14622 VDD.n217 VSS 0.03632f
C14623 VDD.n218 VSS 0.038591f
C14624 VDD.n219 VSS 0.038914f
C14625 VDD.n220 VSS 0.03632f
C14626 VDD.n221 VSS 0.037918f
C14627 VDD.t3589 VSS 0.114531f
C14628 VDD.n222 VSS 0.10977f
C14629 VDD.n223 VSS 0.075189f
C14630 VDD.n224 VSS 0.015962f
C14631 VDD.n225 VSS 0.029939f
C14632 VDD.n226 VSS 0.021976f
C14633 VDD.n227 VSS 0.164845f
C14634 VDD.t143 VSS 0.081164f
C14635 VDD.n228 VSS 0.021976f
C14636 VDD.n229 VSS 0.029982f
C14637 VDD.n230 VSS 0.164845f
C14638 VDD.t185 VSS 0.162311f
C14639 VDD.t230 VSS 0.081164f
C14640 VDD.t224 VSS 0.145418f
C14641 VDD.n231 VSS 0.015962f
C14642 VDD.n232 VSS 0.182618f
C14643 VDD.t196 VSS 0.145418f
C14644 VDD.t150 VSS 0.081164f
C14645 VDD.n233 VSS 0.022391f
C14646 VDD.n234 VSS 0.054109f
C14647 VDD.n235 VSS 0.022391f
C14648 VDD.n236 VSS 0.022391f
C14649 VDD.n237 VSS 0.021976f
C14650 VDD.n238 VSS 0.022392f
C14651 VDD.n239 VSS 0.022391f
C14652 VDD.t133 VSS 0.162311f
C14653 VDD.t97 VSS 0.081164f
C14654 VDD.n240 VSS 0.054109f
C14655 VDD.n241 VSS 0.022391f
C14656 VDD.n242 VSS 0.075888f
C14657 VDD.n243 VSS 0.033567f
C14658 VDD.n244 VSS 0.355421f
C14659 VDD.n245 VSS 0.010237f
C14660 VDD.n246 VSS 0.623036f
C14661 VDD.n247 VSS 0.278708f
C14662 VDD.n248 VSS 0.027576f
C14663 VDD.n249 VSS 0.059971f
C14664 VDD.n250 VSS 0.025802f
C14665 VDD.t3599 VSS 0.114531f
C14666 VDD.n251 VSS 0.108302f
C14667 VDD.n252 VSS 0.064118f
C14668 VDD.n253 VSS 0.038242f
C14669 VDD.t3579 VSS 0.114531f
C14670 VDD.n254 VSS 0.108302f
C14671 VDD.n255 VSS 0.025802f
C14672 VDD.n256 VSS 0.037918f
C14673 VDD.n257 VSS 0.038591f
C14674 VDD.t3601 VSS 0.114531f
C14675 VDD.n258 VSS 0.108302f
C14676 VDD.n259 VSS 0.025802f
C14677 VDD.n260 VSS 0.036993f
C14678 VDD.n261 VSS 0.036993f
C14679 VDD.n262 VSS 0.025802f
C14680 VDD.t3587 VSS 0.114531f
C14681 VDD.n263 VSS 0.108302f
C14682 VDD.n264 VSS 0.038914f
C14683 VDD.n265 VSS 0.038242f
C14684 VDD.t3577 VSS 0.114531f
C14685 VDD.n266 VSS 0.108302f
C14686 VDD.n267 VSS 0.025802f
C14687 VDD.n268 VSS 0.037918f
C14688 VDD.n269 VSS 0.037918f
C14689 VDD.t3591 VSS 0.114531f
C14690 VDD.n270 VSS 0.108302f
C14691 VDD.n271 VSS 0.025802f
C14692 VDD.n272 VSS 0.03632f
C14693 VDD.n273 VSS 0.03632f
C14694 VDD.n274 VSS 0.025802f
C14695 VDD.t3603 VSS 0.114531f
C14696 VDD.n275 VSS 0.108302f
C14697 VDD.n276 VSS 0.038242f
C14698 VDD.n277 VSS 0.038914f
C14699 VDD.t3581 VSS 0.114531f
C14700 VDD.n278 VSS 0.108302f
C14701 VDD.n279 VSS 0.025802f
C14702 VDD.n280 VSS 0.038591f
C14703 VDD.n281 VSS 0.038591f
C14704 VDD.t3585 VSS 0.114531f
C14705 VDD.n282 VSS 0.108302f
C14706 VDD.n283 VSS 0.025802f
C14707 VDD.n284 VSS 0.036993f
C14708 VDD.n285 VSS 0.080834f
C14709 VDD.n286 VSS 0.025802f
C14710 VDD.t3583 VSS 0.114531f
C14711 VDD.n287 VSS 0.108302f
C14712 VDD.n288 VSS -0.022025f
C14713 VDD.n289 VSS 0.085007f
C14714 VDD.n290 VSS 0.053337f
C14715 VDD.n291 VSS 0.099137f
C14716 VDD.n292 VSS 0.296814f
C14717 VDD.t3602 VSS 0.742762f
C14718 VDD.t3580 VSS 0.742762f
C14719 VDD.t3584 VSS 0.742762f
C14720 VDD.t3582 VSS 0.742762f
C14721 VDD.t3595 VSS 0.664711f
C14722 VDD.n293 VSS 0.494814f
C14723 VDD.n294 VSS 0.105003f
C14724 VDD.t3576 VSS 0.742762f
C14725 VDD.t3586 VSS 0.742762f
C14726 VDD.t3600 VSS 0.742762f
C14727 VDD.t3578 VSS 0.637629f
C14728 VDD.t3588 VSS 0.742762f
C14729 VDD.t3598 VSS 0.476515f
C14730 VDD.n295 VSS 0.382761f
C14731 VDD.n296 VSS 0.067469f
C14732 VDD.t63 VSS 0.304195f
C14733 VDD.n297 VSS 0.397216f
C14734 VDD.n298 VSS 0.090637f
C14735 VDD.n299 VSS 0.118436f
C14736 VDD.t59 VSS 0.405242f
C14737 VDD.t60 VSS 0.405242f
C14738 VDD.t71 VSS 0.654091f
C14739 VDD.n300 VSS 0.114991f
C14740 VDD.t67 VSS 0.654091f
C14741 VDD.t61 VSS 0.405242f
C14742 VDD.t57 VSS 0.405242f
C14743 VDD.t70 VSS 0.304195f
C14744 VDD.n301 VSS 0.067469f
C14745 VDD.t1770 VSS 0.135746f
C14746 VDD.n302 VSS 0.017909f
C14747 VDD.n303 VSS 0.017909f
C14748 VDD.n304 VSS 0.151984f
C14749 VDD.n305 VSS 0.067096f
C14750 VDD.n306 VSS 0.05669f
C14751 VDD.n307 VSS 0.046944f
C14752 VDD.n308 VSS 0.047762f
C14753 VDD.n309 VSS 0.05669f
C14754 VDD.n310 VSS 0.058087f
C14755 VDD.n311 VSS 0.057269f
C14756 VDD.n312 VSS 0.078866f
C14757 VDD.n313 VSS 0.104507f
C14758 VDD.n314 VSS 0.03484f
C14759 VDD.n315 VSS 0.057233f
C14760 VDD.n317 VSS 0.103509f
C14761 VDD.n318 VSS 0.01682f
C14762 VDD.n319 VSS 0.017908f
C14763 VDD.n320 VSS 0.013731f
C14764 VDD.n321 VSS 0.017674f
C14765 VDD.n322 VSS 0.100857f
C14766 VDD.n323 VSS 0.367285f
C14767 VDD.t72 VSS 0.728523f
C14768 VDD.t68 VSS 0.405242f
C14769 VDD.t64 VSS 0.405242f
C14770 VDD.t66 VSS 0.304195f
C14771 VDD.n324 VSS 0.133806f
C14772 VDD.n325 VSS 0.057269f
C14773 VDD.n326 VSS 0.05669f
C14774 VDD.n327 VSS 0.022708f
C14775 VDD.n328 VSS 0.133806f
C14776 VDD.t62 VSS 0.304195f
C14777 VDD.t65 VSS 0.405242f
C14778 VDD.t58 VSS 0.405242f
C14779 VDD.t69 VSS 0.728714f
C14780 VDD.n329 VSS 0.483342f
C14781 VDD.n330 VSS 0.04678f
C14782 VDD.n331 VSS 0.046369f
C14783 VDD.n332 VSS 0.159438f
C14784 VDD.n333 VSS 0.213466f
C14785 VDD.n334 VSS 0.447284f
C14786 VDD.n335 VSS 0.225343f
C14787 VDD.t1771 VSS 0.01492f
C14788 VDD.n336 VSS 0.630786f
C14789 VDD.n337 VSS 3.64102f
C14790 VDD.n338 VSS 0.039106f
C14791 VDD.n339 VSS 0.025742f
C14792 VDD.n340 VSS 0.043261f
C14793 VDD.t1208 VSS 0.014212f
C14794 VDD.t2050 VSS 0.021512f
C14795 VDD.n341 VSS 0.029887f
C14796 VDD.n342 VSS 0.037647f
C14797 VDD.t354 VSS 0.014212f
C14798 VDD.n348 VSS 0.018136f
C14799 VDD.n349 VSS 0.036868f
C14800 VDD.t2683 VSS 0.014237f
C14801 VDD.t2947 VSS 0.014748f
C14802 VDD.n350 VSS 0.016089f
C14803 VDD.t1206 VSS 0.012671f
C14804 VDD.n353 VSS 0.074941f
C14805 VDD.t1205 VSS 0.082335f
C14806 VDD.t1203 VSS 0.036272f
C14807 VDD.t1209 VSS 0.036272f
C14808 VDD.t1207 VSS 0.071032f
C14809 VDD.t2049 VSS 0.097155f
C14810 VDD.t2054 VSS 0.263125f
C14811 VDD.n354 VSS 0.015303f
C14812 VDD.n355 VSS 0.013396f
C14813 VDD.n356 VSS 0.024773f
C14814 VDD.n358 VSS 0.015303f
C14815 VDD.n359 VSS 0.036161f
C14816 VDD.n360 VSS 0.018615f
C14817 VDD.n361 VSS 0.018569f
C14818 VDD.n362 VSS 0.263125f
C14819 VDD.n364 VSS 0.019781f
C14820 VDD.n365 VSS 0.025109f
C14821 VDD.n366 VSS 0.016489f
C14822 VDD.n367 VSS 0.018615f
C14823 VDD.n368 VSS 0.263125f
C14824 VDD.n369 VSS 0.018615f
C14825 VDD.n370 VSS 0.025109f
C14826 VDD.n371 VSS 0.019781f
C14827 VDD.n372 VSS 0.035949f
C14828 VDD.n373 VSS 0.015303f
C14829 VDD.n374 VSS 0.015303f
C14830 VDD.n375 VSS 0.219826f
C14831 VDD.n376 VSS 0.035949f
C14832 VDD.n377 VSS 0.021679f
C14833 VDD.n378 VSS 0.024561f
C14834 VDD.n379 VSS 0.015303f
C14835 VDD.n380 VSS 0.021679f
C14836 VDD.n381 VSS 0.024561f
C14837 VDD.n382 VSS 0.015551f
C14838 VDD.n384 VSS 0.013396f
C14839 VDD.t2056 VSS 0.263125f
C14840 VDD.n385 VSS 0.013396f
C14841 VDD.n386 VSS 0.013396f
C14842 VDD.n387 VSS 0.018615f
C14843 VDD.n388 VSS 0.013396f
C14844 VDD.n389 VSS 0.013396f
C14845 VDD.n390 VSS 0.018615f
C14846 VDD.n392 VSS 0.019781f
C14847 VDD.t2051 VSS 0.263125f
C14848 VDD.n397 VSS 0.044122f
C14849 VDD.t2945 VSS 0.061587f
C14850 VDD.t2052 VSS 0.061449f
C14851 VDD.n398 VSS 0.154287f
C14852 VDD.t2057 VSS 0.015015f
C14853 VDD.t2059 VSS 0.014776f
C14854 VDD.n399 VSS 0.12372f
C14855 VDD.n400 VSS 0.100017f
C14856 VDD.n401 VSS 0.045199f
C14857 VDD.n402 VSS 0.018833f
C14858 VDD.n403 VSS 0.018564f
C14859 VDD.n404 VSS 0.146634f
C14860 VDD.n405 VSS 0.037288f
C14861 VDD.t2055 VSS 0.015015f
C14862 VDD.t2058 VSS 0.014776f
C14863 VDD.n406 VSS 0.1215f
C14864 VDD.n407 VSS 0.034552f
C14865 VDD.n408 VSS 0.027442f
C14866 VDD.n409 VSS 0.0862f
C14867 VDD.n410 VSS 0.214484f
C14868 VDD.n411 VSS 0.016444f
C14869 VDD.t2944 VSS 0.263125f
C14870 VDD.n414 VSS 0.263125f
C14871 VDD.n415 VSS 0.036161f
C14872 VDD.n416 VSS 0.022104f
C14873 VDD.n417 VSS 0.022104f
C14874 VDD.n418 VSS 0.024773f
C14875 VDD.n419 VSS 0.015505f
C14876 VDD.n420 VSS 0.015258f
C14877 VDD.n421 VSS 0.175694f
C14878 VDD.n422 VSS 0.140153f
C14879 VDD.t2946 VSS 0.075605f
C14880 VDD.t2636 VSS 0.104309f
C14881 VDD.t357 VSS 0.031978f
C14882 VDD.t2686 VSS 0.031978f
C14883 VDD.t351 VSS 0.031978f
C14884 VDD.t2680 VSS 0.031978f
C14885 VDD.t355 VSS 0.031978f
C14886 VDD.t2684 VSS 0.031978f
C14887 VDD.t353 VSS 0.031978f
C14888 VDD.t2682 VSS 0.092127f
C14889 VDD.n423 VSS 0.071297f
C14890 VDD.n424 VSS 0.023209f
C14891 VDD.n426 VSS 0.022277f
C14892 VDD.n428 VSS 0.011881f
C14893 VDD.n431 VSS 0.015751f
C14894 VDD.n432 VSS 0.010467f
C14895 VDD.n433 VSS 0.013318f
C14896 VDD.t358 VSS 0.012763f
C14897 VDD.n434 VSS 0.011218f
C14898 VDD.n435 VSS 0.026676f
C14899 VDD.n436 VSS 0.232236f
C14900 VDD.n437 VSS 0.221716f
C14901 VDD.n438 VSS 0.03292f
C14902 VDD.n439 VSS 0.019801f
C14903 VDD.n440 VSS 0.019801f
C14904 VDD.n441 VSS 0.019801f
C14905 VDD.n442 VSS 0.019446f
C14906 VDD.n443 VSS 0.067546f
C14907 VDD.n444 VSS 2.35832f
C14908 VDD.n446 VSS 0.011881f
C14909 VDD.t1616 VSS 0.014683f
C14910 VDD.t282 VSS 0.014683f
C14911 VDD.n449 VSS 0.017506f
C14912 VDD.n450 VSS 0.011881f
C14913 VDD.n451 VSS 0.010077f
C14914 VDD.n452 VSS 0.010077f
C14915 VDD.n453 VSS 0.015687f
C14916 VDD.n454 VSS 0.042008f
C14917 VDD.t705 VSS 0.014683f
C14918 VDD.t1151 VSS 0.014683f
C14919 VDD.n457 VSS 0.019839f
C14920 VDD.n459 VSS 0.012144f
C14921 VDD.n462 VSS 0.011881f
C14922 VDD.n463 VSS 0.011881f
C14923 VDD.n467 VSS 0.011881f
C14924 VDD.n468 VSS 0.011881f
C14925 VDD.n471 VSS 0.01031f
C14926 VDD.n472 VSS 0.010077f
C14927 VDD.n473 VSS 0.010077f
C14928 VDD.n475 VSS 0.011881f
C14929 VDD.t704 VSS 0.146946f
C14930 VDD.t702 VSS 0.063956f
C14931 VDD.t706 VSS 0.063956f
C14932 VDD.t708 VSS 0.070428f
C14933 VDD.t2027 VSS 0.065859f
C14934 VDD.t1761 VSS 0.110781f
C14935 VDD.t281 VSS 0.115349f
C14936 VDD.t283 VSS 0.063956f
C14937 VDD.t279 VSS 0.063956f
C14938 VDD.t285 VSS 0.070428f
C14939 VDD.t2887 VSS 0.065859f
C14940 VDD.t1772 VSS 0.085275f
C14941 VDD.t2043 VSS 0.134003f
C14942 VDD.t3094 VSS 0.071189f
C14943 VDD.t1707 VSS 0.071189f
C14944 VDD.t1709 VSS 0.065479f
C14945 VDD.t1705 VSS 0.065479f
C14946 VDD.t1711 VSS 0.108497f
C14947 VDD.t2025 VSS 0.108497f
C14948 VDD.t2956 VSS 0.071189f
C14949 VDD.t1379 VSS 0.071189f
C14950 VDD.t1377 VSS 0.065479f
C14951 VDD.t1383 VSS 0.065479f
C14952 VDD.t1381 VSS 0.089843f
C14953 VDD.n476 VSS 0.127365f
C14954 VDD.t1382 VSS 0.014787f
C14955 VDD.t2547 VSS 0.014787f
C14956 VDD.n478 VSS 0.011881f
C14957 VDD.n481 VSS 0.026075f
C14958 VDD.t2026 VSS 0.013864f
C14959 VDD.t2894 VSS 0.013864f
C14960 VDD.n484 VSS 0.029707f
C14961 VDD.n485 VSS 0.011881f
C14962 VDD.t2362 VSS 0.014787f
C14963 VDD.t1712 VSS 0.014787f
C14964 VDD.t2044 VSS 0.013864f
C14965 VDD.t3706 VSS 0.013864f
C14966 VDD.n487 VSS 0.032563f
C14967 VDD.n488 VSS 0.01221f
C14968 VDD.n491 VSS 0.026075f
C14969 VDD.n494 VSS 0.028639f
C14970 VDD.n496 VSS 0.038332f
C14971 VDD.n497 VSS 0.011881f
C14972 VDD.n498 VSS 0.011881f
C14973 VDD.n500 VSS 0.028059f
C14974 VDD.n503 VSS 0.011881f
C14975 VDD.n504 VSS 0.011881f
C14976 VDD.n507 VSS 0.026075f
C14977 VDD.n509 VSS 0.011881f
C14978 VDD.n510 VSS 0.011881f
C14979 VDD.n511 VSS 0.011881f
C14980 VDD.n513 VSS 0.028059f
C14981 VDD.n515 VSS 0.044176f
C14982 VDD.n516 VSS 0.011881f
C14983 VDD.n517 VSS 0.011881f
C14984 VDD.n518 VSS 0.011881f
C14985 VDD.n520 VSS 0.015687f
C14986 VDD.n523 VSS 0.010719f
C14987 VDD.n524 VSS 0.034682f
C14988 VDD.n526 VSS 0.011881f
C14989 VDD.t2160 VSS 0.014683f
C14990 VDD.t883 VSS 0.014683f
C14991 VDD.n529 VSS 0.017506f
C14992 VDD.n530 VSS 0.011881f
C14993 VDD.n531 VSS 0.010077f
C14994 VDD.n532 VSS 0.010077f
C14995 VDD.n533 VSS 0.015687f
C14996 VDD.n534 VSS 0.042008f
C14997 VDD.t404 VSS 0.014683f
C14998 VDD.t2649 VSS 0.014683f
C14999 VDD.n537 VSS 0.019839f
C15000 VDD.n539 VSS 0.012144f
C15001 VDD.n542 VSS 0.011881f
C15002 VDD.n543 VSS 0.011881f
C15003 VDD.n547 VSS 0.011881f
C15004 VDD.n548 VSS 0.011881f
C15005 VDD.n551 VSS 0.01031f
C15006 VDD.n552 VSS 0.010077f
C15007 VDD.n553 VSS 0.010077f
C15008 VDD.n555 VSS 0.011881f
C15009 VDD.t403 VSS 0.146946f
C15010 VDD.t401 VSS 0.063956f
C15011 VDD.t397 VSS 0.063956f
C15012 VDD.t399 VSS 0.070428f
C15013 VDD.t2036 VSS 0.065859f
C15014 VDD.t2877 VSS 0.110781f
C15015 VDD.t882 VSS 0.115349f
C15016 VDD.t878 VSS 0.063956f
C15017 VDD.t880 VSS 0.063956f
C15018 VDD.t884 VSS 0.070428f
C15019 VDD.t2023 VSS 0.065859f
C15020 VDD.t1962 VSS 0.085275f
C15021 VDD.t1983 VSS 0.134003f
C15022 VDD.t1970 VSS 0.071189f
C15023 VDD.t777 VSS 0.071189f
C15024 VDD.t783 VSS 0.065479f
C15025 VDD.t781 VSS 0.065479f
C15026 VDD.t779 VSS 0.108497f
C15027 VDD.t2889 VSS 0.108497f
C15028 VDD.t3228 VSS 0.071189f
C15029 VDD.t369 VSS 0.071189f
C15030 VDD.t363 VSS 0.065479f
C15031 VDD.t365 VSS 0.065479f
C15032 VDD.t367 VSS 0.089843f
C15033 VDD.n556 VSS 0.127365f
C15034 VDD.t368 VSS 0.014787f
C15035 VDD.t2521 VSS 0.014787f
C15036 VDD.n558 VSS 0.011881f
C15037 VDD.n561 VSS 0.026075f
C15038 VDD.t2890 VSS 0.013864f
C15039 VDD.t3615 VSS 0.013864f
C15040 VDD.n564 VSS 0.029707f
C15041 VDD.n565 VSS 0.011881f
C15042 VDD.t780 VSS 0.014787f
C15043 VDD.t1554 VSS 0.014787f
C15044 VDD.t1984 VSS 0.013864f
C15045 VDD.t2876 VSS 0.013864f
C15046 VDD.n567 VSS 0.032563f
C15047 VDD.n568 VSS 0.01221f
C15048 VDD.n571 VSS 0.026075f
C15049 VDD.n574 VSS 0.028639f
C15050 VDD.n576 VSS 0.038332f
C15051 VDD.n577 VSS 0.011881f
C15052 VDD.n578 VSS 0.011881f
C15053 VDD.n580 VSS 0.028059f
C15054 VDD.n583 VSS 0.011881f
C15055 VDD.n584 VSS 0.011881f
C15056 VDD.n587 VSS 0.026075f
C15057 VDD.n589 VSS 0.011881f
C15058 VDD.n590 VSS 0.011881f
C15059 VDD.n591 VSS 0.011881f
C15060 VDD.n593 VSS 0.028059f
C15061 VDD.n595 VSS 0.044176f
C15062 VDD.n596 VSS 0.011881f
C15063 VDD.n597 VSS 0.011881f
C15064 VDD.n598 VSS 0.011881f
C15065 VDD.n600 VSS 0.015687f
C15066 VDD.n603 VSS 0.010719f
C15067 VDD.n604 VSS 0.015799f
C15068 VDD.n605 VSS 0.508827f
C15069 VDD.n607 VSS 0.011881f
C15070 VDD.t131 VSS 0.010137f
C15071 VDD.t3819 VSS 0.021516f
C15072 VDD.n610 VSS 0.055166f
C15073 VDD.t132 VSS 0.010137f
C15074 VDD.n611 VSS 0.027282f
C15075 VDD.t724 VSS 0.014683f
C15076 VDD.n613 VSS 0.011881f
C15077 VDD.n614 VSS 0.010077f
C15078 VDD.n615 VSS 0.010077f
C15079 VDD.n616 VSS 0.015687f
C15080 VDD.n617 VSS 0.042008f
C15081 VDD.t1375 VSS 0.014683f
C15082 VDD.t1047 VSS 0.014683f
C15083 VDD.n620 VSS 0.019839f
C15084 VDD.n622 VSS 0.012144f
C15085 VDD.n625 VSS 0.011881f
C15086 VDD.n626 VSS 0.011881f
C15087 VDD.n630 VSS 0.011881f
C15088 VDD.n631 VSS 0.011881f
C15089 VDD.n632 VSS 0.013239f
C15090 VDD.n635 VSS 0.010077f
C15091 VDD.n636 VSS 0.051089f
C15092 VDD.n637 VSS 0.011881f
C15093 VDD.t1046 VSS 0.146946f
C15094 VDD.t1044 VSS 0.063956f
C15095 VDD.t1050 VSS 0.063956f
C15096 VDD.t1048 VSS 0.070428f
C15097 VDD.t2922 VSS 0.065859f
C15098 VDD.t1876 VSS 0.110781f
C15099 VDD.t723 VSS 0.092888f
C15100 VDD.t130 VSS 0.031978f
C15101 VDD.t721 VSS 0.054439f
C15102 VDD.t717 VSS 0.063956f
C15103 VDD.t719 VSS 0.070428f
C15104 VDD.t2891 VSS 0.065859f
C15105 VDD.t3093 VSS 0.085275f
C15106 VDD.t1889 VSS 0.134003f
C15107 VDD.t2078 VSS 0.071189f
C15108 VDD.t337 VSS 0.071189f
C15109 VDD.t339 VSS 0.065479f
C15110 VDD.t335 VSS 0.065479f
C15111 VDD.t333 VSS 0.108497f
C15112 VDD.t2918 VSS 0.108497f
C15113 VDD.t3611 VSS 0.071189f
C15114 VDD.t1571 VSS 0.071189f
C15115 VDD.t1577 VSS 0.065479f
C15116 VDD.t1573 VSS 0.065479f
C15117 VDD.t1575 VSS 0.037308f
C15118 VDD.t174 VSS 0.057103f
C15119 VDD.n638 VSS 0.116599f
C15120 VDD.t1576 VSS 0.014734f
C15121 VDD.n639 VSS 0.013562f
C15122 VDD.n640 VSS 0.011881f
C15123 VDD.n642 VSS 0.04808f
C15124 VDD.n643 VSS 0.012787f
C15125 VDD.t175 VSS 0.010822f
C15126 VDD.n644 VSS 0.094896f
C15127 VDD.n645 VSS 0.076512f
C15128 VDD.t3822 VSS 0.056694f
C15129 VDD.n646 VSS 0.028405f
C15130 VDD.n647 VSS 0.080035f
C15131 VDD.t176 VSS 0.01172f
C15132 VDD.n648 VSS 0.127534f
C15133 VDD.n649 VSS 0.011881f
C15134 VDD.n651 VSS 0.013403f
C15135 VDD.t2919 VSS 0.013864f
C15136 VDD.n653 VSS 0.011881f
C15137 VDD.t2320 VSS 0.014787f
C15138 VDD.t334 VSS 0.014787f
C15139 VDD.n654 VSS 0.028059f
C15140 VDD.n659 VSS 0.028639f
C15141 VDD.t2106 VSS 0.013864f
C15142 VDD.t1890 VSS 0.013864f
C15143 VDD.n660 VSS 0.032563f
C15144 VDD.n661 VSS 0.01221f
C15145 VDD.n662 VSS 0.038332f
C15146 VDD.n664 VSS 0.026075f
C15147 VDD.n667 VSS 0.011881f
C15148 VDD.n668 VSS 0.011881f
C15149 VDD.n669 VSS 0.011881f
C15150 VDD.n671 VSS 0.015905f
C15151 VDD.n674 VSS 0.011881f
C15152 VDD.n675 VSS 0.011881f
C15153 VDD.n677 VSS 0.014089f
C15154 VDD.n680 VSS 0.011881f
C15155 VDD.n681 VSS 0.011881f
C15156 VDD.n683 VSS 0.024192f
C15157 VDD.n685 VSS 0.011881f
C15158 VDD.n686 VSS 0.011881f
C15159 VDD.n691 VSS 0.010719f
C15160 VDD.n692 VSS 0.015799f
C15161 VDD.n693 VSS 0.665722f
C15162 VDD.n694 VSS 1.07877f
C15163 VDD.n695 VSS 2.36623f
C15164 VDD.t772 VSS 0.014745f
C15165 VDD.n701 VSS 0.019856f
C15166 VDD.n705 VSS 0.011881f
C15167 VDD.t1920 VSS 0.012528f
C15168 VDD.t819 VSS 0.015994f
C15169 VDD.n706 VSS 0.010205f
C15170 VDD.n708 VSS 0.011881f
C15171 VDD.t813 VSS 0.013927f
C15172 VDD.n710 VSS 0.011863f
C15173 VDD.n711 VSS 0.011881f
C15174 VDD.t2851 VSS 0.085275f
C15175 VDD.t3453 VSS 0.014484f
C15176 VDD.n712 VSS 0.019104f
C15177 VDD.n713 VSS 0.011881f
C15178 VDD.n718 VSS 0.011881f
C15179 VDD.t3438 VSS 0.014219f
C15180 VDD.n721 VSS 0.022117f
C15181 VDD.n722 VSS 0.011881f
C15182 VDD.t3532 VSS 0.01383f
C15183 VDD.n723 VSS 0.013668f
C15184 VDD.n724 VSS 0.018529f
C15185 VDD.n725 VSS 0.011881f
C15186 VDD.n726 VSS 0.010534f
C15187 VDD.t46 VSS 0.014469f
C15188 VDD.t2048 VSS 0.014485f
C15189 VDD.n727 VSS 0.019318f
C15190 VDD.n728 VSS 0.011881f
C15191 VDD.t2732 VSS 0.01449f
C15192 VDD.n730 VSS 0.011881f
C15193 VDD.t444 VSS 0.012563f
C15194 VDD.n731 VSS 0.014135f
C15195 VDD.n732 VSS 0.011881f
C15196 VDD.n733 VSS 0.014537f
C15197 VDD.n736 VSS 0.011881f
C15198 VDD.t3454 VSS 0.033501f
C15199 VDD.t3616 VSS 0.031978f
C15200 VDD.t3470 VSS 0.062433f
C15201 VDD.t3466 VSS 0.041114f
C15202 VDD.t1979 VSS 0.031978f
C15203 VDD.t3526 VSS 0.033501f
C15204 VDD.t1695 VSS 0.031978f
C15205 VDD.t3552 VSS 0.053297f
C15206 VDD.t3529 VSS 0.056342f
C15207 VDD.t3437 VSS 0.031978f
C15208 VDD.t3531 VSS 0.02741f
C15209 VDD.t2966 VSS 0.091366f
C15210 VDD.t1354 VSS 0.072331f
C15211 VDD.t2501 VSS 0.028171f
C15212 VDD.t977 VSS 0.035404f
C15213 VDD.t47 VSS 0.036546f
C15214 VDD.t698 VSS 0.031978f
C15215 VDD.t45 VSS 0.037308f
C15216 VDD.t2502 VSS 0.089843f
C15217 VDD.t3451 VSS 0.073092f
C15218 VDD.t2047 VSS 0.036927f
C15219 VDD.t427 VSS 0.031978f
C15220 VDD.t2731 VSS 0.031978f
C15221 VDD.t924 VSS 0.051774f
C15222 VDD.t2587 VSS 0.070808f
C15223 VDD.t3537 VSS 0.075377f
C15224 VDD.t676 VSS 0.052535f
C15225 VDD.t327 VSS 0.02741f
C15226 VDD.t2305 VSS 0.031978f
C15227 VDD.t561 VSS 0.081468f
C15228 VDD.t328 VSS 0.070808f
C15229 VDD.t443 VSS 0.039211f
C15230 VDD.t3533 VSS 0.035785f
C15231 VDD.t3478 VSS 0.041495f
C15232 VDD.t1441 VSS 0.106974f
C15233 VDD.t1423 VSS 0.08832f
C15234 VDD.n737 VSS 0.043887f
C15235 VDD.n738 VSS 0.010783f
C15236 VDD.n740 VSS 0.011881f
C15237 VDD.n741 VSS 0.011881f
C15238 VDD.t2012 VSS 0.0145f
C15239 VDD.n743 VSS 0.011881f
C15240 VDD.t1106 VSS 0.012563f
C15241 VDD.n744 VSS 0.014135f
C15242 VDD.n745 VSS 0.011881f
C15243 VDD.n746 VSS 0.012976f
C15244 VDD.n749 VSS 0.011881f
C15245 VDD.n750 VSS 0.013668f
C15246 VDD.t1804 VSS 0.012563f
C15247 VDD.n751 VSS 0.011881f
C15248 VDD.t2860 VSS 0.014675f
C15249 VDD.n753 VSS 0.015289f
C15250 VDD.n754 VSS 0.011881f
C15251 VDD.t3717 VSS 0.014219f
C15252 VDD.n755 VSS 0.035607f
C15253 VDD.n756 VSS 0.011881f
C15254 VDD.t2904 VSS 0.014219f
C15255 VDD.n757 VSS 0.026112f
C15256 VDD.n758 VSS 0.011881f
C15257 VDD.n759 VSS 0.024663f
C15258 VDD.n760 VSS 0.044694f
C15259 VDD.n761 VSS 0.011881f
C15260 VDD.n762 VSS 0.013668f
C15261 VDD.t526 VSS 0.012563f
C15262 VDD.t913 VSS 0.014675f
C15263 VDD.n763 VSS 0.029824f
C15264 VDD.n764 VSS 0.011881f
C15265 VDD.t3776 VSS 0.041965f
C15266 VDD.n766 VSS 0.037956f
C15267 VDD.n767 VSS 0.011881f
C15268 VDD.n769 VSS 0.011881f
C15269 VDD.n772 VSS 0.011881f
C15270 VDD.t1806 VSS 0.014219f
C15271 VDD.n774 VSS 0.011881f
C15272 VDD.t2247 VSS 0.010806f
C15273 VDD.n777 VSS 0.012208f
C15274 VDD.n778 VSS 0.011881f
C15275 VDD.n779 VSS 0.013523f
C15276 VDD.n780 VSS 0.011881f
C15277 VDD.t1404 VSS 0.014745f
C15278 VDD.n782 VSS 0.011385f
C15279 VDD.n783 VSS 0.011881f
C15280 VDD.n784 VSS 0.012923f
C15281 VDD.t1466 VSS 0.013927f
C15282 VDD.n786 VSS 0.011881f
C15283 VDD.t3138 VSS 0.085275f
C15284 VDD.n792 VSS 0.011881f
C15285 VDD.n794 VSS 0.011881f
C15286 VDD.n795 VSS 0.013668f
C15287 VDD.n796 VSS 0.011881f
C15288 VDD.n797 VSS 0.011881f
C15289 VDD.t452 VSS 0.014745f
C15290 VDD.n799 VSS 0.011881f
C15291 VDD.n801 VSS 0.012923f
C15292 VDD.t1524 VSS 0.010846f
C15293 VDD.n802 VSS 0.015964f
C15294 VDD.n803 VSS 0.011881f
C15295 VDD.n805 VSS 0.011363f
C15296 VDD.n806 VSS 0.011881f
C15297 VDD.t2601 VSS 0.013927f
C15298 VDD.n808 VSS 0.012081f
C15299 VDD.n809 VSS 0.011881f
C15300 VDD.t2599 VSS 0.015994f
C15301 VDD.n812 VSS 0.011881f
C15302 VDD.t2769 VSS 0.014745f
C15303 VDD.n813 VSS 0.013523f
C15304 VDD.n816 VSS 0.011881f
C15305 VDD.t3626 VSS 0.0145f
C15306 VDD.n817 VSS 0.023826f
C15307 VDD.t2924 VSS 0.073092f
C15308 VDD.n820 VSS 0.011881f
C15309 VDD.n822 VSS 0.012976f
C15310 VDD.n823 VSS 0.012483f
C15311 VDD.n824 VSS 0.011881f
C15312 VDD.n825 VSS 0.013606f
C15313 VDD.n826 VSS 0.015706f
C15314 VDD.n827 VSS 0.011881f
C15315 VDD.n828 VSS 0.011881f
C15316 VDD.n829 VSS 0.012244f
C15317 VDD.n830 VSS 0.011881f
C15318 VDD.n832 VSS 0.011881f
C15319 VDD.n836 VSS 0.011881f
C15320 VDD.n837 VSS 0.011881f
C15321 VDD.t2180 VSS 0.014745f
C15322 VDD.n839 VSS 0.013668f
C15323 VDD.n840 VSS 0.024573f
C15324 VDD.n841 VSS 0.011881f
C15325 VDD.t2135 VSS 0.015901f
C15326 VDD.n842 VSS 0.011881f
C15327 VDD.n843 VSS 0.013668f
C15328 VDD.t408 VSS 0.017003f
C15329 VDD.t262 VSS 0.014714f
C15330 VDD.n844 VSS 0.038996f
C15331 VDD.n845 VSS 0.011881f
C15332 VDD.n846 VSS 0.017519f
C15333 VDD.n847 VSS 0.021056f
C15334 VDD.t147 VSS 0.222704f
C15335 VDD.t3334 VSS 0.091746f
C15336 VDD.t1238 VSS 0.031978f
C15337 VDD.t3332 VSS 0.032739f
C15338 VDD.t1236 VSS 0.036166f
C15339 VDD.t2034 VSS 0.032739f
C15340 VDD.t1234 VSS 0.03312f
C15341 VDD.t1240 VSS 0.069286f
C15342 VDD.t2569 VSS 0.044541f
C15343 VDD.t1991 VSS 0.035404f
C15344 VDD.t835 VSS 0.080706f
C15345 VDD.t1438 VSS 0.014469f
C15346 VDD.n848 VSS 0.017319f
C15347 VDD.n850 VSS 0.011881f
C15348 VDD.t1992 VSS 0.014219f
C15349 VDD.n854 VSS 0.011881f
C15350 VDD.n855 VSS 0.013523f
C15351 VDD.t1239 VSS 0.015761f
C15352 VDD.t3335 VSS 0.014469f
C15353 VDD.n856 VSS 0.017319f
C15354 VDD.t172 VSS 0.010137f
C15355 VDD.t3818 VSS 0.021516f
C15356 VDD.n858 VSS 0.055166f
C15357 VDD.t173 VSS 0.010137f
C15358 VDD.n859 VSS 0.030049f
C15359 VDD.t148 VSS 0.010137f
C15360 VDD.t3796 VSS 0.021516f
C15361 VDD.n861 VSS 0.055166f
C15362 VDD.t149 VSS 0.010137f
C15363 VDD.n862 VSS 0.030049f
C15364 VDD.n863 VSS 0.027374f
C15365 VDD.n864 VSS 0.045507f
C15366 VDD.n866 VSS 0.015826f
C15367 VDD.n868 VSS 0.015061f
C15368 VDD.n870 VSS 0.011881f
C15369 VDD.n871 VSS 0.011881f
C15370 VDD.n873 VSS 0.014892f
C15371 VDD.n875 VSS 0.022117f
C15372 VDD.n877 VSS 0.011881f
C15373 VDD.n878 VSS 0.011881f
C15374 VDD.n879 VSS 0.011881f
C15375 VDD.t256 VSS 0.014219f
C15376 VDD.n881 VSS 0.013668f
C15377 VDD.n882 VSS 0.011881f
C15378 VDD.n883 VSS 0.013104f
C15379 VDD.t2807 VSS 0.014745f
C15380 VDD.n884 VSS 0.011881f
C15381 VDD.n886 VSS 0.011881f
C15382 VDD.n887 VSS 0.013931f
C15383 VDD.n888 VSS 0.01469f
C15384 VDD.n889 VSS 0.013523f
C15385 VDD.t2792 VSS 0.014469f
C15386 VDD.n890 VSS 0.017982f
C15387 VDD.n891 VSS 0.011881f
C15388 VDD.n893 VSS 0.011881f
C15389 VDD.n895 VSS 0.014257f
C15390 VDD.n896 VSS 0.013523f
C15391 VDD.n898 VSS 0.014064f
C15392 VDD.n899 VSS 0.011881f
C15393 VDD.n900 VSS 0.013668f
C15394 VDD.n901 VSS 0.017065f
C15395 VDD.n902 VSS 0.011881f
C15396 VDD.n903 VSS 0.011881f
C15397 VDD.t2218 VSS 0.014745f
C15398 VDD.n905 VSS 0.020999f
C15399 VDD.n907 VSS 0.011881f
C15400 VDD.n908 VSS 0.011881f
C15401 VDD.n909 VSS 0.011881f
C15402 VDD.t1729 VSS 0.014745f
C15403 VDD.n910 VSS 0.020336f
C15404 VDD.n912 VSS 0.015061f
C15405 VDD.n914 VSS 0.011881f
C15406 VDD.n915 VSS 0.011881f
C15407 VDD.n916 VSS 0.011881f
C15408 VDD.t1398 VSS 0.0145f
C15409 VDD.n917 VSS 0.024649f
C15410 VDD.t2558 VSS 0.013749f
C15411 VDD.n918 VSS 0.018467f
C15412 VDD.n920 VSS 0.011881f
C15413 VDD.n921 VSS 0.011881f
C15414 VDD.n923 VSS 0.012435f
C15415 VDD.n925 VSS 0.015061f
C15416 VDD.n927 VSS 0.011881f
C15417 VDD.n928 VSS 0.011881f
C15418 VDD.n929 VSS 0.011881f
C15419 VDD.n931 VSS 0.013668f
C15420 VDD.n932 VSS 0.018529f
C15421 VDD.n934 VSS 0.011881f
C15422 VDD.n935 VSS 0.011881f
C15423 VDD.n936 VSS 0.019467f
C15424 VDD.n938 VSS 0.014066f
C15425 VDD.n939 VSS 0.016065f
C15426 VDD.n941 VSS 0.011881f
C15427 VDD.n942 VSS 0.011881f
C15428 VDD.n943 VSS 0.011881f
C15429 VDD.n944 VSS 0.018529f
C15430 VDD.n946 VSS 0.022117f
C15431 VDD.n948 VSS 0.011881f
C15432 VDD.n949 VSS 0.011881f
C15433 VDD.n950 VSS 0.04473f
C15434 VDD.n951 VSS 0.120098f
C15435 VDD.t1437 VSS 0.059388f
C15436 VDD.t255 VSS 0.031978f
C15437 VDD.t1439 VSS 0.02741f
C15438 VDD.t2962 VSS 0.036166f
C15439 VDD.t1435 VSS 0.08832f
C15440 VDD.t1147 VSS 0.094411f
C15441 VDD.t3516 VSS 0.073092f
C15442 VDD.t1529 VSS 0.047586f
C15443 VDD.t2806 VSS 0.047586f
C15444 VDD.t2808 VSS 0.068144f
C15445 VDD.t2559 VSS 0.089462f
C15446 VDD.t2290 VSS 0.07157f
C15447 VDD.t2865 VSS 0.041114f
C15448 VDD.t1533 VSS 0.036166f
C15449 VDD.t2789 VSS 0.031978f
C15450 VDD.t3422 VSS 0.031978f
C15451 VDD.t2791 VSS 0.085275f
C15452 VDD.t2968 VSS 0.072712f
C15453 VDD.t2557 VSS 0.02741f
C15454 VDD.t1397 VSS 0.07157f
C15455 VDD.t716 VSS 0.07728f
C15456 VDD.t3027 VSS 0.032739f
C15457 VDD.t2088 VSS 0.032739f
C15458 VDD.t3514 VSS 0.036166f
C15459 VDD.t1726 VSS 0.035785f
C15460 VDD.t1728 VSS 0.068905f
C15461 VDD.t3021 VSS 0.071189f
C15462 VDD.t997 VSS 0.066621f
C15463 VDD.t1308 VSS 0.071189f
C15464 VDD.t2217 VSS 0.043399f
C15465 VDD.t3732 VSS 0.031978f
C15466 VDD.t2219 VSS 0.038069f
C15467 VDD.t1531 VSS 0.036166f
C15468 VDD.t3724 VSS 0.059007f
C15469 VDD.t405 VSS 0.053297f
C15470 VDD.t2281 VSS 0.033501f
C15471 VDD.t2373 VSS 0.031978f
C15472 VDD.t999 VSS 0.050251f
C15473 VDD.t3659 VSS 0.068905f
C15474 VDD.t251 VSS 0.096695f
C15475 VDD.t1310 VSS 0.089462f
C15476 VDD.t3134 VSS 0.048348f
C15477 VDD.t3735 VSS 0.031978f
C15478 VDD.t1119 VSS 0.036546f
C15479 VDD.t3015 VSS 0.068905f
C15480 VDD.t2982 VSS 0.078422f
C15481 VDD.t2861 VSS 0.039592f
C15482 VDD.t1307 VSS 0.035023f
C15483 VDD.t1122 VSS 0.032739f
C15484 VDD.t571 VSS 0.037688f
C15485 VDD.t1118 VSS 0.07195f
C15486 VDD.t2988 VSS 0.053297f
C15487 VDD.t2626 VSS 0.037308f
C15488 VDD.t1741 VSS 0.036927f
C15489 VDD.t3355 VSS 0.033501f
C15490 VDD.t1999 VSS 0.074996f
C15491 VDD.t2543 VSS 0.067763f
C15492 VDD.t1743 VSS 0.037688f
C15493 VDD.t1117 VSS 0.058246f
C15494 VDD.t1121 VSS 0.046444f
C15495 VDD.t2179 VSS 0.031978f
C15496 VDD.t2136 VSS 0.031978f
C15497 VDD.t2181 VSS 0.041114f
C15498 VDD.t3420 VSS 0.036166f
C15499 VDD.t2177 VSS 0.031978f
C15500 VDD.t2132 VSS 0.07157f
C15501 VDD.t3558 VSS 0.081848f
C15502 VDD.t2134 VSS 0.036166f
C15503 VDD.t263 VSS 0.034643f
C15504 VDD.t261 VSS 0.073473f
C15505 VDD.t407 VSS 0.053677f
C15506 VDD.n952 VSS 0.03854f
C15507 VDD.n953 VSS 0.024126f
C15508 VDD.n954 VSS 0.011881f
C15509 VDD.n955 VSS 0.011881f
C15510 VDD.n956 VSS 0.011881f
C15511 VDD.n958 VSS 0.037543f
C15512 VDD.n960 VSS 0.010708f
C15513 VDD.n962 VSS 0.011881f
C15514 VDD.n963 VSS 0.011881f
C15515 VDD.n964 VSS 0.011881f
C15516 VDD.n966 VSS 0.020999f
C15517 VDD.t2544 VSS 0.010806f
C15518 VDD.n968 VSS 0.015958f
C15519 VDD.n974 VSS 0.011881f
C15520 VDD.n975 VSS 0.011881f
C15521 VDD.n976 VSS 0.011881f
C15522 VDD.n982 VSS 0.011881f
C15523 VDD.n983 VSS 0.011881f
C15524 VDD.n984 VSS 0.011881f
C15525 VDD.n986 VSS 0.011584f
C15526 VDD.n987 VSS 0.012031f
C15527 VDD.n990 VSS 0.010157f
C15528 VDD.n992 VSS 0.011881f
C15529 VDD.n993 VSS 0.011881f
C15530 VDD.n997 VSS 0.011881f
C15531 VDD.n998 VSS 0.011881f
C15532 VDD.n1001 VSS 0.018529f
C15533 VDD.n1002 VSS 0.011881f
C15534 VDD.n1003 VSS 0.011881f
C15535 VDD.n1004 VSS 0.011881f
C15536 VDD.n1006 VSS 0.012081f
C15537 VDD.n1007 VSS 0.013523f
C15538 VDD.t2996 VSS 0.012563f
C15539 VDD.n1009 VSS 0.011881f
C15540 VDD.n1011 VSS 0.011881f
C15541 VDD.t1446 VSS 0.013611f
C15542 VDD.n1013 VSS 0.017733f
C15543 VDD.n1014 VSS 0.011881f
C15544 VDD.t2813 VSS 0.010846f
C15545 VDD.n1015 VSS 0.015918f
C15546 VDD.n1016 VSS 0.011881f
C15547 VDD.t833 VSS 0.012751f
C15548 VDD.n1020 VSS 0.011385f
C15549 VDD.n1021 VSS 0.011881f
C15550 VDD.t1637 VSS 0.013927f
C15551 VDD.n1024 VSS 0.011881f
C15552 VDD.n1025 VSS 0.011881f
C15553 VDD.t1633 VSS 0.015994f
C15554 VDD.n1031 VSS 0.011881f
C15555 VDD.n1032 VSS 0.011881f
C15556 VDD.n1033 VSS 0.011881f
C15557 VDD.n1034 VSS 0.015472f
C15558 VDD.n1035 VSS 0.011863f
C15559 VDD.n1037 VSS 0.010708f
C15560 VDD.n1039 VSS 0.011881f
C15561 VDD.n1040 VSS 0.011881f
C15562 VDD.n1041 VSS 0.011881f
C15563 VDD.n1046 VSS 0.011881f
C15564 VDD.n1047 VSS 0.011881f
C15565 VDD.n1048 VSS 0.011881f
C15566 VDD.n1052 VSS 0.011101f
C15567 VDD.n1054 VSS 0.011881f
C15568 VDD.n1055 VSS 0.011881f
C15569 VDD.n1056 VSS 0.011881f
C15570 VDD.n1059 VSS 0.015838f
C15571 VDD.n1061 VSS 0.011881f
C15572 VDD.n1062 VSS 0.011881f
C15573 VDD.n1066 VSS 0.014404f
C15574 VDD.n1067 VSS 0.011881f
C15575 VDD.n1068 VSS 0.011881f
C15576 VDD.n1069 VSS 0.011881f
C15577 VDD.t560 VSS 0.014675f
C15578 VDD.n1070 VSS 0.029806f
C15579 VDD.n1072 VSS 0.015061f
C15580 VDD.n1074 VSS 0.011881f
C15581 VDD.n1075 VSS 0.011881f
C15582 VDD.n1076 VSS 0.011881f
C15583 VDD.n1077 VSS 0.044776f
C15584 VDD.n1078 VSS 0.119717f
C15585 VDD.t555 VSS 0.08832f
C15586 VDD.t2098 VSS 0.036166f
C15587 VDD.t557 VSS 0.03312f
C15588 VDD.t559 VSS 0.034643f
C15589 VDD.t2995 VSS 0.07195f
C15590 VDD.t3147 VSS 0.070808f
C15591 VDD.t1906 VSS 0.031978f
C15592 VDD.t2506 VSS 0.031978f
C15593 VDD.t1690 VSS 0.073854f
C15594 VDD.t1445 VSS 0.100121f
C15595 VDD.t902 VSS 0.062814f
C15596 VDD.t2479 VSS 0.043779f
C15597 VDD.t572 VSS 0.037688f
C15598 VDD.t2508 VSS 0.032359f
C15599 VDD.t2984 VSS 0.036166f
C15600 VDD.t1899 VSS 0.04987f
C15601 VDD.t2814 VSS 0.054058f
C15602 VDD.t1855 VSS 0.09365f
C15603 VDD.t834 VSS 0.074996f
C15604 VDD.t2812 VSS 0.031978f
C15605 VDD.t3671 VSS 0.037688f
C15606 VDD.t2505 VSS 0.031978f
C15607 VDD.t3657 VSS 0.032739f
C15608 VDD.t2480 VSS 0.031978f
C15609 VDD.t832 VSS 0.031978f
C15610 VDD.t1628 VSS 0.065859f
C15611 VDD.t1831 VSS 0.046825f
C15612 VDD.t2652 VSS 0.031978f
C15613 VDD.t2481 VSS 0.074615f
C15614 VDD.t2884 VSS 0.074235f
C15615 VDD.t1636 VSS 0.033501f
C15616 VDD.t729 VSS 0.031978f
C15617 VDD.t1630 VSS 0.056342f
C15618 VDD.t1634 VSS 0.063956f
C15619 VDD.t1632 VSS 0.091366f
C15620 VDD.t3625 VSS 0.070047f
C15621 VDD.t1668 VSS 0.070047f
C15622 VDD.t449 VSS 0.074235f
C15623 VDD.t453 VSS 0.063575f
C15624 VDD.t2321 VSS 0.031978f
C15625 VDD.t451 VSS 0.035023f
C15626 VDD.t1285 VSS 0.068144f
C15627 VDD.t1667 VSS 0.090985f
C15628 VDD.t1525 VSS 0.056723f
C15629 VDD.t3274 VSS 0.036927f
C15630 VDD.t1837 VSS 0.036927f
C15631 VDD.t3302 VSS 0.035404f
C15632 VDD.t2339 VSS 0.063956f
C15633 VDD.t1271 VSS 0.039592f
C15634 VDD.t1523 VSS 0.045302f
C15635 VDD.t1666 VSS 0.070428f
C15636 VDD.t1286 VSS 0.046063f
C15637 VDD.t3624 VSS 0.031978f
C15638 VDD.t2596 VSS 0.031978f
C15639 VDD.t1896 VSS 0.041114f
C15640 VDD.t1847 VSS 0.059768f
C15641 VDD.t1670 VSS 0.043018f
C15642 VDD.t240 VSS 0.046825f
C15643 VDD.t3017 VSS 0.063194f
C15644 VDD.t2600 VSS 0.035023f
C15645 VDD.t1652 VSS 0.031978f
C15646 VDD.t2592 VSS 0.056342f
C15647 VDD.t2594 VSS 0.063956f
C15648 VDD.t2598 VSS 0.085655f
C15649 VDD.t2768 VSS 0.085655f
C15650 VDD.t2770 VSS 0.034643f
C15651 VDD.t2571 VSS 0.036166f
C15652 VDD.t2766 VSS 0.10507f
C15653 VDD.t2965 VSS 0.08832f
C15654 VDD.n1079 VSS 0.033972f
C15655 VDD.n1080 VSS 0.024263f
C15656 VDD.n1082 VSS 0.011881f
C15657 VDD.n1083 VSS 0.011881f
C15658 VDD.n1084 VSS 0.011881f
C15659 VDD.n1085 VSS 0.015221f
C15660 VDD.n1086 VSS 0.015061f
C15661 VDD.n1088 VSS 0.020039f
C15662 VDD.n1089 VSS 0.011881f
C15663 VDD.n1090 VSS 0.011881f
C15664 VDD.n1095 VSS 0.011881f
C15665 VDD.n1096 VSS 0.011881f
C15666 VDD.n1098 VSS 0.011863f
C15667 VDD.t241 VSS 0.012528f
C15668 VDD.n1101 VSS 0.010167f
C15669 VDD.n1103 VSS 0.011881f
C15670 VDD.n1104 VSS 0.011881f
C15671 VDD.n1105 VSS 0.011881f
C15672 VDD.n1109 VSS 0.011881f
C15673 VDD.n1110 VSS 0.011881f
C15674 VDD.n1111 VSS 0.011881f
C15675 VDD.n1117 VSS 0.011881f
C15676 VDD.n1118 VSS 0.011881f
C15677 VDD.n1119 VSS 0.011881f
C15678 VDD.n1121 VSS 0.020862f
C15679 VDD.n1122 VSS 0.010349f
C15680 VDD.n1123 VSS 0.017523f
C15681 VDD.n1125 VSS 0.014404f
C15682 VDD.n1126 VSS 0.011881f
C15683 VDD.n1127 VSS 0.011881f
C15684 VDD.n1128 VSS 0.011881f
C15685 VDD.n1131 VSS 0.011881f
C15686 VDD.n1132 VSS 0.011881f
C15687 VDD.t3635 VSS 0.012563f
C15688 VDD.n1133 VSS 0.011812f
C15689 VDD.n1134 VSS 0.011881f
C15690 VDD.n1135 VSS 0.011881f
C15691 VDD.n1138 VSS 0.011101f
C15692 VDD.n1139 VSS 0.011881f
C15693 VDD.t2883 VSS 0.010806f
C15694 VDD.t2412 VSS 0.014469f
C15695 VDD.n1141 VSS 0.011881f
C15696 VDD.n1142 VSS 0.013668f
C15697 VDD.n1144 VSS 0.011881f
C15698 VDD.n1146 VSS 0.011881f
C15699 VDD.t520 VSS 0.014219f
C15700 VDD.n1147 VSS 0.020814f
C15701 VDD.t915 VSS 0.013927f
C15702 VDD.n1148 VSS 0.011881f
C15703 VDD.n1152 VSS 0.011881f
C15704 VDD.t919 VSS 0.015994f
C15705 VDD.t3264 VSS 0.012528f
C15706 VDD.n1154 VSS 0.010182f
C15707 VDD.t1460 VSS 0.015994f
C15708 VDD.n1155 VSS 0.010205f
C15709 VDD.n1158 VSS 0.011881f
C15710 VDD.n1159 VSS 0.011881f
C15711 VDD.n1160 VSS 0.011881f
C15712 VDD.n1163 VSS 0.014405f
C15713 VDD.n1165 VSS 0.011863f
C15714 VDD.n1167 VSS 0.011881f
C15715 VDD.n1168 VSS 0.011881f
C15716 VDD.n1170 VSS 0.011385f
C15717 VDD.n1172 VSS 0.018529f
C15718 VDD.n1173 VSS 0.011881f
C15719 VDD.n1174 VSS 0.011881f
C15720 VDD.n1175 VSS 0.011881f
C15721 VDD.n1177 VSS 0.016565f
C15722 VDD.n1178 VSS 0.012162f
C15723 VDD.n1181 VSS 0.011881f
C15724 VDD.n1182 VSS 0.011881f
C15725 VDD.n1184 VSS 0.018529f
C15726 VDD.n1187 VSS 0.011881f
C15727 VDD.n1188 VSS 0.011881f
C15728 VDD.n1189 VSS 0.011881f
C15729 VDD.n1191 VSS 0.013426f
C15730 VDD.n1192 VSS 0.013261f
C15731 VDD.n1193 VSS 0.014382f
C15732 VDD.n1195 VSS 0.011881f
C15733 VDD.n1196 VSS 0.011881f
C15734 VDD.n1197 VSS 0.011881f
C15735 VDD.n1198 VSS 0.044776f
C15736 VDD.n1199 VSS 0.154741f
C15737 VDD.t865 VSS 0.123344f
C15738 VDD.t3011 VSS 0.067001f
C15739 VDD.t2697 VSS 0.035785f
C15740 VDD.t3634 VSS 0.074615f
C15741 VDD.t1897 VSS 0.097837f
C15742 VDD.t2583 VSS 0.031978f
C15743 VDD.t3269 VSS 0.035023f
C15744 VDD.t3324 VSS 0.067763f
C15745 VDD.t2696 VSS 0.041495f
C15746 VDD.t2107 VSS 0.037308f
C15747 VDD.t2538 VSS 0.04949f
C15748 VDD.t2337 VSS 0.052916f
C15749 VDD.t1845 VSS 0.111923f
C15750 VDD.t2882 VSS 0.089081f
C15751 VDD.t2411 VSS 0.037688f
C15752 VDD.t2699 VSS 0.031978f
C15753 VDD.t2413 VSS 0.032739f
C15754 VDD.t3325 VSS 0.036166f
C15755 VDD.t2777 VSS 0.031978f
C15756 VDD.t920 VSS 0.061291f
C15757 VDD.t1853 VSS 0.051393f
C15758 VDD.t2964 VSS 0.031978f
C15759 VDD.t3326 VSS 0.02741f
C15760 VDD.t519 VSS 0.074235f
C15761 VDD.t914 VSS 0.077661f
C15762 VDD.t2581 VSS 0.031978f
C15763 VDD.t916 VSS 0.035023f
C15764 VDD.t3019 VSS 0.031978f
C15765 VDD.t922 VSS 0.035785f
C15766 VDD.t3263 VSS 0.031978f
C15767 VDD.t918 VSS 0.070808f
C15768 VDD.t1895 VSS 0.086797f
C15769 VDD.t515 VSS 0.050251f
C15770 VDD.t1459 VSS 0.050251f
C15771 VDD.t1463 VSS 0.035023f
C15772 VDD.t3472 VSS 0.057103f
C15773 VDD.t2907 VSS 0.072331f
C15774 VDD.t425 VSS 0.072331f
C15775 VDD.t2011 VSS 0.036546f
C15776 VDD.t1555 VSS 0.02741f
C15777 VDD.t2967 VSS 0.098218f
C15778 VDD.t2306 VSS 0.103548f
C15779 VDD.t1558 VSS 0.054819f
C15780 VDD.t2793 VSS 0.054819f
C15781 VDD.t2298 VSS 0.047967f
C15782 VDD.t1105 VSS 0.031978f
C15783 VDD.t1097 VSS 0.035785f
C15784 VDD.t3474 VSS 0.036927f
C15785 VDD.t2005 VSS 0.035023f
C15786 VDD.t1559 VSS 0.089462f
C15787 VDD.t1717 VSS 0.103548f
C15788 VDD.t1901 VSS 0.036166f
C15789 VDD.t2857 VSS 0.036166f
C15790 VDD.t2859 VSS 0.066621f
C15791 VDD.t1803 VSS 0.070428f
C15792 VDD.t2094 VSS 0.037308f
C15793 VDD.t2296 VSS 0.035023f
C15794 VDD.t1415 VSS 0.10507f
C15795 VDD.t2969 VSS 0.098979f
C15796 VDD.t3716 VSS 0.104309f
C15797 VDD.t212 VSS 0.083752f
C15798 VDD.t2903 VSS 0.034262f
C15799 VDD.t2959 VSS 0.150753f
C15800 VDD.n1200 VSS 0.189764f
C15801 VDD.t1877 VSS 0.085275f
C15802 VDD.t1898 VSS 0.036166f
C15803 VDD.t910 VSS 0.036166f
C15804 VDD.t912 VSS 0.066621f
C15805 VDD.t525 VSS 0.070428f
C15806 VDD.t2092 VSS 0.070808f
C15807 VDD.t1516 VSS 0.035785f
C15808 VDD.t221 VSS 0.07157f
C15809 VDD.t3128 VSS 0.102786f
C15810 VDD.t1675 VSS 0.035023f
C15811 VDD.t3233 VSS 0.036546f
C15812 VDD.t1259 VSS 0.098599f
C15813 VDD.t1518 VSS 0.077661f
C15814 VDD.t1805 VSS 0.035023f
C15815 VDD.t1679 VSS 0.02741f
C15816 VDD.t2963 VSS 0.037688f
C15817 VDD.t1677 VSS 0.07157f
C15818 VDD.t3687 VSS 0.053297f
C15819 VDD.t2248 VSS 0.033501f
C15820 VDD.t2233 VSS 0.036927f
C15821 VDD.t3391 VSS 0.07157f
C15822 VDD.t2579 VSS 0.074996f
C15823 VDD.t2246 VSS 0.036166f
C15824 VDD.t1401 VSS 0.037688f
C15825 VDD.t1674 VSS 0.031978f
C15826 VDD.t1403 VSS 0.032739f
C15827 VDD.t1678 VSS 0.055581f
C15828 VDD.t1461 VSS 0.068144f
C15829 VDD.t3336 VSS 0.041114f
C15830 VDD.t3375 VSS 0.031978f
C15831 VDD.t2235 VSS 0.031978f
C15832 VDD.t1155 VSS 0.031978f
C15833 VDD.t968 VSS 0.063956f
C15834 VDD.t1811 VSS 0.047206f
C15835 VDD.t1465 VSS 0.042257f
C15836 VDD.t1457 VSS 0.06091f
C15837 VDD.n1201 VSS 0.038176f
C15838 VDD.n1202 VSS 0.022866f
C15839 VDD.n1203 VSS 0.011881f
C15840 VDD.n1204 VSS 0.011881f
C15841 VDD.n1205 VSS 0.011881f
C15842 VDD.n1207 VSS 0.011086f
C15843 VDD.n1208 VSS 0.010615f
C15844 VDD.n1210 VSS 0.010708f
C15845 VDD.n1212 VSS 0.011881f
C15846 VDD.n1213 VSS 0.011881f
C15847 VDD.n1214 VSS 0.011881f
C15848 VDD.n1216 VSS 0.020999f
C15849 VDD.n1218 VSS 0.015061f
C15850 VDD.n1220 VSS 0.011881f
C15851 VDD.n1221 VSS 0.011881f
C15852 VDD.n1225 VSS 0.016181f
C15853 VDD.n1226 VSS 0.011881f
C15854 VDD.n1227 VSS 0.011881f
C15855 VDD.n1228 VSS 0.011881f
C15856 VDD.n1231 VSS 0.022117f
C15857 VDD.n1233 VSS 0.011881f
C15858 VDD.n1234 VSS 0.011881f
C15859 VDD.n1236 VSS 0.01782f
C15860 VDD.n1237 VSS 0.013668f
C15861 VDD.t222 VSS 0.010055f
C15862 VDD.n1239 VSS 0.010807f
C15863 VDD.n1240 VSS 0.011881f
C15864 VDD.n1241 VSS 0.011881f
C15865 VDD.n1242 VSS 0.021695f
C15866 VDD.n1243 VSS 0.02557f
C15867 VDD.n1244 VSS 0.016271f
C15868 VDD.t223 VSS 0.010055f
C15869 VDD.n1245 VSS 0.01771f
C15870 VDD.n1246 VSS 0.010807f
C15871 VDD.n1247 VSS 0.011881f
C15872 VDD.n1248 VSS 0.011881f
C15873 VDD.n1249 VSS 0.011881f
C15874 VDD.n1251 VSS 0.018529f
C15875 VDD.n1253 VSS 0.011881f
C15876 VDD.n1254 VSS 0.011881f
C15877 VDD.n1255 VSS 0.011881f
C15878 VDD.n1256 VSS 0.01552f
C15879 VDD.t213 VSS 0.010055f
C15880 VDD.n1257 VSS 0.017919f
C15881 VDD.n1258 VSS 0.023377f
C15882 VDD.t3817 VSS 0.035362f
C15883 VDD.n1259 VSS 0.016265f
C15884 VDD.n1260 VSS 0.053377f
C15885 VDD.n1261 VSS 0.022029f
C15886 VDD.n1262 VSS 0.024663f
C15887 VDD.n1263 VSS 0.011881f
C15888 VDD.n1264 VSS 0.011881f
C15889 VDD.n1265 VSS 0.020579f
C15890 VDD.n1266 VSS 0.035179f
C15891 VDD.n1267 VSS 0.01661f
C15892 VDD.n1268 VSS 0.01661f
C15893 VDD.n1269 VSS 0.011881f
C15894 VDD.n1270 VSS 0.011881f
C15895 VDD.n1271 VSS 0.029153f
C15896 VDD.t214 VSS 0.010055f
C15897 VDD.n1272 VSS 0.01771f
C15898 VDD.n1273 VSS 0.011917f
C15899 VDD.n1275 VSS 0.012081f
C15900 VDD.n1277 VSS 0.011881f
C15901 VDD.n1278 VSS 0.011881f
C15902 VDD.n1279 VSS 0.011881f
C15903 VDD.n1281 VSS 0.029806f
C15904 VDD.n1283 VSS 0.018529f
C15905 VDD.n1284 VSS 0.011881f
C15906 VDD.n1285 VSS 0.011881f
C15907 VDD.n1286 VSS 0.011881f
C15908 VDD.n1288 VSS 0.01365f
C15909 VDD.n1289 VSS 0.01214f
C15910 VDD.n1291 VSS 0.011881f
C15911 VDD.n1292 VSS 0.011881f
C15912 VDD.n1293 VSS 0.011881f
C15913 VDD.n1297 VSS 0.011881f
C15914 VDD.n1298 VSS 0.011881f
C15915 VDD.n1299 VSS 0.011881f
C15916 VDD.n1301 VSS 0.024375f
C15917 VDD.n1302 VSS 0.013273f
C15918 VDD.n1304 VSS 0.015937f
C15919 VDD.n1305 VSS 0.022225f
C15920 VDD.n1306 VSS 0.011881f
C15921 VDD.n1307 VSS 0.011881f
C15922 VDD.n1308 VSS 0.011881f
C15923 VDD.n1310 VSS 0.024168f
C15924 VDD.n1312 VSS 0.011881f
C15925 VDD.n1313 VSS 0.011881f
C15926 VDD.n1314 VSS 0.011881f
C15927 VDD.n1320 VSS 0.011881f
C15928 VDD.n1321 VSS 0.011881f
C15929 VDD.n1322 VSS 0.011881f
C15930 VDD.n1324 VSS 0.022164f
C15931 VDD.n1325 VSS 0.012976f
C15932 VDD.n1326 VSS 0.011958f
C15933 VDD.n1328 VSS 0.011881f
C15934 VDD.n1329 VSS 0.011881f
C15935 VDD.n1330 VSS 0.011881f
C15936 VDD.n1332 VSS 0.017982f
C15937 VDD.n1334 VSS 0.013629f
C15938 VDD.n1336 VSS 0.011881f
C15939 VDD.n1337 VSS 0.011881f
C15940 VDD.n1338 VSS 0.011881f
C15941 VDD.n1341 VSS 0.014169f
C15942 VDD.n1343 VSS 0.011881f
C15943 VDD.n1344 VSS 0.011881f
C15944 VDD.n1348 VSS 0.015655f
C15945 VDD.n1349 VSS 0.011881f
C15946 VDD.n1350 VSS 0.011881f
C15947 VDD.n1354 VSS 0.017774f
C15948 VDD.n1355 VSS 0.011881f
C15949 VDD.n1356 VSS 0.011881f
C15950 VDD.n1357 VSS 0.011881f
C15951 VDD.n1359 VSS 0.011881f
C15952 VDD.n1360 VSS 0.013668f
C15953 VDD.t697 VSS 0.013828f
C15954 VDD.t3708 VSS 0.014421f
C15955 VDD.n1361 VSS 0.011881f
C15956 VDD.t274 VSS 0.014745f
C15957 VDD.t3723 VSS 0.014207f
C15958 VDD.n1362 VSS 0.015995f
C15959 VDD.n1363 VSS 0.011881f
C15960 VDD.n1364 VSS 0.010534f
C15961 VDD.n1365 VSS 0.010684f
C15962 VDD.n1366 VSS 0.016863f
C15963 VDD.n1367 VSS 0.011881f
C15964 VDD.n1368 VSS 0.013668f
C15965 VDD.n1369 VSS 0.018003f
C15966 VDD.n1370 VSS 0.011881f
C15967 VDD.t982 VSS 0.014745f
C15968 VDD.n1371 VSS 0.013668f
C15969 VDD.n1372 VSS 0.017706f
C15970 VDD.t3442 VSS 0.012563f
C15971 VDD.n1373 VSS 0.012671f
C15972 VDD.n1375 VSS 0.011881f
C15973 VDD.n1376 VSS 0.011881f
C15974 VDD.n1378 VSS 0.020336f
C15975 VDD.n1379 VSS 0.019551f
C15976 VDD.n1380 VSS 0.011881f
C15977 VDD.n1381 VSS 0.011881f
C15978 VDD.n1382 VSS 0.011881f
C15979 VDD.n1384 VSS 0.021015f
C15980 VDD.n1386 VSS 0.011881f
C15981 VDD.n1387 VSS 0.011881f
C15982 VDD.n1388 VSS 0.011881f
C15983 VDD.n1391 VSS 0.013629f
C15984 VDD.n1393 VSS 0.011881f
C15985 VDD.n1394 VSS 0.011881f
C15986 VDD.n1396 VSS 0.032809f
C15987 VDD.n1397 VSS 0.017907f
C15988 VDD.n1398 VSS 0.017728f
C15989 VDD.n1399 VSS 0.011881f
C15990 VDD.n1400 VSS 0.011881f
C15991 VDD.n1401 VSS 0.011881f
C15992 VDD.n1403 VSS 0.044136f
C15993 VDD.n1404 VSS 0.119717f
C15994 VDD.t2500 VSS 0.085275f
C15995 VDD.t976 VSS 0.035023f
C15996 VDD.t269 VSS 0.031978f
C15997 VDD.t696 VSS 0.036166f
C15998 VDD.t271 VSS 0.039211f
C15999 VDD.t273 VSS 0.069666f
C16000 VDD.t3707 VSS 0.069666f
C16001 VDD.t3722 VSS 0.035404f
C16002 VDD.t786 VSS 0.040734f
C16003 VDD.t688 VSS 0.073473f
C16004 VDD.t2765 VSS 0.063575f
C16005 VDD.t785 VSS 0.031597f
C16006 VDD.t591 VSS 0.041495f
C16007 VDD.t692 VSS 0.067382f
C16008 VDD.t2990 VSS 0.036166f
C16009 VDD.t2994 VSS 0.033501f
C16010 VDD.t590 VSS 0.065479f
C16011 VDD.t3545 VSS 0.07157f
C16012 VDD.t3714 VSS 0.036166f
C16013 VDD.t983 VSS 0.034643f
C16014 VDD.t981 VSS 0.068905f
C16015 VDD.t3711 VSS 0.068905f
C16016 VDD.t1904 VSS 0.035023f
C16017 VDD.t2203 VSS 0.039211f
C16018 VDD.t773 VSS 0.067763f
C16019 VDD.t3441 VSS 0.031978f
C16020 VDD.t771 VSS 0.035785f
C16021 VDD.t2096 VSS 0.070428f
C16022 VDD.t584 VSS 0.036546f
C16023 VDD.t3450 VSS 0.033501f
C16024 VDD.t1905 VSS 0.086797f
C16025 VDD.t818 VSS 0.070808f
C16026 VDD.t1919 VSS 0.031978f
C16027 VDD.t816 VSS 0.035785f
C16028 VDD.t2100 VSS 0.031978f
C16029 VDD.t814 VSS 0.035023f
C16030 VDD.t1451 VSS 0.031978f
C16031 VDD.t812 VSS 0.053297f
C16032 VDD.t200 VSS 0.222704f
C16033 VDD.t925 VSS 0.120679f
C16034 VDD.t927 VSS 0.068144f
C16035 VDD.t1981 VSS 0.108116f
C16036 VDD.t2449 VSS 0.103928f
C16037 VDD.t2447 VSS 0.068144f
C16038 VDD.t1985 VSS 0.107735f
C16039 VDD.t3747 VSS 0.07195f
C16040 VDD.t311 VSS 0.031978f
C16041 VDD.t1322 VSS 0.031978f
C16042 VDD.t313 VSS 0.036546f
C16043 VDD.t3053 VSS 0.101264f
C16044 VDD.t586 VSS 0.07195f
C16045 VDD.t898 VSS 0.035023f
C16046 VDD.t2773 VSS 0.031978f
C16047 VDD.t900 VSS 0.037688f
C16048 VDD.t1320 VSS 0.036166f
C16049 VDD.t43 VSS 0.053297f
C16050 VDD.t1324 VSS 0.087939f
C16051 VDD.t3363 VSS 0.055961f
C16052 VDD.t1935 VSS 0.0552f
C16053 VDD.t2496 VSS 0.055961f
C16054 VDD.t1263 VSS 0.031978f
C16055 VDD.t2498 VSS 0.037688f
C16056 VDD.t1321 VSS 0.058246f
C16057 VDD.t2774 VSS 0.046063f
C16058 VDD.t2551 VSS 0.031978f
C16059 VDD.t820 VSS 0.036166f
C16060 VDD.t2555 VSS 0.041114f
C16061 VDD.t3373 VSS 0.031978f
C16062 VDD.t2553 VSS 0.031978f
C16063 VDD.t1326 VSS 0.053677f
C16064 VDD.n1405 VSS 0.080433f
C16065 VDD.t2554 VSS 0.014469f
C16066 VDD.n1407 VSS 0.011881f
C16067 VDD.n1408 VSS 0.011881f
C16068 VDD.n1409 VSS 0.013668f
C16069 VDD.t2499 VSS 0.012738f
C16070 VDD.n1410 VSS 0.014651f
C16071 VDD.n1411 VSS 0.011881f
C16072 VDD.t1264 VSS 0.010806f
C16073 VDD.n1414 VSS 0.011101f
C16074 VDD.n1415 VSS 0.011881f
C16075 VDD.n1416 VSS 0.011881f
C16076 VDD.n1417 VSS 0.013668f
C16077 VDD.n1419 VSS 0.011881f
C16078 VDD.t899 VSS 0.014469f
C16079 VDD.n1420 VSS 0.016313f
C16080 VDD.n1422 VSS 0.013668f
C16081 VDD.n1424 VSS 0.011881f
C16082 VDD.n1425 VSS 0.011881f
C16083 VDD.t312 VSS 0.014745f
C16084 VDD.n1426 VSS 0.013668f
C16085 VDD.n1427 VSS 0.013668f
C16086 VDD.n1428 VSS 0.03134f
C16087 VDD.n1429 VSS 0.011881f
C16088 VDD.t2825 VSS 0.014745f
C16089 VDD.t2450 VSS 0.014745f
C16090 VDD.n1430 VSS 0.013668f
C16091 VDD.n1431 VSS 0.013668f
C16092 VDD.n1432 VSS 0.03134f
C16093 VDD.t201 VSS 0.010137f
C16094 VDD.t3808 VSS 0.021516f
C16095 VDD.n1434 VSS 0.055166f
C16096 VDD.t202 VSS 0.010137f
C16097 VDD.n1435 VSS 0.030049f
C16098 VDD.t208 VSS 0.010137f
C16099 VDD.t3814 VSS 0.021516f
C16100 VDD.n1437 VSS 0.055166f
C16101 VDD.t209 VSS 0.010137f
C16102 VDD.n1438 VSS 0.030049f
C16103 VDD.n1439 VSS 0.02678f
C16104 VDD.t1357 VSS 0.014745f
C16105 VDD.t926 VSS 0.014745f
C16106 VDD.n1441 VSS 0.035938f
C16107 VDD.n1443 VSS 0.053216f
C16108 VDD.n1444 VSS 0.011881f
C16109 VDD.n1445 VSS 0.011881f
C16110 VDD.n1447 VSS 0.036601f
C16111 VDD.n1449 VSS 0.011881f
C16112 VDD.n1450 VSS 0.011881f
C16113 VDD.n1451 VSS 0.011881f
C16114 VDD.n1453 VSS 0.020199f
C16115 VDD.n1454 VSS 0.012941f
C16116 VDD.n1455 VSS 0.01782f
C16117 VDD.n1457 VSS 0.011881f
C16118 VDD.n1458 VSS 0.011881f
C16119 VDD.n1459 VSS 0.011881f
C16120 VDD.n1461 VSS 0.018529f
C16121 VDD.n1464 VSS 0.011881f
C16122 VDD.n1465 VSS 0.011881f
C16123 VDD.n1467 VSS 0.016801f
C16124 VDD.n1468 VSS 0.012208f
C16125 VDD.n1470 VSS 0.011881f
C16126 VDD.n1471 VSS 0.011881f
C16127 VDD.n1472 VSS 0.011881f
C16128 VDD.n1474 VSS 0.01766f
C16129 VDD.n1475 VSS 0.010471f
C16130 VDD.n1477 VSS 0.017182f
C16131 VDD.n1479 VSS 0.022477f
C16132 VDD.n1480 VSS 0.011881f
C16133 VDD.n1481 VSS 0.011881f
C16134 VDD.n1483 VSS 0.014405f
C16135 VDD.n1486 VSS 0.011402f
C16136 VDD.n1487 VSS 0.011881f
C16137 VDD.n1497 VSS 0.014542f
C16138 VDD.n1503 VSS 0.778377f
C16139 VDD.t1124 VSS 0.014745f
C16140 VDD.t550 VSS 0.015994f
C16141 VDD.n1510 VSS 0.010205f
C16142 VDD.n1512 VSS 0.011881f
C16143 VDD.t2643 VSS 0.013611f
C16144 VDD.n1515 VSS 0.015838f
C16145 VDD.n1516 VSS 0.011881f
C16146 VDD.t546 VSS 0.013927f
C16147 VDD.t3690 VSS 0.054439f
C16148 VDD.n1518 VSS 0.011881f
C16149 VDD.t3536 VSS 0.012728f
C16150 VDD.n1520 VSS 0.011881f
C16151 VDD.t3254 VSS 0.014121f
C16152 VDD.n1521 VSS 0.020948f
C16153 VDD.n1522 VSS 0.011881f
C16154 VDD.n1524 VSS 0.01373f
C16155 VDD.n1525 VSS 0.011881f
C16156 VDD.t3540 VSS 0.014219f
C16157 VDD.t3003 VSS 0.013964f
C16158 VDD.n1526 VSS 0.017492f
C16159 VDD.n1527 VSS 0.011881f
C16160 VDD.n1529 VSS 0.011881f
C16161 VDD.t2910 VSS 0.014477f
C16162 VDD.n1530 VSS 0.017738f
C16163 VDD.n1531 VSS 0.011881f
C16164 VDD.n1532 VSS 0.024012f
C16165 VDD.t3005 VSS 0.014477f
C16166 VDD.n1533 VSS 0.011881f
C16167 VDD.t3010 VSS 0.01447f
C16168 VDD.t3544 VSS 0.014304f
C16169 VDD.t158 VSS 0.010137f
C16170 VDD.t3781 VSS 0.021516f
C16171 VDD.n1536 VSS 0.055166f
C16172 VDD.t159 VSS 0.010137f
C16173 VDD.n1537 VSS 0.030049f
C16174 VDD.n1538 VSS 0.040326f
C16175 VDD.n1539 VSS 0.011881f
C16176 VDD.t1503 VSS 0.01447f
C16177 VDD.t1508 VSS 0.014207f
C16178 VDD.n1540 VSS 0.010451f
C16179 VDD.n1541 VSS 0.015706f
C16180 VDD.n1542 VSS 0.011881f
C16181 VDD.n1543 VSS 0.011881f
C16182 VDD.t1501 VSS 0.014485f
C16183 VDD.n1544 VSS 0.011881f
C16184 VDD.t1108 VSS 0.014485f
C16185 VDD.t1816 VSS 0.01449f
C16186 VDD.n1545 VSS 0.021272f
C16187 VDD.n1546 VSS 0.011881f
C16188 VDD.t3525 VSS 0.012728f
C16189 VDD.n1549 VSS 0.011881f
C16190 VDD.n1550 VSS 0.011058f
C16191 VDD.n1551 VSS 0.011881f
C16192 VDD.t52 VSS 0.013749f
C16193 VDD.n1553 VSS 0.014257f
C16194 VDD.n1554 VSS 0.011881f
C16195 VDD.t1605 VSS 0.010846f
C16196 VDD.n1556 VSS 0.015301f
C16197 VDD.n1557 VSS 0.011881f
C16198 VDD.t3284 VSS 0.053297f
C16199 VDD.n1559 VSS 0.010783f
C16200 VDD.n1560 VSS 0.015937f
C16201 VDD.n1561 VSS 0.011881f
C16202 VDD.t1110 VSS 0.012563f
C16203 VDD.n1562 VSS 0.014135f
C16204 VDD.n1563 VSS 0.011881f
C16205 VDD.n1565 VSS 0.017313f
C16206 VDD.n1566 VSS 0.011881f
C16207 VDD.n1568 VSS 0.011881f
C16208 VDD.n1569 VSS 0.012923f
C16209 VDD.t1043 VSS 0.015653f
C16210 VDD.n1570 VSS 0.01048f
C16211 VDD.t1868 VSS 0.014504f
C16212 VDD.n1571 VSS 0.011881f
C16213 VDD.t3041 VSS 0.015885f
C16214 VDD.n1572 VSS 0.037012f
C16215 VDD.n1573 VSS 0.011881f
C16216 VDD.t3812 VSS 0.074403f
C16217 VDD.t2750 VSS 0.012931f
C16218 VDD.t170 VSS 0.010055f
C16219 VDD.n1574 VSS 0.01771f
C16220 VDD.n1575 VSS 0.019845f
C16221 VDD.n1576 VSS 0.024263f
C16222 VDD.n1577 VSS 0.011881f
C16223 VDD.n1578 VSS 0.010911f
C16224 VDD.n1579 VSS 0.019199f
C16225 VDD.n1580 VSS 0.011881f
C16226 VDD.n1581 VSS 0.011147f
C16227 VDD.n1582 VSS 0.012614f
C16228 VDD.t89 VSS 0.010055f
C16229 VDD.t3799 VSS 0.042335f
C16230 VDD.n1584 VSS 0.073549f
C16231 VDD.t90 VSS 0.010055f
C16232 VDD.n1585 VSS 0.042203f
C16233 VDD.n1586 VSS 0.026958f
C16234 VDD.n1587 VSS 0.011881f
C16235 VDD.n1588 VSS 0.012073f
C16236 VDD.n1589 VSS 0.011881f
C16237 VDD.n1592 VSS 0.019778f
C16238 VDD.t1483 VSS 0.014485f
C16239 VDD.n1593 VSS 0.012976f
C16240 VDD.t1002 VSS 0.01449f
C16241 VDD.n1594 VSS 0.0215f
C16242 VDD.n1595 VSS 0.011881f
C16243 VDD.t1390 VSS 0.014485f
C16244 VDD.n1596 VSS 0.012233f
C16245 VDD.t2864 VSS 0.014481f
C16246 VDD.t758 VSS 0.035785f
C16247 VDD.t3270 VSS 0.031978f
C16248 VDD.t2625 VSS 0.036546f
C16249 VDD.t962 VSS 0.044921f
C16250 VDD.t308 VSS 0.062433f
C16251 VDD.t1109 VSS 0.061672f
C16252 VDD.t3460 VSS 0.070808f
C16253 VDD.t1549 VSS 0.084513f
C16254 VDD.t2721 VSS 0.081468f
C16255 VDD.t1807 VSS 0.068524f
C16256 VDD.t1823 VSS 0.077661f
C16257 VDD.t1146 VSS 0.043399f
C16258 VDD.t307 VSS 0.034262f
C16259 VDD.t1258 VSS 0.03883f
C16260 VDD.t518 VSS 0.031978f
C16261 VDD.t3306 VSS 0.042637f
C16262 VDD.t1042 VSS 0.036927f
C16263 VDD.t527 VSS 0.073854f
C16264 VDD.t1867 VSS 0.086417f
C16265 VDD.t1257 VSS 0.063956f
C16266 VDD.t1145 VSS 0.103167f
C16267 VDD.t3040 VSS 0.075377f
C16268 VDD.t169 VSS 0.109639f
C16269 VDD.t2749 VSS 0.137429f
C16270 VDD.t523 VSS 0.068905f
C16271 VDD.t3308 VSS 0.0552f
C16272 VDD.t79 VSS 0.112684f
C16273 VDD.t3261 VSS 0.10507f
C16274 VDD.n1597 VSS 0.033972f
C16275 VDD.t2960 VSS 0.06624f
C16276 VDD.t1040 VSS 0.090604f
C16277 VDD.t2935 VSS 0.081848f
C16278 VDD.t3320 VSS 0.072712f
C16279 VDD.t3278 VSS 0.068905f
C16280 VDD.t3182 VSS 0.08261f
C16281 VDD.t166 VSS 0.11573f
C16282 VDD.t88 VSS 0.210902f
C16283 VDD.t1643 VSS 0.172833f
C16284 VDD.t1450 VSS 0.070047f
C16285 VDD.t3107 VSS 0.070808f
C16286 VDD.t1362 VSS 0.038069f
C16287 VDD.t253 VSS 0.035785f
C16288 VDD.t3294 VSS 0.039592f
C16289 VDD.t3620 VSS 0.035023f
C16290 VDD.t277 VSS 0.032739f
C16291 VDD.t3280 VSS 0.070047f
C16292 VDD.t2565 VSS 0.081468f
C16293 VDD.t110 VSS 0.089462f
C16294 VDD.t3630 VSS 0.08832f
C16295 VDD.t1482 VSS 0.036927f
C16296 VDD.t1360 VSS 0.031978f
C16297 VDD.t1001 VSS 0.031978f
C16298 VDD.t731 VSS 0.051774f
C16299 VDD.t803 VSS 0.053297f
C16300 VDD.t1389 VSS 0.053297f
C16301 VDD.t2863 VSS 0.051774f
C16302 VDD.n1598 VSS 0.079654f
C16303 VDD.n1599 VSS 0.011881f
C16304 VDD.t3678 VSS 0.012563f
C16305 VDD.n1601 VSS 0.011881f
C16306 VDD.n1602 VSS 0.02048f
C16307 VDD.n1603 VSS 0.015751f
C16308 VDD.n1604 VSS 0.011881f
C16309 VDD.t3223 VSS 0.013918f
C16310 VDD.n1606 VSS 0.015301f
C16311 VDD.n1607 VSS 0.011881f
C16312 VDD.n1611 VSS 0.015498f
C16313 VDD.n1612 VSS 0.011881f
C16314 VDD.n1613 VSS 0.011783f
C16315 VDD.n1616 VSS 0.012019f
C16316 VDD.n1617 VSS 0.011881f
C16317 VDD.n1620 VSS 0.011881f
C16318 VDD.n1623 VSS 0.011881f
C16319 VDD.n1625 VSS 0.012634f
C16320 VDD.n1626 VSS 0.011881f
C16321 VDD.n1628 VSS 0.011881f
C16322 VDD.t992 VSS 0.010846f
C16323 VDD.t622 VSS 0.013297f
C16324 VDD.n1629 VSS 0.011881f
C16325 VDD.t649 VSS 0.085275f
C16326 VDD.t807 VSS 0.038069f
C16327 VDD.t1302 VSS 0.045683f
C16328 VDD.t1764 VSS 0.064717f
C16329 VDD.t3677 VSS 0.032739f
C16330 VDD.t2867 VSS 0.035785f
C16331 VDD.t3300 VSS 0.063194f
C16332 VDD.t822 VSS 0.106593f
C16333 VDD.t3176 VSS 0.07195f
C16334 VDD.t3222 VSS 0.03312f
C16335 VDD.t3210 VSS 0.065479f
C16336 VDD.t3174 VSS 0.036166f
C16337 VDD.t49 VSS 0.032739f
C16338 VDD.t3206 VSS 0.031978f
C16339 VDD.t2932 VSS 0.032739f
C16340 VDD.t613 VSS 0.036166f
C16341 VDD.t3718 VSS 0.032739f
C16342 VDD.t611 VSS 0.036166f
C16343 VDD.t3 VSS 0.032739f
C16344 VDD.t623 VSS 0.055961f
C16345 VDD.t597 VSS 0.048348f
C16346 VDD.t3145 VSS 0.032739f
C16347 VDD.t625 VSS 0.031978f
C16348 VDD.t1697 VSS 0.032739f
C16349 VDD.t615 VSS 0.050632f
C16350 VDD.t603 VSS 0.065479f
C16351 VDD.t601 VSS 0.051012f
C16352 VDD.t2323 VSS 0.032359f
C16353 VDD.t617 VSS 0.035023f
C16354 VDD.t990 VSS 0.032739f
C16355 VDD.t609 VSS 0.037688f
C16356 VDD.t1699 VSS 0.032739f
C16357 VDD.t605 VSS 0.039592f
C16358 VDD.t627 VSS 0.046444f
C16359 VDD.t2644 VSS 0.032739f
C16360 VDD.t607 VSS 0.036927f
C16361 VDD.t3357 VSS 0.032739f
C16362 VDD.t599 VSS 0.047586f
C16363 VDD.t619 VSS 0.060149f
C16364 VDD.t991 VSS 0.032739f
C16365 VDD.t621 VSS 0.037688f
C16366 VDD.t1700 VSS 0.060149f
C16367 VDD.n1631 VSS 0.039301f
C16368 VDD.n1632 VSS 0.011881f
C16369 VDD.n1636 VSS 0.011881f
C16370 VDD.n1639 VSS 0.011881f
C16371 VDD.n1640 VSS 0.011881f
C16372 VDD.n1643 VSS 0.011881f
C16373 VDD.t3120 VSS 0.012563f
C16374 VDD.n1646 VSS 0.012081f
C16375 VDD.n1647 VSS 0.011881f
C16376 VDD.t1692 VSS 0.013738f
C16377 VDD.n1649 VSS 0.015846f
C16378 VDD.n1650 VSS 0.0111f
C16379 VDD.t390 VSS 0.011212f
C16380 VDD.t392 VSS 0.011298f
C16381 VDD.n1651 VSS 0.014245f
C16382 VDD.n1652 VSS 0.011881f
C16383 VDD.t747 VSS 0.014745f
C16384 VDD.n1653 VSS 0.013523f
C16385 VDD.n1654 VSS 0.015061f
C16386 VDD.n1655 VSS 0.011881f
C16387 VDD.t989 VSS 0.036927f
C16388 VDD.t299 VSS 0.073092f
C16389 VDD.t3404 VSS 0.073092f
C16390 VDD.t2646 VSS 0.053677f
C16391 VDD.t2273 VSS 0.067001f
C16392 VDD.t2380 VSS 0.052535f
C16393 VDD.t303 VSS 0.039211f
C16394 VDD.t301 VSS 0.063956f
C16395 VDD.t305 VSS 0.059007f
C16396 VDD.t1328 VSS 0.031978f
C16397 VDD.t297 VSS 0.04949f
C16398 VDD.t752 VSS 0.095553f
C16399 VDD.t1688 VSS 0.078803f
C16400 VDD.t754 VSS 0.04949f
C16401 VDD.t2519 VSS 0.031978f
C16402 VDD.t2678 VSS 0.081087f
C16403 VDD.t3119 VSS 0.087939f
C16404 VDD.t938 VSS 0.035785f
C16405 VDD.t3013 VSS 0.045302f
C16406 VDD.t830 VSS 0.035023f
C16407 VDD.t2433 VSS 0.079945f
C16408 VDD.t1691 VSS 0.106212f
C16409 VDD.t3109 VSS 0.070047f
C16410 VDD.t2758 VSS 0.041114f
C16411 VDD.t389 VSS 0.044541f
C16412 VDD.t1820 VSS 0.061291f
C16413 VDD.t391 VSS 0.02741f
C16414 VDD.t3244 VSS 0.073473f
C16415 VDD.t746 VSS 0.072712f
C16416 VDD.t2757 VSS 0.031978f
C16417 VDD.t744 VSS 0.031978f
C16418 VDD.t869 VSS 0.036166f
C16419 VDD.t714 VSS 0.085275f
C16420 VDD.n1658 VSS 0.155412f
C16421 VDD.n1659 VSS 0.011881f
C16422 VDD.n1662 VSS 0.011881f
C16423 VDD.t2940 VSS 0.013913f
C16424 VDD.n1664 VSS 0.012351f
C16425 VDD.n1665 VSS 0.011881f
C16426 VDD.n1668 VSS 0.011881f
C16427 VDD.n1669 VSS 0.011881f
C16428 VDD.t634 VSS 0.01406f
C16429 VDD.t2420 VSS 0.012673f
C16430 VDD.n1671 VSS 0.019325f
C16431 VDD.n1672 VSS 0.011881f
C16432 VDD.t3085 VSS 0.014477f
C16433 VDD.n1674 VSS 0.011881f
C16434 VDD.n1675 VSS 0.011881f
C16435 VDD.n1676 VSS 0.013668f
C16436 VDD.t3083 VSS 0.01447f
C16437 VDD.n1677 VSS 0.011881f
C16438 VDD.n1678 VSS 0.011881f
C16439 VDD.t951 VSS 0.014745f
C16440 VDD.t3191 VSS 0.014219f
C16441 VDD.n1679 VSS 0.022117f
C16442 VDD.n1680 VSS 0.011881f
C16443 VDD.n1681 VSS 0.013523f
C16444 VDD.n1682 VSS 0.011881f
C16445 VDD.t2142 VSS 0.014745f
C16446 VDD.n1683 VSS 0.013668f
C16447 VDD.n1684 VSS 0.013668f
C16448 VDD.n1685 VSS 0.03134f
C16449 VDD.n1686 VSS 0.011881f
C16450 VDD.t1275 VSS 0.014745f
C16451 VDD.t1562 VSS 0.014745f
C16452 VDD.t632 VSS 0.014399f
C16453 VDD.n1687 VSS 0.013668f
C16454 VDD.n1688 VSS 0.031565f
C16455 VDD.t91 VSS 0.222704f
C16456 VDD.t1167 VSS 0.120679f
C16457 VDD.t1169 VSS 0.068144f
C16458 VDD.t1165 VSS 0.108116f
C16459 VDD.t2532 VSS 0.072331f
C16460 VDD.t629 VSS 0.031978f
C16461 VDD.t2534 VSS 0.031978f
C16462 VDD.t631 VSS 0.036166f
C16463 VDD.t1801 VSS 0.054058f
C16464 VDD.t3339 VSS 0.127531f
C16465 VDD.t3118 VSS 0.04949f
C16466 VDD.t2667 VSS 0.032739f
C16467 VDD.t3121 VSS 0.047967f
C16468 VDD.t2062 VSS 0.065479f
C16469 VDD.t2065 VSS 0.050251f
C16470 VDD.t2187 VSS 0.062814f
C16471 VDD.t1539 VSS 0.054819f
C16472 VDD.t2939 VSS 0.042257f
C16473 VDD.t2926 VSS 0.065479f
C16474 VDD.t635 VSS 0.037688f
C16475 VDD.t1598 VSS 0.032739f
C16476 VDD.t633 VSS 0.037308f
C16477 VDD.t2417 VSS 0.043018f
C16478 VDD.t2928 VSS 0.067763f
C16479 VDD.t1137 VSS 0.067763f
C16480 VDD.t2419 VSS 0.10507f
C16481 VDD.t2031 VSS 0.072331f
C16482 VDD.t3084 VSS 0.032739f
C16483 VDD.t3082 VSS 0.035404f
C16484 VDD.t948 VSS 0.035404f
C16485 VDD.t950 VSS 0.068905f
C16486 VDD.t2950 VSS 0.064337f
C16487 VDD.t3190 VSS 0.035023f
C16488 VDD.t2041 VSS 0.043779f
C16489 VDD.t2143 VSS 0.068144f
C16490 VDD.t2141 VSS 0.103928f
C16491 VDD.t2029 VSS 0.108116f
C16492 VDD.t1276 VSS 0.068144f
C16493 VDD.t1274 VSS 0.085655f
C16494 VDD.n1689 VSS 0.078512f
C16495 VDD.n1690 VSS 0.011881f
C16496 VDD.t630 VSS 0.014204f
C16497 VDD.t2533 VSS 0.014469f
C16498 VDD.n1691 VSS 0.013668f
C16499 VDD.n1692 VSS 0.013668f
C16500 VDD.n1693 VSS 0.03134f
C16501 VDD.t122 VSS 0.010137f
C16502 VDD.t3791 VSS 0.021516f
C16503 VDD.n1695 VSS 0.055166f
C16504 VDD.t123 VSS 0.010137f
C16505 VDD.n1696 VSS 0.030049f
C16506 VDD.t92 VSS 0.010137f
C16507 VDD.t3782 VSS 0.021516f
C16508 VDD.n1698 VSS 0.055166f
C16509 VDD.t93 VSS 0.010137f
C16510 VDD.n1699 VSS 0.030049f
C16511 VDD.n1700 VSS 0.02678f
C16512 VDD.t1168 VSS 0.014745f
C16513 VDD.t2432 VSS 0.014745f
C16514 VDD.n1702 VSS 0.035938f
C16515 VDD.n1704 VSS 0.053216f
C16516 VDD.n1705 VSS 0.011881f
C16517 VDD.n1706 VSS 0.011881f
C16518 VDD.n1708 VSS 0.017982f
C16519 VDD.n1710 VSS 0.014772f
C16520 VDD.n1712 VSS 0.011881f
C16521 VDD.n1713 VSS 0.011881f
C16522 VDD.n1714 VSS 0.011881f
C16523 VDD.n1715 VSS 0.02392f
C16524 VDD.n1716 VSS 0.035938f
C16525 VDD.n1718 VSS 0.011881f
C16526 VDD.n1719 VSS 0.011881f
C16527 VDD.n1720 VSS 0.011881f
C16528 VDD.n1722 VSS 0.020999f
C16529 VDD.n1724 VSS 0.015061f
C16530 VDD.n1726 VSS 0.011881f
C16531 VDD.n1727 VSS 0.011881f
C16532 VDD.n1729 VSS 0.02061f
C16533 VDD.n1730 VSS 0.016107f
C16534 VDD.n1731 VSS 0.017385f
C16535 VDD.n1732 VSS 0.018287f
C16536 VDD.n1734 VSS 0.016181f
C16537 VDD.n1735 VSS 0.011881f
C16538 VDD.n1736 VSS 0.011881f
C16539 VDD.n1738 VSS 0.014651f
C16540 VDD.n1739 VSS 0.012222f
C16541 VDD.n1740 VSS 0.013667f
C16542 VDD.n1742 VSS 0.011881f
C16543 VDD.n1743 VSS 0.011881f
C16544 VDD.n1748 VSS 0.011881f
C16545 VDD.n1749 VSS 0.011881f
C16546 VDD.n1750 VSS 0.011881f
C16547 VDD.n1752 VSS 0.013584f
C16548 VDD.n1754 VSS 0.011881f
C16549 VDD.n1755 VSS 0.011881f
C16550 VDD.n1756 VSS 0.011881f
C16551 VDD.n1757 VSS 0.025155f
C16552 VDD.n1761 VSS 0.011881f
C16553 VDD.n1762 VSS 0.011881f
C16554 VDD.n1764 VSS 0.020999f
C16555 VDD.n1766 VSS 0.045024f
C16556 VDD.n1767 VSS 0.015831f
C16557 VDD.n1768 VSS 0.015846f
C16558 VDD.n1769 VSS 0.011881f
C16559 VDD.n1771 VSS 0.018754f
C16560 VDD.n1773 VSS 0.011881f
C16561 VDD.n1774 VSS 0.011881f
C16562 VDD.n1778 VSS 0.014135f
C16563 VDD.n1779 VSS 0.011881f
C16564 VDD.n1780 VSS 0.011881f
C16565 VDD.n1781 VSS 0.011881f
C16566 VDD.n1783 VSS 0.013584f
C16567 VDD.t298 VSS 0.015994f
C16568 VDD.n1789 VSS 0.011881f
C16569 VDD.n1790 VSS 0.011881f
C16570 VDD.n1791 VSS 0.011881f
C16571 VDD.t304 VSS 0.013927f
C16572 VDD.n1795 VSS 0.011406f
C16573 VDD.n1797 VSS 0.011881f
C16574 VDD.n1798 VSS 0.011881f
C16575 VDD.n1802 VSS 0.011385f
C16576 VDD.n1803 VSS 0.011881f
C16577 VDD.n1804 VSS 0.011881f
C16578 VDD.n1805 VSS 0.011881f
C16579 VDD.n1806 VSS 0.024904f
C16580 VDD.n1807 VSS 0.016404f
C16581 VDD.n1808 VSS 0.014638f
C16582 VDD.n1809 VSS 0.013577f
C16583 VDD.n1813 VSS 0.011881f
C16584 VDD.n1814 VSS 0.011881f
C16585 VDD.n1815 VSS 0.011881f
C16586 VDD.n1817 VSS 0.014724f
C16587 VDD.n1819 VSS 0.01148f
C16588 VDD.n1821 VSS 0.011881f
C16589 VDD.n1822 VSS 0.011881f
C16590 VDD.n1824 VSS 0.013213f
C16591 VDD.n1829 VSS 0.011881f
C16592 VDD.n1830 VSS 0.011881f
C16593 VDD.n1833 VSS 0.012649f
C16594 VDD.n1834 VSS 0.010467f
C16595 VDD.n1835 VSS 0.011881f
C16596 VDD.n1836 VSS 0.011881f
C16597 VDD.n1837 VSS 0.011881f
C16598 VDD.n1839 VSS 0.021048f
C16599 VDD.n1841 VSS 0.012875f
C16600 VDD.n1843 VSS 0.011881f
C16601 VDD.n1844 VSS 0.011881f
C16602 VDD.n1848 VSS 0.012081f
C16603 VDD.n1850 VSS 0.011881f
C16604 VDD.n1851 VSS 0.011881f
C16605 VDD.n1853 VSS 0.013015f
C16606 VDD.n1854 VSS 0.01741f
C16607 VDD.n1856 VSS 0.011881f
C16608 VDD.n1857 VSS 0.011881f
C16609 VDD.n1858 VSS 0.011881f
C16610 VDD.n1859 VSS 0.041199f
C16611 VDD.n1861 VSS 0.020187f
C16612 VDD.n1862 VSS 0.011881f
C16613 VDD.n1863 VSS 0.011881f
C16614 VDD.n1864 VSS 0.011881f
C16615 VDD.n1866 VSS 0.011958f
C16616 VDD.n1867 VSS 0.018655f
C16617 VDD.t111 VSS 0.010137f
C16618 VDD.t3778 VSS 0.021516f
C16619 VDD.n1869 VSS 0.055166f
C16620 VDD.t112 VSS 0.010137f
C16621 VDD.n1870 VSS 0.030049f
C16622 VDD.n1871 VSS 0.02054f
C16623 VDD.n1872 VSS 0.034122f
C16624 VDD.n1873 VSS 0.019845f
C16625 VDD.n1874 VSS 0.01978f
C16626 VDD.n1875 VSS 0.011881f
C16627 VDD.n1876 VSS 0.014062f
C16628 VDD.n1878 VSS 0.01709f
C16629 VDD.t1363 VSS 0.012563f
C16630 VDD.n1879 VSS 0.012854f
C16631 VDD.n1880 VSS 0.011881f
C16632 VDD.n1881 VSS 0.011881f
C16633 VDD.n1882 VSS 0.011881f
C16634 VDD.t167 VSS 0.011064f
C16635 VDD.t3774 VSS 0.147089f
C16636 VDD.n1886 VSS 0.1075f
C16637 VDD.n1887 VSS 0.012126f
C16638 VDD.n1888 VSS 0.023669f
C16639 VDD.n1889 VSS 0.023938f
C16640 VDD.n1890 VSS 0.023677f
C16641 VDD.n1891 VSS 0.011881f
C16642 VDD.n1893 VSS 0.021342f
C16643 VDD.n1894 VSS 0.012614f
C16644 VDD.n1895 VSS 0.010172f
C16645 VDD.n1896 VSS 0.011881f
C16646 VDD.n1897 VSS 0.011881f
C16647 VDD.n1898 VSS 0.0118f
C16648 VDD.t168 VSS 0.011064f
C16649 VDD.t1041 VSS 0.014825f
C16650 VDD.n1901 VSS 0.013358f
C16651 VDD.n1903 VSS 0.011881f
C16652 VDD.n1904 VSS 0.011881f
C16653 VDD.n1905 VSS 0.01978f
C16654 VDD.t3262 VSS 0.0145f
C16655 VDD.n1906 VSS 0.024123f
C16656 VDD.n1907 VSS 0.010433f
C16657 VDD.t80 VSS 0.010137f
C16658 VDD.t3826 VSS 0.021516f
C16659 VDD.n1909 VSS 0.055166f
C16660 VDD.t81 VSS 0.010137f
C16661 VDD.n1910 VSS 0.030049f
C16662 VDD.n1911 VSS 0.030293f
C16663 VDD.n1912 VSS 0.011038f
C16664 VDD.n1913 VSS 0.019778f
C16665 VDD.n1914 VSS 0.011881f
C16666 VDD.n1915 VSS 0.02936f
C16667 VDD.n1916 VSS 0.100348f
C16668 VDD.n1917 VSS 0.023051f
C16669 VDD.n1918 VSS 0.01661f
C16670 VDD.n1919 VSS 0.011881f
C16671 VDD.n1920 VSS 0.011881f
C16672 VDD.n1921 VSS 0.03017f
C16673 VDD.n1922 VSS 0.031187f
C16674 VDD.t171 VSS 0.010055f
C16675 VDD.n1923 VSS 0.01771f
C16676 VDD.n1924 VSS 0.03017f
C16677 VDD.n1925 VSS 0.011881f
C16678 VDD.n1926 VSS 0.011881f
C16679 VDD.n1927 VSS 0.011881f
C16680 VDD.n1928 VSS 0.026949f
C16681 VDD.n1929 VSS 0.02053f
C16682 VDD.n1930 VSS 0.011027f
C16683 VDD.n1932 VSS 0.011881f
C16684 VDD.n1933 VSS 0.011881f
C16685 VDD.n1934 VSS 0.011881f
C16686 VDD.n1938 VSS 0.011881f
C16687 VDD.n1939 VSS 0.011881f
C16688 VDD.n1940 VSS 0.011881f
C16689 VDD.n1943 VSS 0.015182f
C16690 VDD.n1945 VSS 0.011881f
C16691 VDD.n1946 VSS 0.011881f
C16692 VDD.n1947 VSS 0.011881f
C16693 VDD.n1950 VSS 0.013891f
C16694 VDD.n1952 VSS 0.011881f
C16695 VDD.n1953 VSS 0.011881f
C16696 VDD.n1954 VSS 0.013668f
C16697 VDD.n1955 VSS 0.018529f
C16698 VDD.n1956 VSS 0.011881f
C16699 VDD.n1959 VSS 0.015846f
C16700 VDD.n1961 VSS 0.011881f
C16701 VDD.n1962 VSS 0.010534f
C16702 VDD.n1963 VSS 0.02048f
C16703 VDD.n1965 VSS 0.018233f
C16704 VDD.n1966 VSS 0.011881f
C16705 VDD.n1967 VSS 0.011147f
C16706 VDD.t856 VSS 0.015994f
C16707 VDD.n1968 VSS 0.010205f
C16708 VDD.n1969 VSS 0.011881f
C16709 VDD.n1972 VSS 0.011881f
C16710 VDD.t860 VSS 0.013927f
C16711 VDD.n1973 VSS 0.011863f
C16712 VDD.t743 VSS 0.013749f
C16713 VDD.n1975 VSS 0.01849f
C16714 VDD.n1976 VSS 0.011881f
C16715 VDD.n1977 VSS 0.011881f
C16716 VDD.n1979 VSS 0.010585f
C16717 VDD.n1982 VSS 0.012954f
C16718 VDD.n1984 VSS 0.011881f
C16719 VDD.n1985 VSS 0.011881f
C16720 VDD.n1986 VSS 0.011881f
C16721 VDD.n1990 VSS 0.011062f
C16722 VDD.n1991 VSS 0.014972f
C16723 VDD.n1993 VSS 0.011881f
C16724 VDD.n1994 VSS 0.011881f
C16725 VDD.n1996 VSS 0.01596f
C16726 VDD.n2000 VSS 0.011881f
C16727 VDD.n2001 VSS 0.011881f
C16728 VDD.n2002 VSS 0.011881f
C16729 VDD.n2005 VSS 0.015637f
C16730 VDD.n2006 VSS 0.011845f
C16731 VDD.n2008 VSS 0.011881f
C16732 VDD.n2009 VSS 0.015846f
C16733 VDD.n2010 VSS 0.015831f
C16734 VDD.n2012 VSS 0.034569f
C16735 VDD.t3491 VSS 0.013966f
C16736 VDD.n2014 VSS 0.015084f
C16737 VDD.n2015 VSS 0.026608f
C16738 VDD.n2016 VSS 0.011881f
C16739 VDD.n2017 VSS 0.011881f
C16740 VDD.n2018 VSS 0.011881f
C16741 VDD.n2019 VSS 0.011533f
C16742 VDD.t897 VSS 0.014745f
C16743 VDD.n2020 VSS 0.020107f
C16744 VDD.n2022 VSS 0.011881f
C16745 VDD.n2023 VSS 0.011881f
C16746 VDD.n2024 VSS 0.011881f
C16747 VDD.n2026 VSS 0.022225f
C16748 VDD.n2027 VSS 0.043887f
C16749 VDD.t295 VSS 0.053297f
C16750 VDD.t1859 VSS 0.072331f
C16751 VDD.t1297 VSS 0.036166f
C16752 VDD.t894 VSS 0.032739f
C16753 VDD.t896 VSS 0.034262f
C16754 VDD.t3686 VSS 0.035023f
C16755 VDD.t3267 VSS 0.065479f
C16756 VDD.t756 VSS 0.07195f
C16757 VDD.t2439 VSS 0.072331f
C16758 VDD.t3490 VSS 0.036166f
C16759 VDD.t2986 VSS 0.03845f
C16760 VDD.t2911 VSS 0.067382f
C16761 VDD.t1813 VSS 0.103548f
C16762 VDD.t2755 VSS 0.073092f
C16763 VDD.t2277 VSS 0.03883f
C16764 VDD.t1103 VSS 0.061672f
C16765 VDD.t1925 VSS 0.036546f
C16766 VDD.t2895 VSS 0.032739f
C16767 VDD.t3720 VSS 0.02741f
C16768 VDD.t1261 VSS 0.039592f
C16769 VDD.t3448 VSS 0.070808f
C16770 VDD.t513 VSS 0.04949f
C16771 VDD.t1809 VSS 0.048348f
C16772 VDD.t1101 VSS 0.068905f
C16773 VDD.t521 VSS 0.039972f
C16774 VDD.t855 VSS 0.039972f
C16775 VDD.t857 VSS 0.032739f
C16776 VDD.t2820 VSS 0.031978f
C16777 VDD.t861 VSS 0.063194f
C16778 VDD.t859 VSS 0.06053f
C16779 VDD.t2145 VSS 0.061291f
C16780 VDD.t740 VSS 0.045683f
C16781 VDD.t1183 VSS 0.032359f
C16782 VDD.t1818 VSS 0.031978f
C16783 VDD.t3397 VSS 0.053677f
C16784 VDD.t863 VSS 0.059007f
C16785 VDD.t742 VSS 0.031978f
C16786 VDD.t2331 VSS 0.046825f
C16787 VDD.t2438 VSS 0.039972f
C16788 VDD.t1161 VSS 0.073854f
C16789 VDD.t3248 VSS 0.07195f
C16790 VDD.t3535 VSS 0.070047f
C16791 VDD.t828 VSS 0.065479f
C16792 VDD.t3246 VSS 0.038069f
C16793 VDD.t2138 VSS 0.038069f
C16794 VDD.t2250 VSS 0.063956f
C16795 VDD.t2801 VSS 0.10469f
C16796 VDD.t3253 VSS 0.095173f
C16797 VDD.t1269 VSS 0.032739f
C16798 VDD.t2140 VSS 0.036927f
C16799 VDD.t1304 VSS 0.032739f
C16800 VDD.t2139 VSS 0.02741f
C16801 VDD.t655 VSS 0.038069f
C16802 VDD.t3255 VSS 0.052535f
C16803 VDD.t3048 VSS 0.068524f
C16804 VDD.t3036 VSS 0.034643f
C16805 VDD.t1306 VSS 0.029313f
C16806 VDD.t3539 VSS 0.071189f
C16807 VDD.t3002 VSS 0.076519f
C16808 VDD.t652 VSS 0.034262f
C16809 VDD.t2371 VSS 0.032739f
C16810 VDD.t653 VSS 0.069286f
C16811 VDD.t3000 VSS 0.041114f
C16812 VDD.t324 VSS 0.035785f
C16813 VDD.t2914 VSS 0.065479f
C16814 VDD.t3038 VSS 0.067763f
C16815 VDD.t3528 VSS 0.07195f
C16816 VDD.t1425 VSS 0.068905f
C16817 VDD.t2712 VSS 0.035785f
C16818 VDD.t2909 VSS 0.035785f
C16819 VDD.t2916 VSS 0.10507f
C16820 VDD.t3004 VSS 0.089081f
C16821 VDD.n2028 VSS 0.03854f
C16822 VDD.t3009 VSS 0.053297f
C16823 VDD.t1223 VSS 0.070808f
C16824 VDD.t3428 VSS 0.111161f
C16825 VDD.t3543 VSS 0.08832f
C16826 VDD.t157 VSS 0.02741f
C16827 VDD.t2307 VSS 0.089081f
C16828 VDD.t1502 VSS 0.087178f
C16829 VDD.t853 VSS 0.031978f
C16830 VDD.t1507 VSS 0.02741f
C16831 VDD.t3682 VSS 0.047206f
C16832 VDD.t1149 VSS 0.063575f
C16833 VDD.t1556 VSS 0.058626f
C16834 VDD.t1500 VSS 0.068524f
C16835 VDD.t3492 VSS 0.068524f
C16836 VDD.t2794 VSS 0.035023f
C16837 VDD.t1107 VSS 0.031978f
C16838 VDD.t2280 VSS 0.031978f
C16839 VDD.t1815 VSS 0.07157f
C16840 VDD.t3524 VSS 0.073092f
C16841 VDD.t3097 VSS 0.036546f
C16842 VDD.t2436 VSS 0.067382f
C16843 VDD.t2822 VSS 0.101644f
C16844 VDD.t1490 VSS 0.073473f
C16845 VDD.t51 VSS 0.035023f
C16846 VDD.t2332 VSS 0.065479f
C16847 VDD.t2435 VSS 0.043779f
C16848 VDD.t1515 VSS 0.03845f
C16849 VDD.t3566 VSS 0.047206f
C16850 VDD.t1606 VSS 0.032739f
C16851 VDD.t3343 VSS 0.036927f
C16852 VDD.t3377 VSS 0.09403f
C16853 VDD.t1604 VSS 0.105451f
C16854 VDD.n2029 VSS 0.04425f
C16855 VDD.n2030 VSS 0.024995f
C16856 VDD.n2031 VSS 0.011881f
C16857 VDD.n2032 VSS 0.011881f
C16858 VDD.n2033 VSS 0.011881f
C16859 VDD.n2038 VSS 0.011881f
C16860 VDD.n2039 VSS 0.011881f
C16861 VDD.n2042 VSS 0.019222f
C16862 VDD.n2043 VSS 0.011881f
C16863 VDD.n2044 VSS 0.011881f
C16864 VDD.n2045 VSS 0.011881f
C16865 VDD.n2047 VSS 0.01782f
C16866 VDD.n2048 VSS 0.012895f
C16867 VDD.n2049 VSS 0.013652f
C16868 VDD.n2050 VSS 0.011881f
C16869 VDD.n2051 VSS 0.011881f
C16870 VDD.n2052 VSS 0.011881f
C16871 VDD.n2054 VSS 0.020187f
C16872 VDD.n2055 VSS 0.020187f
C16873 VDD.t1557 VSS 0.014214f
C16874 VDD.n2057 VSS 0.018324f
C16875 VDD.n2059 VSS 0.011881f
C16876 VDD.n2060 VSS 0.011881f
C16877 VDD.n2062 VSS 0.015995f
C16878 VDD.n2064 VSS 0.016907f
C16879 VDD.n2065 VSS 0.01978f
C16880 VDD.n2066 VSS 0.019845f
C16881 VDD.n2067 VSS 0.019778f
C16882 VDD.n2069 VSS 0.01814f
C16883 VDD.n2070 VSS 0.016152f
C16884 VDD.n2071 VSS 0.011881f
C16885 VDD.n2072 VSS 0.011881f
C16886 VDD.n2073 VSS 0.011881f
C16887 VDD.n2074 VSS 0.01783f
C16888 VDD.t2917 VSS 0.01447f
C16889 VDD.n2075 VSS 0.016427f
C16890 VDD.t2713 VSS 0.01449f
C16891 VDD.n2076 VSS 0.02102f
C16892 VDD.n2077 VSS 0.011881f
C16893 VDD.n2078 VSS 0.011881f
C16894 VDD.n2079 VSS 0.011881f
C16895 VDD.t1426 VSS 0.014485f
C16896 VDD.n2080 VSS 0.019753f
C16897 VDD.t3039 VSS 0.01311f
C16898 VDD.n2081 VSS 0.023876f
C16899 VDD.n2087 VSS 0.011881f
C16900 VDD.n2088 VSS 0.011881f
C16901 VDD.n2089 VSS 0.011881f
C16902 VDD.t2372 VSS 0.013966f
C16903 VDD.n2091 VSS 0.018794f
C16904 VDD.n2093 VSS 0.011881f
C16905 VDD.n2094 VSS 0.011881f
C16906 VDD.n2096 VSS 0.0215f
C16907 VDD.t3037 VSS 0.01311f
C16908 VDD.n2097 VSS 0.024402f
C16909 VDD.n2099 VSS 0.011881f
C16910 VDD.n2100 VSS 0.011881f
C16911 VDD.n2101 VSS 0.011881f
C16912 VDD.n2103 VSS 0.010601f
C16913 VDD.n2104 VSS 0.019192f
C16914 VDD.n2106 VSS 0.011881f
C16915 VDD.n2107 VSS 0.011881f
C16916 VDD.n2108 VSS 0.011881f
C16917 VDD.t3247 VSS 0.014485f
C16918 VDD.n2111 VSS 0.02085f
C16919 VDD.n2112 VSS 0.011881f
C16920 VDD.n2113 VSS 0.011881f
C16921 VDD.n2114 VSS 0.011881f
C16922 VDD.t829 VSS 0.014435f
C16923 VDD.n2115 VSS 0.031845f
C16924 VDD.n2118 VSS 0.018529f
C16925 VDD.n2119 VSS 0.011881f
C16926 VDD.n2120 VSS 0.011881f
C16927 VDD.n2121 VSS 0.011881f
C16928 VDD.n2122 VSS 0.010736f
C16929 VDD.n2123 VSS 0.016889f
C16930 VDD.n2124 VSS 0.011881f
C16931 VDD.n2125 VSS 0.011881f
C16932 VDD.t3542 VSS 0.012728f
C16933 VDD.n2127 VSS 0.014315f
C16934 VDD.n2128 VSS 0.011881f
C16935 VDD.t6 VSS 0.013749f
C16936 VDD.t2631 VSS 0.014194f
C16937 VDD.n2130 VSS 0.012328f
C16938 VDD.n2131 VSS 0.015831f
C16939 VDD.t2998 VSS 0.01383f
C16940 VDD.n2132 VSS 0.010601f
C16941 VDD.n2134 VSS 0.011881f
C16942 VDD.n2135 VSS 0.010127f
C16943 VDD.n2136 VSS 0.017108f
C16944 VDD.n2137 VSS 0.014066f
C16945 VDD.n2138 VSS 0.013523f
C16946 VDD.n2139 VSS 0.012275f
C16947 VDD.n2140 VSS 0.014169f
C16948 VDD.n2143 VSS 0.011881f
C16949 VDD.n2145 VSS 0.016065f
C16950 VDD.n2148 VSS 0.011881f
C16951 VDD.n2149 VSS 0.011881f
C16952 VDD.n2150 VSS 0.015846f
C16953 VDD.n2152 VSS 0.033361f
C16954 VDD.n2154 VSS 0.015846f
C16955 VDD.n2155 VSS 0.011881f
C16956 VDD.n2157 VSS 0.017774f
C16957 VDD.n2158 VSS 0.01785f
C16958 VDD.n2159 VSS 0.011881f
C16959 VDD.n2160 VSS 0.011881f
C16960 VDD.n2161 VSS 0.011881f
C16961 VDD.n2163 VSS 0.017733f
C16962 VDD.n2166 VSS 0.011881f
C16963 VDD.n2167 VSS 0.011881f
C16964 VDD.n2168 VSS 0.011881f
C16965 VDD.n2170 VSS 0.025155f
C16966 VDD.n2171 VSS 0.033972f
C16967 VDD.t978 VSS 0.047967f
C16968 VDD.t3550 VSS 0.073854f
C16969 VDD.t2165 VSS 0.075377f
C16970 VDD.t2493 VSS 0.070047f
C16971 VDD.t654 VSS 0.036166f
C16972 VDD.t826 VSS 0.031978f
C16973 VDD.t3523 VSS 0.032739f
C16974 VDD.t3250 VSS 0.037308f
C16975 VDD.t3507 VSS 0.066621f
C16976 VDD.t3541 VSS 0.070808f
C16977 VDD.t3006 VSS 0.037308f
C16978 VDD.t5 VSS 0.035404f
C16979 VDD.t2494 VSS 0.072331f
C16980 VDD.t2630 VSS 0.096315f
C16981 VDD.t1038 VSS 0.07157f
C16982 VDD.t2997 VSS 0.036927f
C16983 VDD.t3680 VSS 0.036166f
C16984 VDD.t1036 VSS 0.02741f
C16985 VDD.t1037 VSS 0.044921f
C16986 VDD.t3458 VSS 0.067763f
C16987 VDD.t684 VSS 0.074235f
C16988 VDD.t3518 VSS 0.07728f
C16989 VDD.t1253 VSS 0.053297f
C16990 VDD.t2741 VSS 0.031978f
C16991 VDD.t690 VSS 0.036166f
C16992 VDD.t1125 VSS 0.048348f
C16993 VDD.t1123 VSS 0.10507f
C16994 VDD.t1902 VSS 0.088701f
C16995 VDD.t549 VSS 0.032739f
C16996 VDD.t1913 VSS 0.031978f
C16997 VDD.t551 VSS 0.032359f
C16998 VDD.t2639 VSS 0.031978f
C16999 VDD.t553 VSS 0.046444f
C17000 VDD.t545 VSS 0.057103f
C17001 VDD.t2642 VSS 0.074235f
C17002 VDD.t543 VSS 0.054058f
C17003 VDD.t177 VSS 0.222704f
C17004 VDD.t287 VSS 0.120679f
C17005 VDD.t289 VSS 0.068144f
C17006 VDD.t1762 VSS 0.108116f
C17007 VDD.t2213 VSS 0.103928f
C17008 VDD.t2215 VSS 0.034643f
C17009 VDD.t3741 VSS 0.034643f
C17010 VDD.t2688 VSS 0.033501f
C17011 VDD.t3051 VSS 0.101644f
C17012 VDD.t582 VSS 0.106593f
C17013 VDD.t3745 VSS 0.035023f
C17014 VDD.t2327 VSS 0.031978f
C17015 VDD.t1600 VSS 0.037688f
C17016 VDD.t2691 VSS 0.087559f
C17017 VDD.t1453 VSS 0.067382f
C17018 VDD.t2577 VSS 0.036927f
C17019 VDD.t3369 VSS 0.035023f
C17020 VDD.t542 VSS 0.04987f
C17021 VDD.t1603 VSS 0.062814f
C17022 VDD.t2421 VSS 0.053297f
C17023 VDD.t447 VSS 0.037688f
C17024 VDD.t2690 VSS 0.036927f
C17025 VDD.t3389 VSS 0.032739f
C17026 VDD.t2328 VSS 0.037308f
C17027 VDD.t2739 VSS 0.069666f
C17028 VDD.t445 VSS 0.041114f
C17029 VDD.t3381 VSS 0.035404f
C17030 VDD.t2329 VSS 0.034262f
C17031 VDD.t1602 VSS 0.035023f
C17032 VDD.t541 VSS 0.064717f
C17033 VDD.t547 VSS 0.046825f
C17034 VDD.t2737 VSS 0.041114f
C17035 VDD.t3399 VSS 0.053297f
C17036 VDD.n2172 VSS 0.038176f
C17037 VDD.n2174 VSS 0.010585f
C17038 VDD.n2175 VSS 0.011881f
C17039 VDD.t2738 VSS 0.015916f
C17040 VDD.n2177 VSS 0.011881f
C17041 VDD.t446 VSS 0.010806f
C17042 VDD.n2180 VSS 0.01191f
C17043 VDD.t2422 VSS 0.010846f
C17044 VDD.n2182 VSS 0.015964f
C17045 VDD.n2183 VSS 0.011881f
C17046 VDD.n2185 VSS 0.011881f
C17047 VDD.n2187 VSS 0.011881f
C17048 VDD.n2190 VSS 0.011881f
C17049 VDD.n2192 VSS 0.013523f
C17050 VDD.t2214 VSS 0.014745f
C17051 VDD.n2193 VSS 0.011881f
C17052 VDD.n2194 VSS 0.013668f
C17053 VDD.n2195 VSS 0.013668f
C17054 VDD.n2196 VSS 0.03134f
C17055 VDD.t231 VSS 0.010137f
C17056 VDD.t3821 VSS 0.021516f
C17057 VDD.n2198 VSS 0.055166f
C17058 VDD.t232 VSS 0.010137f
C17059 VDD.n2199 VSS 0.030049f
C17060 VDD.t178 VSS 0.010137f
C17061 VDD.t3803 VSS 0.021516f
C17062 VDD.n2201 VSS 0.055166f
C17063 VDD.t179 VSS 0.010137f
C17064 VDD.n2202 VSS 0.030049f
C17065 VDD.n2203 VSS 0.02678f
C17066 VDD.t459 VSS 0.014745f
C17067 VDD.t288 VSS 0.014745f
C17068 VDD.n2205 VSS 0.035938f
C17069 VDD.n2207 VSS 0.053216f
C17070 VDD.n2208 VSS 0.011881f
C17071 VDD.n2209 VSS 0.011881f
C17072 VDD.n2211 VSS 0.020999f
C17073 VDD.n2213 VSS 0.015015f
C17074 VDD.n2216 VSS 0.011881f
C17075 VDD.n2217 VSS 0.011881f
C17076 VDD.n2218 VSS 0.011881f
C17077 VDD.n2220 VSS 0.011012f
C17078 VDD.n2221 VSS 0.014267f
C17079 VDD.n2222 VSS 0.011881f
C17080 VDD.n2223 VSS 0.011881f
C17081 VDD.n2224 VSS 0.011881f
C17082 VDD.n2226 VSS 0.010074f
C17083 VDD.n2227 VSS 0.010964f
C17084 VDD.n2230 VSS 0.011881f
C17085 VDD.n2231 VSS 0.011881f
C17086 VDD.n2232 VSS 0.011881f
C17087 VDD.n2234 VSS 0.011101f
C17088 VDD.n2237 VSS 0.011881f
C17089 VDD.n2238 VSS 0.011881f
C17090 VDD.n2239 VSS 0.011881f
C17091 VDD.n2241 VSS 0.010708f
C17092 VDD.n2243 VSS 0.023734f
C17093 VDD.n2244 VSS 0.011881f
C17094 VDD.n2245 VSS 0.011881f
C17095 VDD.n2246 VSS 0.011881f
C17096 VDD.n2247 VSS 0.023117f
C17097 VDD.n2250 VSS 0.011863f
C17098 VDD.n2252 VSS 0.011881f
C17099 VDD.n2253 VSS 0.011881f
C17100 VDD.n2257 VSS 0.014257f
C17101 VDD.n2268 VSS 0.020999f
C17102 VDD.n2274 VSS 0.500541f
C17103 VDD.n2284 VSS 0.011881f
C17104 VDD.n2285 VSS 0.014361f
C17105 VDD.n2286 VSS 0.011267f
C17106 VDD.n2287 VSS 0.011881f
C17107 VDD.n2288 VSS 0.013931f
C17108 VDD.n2289 VSS 0.012343f
C17109 VDD.n2290 VSS 0.011881f
C17110 VDD.t1176 VSS 0.015709f
C17111 VDD.n2291 VSS 0.020097f
C17112 VDD.t2993 VSS 0.014219f
C17113 VDD.n2292 VSS 0.022117f
C17114 VDD.n2293 VSS 0.023669f
C17115 VDD.n2295 VSS 0.025888f
C17116 VDD.t330 VSS 0.010817f
C17117 VDD.n2296 VSS 0.011881f
C17118 VDD.t3779 VSS 0.075443f
C17119 VDD.t145 VSS 0.010055f
C17120 VDD.n2297 VSS 0.126327f
C17121 VDD.n2298 VSS 0.033189f
C17122 VDD.t146 VSS 0.010055f
C17123 VDD.n2300 VSS 0.01771f
C17124 VDD.n2301 VSS 0.011881f
C17125 VDD.n2304 VSS 0.011881f
C17126 VDD.n2307 VSS 0.011881f
C17127 VDD.n2308 VSS 0.013523f
C17128 VDD.n2309 VSS 0.015015f
C17129 VDD.t1158 VSS 0.014745f
C17130 VDD.n2310 VSS 0.013668f
C17131 VDD.n2311 VSS 0.013668f
C17132 VDD.n2312 VSS 0.03134f
C17133 VDD.t77 VSS 0.010137f
C17134 VDD.t3795 VSS 0.021516f
C17135 VDD.n2314 VSS 0.055166f
C17136 VDD.t78 VSS 0.010137f
C17137 VDD.n2315 VSS 0.030049f
C17138 VDD.t186 VSS 0.010137f
C17139 VDD.t3801 VSS 0.021516f
C17140 VDD.n2317 VSS 0.055166f
C17141 VDD.t187 VSS 0.010137f
C17142 VDD.n2318 VSS 0.030049f
C17143 VDD.n2319 VSS 0.02678f
C17144 VDD.t260 VSS 0.014745f
C17145 VDD.t2167 VSS 0.014745f
C17146 VDD.n2321 VSS 0.035938f
C17147 VDD.n2323 VSS 0.053216f
C17148 VDD.n2324 VSS 0.011881f
C17149 VDD.n2325 VSS 0.011881f
C17150 VDD.n2327 VSS 0.020999f
C17151 VDD.n2329 VSS 0.011881f
C17152 VDD.n2330 VSS 0.011881f
C17153 VDD.n2334 VSS 0.011881f
C17154 VDD.n2335 VSS 0.011881f
C17155 VDD.n2336 VSS 0.015495f
C17156 VDD.n2338 VSS 0.011917f
C17157 VDD.n2339 VSS 0.011881f
C17158 VDD.n2340 VSS 0.011881f
C17159 VDD.n2341 VSS 0.03017f
C17160 VDD.n2342 VSS 0.023899f
C17161 VDD.n2343 VSS 0.023127f
C17162 VDD.n2344 VSS 0.017288f
C17163 VDD.n2345 VSS 0.023677f
C17164 VDD.n2346 VSS 0.023938f
C17165 VDD.n2347 VSS 0.036541f
C17166 VDD.n2351 VSS 0.011881f
C17167 VDD.n2352 VSS 0.011881f
C17168 VDD.n2354 VSS 0.010708f
C17169 VDD.n2357 VSS 0.011881f
C17170 VDD.n2358 VSS 0.011881f
C17171 VDD.t37 VSS 0.062814f
C17172 VDD.n2362 VSS 0.012066f
C17173 VDD.n2363 VSS 0.011881f
C17174 VDD.n2364 VSS 0.010563f
C17175 VDD.n2367 VSS 0.015126f
C17176 VDD.n2368 VSS 0.011881f
C17177 VDD.n2369 VSS 0.010783f
C17178 VDD.n2370 VSS 0.014062f
C17179 VDD.n2371 VSS 0.011881f
C17180 VDD.n2375 VSS 0.018262f
C17181 VDD.n2376 VSS 0.011881f
C17182 VDD.n2378 VSS 0.011881f
C17183 VDD.n2379 VSS 0.011147f
C17184 VDD.t434 VSS 0.013682f
C17185 VDD.t322 VSS 0.01447f
C17186 VDD.n2380 VSS 0.01757f
C17187 VDD.n2381 VSS 0.011881f
C17188 VDD.t563 VSS 0.01449f
C17189 VDD.n2383 VSS 0.011881f
C17190 VDD.t316 VSS 0.014212f
C17191 VDD.t2260 VSS 0.012962f
C17192 VDD.n2384 VSS 0.031771f
C17193 VDD.n2385 VSS 0.011881f
C17194 VDD.n2386 VSS 0.010543f
C17195 VDD.n2387 VSS 0.011881f
C17196 VDD.t1315 VSS 0.012738f
C17197 VDD.n2389 VSS 0.014011f
C17198 VDD.n2390 VSS 0.011881f
C17199 VDD.t1112 VSS 0.013828f
C17200 VDD.t1114 VSS 0.012728f
C17201 VDD.n2391 VSS 0.011881f
C17202 VDD.n2393 VSS 0.018529f
C17203 VDD.n2394 VSS 0.011881f
C17204 VDD.n2395 VSS 0.010127f
C17205 VDD.n2397 VSS 0.011881f
C17206 VDD.t1096 VSS 0.012563f
C17207 VDD.t1506 VSS 0.013789f
C17208 VDD.n2398 VSS 0.025097f
C17209 VDD.n2399 VSS 0.011881f
C17210 VDD.t2446 VSS 0.014194f
C17211 VDD.n2400 VSS 0.011881f
C17212 VDD.t3205 VSS 0.014068f
C17213 VDD.n2402 VSS 0.012875f
C17214 VDD.n2403 VSS 0.011881f
C17215 VDD.n2405 VSS 0.011867f
C17216 VDD.n2406 VSS 0.011881f
C17217 VDD.t3342 VSS 0.014214f
C17218 VDD.n2409 VSS 0.012066f
C17219 VDD.n2410 VSS 0.011881f
C17220 VDD.t3561 VSS 0.014212f
C17221 VDD.n2413 VSS 0.014646f
C17222 VDD.n2414 VSS 0.011881f
C17223 VDD.t493 VSS 0.036927f
C17224 VDD.n2416 VSS 0.012066f
C17225 VDD.n2418 VSS 0.014722f
C17226 VDD.n2419 VSS 0.011881f
C17227 VDD.n2423 VSS 0.011881f
C17228 VDD.n2427 VSS 0.016408f
C17229 VDD.n2428 VSS 0.011881f
C17230 VDD.t3695 VSS 0.014068f
C17231 VDD.n2429 VSS 0.011881f
C17232 VDD.t310 VSS 0.01449f
C17233 VDD.t2426 VSS 0.012672f
C17234 VDD.n2431 VSS 0.019325f
C17235 VDD.n2432 VSS 0.011881f
C17236 VDD.t1866 VSS 0.014212f
C17237 VDD.t510 VSS 0.01447f
C17238 VDD.n2434 VSS 0.011881f
C17239 VDD.n2435 VSS 0.011881f
C17240 VDD.t512 VSS 0.014477f
C17241 VDD.t1410 VSS 0.01449f
C17242 VDD.n2436 VSS 0.011881f
C17243 VDD.n2437 VSS 0.013378f
C17244 VDD.n2438 VSS 0.011881f
C17245 VDD.t2835 VSS 0.014212f
C17246 VDD.t3113 VSS 0.014498f
C17247 VDD.n2439 VSS 0.024723f
C17248 VDD.n2440 VSS 0.011881f
C17249 VDD.t2615 VSS 0.012672f
C17250 VDD.n2442 VSS 0.011881f
C17251 VDD.t3608 VSS 0.01449f
C17252 VDD.n2444 VSS 0.011881f
C17253 VDD.t2351 VSS 0.01445f
C17254 VDD.t3648 VSS 0.014458f
C17255 VDD.n2445 VSS 0.040246f
C17256 VDD.n2446 VSS 0.011881f
C17257 VDD.t3637 VSS 0.01447f
C17258 VDD.t1282 VSS 0.014485f
C17259 VDD.t3628 VSS 0.014477f
C17260 VDD.n2447 VSS 0.011881f
C17261 VDD.t1750 VSS 0.014214f
C17262 VDD.n2448 VSS 0.017968f
C17263 VDD.n2449 VSS 0.011881f
C17264 VDD.t3772 VSS 0.041965f
C17265 VDD.t346 VSS 0.014214f
C17266 VDD.n2450 VSS 0.026838f
C17267 VDD.n2451 VSS 0.011881f
C17268 VDD.t2190 VSS 0.014485f
C17269 VDD.t237 VSS 0.013966f
C17270 VDD.t2232 VSS 0.01449f
C17271 VDD.n2452 VSS 0.011881f
C17272 VDD.n2453 VSS 0.011881f
C17273 VDD.n2455 VSS 0.014361f
C17274 VDD.n2457 VSS 0.011881f
C17275 VDD.n2458 VSS 0.011881f
C17276 VDD.t1301 VSS 0.013966f
C17277 VDD.n2461 VSS 0.011881f
C17278 VDD.n2463 VSS 0.011064f
C17279 VDD.n2464 VSS 0.018905f
C17280 VDD.n2465 VSS 0.011881f
C17281 VDD.n2467 VSS 0.011881f
C17282 VDD.t1449 VSS 0.01449f
C17283 VDD.t3759 VSS 0.014485f
C17284 VDD.n2468 VSS 0.02085f
C17285 VDD.n2469 VSS 0.011881f
C17286 VDD.n2470 VSS 0.011147f
C17287 VDD.n2471 VSS 0.01596f
C17288 VDD.t1638 VSS 0.053297f
C17289 VDD.n2473 VSS 0.011417f
C17290 VDD.n2475 VSS 0.011881f
C17291 VDD.t986 VSS 0.015916f
C17292 VDD.n2476 VSS 0.024603f
C17293 VDD.n2477 VSS 0.011881f
C17294 VDD.n2478 VSS 0.010534f
C17295 VDD.n2481 VSS 0.011881f
C17296 VDD.t2788 VSS 0.010846f
C17297 VDD.n2482 VSS 0.015232f
C17298 VDD.n2483 VSS 0.010736f
C17299 VDD.n2484 VSS 0.011881f
C17300 VDD.n2485 VSS 0.021015f
C17301 VDD.n2486 VSS 0.011881f
C17302 VDD.n2488 VSS 0.011881f
C17303 VDD.t1485 VSS 0.014477f
C17304 VDD.n2489 VSS 0.018218f
C17305 VDD.t1544 VSS 0.015219f
C17306 VDD.n2490 VSS 0.011881f
C17307 VDD.n2491 VSS 0.013931f
C17308 VDD.t1488 VSS 0.014204f
C17309 VDD.t868 VSS 0.014219f
C17310 VDD.n2492 VSS 0.021226f
C17311 VDD.n2493 VSS 0.011881f
C17312 VDD.t3734 VSS 0.0145f
C17313 VDD.n2494 VSS 0.023986f
C17314 VDD.t188 VSS 0.222704f
C17315 VDD.t393 VSS 0.120679f
C17316 VDD.t395 VSS 0.068144f
C17317 VDD.t1891 VSS 0.108116f
C17318 VDD.t595 VSS 0.08832f
C17319 VDD.t140 VSS 0.031978f
C17320 VDD.t593 VSS 0.051774f
C17321 VDD.t1965 VSS 0.054439f
C17322 VDD.t1227 VSS 0.014745f
C17323 VDD.n2495 VSS 0.019581f
C17324 VDD.n2496 VSS 0.011881f
C17325 VDD.n2497 VSS 0.011578f
C17326 VDD.n2498 VSS 0.011881f
C17327 VDD.t3771 VSS 0.05912f
C17328 VDD.t3137 VSS 0.014204f
C17329 VDD.n2499 VSS 0.013685f
C17330 VDD.t128 VSS 0.010055f
C17331 VDD.n2500 VSS 0.017032f
C17332 VDD.t3150 VSS 0.014207f
C17333 VDD.n2502 VSS 0.024333f
C17334 VDD.n2503 VSS 0.011881f
C17335 VDD.n2505 VSS 0.011881f
C17336 VDD.n2508 VSS 0.011881f
C17337 VDD.t1182 VSS 0.010806f
C17338 VDD.n2511 VSS 0.012162f
C17339 VDD.n2512 VSS 0.011881f
C17340 VDD.t2152 VSS 0.014469f
C17341 VDD.n2513 VSS 0.016565f
C17342 VDD.n2515 VSS 0.013668f
C17343 VDD.n2516 VSS 0.011881f
C17344 VDD.t2672 VSS 0.015916f
C17345 VDD.n2517 VSS 0.023711f
C17346 VDD.n2518 VSS 0.011881f
C17347 VDD.n2519 VSS 0.011881f
C17348 VDD.n2520 VSS 0.011881f
C17349 VDD.n2522 VSS 0.010708f
C17350 VDD.n2525 VSS 0.011385f
C17351 VDD.n2526 VSS 0.011881f
C17352 VDD.n2527 VSS 0.011881f
C17353 VDD.n2528 VSS 0.011881f
C17354 VDD.n2529 VSS 0.018529f
C17355 VDD.n2532 VSS 0.011881f
C17356 VDD.n2533 VSS 0.011881f
C17357 VDD.n2539 VSS 0.011881f
C17358 VDD.n2540 VSS 0.011881f
C17359 VDD.n2541 VSS 0.011881f
C17360 VDD.n2546 VSS 0.011881f
C17361 VDD.n2547 VSS 0.011881f
C17362 VDD.n2549 VSS 0.011917f
C17363 VDD.t129 VSS 0.010055f
C17364 VDD.n2550 VSS 0.01771f
C17365 VDD.n2551 VSS 0.014915f
C17366 VDD.n2552 VSS 0.011881f
C17367 VDD.n2553 VSS 0.011881f
C17368 VDD.n2554 VSS 0.030848f
C17369 VDD.n2555 VSS 0.015933f
C17370 VDD.n2556 VSS 0.029485f
C17371 VDD.n2557 VSS 0.079913f
C17372 VDD.n2558 VSS 0.011881f
C17373 VDD.n2559 VSS 0.011881f
C17374 VDD.n2560 VSS 0.011881f
C17375 VDD.n2562 VSS 0.013668f
C17376 VDD.n2563 VSS 0.017774f
C17377 VDD.n2565 VSS 0.017065f
C17378 VDD.n2566 VSS 0.011881f
C17379 VDD.n2567 VSS 0.011881f
C17380 VDD.n2568 VSS 0.019778f
C17381 VDD.t141 VSS 0.010137f
C17382 VDD.t3810 VSS 0.021516f
C17383 VDD.n2570 VSS 0.055166f
C17384 VDD.t142 VSS 0.010137f
C17385 VDD.n2571 VSS 0.030049f
C17386 VDD.n2572 VSS 0.019845f
C17387 VDD.n2573 VSS 0.013523f
C17388 VDD.t596 VSS 0.014469f
C17389 VDD.n2574 VSS 0.031602f
C17390 VDD.n2575 VSS 0.013668f
C17391 VDD.n2576 VSS 0.013668f
C17392 VDD.n2577 VSS 0.03134f
C17393 VDD.t189 VSS 0.010137f
C17394 VDD.t3827 VSS 0.021516f
C17395 VDD.n2579 VSS 0.055166f
C17396 VDD.t190 VSS 0.010137f
C17397 VDD.n2580 VSS 0.030049f
C17398 VDD.t210 VSS 0.010137f
C17399 VDD.t3807 VSS 0.021516f
C17400 VDD.n2582 VSS 0.055166f
C17401 VDD.t211 VSS 0.010137f
C17402 VDD.n2583 VSS 0.030049f
C17403 VDD.n2584 VSS 0.02678f
C17404 VDD.t578 VSS 0.014745f
C17405 VDD.t394 VSS 0.014745f
C17406 VDD.n2586 VSS 0.035938f
C17407 VDD.n2588 VSS 0.053216f
C17408 VDD.n2589 VSS 0.011881f
C17409 VDD.n2590 VSS 0.01978f
C17410 VDD.n2592 VSS 0.017356f
C17411 VDD.n2593 VSS 0.023851f
C17412 VDD.n2594 VSS 0.078132f
C17413 VDD.t2242 VSS 0.053677f
C17414 VDD.t1226 VSS 0.032359f
C17415 VDD.t1228 VSS 0.03312f
C17416 VDD.t3574 VSS 0.036166f
C17417 VDD.t347 VSS 0.107355f
C17418 VDD.t3136 VSS 0.104309f
C17419 VDD.t3149 VSS 0.068524f
C17420 VDD.t127 VSS 0.072331f
C17421 VDD.t3140 VSS 0.067763f
C17422 VDD.t1647 VSS 0.113446f
C17423 VDD.t3345 VSS 0.101644f
C17424 VDD.t2781 VSS 0.045302f
C17425 VDD.t2427 VSS 0.035023f
C17426 VDD.t2415 VSS 0.047586f
C17427 VDD.t1646 VSS 0.08832f
C17428 VDD.t2429 VSS 0.053297f
C17429 VDD.t2604 VSS 0.039592f
C17430 VDD.t3349 VSS 0.046825f
C17431 VDD.t1255 VSS 0.074996f
C17432 VDD.t1181 VSS 0.079184f
C17433 VDD.t2151 VSS 0.037688f
C17434 VDD.t1649 VSS 0.031978f
C17435 VDD.t2149 VSS 0.032739f
C17436 VDD.t2416 VSS 0.036166f
C17437 VDD.t1541 VSS 0.031978f
C17438 VDD.t2673 VSS 0.061291f
C17439 VDD.t3426 VSS 0.073092f
C17440 VDD.t2702 VSS 0.080326f
C17441 VDD.t1309 VSS 0.075757f
C17442 VDD.t3733 VSS 0.033501f
C17443 VDD.t2671 VSS 0.059388f
C17444 VDD.t1960 VSS 0.106593f
C17445 VDD.t985 VSS 0.07157f
C17446 VDD.t3522 VSS 0.037688f
C17447 VDD.t2854 VSS 0.063956f
C17448 VDD.t849 VSS 0.04416f
C17449 VDD.t2199 VSS 0.034643f
C17450 VDD.t3673 VSS 0.031978f
C17451 VDD.t3351 VSS 0.037308f
C17452 VDD.t850 VSS 0.041114f
C17453 VDD.t987 VSS 0.04949f
C17454 VDD.t2198 VSS 0.056342f
C17455 VDD.t2369 VSS 0.032739f
C17456 VDD.t2658 VSS 0.037308f
C17457 VDD.t3675 VSS 0.037688f
C17458 VDD.t2787 VSS 0.036166f
C17459 VDD.t244 VSS 0.054819f
C17460 VDD.t2368 VSS 0.047586f
C17461 VDD.t3406 VSS 0.057103f
C17462 VDD.t2201 VSS 0.051393f
C17463 VDD.t3122 VSS 0.053297f
C17464 VDD.t2655 VSS 0.07157f
C17465 VDD.t3186 VSS 0.037688f
C17466 VDD.t2197 VSS 0.037308f
C17467 VDD.t2745 VSS 0.035023f
C17468 VDD.t293 VSS 0.036546f
C17469 VDD.t2747 VSS 0.096315f
C17470 VDD.t1535 VSS 0.067763f
C17471 VDD.t2656 VSS 0.031978f
C17472 VDD.t1543 VSS 0.031978f
C17473 VDD.t3142 VSS 0.077661f
C17474 VDD.t1484 VSS 0.08832f
C17475 VDD.t2675 VSS 0.031978f
C17476 VDD.t1487 VSS 0.041114f
C17477 VDD.t2930 VSS 0.057103f
C17478 VDD.t3200 VSS 0.053297f
C17479 VDD.t867 VSS 0.048728f
C17480 VDD.t3090 VSS 0.045683f
C17481 VDD.n2595 VSS 0.078132f
C17482 VDD.n2596 VSS 0.024538f
C17483 VDD.n2597 VSS 0.012298f
C17484 VDD.n2599 VSS 0.011881f
C17485 VDD.n2600 VSS 0.011881f
C17486 VDD.n2603 VSS 0.013812f
C17487 VDD.n2604 VSS 0.014599f
C17488 VDD.n2606 VSS 0.011881f
C17489 VDD.n2607 VSS 0.011881f
C17490 VDD.n2608 VSS 0.011881f
C17491 VDD.n2609 VSS 0.024257f
C17492 VDD.n2611 VSS 0.013449f
C17493 VDD.n2613 VSS 0.012779f
C17494 VDD.n2614 VSS 0.014394f
C17495 VDD.n2617 VSS 0.011881f
C17496 VDD.n2618 VSS 0.011881f
C17497 VDD.n2619 VSS 0.011881f
C17498 VDD.n2620 VSS 0.011028f
C17499 VDD.n2621 VSS 0.010601f
C17500 VDD.n2622 VSS 0.01554f
C17501 VDD.n2624 VSS 0.011881f
C17502 VDD.n2625 VSS 0.011881f
C17503 VDD.n2626 VSS 0.011881f
C17504 VDD.n2629 VSS 0.011101f
C17505 VDD.n2632 VSS 0.011881f
C17506 VDD.n2633 VSS 0.011881f
C17507 VDD.n2634 VSS 0.011881f
C17508 VDD.n2635 VSS 0.016729f
C17509 VDD.n2638 VSS 0.011881f
C17510 VDD.n2639 VSS 0.011881f
C17511 VDD.n2641 VSS 0.013629f
C17512 VDD.n2643 VSS 0.010708f
C17513 VDD.n2645 VSS 0.011881f
C17514 VDD.n2646 VSS 0.011881f
C17515 VDD.n2647 VSS 0.011881f
C17516 VDD.n2650 VSS 0.02494f
C17517 VDD.n2651 VSS 0.011881f
C17518 VDD.n2652 VSS 0.011881f
C17519 VDD.t3670 VSS 0.012563f
C17520 VDD.n2654 VSS 0.011881f
C17521 VDD.t2844 VSS 0.014485f
C17522 VDD.n2655 VSS 0.010736f
C17523 VDD.n2656 VSS 0.011881f
C17524 VDD.t806 VSS 0.01449f
C17525 VDD.n2658 VSS 0.011385f
C17526 VDD.n2659 VSS 0.011881f
C17527 VDD.n2662 VSS 0.011064f
C17528 VDD.n2663 VSS 0.018196f
C17529 VDD.n2664 VSS 0.011881f
C17530 VDD.t56 VSS 0.012707f
C17531 VDD.t2839 VSS 0.014477f
C17532 VDD.t2846 VSS 0.014204f
C17533 VDD.n2665 VSS 0.014772f
C17534 VDD.n2666 VSS 0.011881f
C17535 VDD.t2164 VSS 0.012673f
C17536 VDD.n2670 VSS 0.011881f
C17537 VDD.n2673 VSS 0.011881f
C17538 VDD.n2674 VSS 0.010911f
C17539 VDD.n2675 VSS 0.014361f
C17540 VDD.n2676 VSS 0.011881f
C17541 VDD.n2678 VSS 0.011267f
C17542 VDD.n2680 VSS 0.013817f
C17543 VDD.n2682 VSS 0.011881f
C17544 VDD.n2683 VSS 0.011881f
C17545 VDD.n2684 VSS 0.011881f
C17546 VDD.n2689 VSS 0.011881f
C17547 VDD.n2690 VSS 0.011881f
C17548 VDD.n2693 VSS 0.019325f
C17549 VDD.n2695 VSS 0.011881f
C17550 VDD.n2696 VSS 0.011881f
C17551 VDD.n2698 VSS 0.018447f
C17552 VDD.n2699 VSS 0.011907f
C17553 VDD.n2700 VSS 0.011881f
C17554 VDD.n2701 VSS 0.011881f
C17555 VDD.n2702 VSS 0.011881f
C17556 VDD.n2706 VSS 0.010327f
C17557 VDD.n2708 VSS 0.011881f
C17558 VDD.n2709 VSS 0.011881f
C17559 VDD.n2710 VSS 0.011881f
C17560 VDD.n2712 VSS 0.021615f
C17561 VDD.n2713 VSS 0.015746f
C17562 VDD.n2714 VSS 0.020118f
C17563 VDD.n2715 VSS 0.011881f
C17564 VDD.n2716 VSS 0.011881f
C17565 VDD.n2717 VSS 0.011881f
C17566 VDD.n2720 VSS 0.029776f
C17567 VDD.n2721 VSS 0.011881f
C17568 VDD.n2722 VSS 0.011881f
C17569 VDD.n2723 VSS 0.011881f
C17570 VDD.n2724 VSS 0.022317f
C17571 VDD.n2725 VSS 0.041222f
C17572 VDD.t3292 VSS 0.054058f
C17573 VDD.t3669 VSS 0.070047f
C17574 VDD.t1520 VSS 0.070808f
C17575 VDD.t1000 VSS 0.068524f
C17576 VDD.t3111 VSS 0.035023f
C17577 VDD.t2504 VSS 0.030455f
C17578 VDD.t2853 VSS 0.063575f
C17579 VDD.t1957 VSS 0.041114f
C17580 VDD.t2843 VSS 0.036927f
C17581 VDD.t805 VSS 0.032359f
C17582 VDD.t750 VSS 0.073092f
C17583 VDD.t3643 VSS 0.09936f
C17584 VDD.t1003 VSS 0.036546f
C17585 VDD.t3025 VSS 0.036546f
C17586 VDD.t3664 VSS 0.036546f
C17587 VDD.t847 VSS 0.036546f
C17588 VDD.t3105 VSS 0.031978f
C17589 VDD.t3548 VSS 0.035785f
C17590 VDD.t3726 VSS 0.031978f
C17591 VDD.t42 VSS 0.037688f
C17592 VDD.t1387 VSS 0.07157f
C17593 VDD.t55 VSS 0.072712f
C17594 VDD.t2838 VSS 0.069286f
C17595 VDD.t2845 VSS 0.034262f
C17596 VDD.t2163 VSS 0.070047f
C17597 VDD.t3124 VSS 0.087559f
C17598 VDD.t1287 VSS 0.033501f
C17599 VDD.t1431 VSS 0.036546f
C17600 VDD.t979 VSS 0.037308f
C17601 VDD.t3661 VSS 0.02741f
C17602 VDD.t3110 VSS 0.094411f
C17603 VDD.t648 VSS 0.112684f
C17604 VDD.t2717 VSS 0.039211f
C17605 VDD.t1292 VSS 0.040734f
C17606 VDD.t3114 VSS 0.041495f
C17607 VDD.t533 VSS 0.031978f
C17608 VDD.t1370 VSS 0.053297f
C17609 VDD.t505 VSS 0.062433f
C17610 VDD.t1973 VSS 0.032739f
C17611 VDD.t489 VSS 0.035785f
C17612 VDD.t503 VSS 0.03312f
C17613 VDD.t1650 VSS 0.032739f
C17614 VDD.t507 VSS 0.065098f
C17615 VDD.t483 VSS 0.052916f
C17616 VDD.t1294 VSS 0.032739f
C17617 VDD.t479 VSS 0.036166f
C17618 VDD.t2205 VSS 0.032739f
C17619 VDD.t3696 VSS 0.041876f
C17620 VDD.t3698 VSS 0.062433f
C17621 VDD.t265 VSS 0.032739f
C17622 VDD.t3700 VSS 0.035785f
C17623 VDD.t3694 VSS 0.03312f
C17624 VDD.t267 VSS 0.07195f
C17625 VDD.t2425 VSS 0.073092f
C17626 VDD.t309 VSS 0.033501f
C17627 VDD.t1865 VSS 0.06624f
C17628 VDD.t3265 VSS 0.067763f
C17629 VDD.t2423 VSS 0.038069f
C17630 VDD.t509 VSS 0.036546f
C17631 VDD.t511 VSS 0.032739f
C17632 VDD.t966 VSS 0.073854f
C17633 VDD.t1409 VSS 0.10507f
C17634 VDD.t2834 VSS 0.068524f
C17635 VDD.t3704 VSS 0.077661f
C17636 VDD.t3047 VSS 0.068524f
C17637 VDD.t3112 VSS 0.063956f
C17638 VDD.t2614 VSS 0.07157f
C17639 VDD.t3042 VSS 0.067001f
C17640 VDD.t3607 VSS 0.032739f
C17641 VDD.t3618 VSS 0.034262f
C17642 VDD.t2612 VSS 0.070808f
C17643 VDD.t3310 VSS 0.040353f
C17644 VDD.t2350 VSS 0.035023f
C17645 VDD.t3647 VSS 0.050251f
C17646 VDD.n2726 VSS 0.078893f
C17647 VDD.t3636 VSS 0.086036f
C17648 VDD.t3627 VSS 0.034262f
C17649 VDD.t1281 VSS 0.034262f
C17650 VDD.t1749 VSS 0.104309f
C17651 VDD.t163 VSS 0.073092f
C17652 VDD.t1975 VSS 0.032739f
C17653 VDD.t345 VSS 0.10507f
C17654 VDD.t2189 VSS 0.073473f
C17655 VDD.t236 VSS 0.031978f
C17656 VDD.t2231 VSS 0.072331f
C17657 VDD.t1641 VSS 0.073092f
C17658 VDD.t2229 VSS 0.032739f
C17659 VDD.t249 VSS 0.03312f
C17660 VDD.t3679 VSS 0.041114f
C17661 VDD.t1298 VSS 0.035023f
C17662 VDD.t1289 VSS 0.039211f
C17663 VDD.t1640 VSS 0.072331f
C17664 VDD.t1300 VSS 0.081468f
C17665 VDD.t647 VSS 0.049109f
C17666 VDD.t2715 VSS 0.050632f
C17667 VDD.t650 VSS 0.036546f
C17668 VDD.t1290 VSS 0.032739f
C17669 VDD.t3116 VSS 0.052155f
C17670 VDD.t3689 VSS 0.067763f
C17671 VDD.t1296 VSS 0.037308f
C17672 VDD.t2849 VSS 0.039972f
C17673 VDD.t3730 VSS 0.073473f
C17674 VDD.t242 VSS 0.072331f
C17675 VDD.t1364 VSS 0.067763f
C17676 VDD.t1448 VSS 0.036546f
C17677 VDD.t804 VSS 0.031978f
C17678 VDD.t3758 VSS 0.108116f
C17679 VDD.t238 VSS 0.08832f
C17680 VDD.n2727 VSS 0.043125f
C17681 VDD.n2728 VSS 0.022751f
C17682 VDD.n2730 VSS 0.011881f
C17683 VDD.n2731 VSS 0.011881f
C17684 VDD.n2732 VSS 0.011881f
C17685 VDD.n2734 VSS 0.021089f
C17686 VDD.n2735 VSS 0.013228f
C17687 VDD.n2737 VSS 0.011881f
C17688 VDD.n2738 VSS 0.011881f
C17689 VDD.n2739 VSS 0.011881f
C17690 VDD.n2742 VSS 0.011121f
C17691 VDD.n2743 VSS 0.011881f
C17692 VDD.n2744 VSS 0.011881f
C17693 VDD.n2746 VSS 0.018794f
C17694 VDD.n2749 VSS 0.011881f
C17695 VDD.n2750 VSS 0.011881f
C17696 VDD.n2751 VSS 0.011881f
C17697 VDD.n2753 VSS 0.010375f
C17698 VDD.n2754 VSS 0.011464f
C17699 VDD.n2755 VSS 0.020792f
C17700 VDD.n2756 VSS 0.017651f
C17701 VDD.n2757 VSS 0.019985f
C17702 VDD.n2758 VSS 0.011881f
C17703 VDD.n2759 VSS 0.011881f
C17704 VDD.t164 VSS 0.010055f
C17705 VDD.n2762 VSS 0.037956f
C17706 VDD.n2763 VSS 0.02339f
C17707 VDD.t1976 VSS 0.014212f
C17708 VDD.t165 VSS 0.010055f
C17709 VDD.n2764 VSS 0.017032f
C17710 VDD.n2765 VSS 0.030304f
C17711 VDD.n2766 VSS 0.016102f
C17712 VDD.n2767 VSS 0.011881f
C17713 VDD.n2768 VSS 0.011881f
C17714 VDD.n2769 VSS 0.01046f
C17715 VDD.n2770 VSS 0.018193f
C17716 VDD.n2771 VSS 0.019707f
C17717 VDD.n2772 VSS 0.016244f
C17718 VDD.n2773 VSS 0.011881f
C17719 VDD.n2774 VSS 0.011881f
C17720 VDD.n2775 VSS 0.011881f
C17721 VDD.n2777 VSS 0.0296f
C17722 VDD.n2778 VSS 0.021455f
C17723 VDD.n2780 VSS 0.019325f
C17724 VDD.t3043 VSS 0.014212f
C17725 VDD.n2781 VSS 0.017191f
C17726 VDD.n2783 VSS 0.011881f
C17727 VDD.n2784 VSS 0.011881f
C17728 VDD.n2785 VSS 0.011881f
C17729 VDD.n2788 VSS 0.017831f
C17730 VDD.n2790 VSS 0.011881f
C17731 VDD.n2791 VSS 0.011881f
C17732 VDD.n2793 VSS 0.021683f
C17733 VDD.n2794 VSS 0.017418f
C17734 VDD.n2795 VSS 0.012405f
C17735 VDD.n2796 VSS 0.016793f
C17736 VDD.n2797 VSS 0.017442f
C17737 VDD.n2799 VSS 0.011881f
C17738 VDD.n2800 VSS 0.011881f
C17739 VDD.n2802 VSS 0.021546f
C17740 VDD.n2803 VSS 0.018105f
C17741 VDD.n2807 VSS 0.011881f
C17742 VDD.n2808 VSS 0.011881f
C17743 VDD.n2809 VSS 0.011881f
C17744 VDD.n2811 VSS 0.012736f
C17745 VDD.n2813 VSS 0.010876f
C17746 VDD.n2815 VSS 0.013213f
C17747 VDD.n2817 VSS 0.011881f
C17748 VDD.n2818 VSS 0.011881f
C17749 VDD.n2819 VSS 0.011881f
C17750 VDD.n2821 VSS 0.024658f
C17751 VDD.n2823 VSS 0.011881f
C17752 VDD.n2824 VSS 0.011881f
C17753 VDD.n2827 VSS 0.013876f
C17754 VDD.n2828 VSS 0.011881f
C17755 VDD.t492 VSS 0.013297f
C17756 VDD.n2829 VSS 0.015855f
C17757 VDD.n2830 VSS 0.011881f
C17758 VDD.n2831 VSS 0.010602f
C17759 VDD.n2832 VSS 0.011474f
C17760 VDD.n2833 VSS 0.011881f
C17761 VDD.n2834 VSS 0.010736f
C17762 VDD.n2835 VSS 0.015746f
C17763 VDD.t2831 VSS 0.01449f
C17764 VDD.n2836 VSS 0.011881f
C17765 VDD.n2839 VSS 0.011881f
C17766 VDD.n2841 VSS 0.011912f
C17767 VDD.n2844 VSS 0.014694f
C17768 VDD.n2845 VSS 0.011912f
C17769 VDD.n2846 VSS 0.014361f
C17770 VDD.n2847 VSS 0.010174f
C17771 VDD.n2849 VSS 0.011881f
C17772 VDD.n2850 VSS 0.011912f
C17773 VDD.n2851 VSS 0.011881f
C17774 VDD.n2853 VSS 0.014694f
C17775 VDD.n2855 VSS 0.01215f
C17776 VDD.n2857 VSS 0.011881f
C17777 VDD.n2858 VSS 0.011881f
C17778 VDD.t1025 VSS 0.013297f
C17779 VDD.n2860 VSS 0.016564f
C17780 VDD.t3102 VSS 0.014485f
C17781 VDD.n2861 VSS 0.02005f
C17782 VDD.n2862 VSS 0.011881f
C17783 VDD.n2863 VSS 0.011881f
C17784 VDD.n2864 VSS 0.011881f
C17785 VDD.n2865 VSS 0.021432f
C17786 VDD.n2868 VSS 0.011881f
C17787 VDD.n2869 VSS 0.011881f
C17788 VDD.n2870 VSS 0.011881f
C17789 VDD.n2871 VSS 0.02026f
C17790 VDD.t530 VSS 0.01455f
C17791 VDD.n2873 VSS 0.023997f
C17792 VDD.n2874 VSS 0.011881f
C17793 VDD.n2875 VSS 0.011881f
C17794 VDD.n2876 VSS 0.011881f
C17795 VDD.n2877 VSS 0.010684f
C17796 VDD.n2878 VSS 0.015537f
C17797 VDD.n2880 VSS 0.013924f
C17798 VDD.t3568 VSS 0.014498f
C17799 VDD.n2881 VSS 0.023522f
C17800 VDD.n2882 VSS 0.011881f
C17801 VDD.n2883 VSS 0.011881f
C17802 VDD.n2884 VSS 0.011881f
C17803 VDD.n2886 VSS 0.01148f
C17804 VDD.n2888 VSS 0.013439f
C17805 VDD.n2890 VSS 0.011881f
C17806 VDD.n2891 VSS 0.011881f
C17807 VDD.n2892 VSS 0.011881f
C17808 VDD.n2893 VSS 0.02342f
C17809 VDD.n2894 VSS 0.038938f
C17810 VDD.t477 VSS 0.06091f
C17811 VDD.t485 VSS 0.065098f
C17812 VDD.t497 VSS 0.062433f
C17813 VDD.t3045 VSS 0.032739f
C17814 VDD.t481 VSS 0.035785f
C17815 VDD.t499 VSS 0.038069f
C17816 VDD.t2279 VSS 0.032739f
C17817 VDD.t487 VSS 0.060149f
C17818 VDD.t495 VSS 0.065479f
C17819 VDD.t501 VSS 0.040353f
C17820 VDD.t874 VSS 0.032739f
C17821 VDD.t491 VSS 0.037308f
C17822 VDD.t964 VSS 0.048728f
C17823 VDD.t2004 VSS 0.063956f
C17824 VDD.t1959 VSS 0.030074f
C17825 VDD.t529 VSS 0.030074f
C17826 VDD.t3565 VSS 0.068524f
C17827 VDD.t3286 VSS 0.042257f
C17828 VDD.t1878 VSS 0.041114f
C17829 VDD.t956 VSS 0.07157f
C17830 VDD.t2 VSS 0.059007f
C17831 VDD.t2913 VSS 0.063575f
C17832 VDD.t970 VSS 0.042637f
C17833 VDD.t2830 VSS 0.037308f
C17834 VDD.t0 VSS 0.031978f
C17835 VDD.t3101 VSS 0.079564f
C17836 VDD.t1024 VSS 0.089081f
C17837 VDD.t2333 VSS 0.032739f
C17838 VDD.t1010 VSS 0.036546f
C17839 VDD.t2832 VSS 0.032739f
C17840 VDD.t1004 VSS 0.02741f
C17841 VDD.t2679 VSS 0.032739f
C17842 VDD.t1022 VSS 0.056342f
C17843 VDD.t1028 VSS 0.057865f
C17844 VDD.t1882 VSS 0.032739f
C17845 VDD.t1026 VSS 0.039211f
C17846 VDD.t2335 VSS 0.032739f
C17847 VDD.t1030 VSS 0.033881f
C17848 VDD.t1006 VSS 0.040353f
C17849 VDD.t3493 VSS 0.032359f
C17850 VDD.t1016 VSS 0.053297f
C17851 VDD.t11 VSS 0.051774f
C17852 VDD.t387 VSS 0.032739f
C17853 VDD.t35 VSS 0.041114f
C17854 VDD.t2775 VSS 0.032739f
C17855 VDD.t3214 VSS 0.038069f
C17856 VDD.t3172 VSS 0.035785f
C17857 VDD.t326 VSS 0.030455f
C17858 VDD.t686 VSS 0.029694f
C17859 VDD.t3226 VSS 0.035023f
C17860 VDD.t3224 VSS 0.070047f
C17861 VDD.t565 VSS 0.074996f
C17862 VDD.t3468 VSS 0.038069f
C17863 VDD.t666 VSS 0.03312f
C17864 VDD.t672 VSS 0.035404f
C17865 VDD.t1929 VSS 0.032739f
C17866 VDD.t670 VSS 0.036546f
C17867 VDD.t439 VSS 0.032739f
C17868 VDD.t668 VSS 0.036546f
C17869 VDD.t564 VSS 0.036546f
C17870 VDD.t1967 VSS 0.133241f
C17871 VDD.t3462 VSS 0.126008f
C17872 VDD.t1567 VSS 0.031978f
C17873 VDD.t3456 VSS 0.040734f
C17874 VDD.t2899 VSS 0.031978f
C17875 VDD.t435 VSS 0.031978f
C17876 VDD.t441 VSS 0.031978f
C17877 VDD.t433 VSS 0.036927f
C17878 VDD.t1911 VSS 0.079945f
C17879 VDD.t321 VSS 0.079184f
C17880 VDD.t317 VSS 0.104309f
C17881 VDD.t1826 VSS 0.073854f
C17882 VDD.t562 VSS 0.02741f
C17883 VDD.t2896 VSS 0.031978f
C17884 VDD.t315 VSS 0.129435f
C17885 VDD.n2895 VSS 0.147798f
C17886 VDD.t2259 VSS 0.04987f
C17887 VDD.t2905 VSS 0.068905f
C17888 VDD.t2017 VSS 0.03883f
C17889 VDD.t2743 VSS 0.038069f
C17890 VDD.t1312 VSS 0.068144f
C17891 VDD.t1314 VSS 0.033501f
C17892 VDD.t1819 VSS 0.033501f
C17893 VDD.t2261 VSS 0.063956f
C17894 VDD.t852 VSS 0.042637f
C17895 VDD.t1111 VSS 0.042637f
C17896 VDD.t2898 VSS 0.06091f
C17897 VDD.t1113 VSS 0.031978f
C17898 VDD.t1262 VSS 0.036546f
C17899 VDD.t2901 VSS 0.068905f
C17900 VDD.t2147 VSS 0.055961f
C17901 VDD.t1099 VSS 0.058626f
C17902 VDD.t3288 VSS 0.052155f
C17903 VDD.t1115 VSS 0.044921f
C17904 VDD.t854 VSS 0.035023f
C17905 VDD.t1480 VSS 0.036166f
C17906 VDD.t1505 VSS 0.035785f
C17907 VDD.t1095 VSS 0.07157f
C17908 VDD.t2445 VSS 0.070808f
C17909 VDD.t3044 VSS 0.035023f
C17910 VDD.t3606 VSS 0.068905f
C17911 VDD.t3204 VSS 0.069666f
C17912 VDD.t3218 VSS 0.065479f
C17913 VDD.t3208 VSS 0.050632f
C17914 VDD.t3569 VSS 0.032739f
C17915 VDD.t3220 VSS 0.031978f
C17916 VDD.t1791 VSS 0.032739f
C17917 VDD.t1008 VSS 0.041114f
C17918 VDD.t1272 VSS 0.032739f
C17919 VDD.t1018 VSS 0.039972f
C17920 VDD.t1012 VSS 0.065479f
C17921 VDD.t1014 VSS 0.04987f
C17922 VDD.t3341 VSS 0.032739f
C17923 VDD.t1032 VSS 0.031978f
C17924 VDD.t3560 VSS 0.032739f
C17925 VDD.t1034 VSS 0.049109f
C17926 VDD.t1020 VSS 0.036927f
C17927 VDD.n2896 VSS 0.038938f
C17928 VDD.n2897 VSS 0.02342f
C17929 VDD.n2898 VSS 0.011995f
C17930 VDD.n2899 VSS 0.01662f
C17931 VDD.n2902 VSS 0.011881f
C17932 VDD.n2903 VSS 0.011881f
C17933 VDD.n2905 VSS 0.019116f
C17934 VDD.n2907 VSS 0.013218f
C17935 VDD.n2908 VSS 0.014074f
C17936 VDD.n2909 VSS 0.015973f
C17937 VDD.n2911 VSS 0.011881f
C17938 VDD.n2912 VSS 0.011881f
C17939 VDD.n2915 VSS 0.012435f
C17940 VDD.n2917 VSS 0.011881f
C17941 VDD.n2918 VSS 0.011881f
C17942 VDD.n2920 VSS 0.018605f
C17943 VDD.n2922 VSS 0.012328f
C17944 VDD.n2924 VSS 0.011881f
C17945 VDD.n2925 VSS 0.011881f
C17946 VDD.n2926 VSS 0.011881f
C17947 VDD.n2928 VSS 0.015182f
C17948 VDD.n2930 VSS 0.017108f
C17949 VDD.n2932 VSS 0.011881f
C17950 VDD.n2933 VSS 0.011881f
C17951 VDD.n2934 VSS 0.011881f
C17952 VDD.n2936 VSS 0.015116f
C17953 VDD.n2938 VSS 0.01873f
C17954 VDD.n2939 VSS 0.011881f
C17955 VDD.n2940 VSS 0.011881f
C17956 VDD.n2941 VSS 0.011881f
C17957 VDD.n2943 VSS 0.018345f
C17958 VDD.n2944 VSS 0.014686f
C17959 VDD.n2946 VSS 0.011881f
C17960 VDD.n2947 VSS 0.011881f
C17961 VDD.n2948 VSS 0.011881f
C17962 VDD.n2951 VSS 0.017831f
C17963 VDD.t2897 VSS 0.014219f
C17964 VDD.n2952 VSS 0.022117f
C17965 VDD.n2954 VSS 0.011881f
C17966 VDD.n2955 VSS 0.011881f
C17967 VDD.n2956 VSS 0.011881f
C17968 VDD.n2957 VSS 0.021683f
C17969 VDD.t318 VSS 0.014477f
C17970 VDD.n2958 VSS 0.018218f
C17971 VDD.n2960 VSS 0.011881f
C17972 VDD.n2961 VSS 0.011881f
C17973 VDD.n2962 VSS 0.011881f
C17974 VDD.n2964 VSS 0.011947f
C17975 VDD.n2965 VSS 0.015548f
C17976 VDD.n2968 VSS 0.010911f
C17977 VDD.n2969 VSS 0.013589f
C17978 VDD.n2972 VSS 0.011881f
C17979 VDD.n2973 VSS 0.011881f
C17980 VDD.n2974 VSS 0.011881f
C17981 VDD.t3463 VSS 0.014485f
C17982 VDD.n2975 VSS 0.02085f
C17983 VDD.n2978 VSS 0.011881f
C17984 VDD.n2979 VSS 0.011881f
C17985 VDD.n2980 VSS 0.011881f
C17986 VDD.n2982 VSS 0.010304f
C17987 VDD.t667 VSS 0.015761f
C17988 VDD.n2985 VSS 0.015688f
C17989 VDD.n2987 VSS 0.011881f
C17990 VDD.n2988 VSS 0.011881f
C17991 VDD.t3225 VSS 0.014068f
C17992 VDD.n2990 VSS 0.017988f
C17993 VDD.t687 VSS 0.01455f
C17994 VDD.n2991 VSS 0.022785f
C17995 VDD.n2992 VSS 0.011881f
C17996 VDD.n2993 VSS 0.011881f
C17997 VDD.n2994 VSS 0.011881f
C17998 VDD.n2996 VSS 0.012736f
C17999 VDD.n2999 VSS 0.013218f
C18000 VDD.n3001 VSS 0.011881f
C18001 VDD.n3002 VSS 0.011881f
C18002 VDD.n3003 VSS 0.011881f
C18003 VDD.t679 VSS 0.0127f
C18004 VDD.n3006 VSS 0.011115f
C18005 VDD.n3007 VSS 0.011881f
C18006 VDD.t384 VSS 0.01447f
C18007 VDD.n3009 VSS 0.013391f
C18008 VDD.n3010 VSS 0.011912f
C18009 VDD.t380 VSS 0.014477f
C18010 VDD.n3012 VSS 0.014705f
C18011 VDD.t3440 VSS 0.01449f
C18012 VDD.n3013 VSS 0.017993f
C18013 VDD.n3016 VSS 0.01215f
C18014 VDD.n3017 VSS 0.011881f
C18015 VDD.n3018 VSS 0.011881f
C18016 VDD.n3019 VSS 0.011881f
C18017 VDD.t3793 VSS 0.041965f
C18018 VDD.t20 VSS 0.013232f
C18019 VDD.n3020 VSS 0.01661f
C18020 VDD.n3021 VSS 0.011881f
C18021 VDD.t975 VSS 0.014286f
C18022 VDD.n3022 VSS 0.033371f
C18023 VDD.t235 VSS 0.010055f
C18024 VDD.n3023 VSS 0.016693f
C18025 VDD.t2531 VSS 0.01449f
C18026 VDD.n3024 VSS 0.011881f
C18027 VDD.n3025 VSS 0.010602f
C18028 VDD.t2104 VSS 0.014485f
C18029 VDD.n3026 VSS 0.011881f
C18030 VDD.n3027 VSS 0.010684f
C18031 VDD.n3029 VSS 0.016863f
C18032 VDD.n3031 VSS 0.011881f
C18033 VDD.n3033 VSS 0.020096f
C18034 VDD.n3034 VSS 0.010856f
C18035 VDD.n3035 VSS 0.021333f
C18036 VDD.n3036 VSS 0.011038f
C18037 VDD.n3037 VSS 0.011881f
C18038 VDD.n3038 VSS 0.011881f
C18039 VDD.n3039 VSS 0.011881f
C18040 VDD.n3040 VSS 0.018305f
C18041 VDD.n3041 VSS 0.019645f
C18042 VDD.n3042 VSS 0.035244f
C18043 VDD.t234 VSS 0.010055f
C18044 VDD.n3044 VSS 0.011038f
C18045 VDD.t701 VSS 0.01443f
C18046 VDD.n3045 VSS 0.018713f
C18047 VDD.n3046 VSS 0.011881f
C18048 VDD.n3047 VSS 0.011881f
C18049 VDD.n3049 VSS 0.013089f
C18050 VDD.n3051 VSS 0.013517f
C18051 VDD.n3053 VSS 0.01108f
C18052 VDD.n3055 VSS 0.011881f
C18053 VDD.n3056 VSS 0.011881f
C18054 VDD.n3058 VSS 0.012066f
C18055 VDD.n3059 VSS 0.016338f
C18056 VDD.n3061 VSS 0.011881f
C18057 VDD.n3062 VSS 0.011881f
C18058 VDD.n3063 VSS 0.023326f
C18059 VDD.n3064 VSS 0.038938f
C18060 VDD.t33 VSS 0.035404f
C18061 VDD.t21 VSS 0.051012f
C18062 VDD.t437 VSS 0.032739f
C18063 VDD.t13 VSS 0.036166f
C18064 VDD.t680 VSS 0.032739f
C18065 VDD.t31 VSS 0.031978f
C18066 VDD.t678 VSS 0.032739f
C18067 VDD.t9 VSS 0.04416f
C18068 VDD.t15 VSS 0.06053f
C18069 VDD.t383 VSS 0.032739f
C18070 VDD.t27 VSS 0.031978f
C18071 VDD.t379 VSS 0.032739f
C18072 VDD.t29 VSS 0.038069f
C18073 VDD.t17 VSS 0.065479f
C18074 VDD.t25 VSS 0.035785f
C18075 VDD.t3439 VSS 0.032739f
C18076 VDD.t23 VSS 0.031978f
C18077 VDD.t700 VSS 0.032739f
C18078 VDD.t7 VSS 0.063194f
C18079 VDD.t19 VSS 0.075377f
C18080 VDD.t233 VSS 0.078803f
C18081 VDD.t974 VSS 0.063575f
C18082 VDD.t1251 VSS 0.068524f
C18083 VDD.t3464 VSS 0.043779f
C18084 VDD.t2530 VSS 0.034643f
C18085 VDD.t2103 VSS 0.03845f
C18086 VDD.t694 VSS 0.072712f
C18087 VDD.t2700 VSS 0.103548f
C18088 VDD.t381 VSS 0.051393f
C18089 VDD.t3654 VSS 0.036166f
C18090 VDD.t3710 VSS 0.036546f
C18091 VDD.t2735 VSS 0.02741f
C18092 VDD.t2779 VSS 0.02741f
C18093 VDD.t1883 VSS 0.07157f
C18094 VDD.t3444 VSS 0.081468f
C18095 VDD.t2264 VSS 0.063575f
C18096 VDD.t3652 VSS 0.080706f
C18097 VDD.t1230 VSS 0.059768f
C18098 VDD.t2262 VSS 0.053297f
C18099 VDD.t76 VSS 0.222704f
C18100 VDD.t259 VSS 0.120679f
C18101 VDD.t257 VSS 0.068144f
C18102 VDD.t1163 VSS 0.108116f
C18103 VDD.t1157 VSS 0.103928f
C18104 VDD.t1159 VSS 0.034643f
C18105 VDD.t3749 VSS 0.034643f
C18106 VDD.t1318 VSS 0.033501f
C18107 VDD.t3488 VSS 0.073092f
C18108 VDD.t2634 VSS 0.100121f
C18109 VDD.t645 VSS 0.033501f
C18110 VDD.t3091 VSS 0.035023f
C18111 VDD.t2491 VSS 0.067763f
C18112 VDD.t1317 VSS 0.090985f
C18113 VDD.t331 VSS 0.090223f
C18114 VDD.t3365 VSS 0.054819f
C18115 VDD.t144 VSS 0.074996f
C18116 VDD.t329 VSS 0.094792f
C18117 VDD.t1316 VSS 0.070428f
C18118 VDD.t2492 VSS 0.064717f
C18119 VDD.t1177 VSS 0.073092f
C18120 VDD.t3393 VSS 0.057484f
C18121 VDD.t2992 VSS 0.031978f
C18122 VDD.t2719 VSS 0.02741f
C18123 VDD.t2961 VSS 0.081848f
C18124 VDD.t1175 VSS 0.085275f
C18125 VDD.t1249 VSS 0.047206f
C18126 VDD.t1795 VSS 0.038069f
C18127 VDD.n3065 VSS 0.047313f
C18128 VDD.n3066 VSS 0.023232f
C18129 VDD.n3067 VSS 0.01469f
C18130 VDD.n3069 VSS 0.011881f
C18131 VDD.n3070 VSS 0.011881f
C18132 VDD.n3073 VSS 0.021015f
C18133 VDD.n3074 VSS 0.011881f
C18134 VDD.n3090 VSS 0.500541f
C18135 VDD.n3097 VSS 0.022244f
C18136 VDD.n3100 VSS 0.011881f
C18137 VDD.t2452 VSS 0.015994f
C18138 VDD.n3101 VSS 0.010205f
C18139 VDD.n3103 VSS 0.014361f
C18140 VDD.n3104 VSS 0.011267f
C18141 VDD.n3105 VSS 0.011881f
C18142 VDD.t2456 VSS 0.013927f
C18143 VDD.n3107 VSS 0.011881f
C18144 VDD.n3108 VSS 0.011147f
C18145 VDD.n3111 VSS 0.015663f
C18146 VDD.t161 VSS 0.010137f
C18147 VDD.t3769 VSS 0.021516f
C18148 VDD.n3113 VSS 0.055166f
C18149 VDD.t162 VSS 0.010137f
C18150 VDD.n3114 VSS 0.030049f
C18151 VDD.t3348 VSS 0.010842f
C18152 VDD.n3116 VSS 0.018988f
C18153 VDD.n3117 VSS 0.023013f
C18154 VDD.n3118 VSS 0.011881f
C18155 VDD.t3809 VSS 0.074403f
C18156 VDD.n3119 VSS 0.018814f
C18157 VDD.n3120 VSS 0.011881f
C18158 VDD.n3121 VSS 0.022101f
C18159 VDD.n3123 VSS 0.023316f
C18160 VDD.n3124 VSS 0.011881f
C18161 VDD.t121 VSS 0.010055f
C18162 VDD.n3125 VSS 0.017371f
C18163 VDD.n3126 VSS 0.013668f
C18164 VDD.n3127 VSS 0.011881f
C18165 VDD.n3128 VSS 0.013668f
C18166 VDD.t1733 VSS 0.014745f
C18167 VDD.t2525 VSS 0.014745f
C18168 VDD.n3129 VSS 0.036601f
C18169 VDD.n3130 VSS 0.011881f
C18170 VDD.n3131 VSS 0.013668f
C18171 VDD.n3132 VSS 0.013668f
C18172 VDD.t1406 VSS 0.014745f
C18173 VDD.t2567 VSS 0.014745f
C18174 VDD.n3133 VSS 0.035938f
C18175 VDD.t155 VSS 0.010137f
C18176 VDD.t3813 VSS 0.021516f
C18177 VDD.n3135 VSS 0.055166f
C18178 VDD.t156 VSS 0.010137f
C18179 VDD.n3136 VSS 0.030049f
C18180 VDD.t228 VSS 0.010137f
C18181 VDD.t3777 VSS 0.021516f
C18182 VDD.n3138 VSS 0.055166f
C18183 VDD.t229 VSS 0.010137f
C18184 VDD.n3139 VSS 0.030049f
C18185 VDD.n3140 VSS 0.02678f
C18186 VDD.n3142 VSS 0.053216f
C18187 VDD.n3144 VSS 0.03134f
C18188 VDD.n3146 VSS 0.011881f
C18189 VDD.n3147 VSS 0.011881f
C18190 VDD.n3148 VSS 0.011881f
C18191 VDD.n3150 VSS 0.03134f
C18192 VDD.n3152 VSS 0.011917f
C18193 VDD.n3153 VSS 0.011881f
C18194 VDD.n3154 VSS 0.011881f
C18195 VDD.n3155 VSS 0.015933f
C18196 VDD.n3156 VSS 0.031187f
C18197 VDD.n3157 VSS 0.027967f
C18198 VDD.n3158 VSS 0.011881f
C18199 VDD.n3159 VSS 0.011881f
C18200 VDD.n3160 VSS 0.011881f
C18201 VDD.n3161 VSS 0.023051f
C18202 VDD.n3162 VSS 0.100348f
C18203 VDD.n3163 VSS 0.022712f
C18204 VDD.t120 VSS 0.010055f
C18205 VDD.n3164 VSS 0.01771f
C18206 VDD.n3165 VSS 0.011038f
C18207 VDD.n3166 VSS 0.023665f
C18208 VDD.n3167 VSS 0.023955f
C18209 VDD.n3168 VSS 0.023665f
C18210 VDD.n3170 VSS 0.011062f
C18211 VDD.n3171 VSS 0.014972f
C18212 VDD.n3174 VSS 0.011881f
C18213 VDD.n3175 VSS 0.011881f
C18214 VDD.n3176 VSS 0.011881f
C18215 VDD.t1872 VSS 0.101644f
C18216 VDD.n3180 VSS 0.011881f
C18217 VDD.n3183 VSS 0.011881f
C18218 VDD.n3186 VSS 0.011881f
C18219 VDD.t2226 VSS 0.01592f
C18220 VDD.n3187 VSS 0.018274f
C18221 VDD.n3188 VSS 0.011881f
C18222 VDD.n3190 VSS 0.017713f
C18223 VDD.n3191 VSS 0.011881f
C18224 VDD.n3192 VSS 0.014066f
C18225 VDD.n3193 VSS 0.016065f
C18226 VDD.n3194 VSS 0.011881f
C18227 VDD.n3195 VSS 0.017819f
C18228 VDD.n3196 VSS 0.011881f
C18229 VDD.t2693 VSS 0.014745f
C18230 VDD.n3197 VSS 0.019856f
C18231 VDD.t1894 VSS 0.014485f
C18232 VDD.n3198 VSS 0.011881f
C18233 VDD.t1337 VSS 0.014745f
C18234 VDD.n3199 VSS 0.020336f
C18235 VDD.t469 VSS 0.058246f
C18236 VDD.n3201 VSS 0.011038f
C18237 VDD.n3202 VSS 0.011881f
C18238 VDD.t3788 VSS 0.05912f
C18239 VDD.n3203 VSS 0.066015f
C18240 VDD.n3204 VSS 0.011881f
C18241 VDD.n3205 VSS 0.014361f
C18242 VDD.n3206 VSS 0.011267f
C18243 VDD.n3207 VSS 0.011881f
C18244 VDD.n3208 VSS 0.011881f
C18245 VDD.n3209 VSS 0.010602f
C18246 VDD.n3211 VSS 0.011881f
C18247 VDD.t973 VSS 0.01455f
C18248 VDD.n3213 VSS 0.011881f
C18249 VDD.n3214 VSS 0.011064f
C18250 VDD.t961 VSS 0.014485f
C18251 VDD.n3215 VSS 0.011881f
C18252 VDD.n3216 VSS 0.011881f
C18253 VDD.t3564 VSS 0.01449f
C18254 VDD.n3218 VSS 0.011881f
C18255 VDD.n3220 VSS 0.011881f
C18256 VDD.t344 VSS 0.014218f
C18257 VDD.t2623 VSS 0.01449f
C18258 VDD.n3221 VSS 0.011881f
C18259 VDD.n3222 VSS 0.011881f
C18260 VDD.n3224 VSS 0.011881f
C18261 VDD.t40 VSS 0.0552f
C18262 VDD.t2365 VSS 0.012966f
C18263 VDD.n3229 VSS 0.011775f
C18264 VDD.n3230 VSS 0.011881f
C18265 VDD.n3234 VSS 0.016465f
C18266 VDD.n3235 VSS 0.011881f
C18267 VDD.n3236 VSS 0.011881f
C18268 VDD.n3239 VSS 0.018025f
C18269 VDD.n3240 VSS 0.011881f
C18270 VDD.t839 VSS 0.012738f
C18271 VDD.n3243 VSS 0.016786f
C18272 VDD.n3244 VSS 0.011881f
C18273 VDD.n3246 VSS 0.011881f
C18274 VDD.n3249 VSS 0.01397f
C18275 VDD.n3250 VSS 0.011881f
C18276 VDD.n3251 VSS 0.011064f
C18277 VDD.n3253 VSS 0.010327f
C18278 VDD.n3254 VSS 0.011881f
C18279 VDD.n3256 VSS 0.011881f
C18280 VDD.t996 VSS 0.010806f
C18281 VDD.t2486 VSS 0.0127f
C18282 VDD.n3258 VSS 0.024492f
C18283 VDD.n3259 VSS 0.011881f
C18284 VDD.n3261 VSS 0.011881f
C18285 VDD.n3262 VSS 0.010708f
C18286 VDD.n3263 VSS 0.011881f
C18287 VDD.n3264 VSS 0.010534f
C18288 VDD.t802 VSS 0.015709f
C18289 VDD.t3171 VSS 0.014068f
C18290 VDD.n3265 VSS 0.017805f
C18291 VDD.n3266 VSS 0.011881f
C18292 VDD.n3270 VSS 0.022409f
C18293 VDD.n3271 VSS 0.011881f
C18294 VDD.n3274 VSS 0.013213f
C18295 VDD.n3275 VSS 0.011881f
C18296 VDD.t540 VSS 0.010806f
C18297 VDD.n3278 VSS 0.012268f
C18298 VDD.n3279 VSS 0.011881f
C18299 VDD.n3282 VSS 0.011881f
C18300 VDD.n3285 VSS 0.011881f
C18301 VDD.t2347 VSS 0.015916f
C18302 VDD.n3288 VSS 0.023614f
C18303 VDD.n3289 VSS 0.011881f
C18304 VDD.t1060 VSS 0.013297f
C18305 VDD.t2301 VSS 0.036927f
C18306 VDD.n3293 VSS 0.011881f
C18307 VDD.n3295 VSS 0.011881f
C18308 VDD.t770 VSS 0.015709f
C18309 VDD.n3296 VSS 0.014361f
C18310 VDD.n3297 VSS 0.011267f
C18311 VDD.n3298 VSS 0.011881f
C18312 VDD.n3301 VSS 0.011881f
C18313 VDD.t2478 VSS 0.010846f
C18314 VDD.n3304 VSS 0.011881f
C18315 VDD.n3305 VSS 0.016271f
C18316 VDD.t1740 VSS 0.015709f
C18317 VDD.n3306 VSS 0.029206f
C18318 VDD.n3307 VSS 0.032511f
C18319 VDD.t3820 VSS 0.075443f
C18320 VDD.n3308 VSS 0.126327f
C18321 VDD.t226 VSS 0.010055f
C18322 VDD.n3309 VSS 0.025888f
C18323 VDD.t74 VSS 0.010137f
C18324 VDD.t3789 VSS 0.021516f
C18325 VDD.n3311 VSS 0.055166f
C18326 VDD.t75 VSS 0.010137f
C18327 VDD.n3312 VSS 0.029585f
C18328 VDD.n3313 VSS 0.033748f
C18329 VDD.n3314 VSS 0.011881f
C18330 VDD.n3315 VSS 0.013668f
C18331 VDD.n3316 VSS 0.013668f
C18332 VDD.t1333 VSS 0.014745f
C18333 VDD.t1434 VSS 0.014745f
C18334 VDD.n3317 VSS 0.035938f
C18335 VDD.n3318 VSS 0.019845f
C18336 VDD.t107 VSS 0.222704f
C18337 VDD.t473 VSS 0.120679f
C18338 VDD.t475 VSS 0.068144f
C18339 VDD.t3099 VSS 0.108116f
C18340 VDD.t2286 VSS 0.08832f
C18341 VDD.t218 VSS 0.031978f
C18342 VDD.t2284 VSS 0.051774f
C18343 VDD.t2045 VSS 0.054439f
C18344 VDD.t767 VSS 0.048348f
C18345 VDD.t3164 VSS 0.041114f
C18346 VDD.t3424 VSS 0.031978f
C18347 VDD.t2473 VSS 0.031978f
C18348 VDD.t2303 VSS 0.101644f
C18349 VDD.t872 VSS 0.081848f
C18350 VDD.t769 VSS 0.035023f
C18351 VDD.t2611 VSS 0.067763f
C18352 VDD.t2475 VSS 0.041495f
C18353 VDD.t2489 VSS 0.045302f
C18354 VDD.t2063 VSS 0.04949f
C18355 VDD.t1247 VSS 0.039211f
C18356 VDD.t3666 VSS 0.036927f
C18357 VDD.t3408 VSS 0.080706f
C18358 VDD.t2477 VSS 0.075757f
C18359 VDD.t1054 VSS 0.028171f
C18360 VDD.t1751 VSS 0.036927f
C18361 VDD.t2476 VSS 0.036546f
C18362 VDD.t2060 VSS 0.032739f
C18363 VDD.t2610 VSS 0.037688f
C18364 VDD.t1737 VSS 0.073092f
C18365 VDD.t3361 VSS 0.073092f
C18366 VDD.t1735 VSS 0.113826f
C18367 VDD.t1739 VSS 0.08261f
C18368 VDD.t225 VSS 0.08832f
C18369 VDD.t73 VSS 0.175879f
C18370 VDD.t2086 VSS 0.124486f
C18371 VDD.t1330 VSS 0.068144f
C18372 VDD.t1332 VSS 0.085655f
C18373 VDD.n3319 VSS 0.078512f
C18374 VDD.t219 VSS 0.010137f
C18375 VDD.t3802 VSS 0.021516f
C18376 VDD.n3321 VSS 0.055166f
C18377 VDD.t220 VSS 0.010137f
C18378 VDD.n3322 VSS 0.030049f
C18379 VDD.n3323 VSS 0.013523f
C18380 VDD.t2287 VSS 0.014469f
C18381 VDD.n3324 VSS 0.031602f
C18382 VDD.n3325 VSS 0.013668f
C18383 VDD.n3326 VSS 0.013668f
C18384 VDD.n3327 VSS 0.03134f
C18385 VDD.t108 VSS 0.010137f
C18386 VDD.t3797 VSS 0.021516f
C18387 VDD.n3329 VSS 0.055166f
C18388 VDD.t109 VSS 0.010137f
C18389 VDD.n3330 VSS 0.030049f
C18390 VDD.t206 VSS 0.010137f
C18391 VDD.t3816 VSS 0.021516f
C18392 VDD.n3332 VSS 0.055166f
C18393 VDD.t207 VSS 0.010137f
C18394 VDD.n3333 VSS 0.030049f
C18395 VDD.n3334 VSS 0.02678f
C18396 VDD.t2212 VSS 0.014745f
C18397 VDD.t474 VSS 0.014745f
C18398 VDD.n3336 VSS 0.035938f
C18399 VDD.n3338 VSS 0.053216f
C18400 VDD.n3339 VSS 0.011881f
C18401 VDD.n3340 VSS 0.01978f
C18402 VDD.n3342 VSS 0.017356f
C18403 VDD.n3343 VSS 0.023851f
C18404 VDD.n3344 VSS 0.019778f
C18405 VDD.n3345 VSS 0.011881f
C18406 VDD.n3346 VSS 0.011881f
C18407 VDD.n3348 VSS 0.03134f
C18408 VDD.n3350 VSS 0.023665f
C18409 VDD.n3351 VSS 0.023955f
C18410 VDD.n3352 VSS 0.023665f
C18411 VDD.n3353 VSS 0.011881f
C18412 VDD.n3354 VSS 0.021526f
C18413 VDD.n3355 VSS 0.022727f
C18414 VDD.n3356 VSS 0.024238f
C18415 VDD.t227 VSS 0.010055f
C18416 VDD.n3357 VSS 0.01771f
C18417 VDD.n3359 VSS 0.014367f
C18418 VDD.n3361 VSS 0.011881f
C18419 VDD.n3362 VSS 0.011881f
C18420 VDD.n3363 VSS 0.011881f
C18421 VDD.n3367 VSS 0.015964f
C18422 VDD.n3368 VSS 0.011881f
C18423 VDD.n3369 VSS 0.011881f
C18424 VDD.n3370 VSS 0.011881f
C18425 VDD.n3372 VSS 0.011101f
C18426 VDD.n3375 VSS 0.011881f
C18427 VDD.n3376 VSS 0.011881f
C18428 VDD.n3379 VSS 0.021309f
C18429 VDD.n3381 VSS 0.011881f
C18430 VDD.n3382 VSS 0.011881f
C18431 VDD.n3384 VSS 0.010708f
C18432 VDD.n3391 VSS 0.011881f
C18433 VDD.n3392 VSS 0.011881f
C18434 VDD.n3393 VSS 0.011881f
C18435 VDD.t2387 VSS 0.015709f
C18436 VDD.n3394 VSS 0.021309f
C18437 VDD.t2121 VSS 0.010806f
C18438 VDD.n3396 VSS 0.010826f
C18439 VDD.n3397 VSS 0.011881f
C18440 VDD.n3399 VSS 0.011881f
C18441 VDD.n3402 VSS 0.011881f
C18442 VDD.t1394 VSS 0.014477f
C18443 VDD.n3405 VSS 0.011881f
C18444 VDD.t1400 VSS 0.014204f
C18445 VDD.n3406 VSS 0.014772f
C18446 VDD.n3408 VSS 0.013261f
C18447 VDD.n3409 VSS 0.011064f
C18448 VDD.n3410 VSS 0.011881f
C18449 VDD.t1347 VSS 0.014194f
C18450 VDD.t1825 VSS 0.01383f
C18451 VDD.n3411 VSS 0.016273f
C18452 VDD.n3412 VSS 0.011881f
C18453 VDD.t2186 VSS 0.0127f
C18454 VDD.n3414 VSS 0.010162f
C18455 VDD.n3415 VSS 0.015637f
C18456 VDD.n3416 VSS 0.011881f
C18457 VDD.n3417 VSS 0.011881f
C18458 VDD.n3420 VSS 0.018848f
C18459 VDD.n3422 VSS 0.011881f
C18460 VDD.n3423 VSS 0.011881f
C18461 VDD.n3424 VSS 0.011881f
C18462 VDD.n3426 VSS 0.012328f
C18463 VDD.n3429 VSS 0.01309f
C18464 VDD.n3430 VSS 0.011881f
C18465 VDD.n3431 VSS 0.011881f
C18466 VDD.n3432 VSS 0.011881f
C18467 VDD.n3433 VSS 0.018196f
C18468 VDD.n3437 VSS 0.011881f
C18469 VDD.n3438 VSS 0.011881f
C18470 VDD.n3439 VSS 0.011881f
C18471 VDD.n3440 VSS 0.018882f
C18472 VDD.n3442 VSS 0.010843f
C18473 VDD.n3444 VSS 0.011881f
C18474 VDD.n3445 VSS 0.011881f
C18475 VDD.t3323 VSS 0.010846f
C18476 VDD.n3448 VSS 0.022439f
C18477 VDD.n3449 VSS 0.011881f
C18478 VDD.n3450 VSS 0.011881f
C18479 VDD.n3451 VSS 0.011881f
C18480 VDD.n3456 VSS 0.011881f
C18481 VDD.n3457 VSS 0.011881f
C18482 VDD.n3459 VSS 0.010708f
C18483 VDD.n3461 VSS 0.012208f
C18484 VDD.n3463 VSS 0.011881f
C18485 VDD.n3464 VSS 0.011881f
C18486 VDD.n3465 VSS 0.011881f
C18487 VDD.n3466 VSS 0.025155f
C18488 VDD.n3467 VSS 0.039301f
C18489 VDD.t2463 VSS 0.053297f
C18490 VDD.t2386 VSS 0.037688f
C18491 VDD.t2120 VSS 0.081848f
C18492 VDD.t2616 VSS 0.074996f
C18493 VDD.t3418 VSS 0.031978f
C18494 VDD.t3416 VSS 0.036927f
C18495 VDD.t2122 VSS 0.041114f
C18496 VDD.t2384 VSS 0.053297f
C18497 VDD.t2464 VSS 0.031978f
C18498 VDD.t2344 VSS 0.037688f
C18499 VDD.t2302 VSS 0.032739f
C18500 VDD.t2340 VSS 0.035023f
C18501 VDD.t1413 VSS 0.037688f
C18502 VDD.t3322 VSS 0.082229f
C18503 VDD.t3410 VSS 0.094411f
C18504 VDD.t2461 VSS 0.036927f
C18505 VDD.t1563 VSS 0.031978f
C18506 VDD.t3153 VSS 0.053297f
C18507 VDD.t2343 VSS 0.072331f
C18508 VDD.t1393 VSS 0.037688f
C18509 VDD.t2345 VSS 0.031978f
C18510 VDD.t1399 VSS 0.035023f
C18511 VDD.t2785 VSS 0.072712f
C18512 VDD.t3520 VSS 0.101644f
C18513 VDD.t2341 VSS 0.037688f
C18514 VDD.t2378 VSS 0.031978f
C18515 VDD.t3155 VSS 0.035785f
C18516 VDD.t1193 VSS 0.041876f
C18517 VDD.t1693 VSS 0.06624f
C18518 VDD.t1346 VSS 0.036546f
C18519 VDD.t3764 VSS 0.07157f
C18520 VDD.t1824 VSS 0.098599f
C18521 VDD.t2271 VSS 0.036166f
C18522 VDD.t1522 VSS 0.036166f
C18523 VDD.t2183 VSS 0.044921f
C18524 VDD.t1793 VSS 0.031978f
C18525 VDD.t2185 VSS 0.038069f
C18526 VDD.t1955 VSS 0.053297f
C18527 VDD.t2364 VSS 0.034643f
C18528 VDD.t2366 VSS 0.034262f
C18529 VDD.t3632 VSS 0.032739f
C18530 VDD.t3501 VSS 0.035404f
C18531 VDD.t3312 VSS 0.032739f
C18532 VDD.t3503 VSS 0.057865f
C18533 VDD.t2951 VSS 0.075377f
C18534 VDD.t1644 VSS 0.047206f
C18535 VDD.t1724 VSS 0.032739f
C18536 VDD.t1645 VSS 0.031978f
C18537 VDD.t3194 VSS 0.032739f
C18538 VDD.t1368 VSS 0.065098f
C18539 VDD.t1366 VSS 0.039211f
C18540 VDD.t643 VSS 0.042637f
C18541 VDD.t247 VSS 0.070047f
C18542 VDD.t838 VSS 0.035404f
C18543 VDD.t3318 VSS 0.031978f
C18544 VDD.t836 VSS 0.057865f
C18545 VDD.t2941 VSS 0.036166f
C18546 VDD.t1997 VSS 0.047206f
C18547 VDD.t1745 VSS 0.070428f
C18548 VDD.t3196 VSS 0.068524f
C18549 VDD.t3157 VSS 0.068524f
C18550 VDD.t1624 VSS 0.035404f
C18551 VDD.t2299 VSS 0.041114f
C18552 VDD.t3290 VSS 0.073473f
C18553 VDD.t3622 VSS 0.06053f
C18554 VDD.t291 VSS 0.036546f
C18555 VDD.t3304 VSS 0.035023f
C18556 VDD.t994 VSS 0.036546f
C18557 VDD.t1447 VSS 0.037688f
C18558 VDD.t1626 VSS 0.077661f
C18559 VDD.t2155 VSS 0.074235f
C18560 VDD.t3086 VSS 0.036927f
C18561 VDD.t1843 VSS 0.036166f
C18562 VDD.t2487 VSS 0.052155f
C18563 VDD.t2485 VSS 0.054819f
C18564 VDD.t995 VSS 0.053297f
C18565 VDD.n3468 VSS 0.04425f
C18566 VDD.t1627 VSS 0.039972f
C18567 VDD.t993 VSS 0.046063f
C18568 VDD.t245 VSS 0.031978f
C18569 VDD.t799 VSS 0.059768f
C18570 VDD.t1839 VSS 0.052916f
C18571 VDD.t579 VSS 0.031978f
C18572 VDD.t797 VSS 0.02741f
C18573 VDD.t3629 VSS 0.043399f
C18574 VDD.t1358 VSS 0.073473f
C18575 VDD.t580 VSS 0.03845f
C18576 VDD.t801 VSS 0.072712f
C18577 VDD.t3166 VSS 0.07195f
C18578 VDD.t3170 VSS 0.031978f
C18579 VDD.t536 VSS 0.032739f
C18580 VDD.t3216 VSS 0.033881f
C18581 VDD.t3212 VSS 0.065479f
C18582 VDD.t3168 VSS 0.065479f
C18583 VDD.t1087 VSS 0.035023f
C18584 VDD.t3505 VSS 0.032739f
C18585 VDD.t1075 VSS 0.035023f
C18586 VDD.t2483 VSS 0.032739f
C18587 VDD.t1067 VSS 0.037688f
C18588 VDD.t535 VSS 0.032739f
C18589 VDD.t1089 VSS 0.053297f
C18590 VDD.t2816 VSS 0.032739f
C18591 VDD.t1073 VSS 0.035404f
C18592 VDD.t1071 VSS 0.034262f
C18593 VDD.t3412 VSS 0.032739f
C18594 VDD.t1069 VSS 0.063956f
C18595 VDD.t1079 VSS 0.043779f
C18596 VDD.t539 VSS 0.032359f
C18597 VDD.t1065 VSS 0.037688f
C18598 VDD.t538 VSS 0.032739f
C18599 VDD.t1077 VSS 0.032739f
C18600 VDD.t2484 VSS 0.032739f
C18601 VDD.t1061 VSS 0.031978f
C18602 VDD.t2348 VSS 0.032739f
C18603 VDD.t1083 VSS 0.041114f
C18604 VDD.t3353 VSS 0.032739f
C18605 VDD.t1085 VSS 0.031978f
C18606 VDD.t2818 VSS 0.032739f
C18607 VDD.t1063 VSS 0.042257f
C18608 VDD.t1081 VSS 0.065479f
C18609 VDD.t1059 VSS 0.039592f
C18610 VDD.t2346 VSS 0.060149f
C18611 VDD.n3469 VSS 0.096024f
C18612 VDD.n3470 VSS 0.024904f
C18613 VDD.n3471 VSS 0.015764f
C18614 VDD.n3472 VSS 0.011881f
C18615 VDD.n3473 VSS 0.011881f
C18616 VDD.n3474 VSS 0.011881f
C18617 VDD.n3476 VSS 0.010528f
C18618 VDD.n3479 VSS 0.011785f
C18619 VDD.n3480 VSS 0.011881f
C18620 VDD.n3481 VSS 0.011881f
C18621 VDD.n3483 VSS 0.014724f
C18622 VDD.n3485 VSS 0.01148f
C18623 VDD.n3487 VSS 0.011881f
C18624 VDD.n3488 VSS 0.011881f
C18625 VDD.n3490 VSS 0.013213f
C18626 VDD.n3492 VSS 0.011207f
C18627 VDD.n3494 VSS 0.011881f
C18628 VDD.n3495 VSS 0.011881f
C18629 VDD.n3498 VSS 0.013213f
C18630 VDD.n3500 VSS 0.011881f
C18631 VDD.n3501 VSS 0.011881f
C18632 VDD.n3502 VSS 0.011881f
C18633 VDD.n3504 VSS 0.015309f
C18634 VDD.n3505 VSS 0.012941f
C18635 VDD.n3506 VSS 0.011881f
C18636 VDD.n3507 VSS 0.011881f
C18637 VDD.n3508 VSS 0.011881f
C18638 VDD.n3510 VSS 0.021309f
C18639 VDD.n3512 VSS 0.013629f
C18640 VDD.n3514 VSS 0.011881f
C18641 VDD.n3515 VSS 0.011881f
C18642 VDD.n3517 VSS 0.011385f
C18643 VDD.n3519 VSS 0.020351f
C18644 VDD.n3520 VSS 0.011881f
C18645 VDD.n3521 VSS 0.011881f
C18646 VDD.n3522 VSS 0.011881f
C18647 VDD.n3525 VSS 0.012071f
C18648 VDD.n3529 VSS 0.016366f
C18649 VDD.n3530 VSS 0.011881f
C18650 VDD.n3531 VSS 0.011881f
C18651 VDD.n3532 VSS 0.011881f
C18652 VDD.n3536 VSS 0.011881f
C18653 VDD.n3537 VSS 0.011881f
C18654 VDD.n3541 VSS 0.018196f
C18655 VDD.n3542 VSS 0.011881f
C18656 VDD.n3543 VSS 0.011881f
C18657 VDD.n3544 VSS 0.011881f
C18658 VDD.n3546 VSS 0.013384f
C18659 VDD.n3548 VSS 0.016663f
C18660 VDD.n3549 VSS 0.011881f
C18661 VDD.n3550 VSS 0.011881f
C18662 VDD.n3552 VSS 0.013828f
C18663 VDD.n3553 VSS 0.01174f
C18664 VDD.n3554 VSS 0.011881f
C18665 VDD.n3555 VSS 0.011881f
C18666 VDD.n3556 VSS 0.011881f
C18667 VDD.n3558 VSS 0.013384f
C18668 VDD.t3504 VSS 0.01383f
C18669 VDD.n3560 VSS 0.014494f
C18670 VDD.n3562 VSS 0.011881f
C18671 VDD.n3563 VSS 0.011881f
C18672 VDD.n3565 VSS 0.017065f
C18673 VDD.n3566 VSS 0.011397f
C18674 VDD.n3567 VSS 0.011881f
C18675 VDD.n3568 VSS 0.011881f
C18676 VDD.n3569 VSS 0.011881f
C18677 VDD.n3570 VSS 0.012244f
C18678 VDD.n3571 VSS 0.012328f
C18679 VDD.t1870 VSS 0.01449f
C18680 VDD.n3572 VSS 0.011881f
C18681 VDD.n3573 VSS 0.014361f
C18682 VDD.n3576 VSS 0.011881f
C18683 VDD.n3578 VSS 0.010602f
C18684 VDD.n3579 VSS 0.012f
C18685 VDD.n3580 VSS 0.011881f
C18686 VDD.t3277 VSS 0.01447f
C18687 VDD.n3581 VSS 0.01693f
C18688 VDD.n3582 VSS 0.011881f
C18689 VDD.n3583 VSS 0.012244f
C18690 VDD.n3584 VSS 0.012283f
C18691 VDD.n3586 VSS 0.011881f
C18692 VDD.n3587 VSS 0.014361f
C18693 VDD.n3590 VSS 0.011881f
C18694 VDD.n3591 VSS 0.011881f
C18695 VDD.n3592 VSS 0.011881f
C18696 VDD.n3593 VSS 0.013759f
C18697 VDD.n3594 VSS 0.019212f
C18698 VDD.n3596 VSS 0.011267f
C18699 VDD.n3598 VSS 0.011881f
C18700 VDD.n3599 VSS 0.011881f
C18701 VDD.n3600 VSS 0.011881f
C18702 VDD.n3601 VSS 0.018619f
C18703 VDD.t955 VSS 0.012738f
C18704 VDD.n3603 VSS 0.014262f
C18705 VDD.n3604 VSS 0.011881f
C18706 VDD.n3605 VSS 0.011881f
C18707 VDD.n3606 VSS 0.011881f
C18708 VDD.t3273 VSS 0.014477f
C18709 VDD.n3608 VSS 0.018882f
C18710 VDD.n3610 VSS 0.011881f
C18711 VDD.n3611 VSS 0.011881f
C18712 VDD.n3612 VSS 0.011881f
C18713 VDD.t1581 VSS 0.01455f
C18714 VDD.n3616 VSS 0.024248f
C18715 VDD.n3617 VSS 0.011881f
C18716 VDD.n3618 VSS 0.011881f
C18717 VDD.n3619 VSS 0.011881f
C18718 VDD.n3620 VSS 0.013759f
C18719 VDD.n3621 VSS 0.019212f
C18720 VDD.n3624 VSS 0.011881f
C18721 VDD.n3625 VSS 0.011881f
C18722 VDD.n3626 VSS 0.011881f
C18723 VDD.n3627 VSS 0.021935f
C18724 VDD.t3315 VSS 0.014485f
C18725 VDD.n3629 VSS 0.02085f
C18726 VDD.n3630 VSS 0.011881f
C18727 VDD.n3631 VSS 0.011881f
C18728 VDD.n3632 VSS 0.011881f
C18729 VDD.n3633 VSS 0.024629f
C18730 VDD.n3634 VSS 0.148179f
C18731 VDD.t3314 VSS 0.088701f
C18732 VDD.t1579 VSS 0.031978f
C18733 VDD.t1869 VSS 0.032739f
C18734 VDD.t1225 VSS 0.040734f
C18735 VDD.t1279 VSS 0.07195f
C18736 VDD.t1199 VSS 0.045683f
C18737 VDD.t3023 VSS 0.041495f
C18738 VDD.t2706 VSS 0.036546f
C18739 VDD.t2628 VSS 0.039211f
C18740 VDD.t2714 VSS 0.048348f
C18741 VDD.t2602 VSS 0.081468f
C18742 VDD.t1888 VSS 0.07728f
C18743 VDD.t1580 VSS 0.02741f
C18744 VDD.t2708 VSS 0.02741f
C18745 VDD.t1875 VSS 0.036546f
C18746 VDD.t2704 VSS 0.041114f
C18747 VDD.t3296 VSS 0.059007f
C18748 VDD.t3316 VSS 0.106974f
C18749 VDD.t3272 VSS 0.097837f
C18750 VDD.t3276 VSS 0.104309f
C18751 VDD.t954 VSS 0.072712f
C18752 VDD.t1278 VSS 0.031978f
C18753 VDD.t952 VSS 0.032739f
C18754 VDD.t39 VSS 0.036166f
C18755 VDD.t1863 VSS 0.039592f
C18756 VDD.t531 VSS 0.050251f
C18757 VDD.t3029 VSS 0.067382f
C18758 VDD.t765 VSS 0.036546f
C18759 VDD.t2665 VSS 0.041495f
C18760 VDD.t1701 VSS 0.048348f
C18761 VDD.t1129 VSS 0.039211f
C18762 VDD.t764 VSS 0.098979f
C18763 VDD.t3641 VSS 0.108877f
C18764 VDD.t1747 VSS 0.029694f
C18765 VDD.t2573 VSS 0.09936f
C18766 VDD.t197 VSS 0.101644f
C18767 VDD.t2751 VSS 0.069286f
C18768 VDD.t3130 VSS 0.138571f
C18769 VDD.t841 VSS 0.148088f
C18770 VDD.t1141 VSS 0.063575f
C18771 VDD.t1492 VSS 0.039211f
C18772 VDD.t1885 VSS 0.041114f
C18773 VDD.t1348 VSS 0.065098f
C18774 VDD.t755 VSS 0.057484f
C18775 VDD.t840 VSS 0.02741f
C18776 VDD.t972 VSS 0.02741f
C18777 VDD.t1143 VSS 0.052916f
C18778 VDD.t1139 VSS 0.055961f
C18779 VDD.t2590 VSS 0.057103f
C18780 VDD.t3298 VSS 0.069666f
C18781 VDD.t960 VSS 0.035785f
C18782 VDD.t516 VSS 0.031978f
C18783 VDD.t3563 VSS 0.036546f
C18784 VDD.t958 VSS 0.044921f
C18785 VDD.t2624 VSS 0.134764f
C18786 VDD.t343 VSS 0.125628f
C18787 VDD.t3562 VSS 0.031978f
C18788 VDD.t2622 VSS 0.041114f
C18789 VDD.t876 VSS 0.125628f
C18790 VDD.t1703 VSS 0.123344f
C18791 VDD.n3635 VSS 0.043108f
C18792 VDD.n3636 VSS 0.024103f
C18793 VDD.n3637 VSS 0.011881f
C18794 VDD.n3638 VSS 0.011881f
C18795 VDD.n3639 VSS 0.011881f
C18796 VDD.n3641 VSS 0.015843f
C18797 VDD.n3642 VSS 0.021638f
C18798 VDD.n3644 VSS 0.021505f
C18799 VDD.t3243 VSS 0.014212f
C18800 VDD.n3645 VSS 0.017831f
C18801 VDD.n3647 VSS 0.011881f
C18802 VDD.n3648 VSS 0.011881f
C18803 VDD.n3649 VSS 0.011881f
C18804 VDD.n3651 VSS 0.021089f
C18805 VDD.n3652 VSS 0.012748f
C18806 VDD.n3653 VSS 0.019707f
C18807 VDD.n3654 VSS 0.018242f
C18808 VDD.n3657 VSS 0.023196f
C18809 VDD.n3658 VSS 0.011881f
C18810 VDD.n3659 VSS 0.011881f
C18811 VDD.n3660 VSS 0.011881f
C18812 VDD.n3662 VSS 0.012f
C18813 VDD.n3665 VSS 0.011881f
C18814 VDD.n3666 VSS 0.011881f
C18815 VDD.n3670 VSS 0.023316f
C18816 VDD.t198 VSS 0.010055f
C18817 VDD.n3671 VSS 0.017371f
C18818 VDD.n3672 VSS 0.011917f
C18819 VDD.n3673 VSS 0.011881f
C18820 VDD.n3674 VSS 0.011881f
C18821 VDD.n3675 VSS 0.011881f
C18822 VDD.n3676 VSS 0.031187f
C18823 VDD.n3677 VSS 0.027967f
C18824 VDD.n3678 VSS 0.022101f
C18825 VDD.t199 VSS 0.010055f
C18826 VDD.n3679 VSS 0.01771f
C18827 VDD.n3680 VSS 0.017797f
C18828 VDD.n3681 VSS 0.011881f
C18829 VDD.n3682 VSS 0.011881f
C18830 VDD.n3683 VSS 0.011881f
C18831 VDD.n3684 VSS 0.014361f
C18832 VDD.t472 VSS 0.010846f
C18833 VDD.n3685 VSS 0.015964f
C18834 VDD.n3686 VSS 0.011881f
C18835 VDD.n3688 VSS 0.010333f
C18836 VDD.n3689 VSS 0.011881f
C18837 VDD.t2014 VSS 0.014414f
C18838 VDD.n3693 VSS 0.011881f
C18839 VDD.n3696 VSS 0.011881f
C18840 VDD.n3697 VSS 0.014066f
C18841 VDD.n3698 VSS 0.016065f
C18842 VDD.n3699 VSS 0.011881f
C18843 VDD.n3701 VSS 0.014498f
C18844 VDD.n3702 VSS 0.011881f
C18845 VDD.n3703 VSS 0.010563f
C18846 VDD.n3704 VSS 0.013523f
C18847 VDD.n3705 VSS 0.011881f
C18848 VDD.n3706 VSS 0.011881f
C18849 VDD.n3708 VSS 0.015061f
C18850 VDD.n3711 VSS 0.011881f
C18851 VDD.n3712 VSS 0.011881f
C18852 VDD.n3713 VSS 0.011881f
C18853 VDD.t342 VSS 0.01455f
C18854 VDD.n3714 VSS 0.033274f
C18855 VDD.n3717 VSS 0.011881f
C18856 VDD.n3718 VSS 0.011881f
C18857 VDD.n3721 VSS 0.013652f
C18858 VDD.n3723 VSS 0.011881f
C18859 VDD.n3724 VSS 0.011881f
C18860 VDD.t2016 VSS 0.014429f
C18861 VDD.t934 VSS 0.014483f
C18862 VDD.n3727 VSS 0.032636f
C18863 VDD.n3728 VSS 0.011881f
C18864 VDD.n3729 VSS 0.011881f
C18865 VDD.n3730 VSS 0.011881f
C18866 VDD.t932 VSS 0.015916f
C18867 VDD.n3731 VSS 0.038286f
C18868 VDD.n3733 VSS 0.010708f
C18869 VDD.n3735 VSS 0.011881f
C18870 VDD.n3736 VSS 0.011881f
C18871 VDD.n3737 VSS 0.011881f
C18872 VDD.n3741 VSS 0.011881f
C18873 VDD.n3742 VSS 0.011881f
C18874 VDD.n3743 VSS 0.011881f
C18875 VDD.n3745 VSS 0.011267f
C18876 VDD.n3748 VSS 0.011101f
C18877 VDD.n3750 VSS 0.011881f
C18878 VDD.n3751 VSS 0.011881f
C18879 VDD.n3752 VSS 0.011881f
C18880 VDD.n3753 VSS 0.025079f
C18881 VDD.n3754 VSS 0.04425f
C18882 VDD.t2753 VSS 0.067763f
C18883 VDD.t2733 VSS 0.090223f
C18884 VDD.t2978 VSS 0.055581f
C18885 VDD.t2382 VSS 0.060149f
C18886 VDD.t2007 VSS 0.056342f
C18887 VDD.t471 VSS 0.039211f
C18888 VDD.t1489 VSS 0.037688f
C18889 VDD.t2754 VSS 0.046063f
C18890 VDD.t470 VSS 0.064717f
C18891 VDD.t929 VSS 0.035404f
C18892 VDD.t1504 VSS 0.030836f
C18893 VDD.t1565 VSS 0.037688f
C18894 VDD.t2974 VSS 0.036546f
C18895 VDD.t2002 VSS 0.031978f
C18896 VDD.t2585 VSS 0.087559f
C18897 VDD.t931 VSS 0.084132f
C18898 VDD.t2013 VSS 0.031978f
C18899 VDD.t933 VSS 0.031978f
C18900 VDD.t2015 VSS 0.092127f
C18901 VDD.t361 VSS 0.126389f
C18902 VDD.t2729 VSS 0.063956f
C18903 VDD.t3483 VSS 0.029694f
C18904 VDD.t1498 VSS 0.034262f
C18905 VDD.t1787 VSS 0.073092f
C18906 VDD.t1135 VSS 0.047206f
C18907 VDD.t1880 VSS 0.045302f
C18908 VDD.t359 VSS 0.080706f
C18909 VDD.t588 VSS 0.043399f
C18910 VDD.t341 VSS 0.029313f
C18911 VDD.t3258 VSS 0.068524f
C18912 VDD.t3476 VSS 0.042257f
C18913 VDD.t1857 VSS 0.037308f
C18914 VDD.t1334 VSS 0.039972f
C18915 VDD.t423 VSS 0.031978f
C18916 VDD.t1336 VSS 0.081848f
C18917 VDD.t429 VSS 0.081468f
C18918 VDD.t3241 VSS 0.036166f
C18919 VDD.t1127 VSS 0.063956f
C18920 VDD.t375 VSS 0.085275f
C18921 VDD.t385 VSS 0.084894f
C18922 VDD.t2826 VSS 0.041114f
C18923 VDD.t3691 VSS 0.036927f
C18924 VDD.t3684 VSS 0.066621f
C18925 VDD.t2828 VSS 0.070808f
C18926 VDD.t3337 VSS 0.03845f
C18927 VDD.t3486 VSS 0.073854f
C18928 VDD.t1817 VSS 0.072712f
C18929 VDD.t2225 VSS 0.032359f
C18930 VDD.t2292 VSS 0.032739f
C18931 VDD.t2221 VSS 0.032739f
C18932 VDD.t1569 VSS 0.032739f
C18933 VDD.t2223 VSS 0.034262f
C18934 VDD.t2227 VSS 0.069286f
C18935 VDD.t3282 VSS 0.039592f
C18936 VDD.t760 VSS 0.040353f
C18937 VDD.t431 VSS 0.073473f
C18938 VDD.t3443 VSS 0.048348f
C18939 VDD.t2725 VSS 0.02741f
C18940 VDD.t759 VSS 0.041114f
C18941 VDD.t1781 VSS 0.057865f
C18942 VDD.t319 VSS 0.045683f
C18943 VDD.t1915 VSS 0.085275f
C18944 VDD.t3728 VSS 0.107735f
C18945 VDD.t2694 VSS 0.068144f
C18946 VDD.t2692 VSS 0.033881f
C18947 VDD.t1893 VSS 0.033881f
C18948 VDD.t2388 VSS 0.086797f
C18949 VDD.n3755 VSS 0.115059f
C18950 VDD.n3756 VSS 0.023851f
C18951 VDD.t2389 VSS 0.01449f
C18952 VDD.n3757 VSS 0.02086f
C18953 VDD.n3758 VSS 0.011881f
C18954 VDD.n3759 VSS 0.011881f
C18955 VDD.n3760 VSS 0.011881f
C18956 VDD.n3761 VSS 0.019387f
C18957 VDD.n3762 VSS 0.013668f
C18958 VDD.n3763 VSS 0.017866f
C18959 VDD.n3765 VSS 0.011881f
C18960 VDD.n3766 VSS 0.011881f
C18961 VDD.n3768 VSS 0.012435f
C18962 VDD.n3771 VSS 0.011881f
C18963 VDD.n3772 VSS 0.011881f
C18964 VDD.n3775 VSS 0.010736f
C18965 VDD.n3776 VSS 0.016317f
C18966 VDD.n3777 VSS 0.011881f
C18967 VDD.n3778 VSS 0.011881f
C18968 VDD.n3779 VSS 0.011881f
C18969 VDD.n3783 VSS 0.023899f
C18970 VDD.n3785 VSS 0.011881f
C18971 VDD.n3786 VSS 0.011881f
C18972 VDD.n3787 VSS 0.011881f
C18973 VDD.t3487 VSS 0.013749f
C18974 VDD.n3788 VSS 0.019132f
C18975 VDD.t3685 VSS 0.01447f
C18976 VDD.n3792 VSS 0.017588f
C18977 VDD.n3793 VSS 0.011881f
C18978 VDD.n3794 VSS 0.011881f
C18979 VDD.n3795 VSS 0.011881f
C18980 VDD.t3692 VSS 0.014373f
C18981 VDD.n3796 VSS 0.02836f
C18982 VDD.n3799 VSS 0.011881f
C18983 VDD.n3800 VSS 0.011881f
C18984 VDD.n3806 VSS 0.011881f
C18985 VDD.n3807 VSS 0.011881f
C18986 VDD.n3808 VSS 0.011881f
C18987 VDD.n3809 VSS 0.014361f
C18988 VDD.n3810 VSS 0.011267f
C18989 VDD.n3811 VSS 0.011881f
C18990 VDD.t374 VSS 0.014485f
C18991 VDD.t3260 VSS 0.01449f
C18992 VDD.n3812 VSS 0.021089f
C18993 VDD.n3813 VSS 0.011881f
C18994 VDD.n3815 VSS 0.010911f
C18995 VDD.n3816 VSS 0.010783f
C18996 VDD.n3818 VSS 0.011881f
C18997 VDD.n3819 VSS 0.011427f
C18998 VDD.n3820 VSS 0.016823f
C18999 VDD.n3823 VSS 0.011881f
C19000 VDD.n3825 VSS 0.014537f
C19001 VDD.n3826 VSS 0.011064f
C19002 VDD.n3827 VSS 0.027891f
C19003 VDD.t3768 VSS 0.041965f
C19004 VDD.n3829 VSS 0.015593f
C19005 VDD.n3830 VSS 0.037956f
C19006 VDD.t125 VSS 0.010055f
C19007 VDD.n3832 VSS 0.011917f
C19008 VDD.n3834 VSS 0.011881f
C19009 VDD.n3835 VSS 0.011881f
C19010 VDD.n3836 VSS 0.011881f
C19011 VDD.n3838 VSS 0.013891f
C19012 VDD.n3840 VSS 0.011881f
C19013 VDD.n3841 VSS 0.011881f
C19014 VDD.n3842 VSS 0.011881f
C19015 VDD.n3847 VSS 0.011881f
C19016 VDD.n3848 VSS 0.011881f
C19017 VDD.n3849 VSS 0.011881f
C19018 VDD.n3851 VSS 0.014565f
C19019 VDD.n3852 VSS 0.01368f
C19020 VDD.n3854 VSS 0.013228f
C19021 VDD.n3855 VSS 0.011881f
C19022 VDD.n3856 VSS 0.011881f
C19023 VDD.n3857 VSS 0.011881f
C19024 VDD.n3859 VSS 0.02085f
C19025 VDD.n3861 VSS 0.011881f
C19026 VDD.n3862 VSS 0.011881f
C19027 VDD.n3864 VSS 0.025155f
C19028 VDD.n3865 VSS 0.045773f
C19029 VDD.t377 VSS 0.051774f
C19030 VDD.t1385 VSS 0.113065f
C19031 VDD.t373 VSS 0.098218f
C19032 VDD.t3763 VSS 0.031978f
C19033 VDD.t3259 VSS 0.036546f
C19034 VDD.t1797 VSS 0.067763f
C19035 VDD.t824 VSS 0.06091f
C19036 VDD.t2588 VSS 0.035785f
C19037 VDD.t53 VSS 0.040734f
C19038 VDD.t3435 VSS 0.037688f
C19039 VDD.t2471 VSS 0.031978f
C19040 VDD.t371 VSS 0.06053f
C19041 VDD.t3712 VSS 0.065859f
C19042 VDD.t1417 VSS 0.065479f
C19043 VDD.t1421 VSS 0.063956f
C19044 VDD.t3008 VSS 0.042637f
C19045 VDD.t3762 VSS 0.051774f
C19046 VDD.t2090 VSS 0.06624f
C19047 VDD.t3640 VSS 0.036546f
C19048 VDD.t2723 VSS 0.039211f
C19049 VDD.t1419 VSS 0.035785f
C19050 VDD.t727 VSS 0.041114f
C19051 VDD.t3508 VSS 0.038069f
C19052 VDD.t349 VSS 0.089462f
C19053 VDD.t3510 VSS 0.105832f
C19054 VDD.t124 VSS 0.036546f
C19055 VDD.t2880 VSS 0.047206f
C19056 VDD.t3252 VSS 0.102786f
C19057 VDD.t2451 VSS 0.081468f
C19058 VDD.t3638 VSS 0.031978f
C19059 VDD.t2459 VSS 0.039211f
C19060 VDD.t3512 VSS 0.031978f
C19061 VDD.t2457 VSS 0.041495f
C19062 VDD.t2810 VSS 0.031978f
C19063 VDD.t2455 VSS 0.053297f
C19064 VDD.t154 VSS 0.222704f
C19065 VDD.t1405 VSS 0.120679f
C19066 VDD.t1407 VSS 0.068144f
C19067 VDD.t2761 VSS 0.108116f
C19068 VDD.t1732 VSS 0.103928f
C19069 VDD.t1730 VSS 0.068144f
C19070 VDD.t2021 VSS 0.107735f
C19071 VDD.t3743 VSS 0.103548f
C19072 VDD.t1586 VSS 0.104309f
C19073 VDD.t119 VSS 0.101644f
C19074 VDD.t2352 VSS 0.064337f
C19075 VDD.t1590 VSS 0.072712f
C19076 VDD.t1588 VSS 0.090985f
C19077 VDD.t2710 VSS 0.090223f
C19078 VDD.t3371 VSS 0.037308f
C19079 VDD.t160 VSS 0.074996f
C19080 VDD.t3347 VSS 0.107355f
C19081 VDD.t725 VSS 0.037688f
C19082 VDD.t1589 VSS 0.037688f
C19083 VDD.t1591 VSS 0.035785f
C19084 VDD.t1927 VSS 0.031978f
C19085 VDD.t2453 VSS 0.031978f
C19086 VDD.t682 VSS 0.039972f
C19087 VDD.t3446 VSS 0.038069f
C19088 VDD.t3395 VSS 0.03312f
C19089 VDD.t1455 VSS 0.062053f
C19090 VDD.n3866 VSS 0.080433f
C19091 VDD.n3867 VSS 0.022477f
C19092 VDD.n3868 VSS 0.011863f
C19093 VDD.n3870 VSS 0.011881f
C19094 VDD.n3871 VSS 0.011881f
C19095 VDD.n3876 VSS 0.011881f
C19096 VDD.n3885 VSS 0.011917f
C19097 VDD.t126 VSS 0.010055f
C19098 VDD.n3886 VSS 0.01771f
C19099 VDD.n3887 VSS 0.022373f
C19100 VDD.n3893 VSS 0.500541f
C19101 VDD.n3903 VSS 0.011881f
C19102 VDD.t3784 VSS 0.041965f
C19103 VDD.n3904 VSS 0.014361f
C19104 VDD.n3905 VSS 0.023739f
C19105 VDD.n3906 VSS 0.011881f
C19106 VDD.t96 VSS 0.010055f
C19107 VDD.n3907 VSS 0.017371f
C19108 VDD.t3496 VSS 0.014477f
C19109 VDD.n3909 VSS 0.027503f
C19110 VDD.t3498 VSS 0.014204f
C19111 VDD.n3910 VSS 0.013931f
C19112 VDD.n3911 VSS 0.014599f
C19113 VDD.n3912 VSS 0.013812f
C19114 VDD.n3914 VSS 0.028154f
C19115 VDD.n3916 VSS 0.031187f
C19116 VDD.n3917 VSS 0.011881f
C19117 VDD.t1174 VSS 0.01469f
C19118 VDD.n3918 VSS 0.013668f
C19119 VDD.n3919 VSS 0.034187f
C19120 VDD.n3920 VSS 0.011881f
C19121 VDD.n3921 VSS 0.013668f
C19122 VDD.t3331 VSS 0.01469f
C19123 VDD.t844 VSS 0.01469f
C19124 VDD.n3922 VSS 0.013668f
C19125 VDD.n3923 VSS 0.034187f
C19126 VDD.n3924 VSS 0.011881f
C19127 VDD.t574 VSS 0.014703f
C19128 VDD.n3928 VSS 0.011881f
C19129 VDD.n3929 VSS 0.013523f
C19130 VDD.t420 VSS 0.015761f
C19131 VDD.t1134 VSS 0.014469f
C19132 VDD.n3930 VSS 0.017319f
C19133 VDD.t138 VSS 0.010137f
C19134 VDD.t3767 VSS 0.021516f
C19135 VDD.n3932 VSS 0.055166f
C19136 VDD.t139 VSS 0.010137f
C19137 VDD.n3933 VSS 0.030049f
C19138 VDD.t183 VSS 0.010137f
C19139 VDD.t3806 VSS 0.021516f
C19140 VDD.n3935 VSS 0.055166f
C19141 VDD.t184 VSS 0.010137f
C19142 VDD.n3936 VSS 0.030049f
C19143 VDD.n3937 VSS 0.027374f
C19144 VDD.n3938 VSS 0.045507f
C19145 VDD.n3940 VSS 0.015826f
C19146 VDD.n3942 VSS 0.015061f
C19147 VDD.n3944 VSS 0.011881f
C19148 VDD.n3945 VSS 0.011881f
C19149 VDD.n3947 VSS 0.033907f
C19150 VDD.n3949 VSS 0.011881f
C19151 VDD.n3950 VSS 0.011881f
C19152 VDD.n3951 VSS 0.011881f
C19153 VDD.n3953 VSS 0.034187f
C19154 VDD.n3955 VSS 0.011881f
C19155 VDD.n3956 VSS 0.011881f
C19156 VDD.n3957 VSS 0.011881f
C19157 VDD.n3959 VSS 0.013536f
C19158 VDD.n3960 VSS 0.018903f
C19159 VDD.t205 VSS 0.010055f
C19160 VDD.n3962 VSS 0.01771f
C19161 VDD.n3963 VSS 0.03017f
C19162 VDD.n3964 VSS 0.011881f
C19163 VDD.n3965 VSS 0.011881f
C19164 VDD.n3966 VSS 0.027508f
C19165 VDD.n3967 VSS 0.03855f
C19166 VDD.n3968 VSS 0.033189f
C19167 VDD.t3790 VSS 0.075443f
C19168 VDD.n3969 VSS 0.126327f
C19169 VDD.t204 VSS 0.010055f
C19170 VDD.n3970 VSS 0.025888f
C19171 VDD.n3971 VSS 0.022914f
C19172 VDD.t3811 VSS 0.0416f
C19173 VDD.t192 VSS 0.010055f
C19174 VDD.n3972 VSS 0.010971f
C19175 VDD.n3973 VSS 0.024377f
C19176 VDD.n3974 VSS 0.027704f
C19177 VDD.t193 VSS 0.010055f
C19178 VDD.n3975 VSS 0.021153f
C19179 VDD.n3976 VSS 0.051708f
C19180 VDD.n3979 VSS 0.011881f
C19181 VDD.n3980 VSS 0.011881f
C19182 VDD.n3981 VSS 0.011881f
C19183 VDD.n3982 VSS 0.018218f
C19184 VDD.t940 VSS 0.053297f
C19185 VDD.n3984 VSS 0.010543f
C19186 VDD.n3985 VSS 0.014731f
C19187 VDD.n3986 VSS 0.011881f
C19188 VDD.t943 VSS 0.012972f
C19189 VDD.n3988 VSS 0.011881f
C19190 VDD.n3991 VSS 0.011812f
C19191 VDD.n3992 VSS 0.011881f
C19192 VDD.n3993 VSS 0.014361f
C19193 VDD.n3995 VSS 0.011881f
C19194 VDD.n3996 VSS 0.011881f
C19195 VDD.t2784 VSS 0.010846f
C19196 VDD.n3999 VSS 0.011881f
C19197 VDD.t1620 VSS 0.01447f
C19198 VDD.t1618 VSS 0.014477f
C19199 VDD.n4001 VSS 0.011881f
C19200 VDD.n4003 VSS 0.019845f
C19201 VDD.t2396 VSS 0.015761f
C19202 VDD.n4005 VSS 0.022693f
C19203 VDD.t114 VSS 0.010137f
C19204 VDD.t3773 VSS 0.021516f
C19205 VDD.n4007 VSS 0.055166f
C19206 VDD.t115 VSS 0.010137f
C19207 VDD.n4008 VSS 0.030049f
C19208 VDD.t1713 VSS 0.036927f
C19209 VDD.t3033 VSS 0.033881f
C19210 VDD.t942 VSS 0.039592f
C19211 VDD.t1923 VSS 0.046825f
C19212 VDD.t1871 VSS 0.098599f
C19213 VDD.t3739 VSS 0.081468f
C19214 VDD.t2999 VSS 0.031978f
C19215 VDD.t2797 VSS 0.02741f
C19216 VDD.t1513 VSS 0.054058f
C19217 VDD.t1917 VSS 0.084132f
C19218 VDD.t748 VSS 0.08261f
C19219 VDD.t1684 VSS 0.041495f
C19220 VDD.t664 VSS 0.037688f
C19221 VDD.t2799 VSS 0.041495f
C19222 VDD.t2608 VSS 0.04949f
C19223 VDD.t1884 VSS 0.043018f
C19224 VDD.t2325 VSS 0.040734f
C19225 VDD.t3385 VSS 0.077661f
C19226 VDD.t1479 VSS 0.068144f
C19227 VDD.t2509 VSS 0.034262f
C19228 VDD.t2783 VSS 0.036546f
C19229 VDD.t2606 VSS 0.037688f
C19230 VDD.t2800 VSS 0.040734f
C19231 VDD.t1685 VSS 0.064717f
C19232 VDD.t1055 VSS 0.049109f
C19233 VDD.t1619 VSS 0.041114f
C19234 VDD.t3379 VSS 0.031978f
C19235 VDD.t1617 VSS 0.031978f
C19236 VDD.t1686 VSS 0.072712f
C19237 VDD.t1621 VSS 0.081848f
C19238 VDD.t1057 VSS 0.036546f
C19239 VDD.t2397 VSS 0.036166f
C19240 VDD.t2393 VSS 0.065479f
C19241 VDD.t2399 VSS 0.052155f
C19242 VDD.t113 VSS 0.032739f
C19243 VDD.t2395 VSS 0.070047f
C19244 VDD.n4010 VSS 0.123143f
C19245 VDD.n4011 VSS 0.011881f
C19246 VDD.n4012 VSS 0.014498f
C19247 VDD.n4014 VSS 0.011812f
C19248 VDD.n4015 VSS 0.011881f
C19249 VDD.t102 VSS 0.010137f
C19250 VDD.t3815 VSS 0.021516f
C19251 VDD.n4019 VSS 0.055166f
C19252 VDD.t103 VSS 0.010137f
C19253 VDD.n4020 VSS 0.030049f
C19254 VDD.t1190 VSS 0.010815f
C19255 VDD.n4022 VSS 0.019545f
C19256 VDD.n4023 VSS 0.019504f
C19257 VDD.n4024 VSS 0.011881f
C19258 VDD.t1345 VSS 0.01592f
C19259 VDD.n4026 VSS 0.011881f
C19260 VDD.n4027 VSS 0.011881f
C19261 VDD.n4031 VSS 0.011881f
C19262 VDD.t1497 VSS 0.015916f
C19263 VDD.t2442 VSS 0.01447f
C19264 VDD.n4032 VSS 0.017524f
C19265 VDD.n4033 VSS 0.011881f
C19266 VDD.t2444 VSS 0.014477f
C19267 VDD.t2239 VSS 0.014477f
C19268 VDD.n4034 VSS 0.011881f
C19269 VDD.t2237 VSS 0.01447f
C19270 VDD.n4035 VSS 0.01757f
C19271 VDD.n4036 VSS 0.011881f
C19272 VDD.t2515 VSS 0.070047f
C19273 VDD.t2516 VSS 0.014483f
C19274 VDD.n4040 VSS 0.01953f
C19275 VDD.n4041 VSS 0.011881f
C19276 VDD.n4042 VSS 0.013931f
C19277 VDD.t2512 VSS 0.015709f
C19278 VDD.n4044 VSS 0.011881f
C19279 VDD.n4046 VSS 0.031187f
C19280 VDD.n4047 VSS 0.023955f
C19281 VDD.t3823 VSS 0.075443f
C19282 VDD.n4048 VSS 0.126327f
C19283 VDD.t570 VSS 0.010806f
C19284 VDD.n4050 VSS 0.021502f
C19285 VDD.n4051 VSS 0.013652f
C19286 VDD.n4052 VSS 0.011881f
C19287 VDD.n4053 VSS 0.014066f
C19288 VDD.n4054 VSS 0.011881f
C19289 VDD.n4056 VSS 0.011881f
C19290 VDD.n4060 VSS 0.011881f
C19291 VDD.n4061 VSS 0.011881f
C19292 VDD.t462 VSS 0.01592f
C19293 VDD.n4063 VSS 0.019778f
C19294 VDD.t216 VSS 0.010137f
C19295 VDD.t3800 VSS 0.021516f
C19296 VDD.n4065 VSS 0.055166f
C19297 VDD.t217 VSS 0.010137f
C19298 VDD.n4066 VSS 0.030049f
C19299 VDD.n4067 VSS 0.019845f
C19300 VDD.n4068 VSS 0.011038f
C19301 VDD.t1232 VSS 0.031978f
C19302 VDD.t2511 VSS 0.041114f
C19303 VDD.t1799 VSS 0.054819f
C19304 VDD.t1873 VSS 0.059007f
C19305 VDD.t2653 VSS 0.059007f
C19306 VDD.t1827 VSS 0.073092f
C19307 VDD.t2513 VSS 0.073092f
C19308 VDD.t2295 VSS 0.064717f
C19309 VDD.t713 VSS 0.057484f
C19310 VDD.t151 VSS 0.037688f
C19311 VDD.t569 VSS 0.087939f
C19312 VDD.t1841 VSS 0.111923f
C19313 VDD.t275 VSS 0.090223f
C19314 VDD.t710 VSS 0.064717f
C19315 VDD.t3751 VSS 0.037688f
C19316 VDD.t2294 VSS 0.031978f
C19317 VDD.t1789 VSS 0.035023f
C19318 VDD.t1582 VSS 0.041114f
C19319 VDD.t2545 VSS 0.100502f
C19320 VDD.t2517 VSS 0.089843f
C19321 VDD.t711 VSS 0.03312f
C19322 VDD.t3162 VSS 0.035404f
C19323 VDD.t465 VSS 0.036166f
C19324 VDD.t463 VSS 0.065479f
C19325 VDD.t467 VSS 0.035404f
C19326 VDD.t3159 VSS 0.032739f
C19327 VDD.t461 VSS 0.031978f
C19328 VDD.t639 VSS 0.091746f
C19329 VDD.t215 VSS 0.101644f
C19330 VDD.t1201 VSS 0.046825f
C19331 VDD.t1444 VSS 0.058246f
C19332 VDD.n4069 VSS 0.04425f
C19333 VDD.n4070 VSS 0.011881f
C19334 VDD.t1428 VSS 0.010806f
C19335 VDD.n4072 VSS 0.025697f
C19336 VDD.n4073 VSS 0.011881f
C19337 VDD.t3804 VSS 0.05912f
C19338 VDD.t3757 VSS 0.01447f
C19339 VDD.n4074 VSS 0.016701f
C19340 VDD.n4075 VSS 0.011881f
C19341 VDD.t3755 VSS 0.014477f
C19342 VDD.t2805 VSS 0.015916f
C19343 VDD.n4077 VSS 0.024603f
C19344 VDD.n4078 VSS 0.011881f
C19345 VDD.n4080 VSS 0.011881f
C19346 VDD.n4081 VSS 0.010841f
C19347 VDD.n4083 VSS 0.011881f
C19348 VDD.n4084 VSS 0.014361f
C19349 VDD.t790 VSS 0.013903f
C19350 VDD.n4085 VSS 0.016738f
C19351 VDD.n4086 VSS 0.011881f
C19352 VDD.t83 VSS 0.010137f
C19353 VDD.t3780 VSS 0.021516f
C19354 VDD.n4089 VSS 0.055166f
C19355 VDD.t84 VSS 0.010137f
C19356 VDD.n4090 VSS 0.030049f
C19357 VDD.n4092 VSS 0.02676f
C19358 VDD.n4093 VSS 0.011881f
C19359 VDD.t2126 VSS 0.063194f
C19360 VDD.t891 VSS 0.014483f
C19361 VDD.n4095 VSS 0.018959f
C19362 VDD.t2127 VSS 0.015869f
C19363 VDD.t2254 VSS 0.014892f
C19364 VDD.n4096 VSS 0.038735f
C19365 VDD.t3181 VSS 0.0144f
C19366 VDD.n4097 VSS 0.011881f
C19367 VDD.t2252 VSS 0.012721f
C19368 VDD.n4100 VSS 0.018262f
C19369 VDD.n4101 VSS 0.011881f
C19370 VDD.t2174 VSS 0.01592f
C19371 VDD.n4104 VSS 0.011303f
C19372 VDD.n4105 VSS 0.011881f
C19373 VDD.n4108 VSS 0.011881f
C19374 VDD.t458 VSS 0.014745f
C19375 VDD.n4110 VSS 0.020519f
C19376 VDD.n4111 VSS 0.011881f
C19377 VDD.t2377 VSS 0.012972f
C19378 VDD.n4112 VSS 0.013668f
C19379 VDD.n4113 VSS 0.011881f
C19380 VDD.n4114 VSS 0.010543f
C19381 VDD.n4116 VSS 0.011881f
C19382 VDD.t1546 VSS 0.012958f
C19383 VDD.t1412 VSS 0.013749f
C19384 VDD.n4117 VSS 0.010543f
C19385 VDD.n4118 VSS 0.01464f
C19386 VDD.n4119 VSS 0.011881f
C19387 VDD.n4122 VSS 0.011881f
C19388 VDD.n4123 VSS 0.0447f
C19389 VDD.n4124 VSS 0.011881f
C19390 VDD.n4126 VSS 0.027967f
C19391 VDD.n4127 VSS 0.011881f
C19392 VDD.t3775 VSS 0.074403f
C19393 VDD.t135 VSS 0.010055f
C19394 VDD.n4128 VSS 0.01771f
C19395 VDD.n4129 VSS 0.011881f
C19396 VDD.n4132 VSS 0.010815f
C19397 VDD.n4133 VSS 0.011881f
C19398 VDD.t2856 VSS 0.010846f
C19399 VDD.n4136 VSS 0.011881f
C19400 VDD.n4137 VSS 0.011881f
C19401 VDD.n4139 VSS 0.010708f
C19402 VDD.n4140 VSS 0.011881f
C19403 VDD.t1510 VSS 0.015916f
C19404 VDD.n4142 VSS 0.011881f
C19405 VDD.n4143 VSS 0.011881f
C19406 VDD.t1268 VSS 0.014745f
C19407 VDD.n4144 VSS 0.013668f
C19408 VDD.n4145 VSS 0.018529f
C19409 VDD.n4146 VSS 0.011881f
C19410 VDD.n4147 VSS 0.013668f
C19411 VDD.n4148 VSS 0.011881f
C19412 VDD.t2268 VSS 0.014745f
C19413 VDD.n4150 VSS 0.011881f
C19414 VDD.t104 VSS 0.222704f
C19415 VDD.t946 VSS 0.120679f
C19416 VDD.t944 VSS 0.068144f
C19417 VDD.t1977 VSS 0.107735f
C19418 VDD.t3572 VSS 0.07195f
C19419 VDD.t1680 VSS 0.032359f
C19420 VDD.t1682 VSS 0.03312f
C19421 VDD.t674 VSS 0.036166f
C19422 VDD.t2836 VSS 0.053297f
C19423 VDD.t2253 VSS 0.032739f
C19424 VDD.t2128 VSS 0.031978f
C19425 VDD.t2251 VSS 0.032739f
C19426 VDD.t2124 VSS 0.059768f
C19427 VDD.t2130 VSS 0.044541f
C19428 VDD.t2943 VSS 0.036546f
C19429 VDD.t1851 VSS 0.034643f
C19430 VDD.t2934 VSS 0.041876f
C19431 VDD.t3188 VSS 0.063956f
C19432 VDD.t3178 VSS 0.033501f
C19433 VDD.t2173 VSS 0.034262f
C19434 VDD.t2169 VSS 0.065479f
C19435 VDD.t2171 VSS 0.040353f
C19436 VDD.t3184 VSS 0.032739f
C19437 VDD.t2175 VSS 0.031978f
C19438 VDD.t3192 VSS 0.036546f
C19439 VDD.t1596 VSS 0.031978f
C19440 VDD.t2937 VSS 0.034262f
C19441 VDD.t2948 VSS 0.10507f
C19442 VDD.t457 VSS 0.10507f
C19443 VDD.t455 VSS 0.034262f
C19444 VDD.t2376 VSS 0.034262f
C19445 VDD.t3667 VSS 0.033881f
C19446 VDD.t1395 VSS 0.036927f
C19447 VDD.t3103 VSS 0.142378f
C19448 VDD.t1411 VSS 0.141236f
C19449 VDD.t1545 VSS 0.065859f
C19450 VDD.t1594 VSS 0.037688f
C19451 VDD.t871 VSS 0.036927f
C19452 VDD.t1537 VSS 0.032359f
C19453 VDD.t2663 VSS 0.033881f
C19454 VDD.t2066 VSS 0.070428f
C19455 VDD.t2795 VSS 0.071189f
C19456 VDD.t2873 VSS 0.086797f
C19457 VDD.n4151 VSS 0.119717f
C19458 VDD.t3151 VSS 0.085275f
C19459 VDD.t1196 VSS 0.104309f
C19460 VDD.t134 VSS 0.101644f
C19461 VDD.t2288 VSS 0.064337f
C19462 VDD.t1350 VSS 0.072712f
C19463 VDD.t1198 VSS 0.090985f
C19464 VDD.t2563 VSS 0.073854f
C19465 VDD.t2661 VSS 0.036927f
C19466 VDD.t1833 VSS 0.036166f
C19467 VDD.t2659 VSS 0.074996f
C19468 VDD.t2855 VSS 0.07157f
C19469 VDD.t1391 VSS 0.037688f
C19470 VDD.t1195 VSS 0.036166f
C19471 VDD.t1993 VSS 0.032739f
C19472 VDD.t1351 VSS 0.04987f
C19473 VDD.t1511 VSS 0.067382f
C19474 VDD.t2401 VSS 0.041114f
C19475 VDD.t1849 VSS 0.036166f
C19476 VDD.t1861 VSS 0.031978f
C19477 VDD.t1352 VSS 0.083371f
C19478 VDD.t1509 VSS 0.083371f
C19479 VDD.t1052 VSS 0.035023f
C19480 VDD.t2871 VSS 0.070428f
C19481 VDD.t1267 VSS 0.068905f
C19482 VDD.t1265 VSS 0.068144f
C19483 VDD.t1989 VSS 0.072712f
C19484 VDD.t1283 VSS 0.07157f
C19485 VDD.t1527 VSS 0.036166f
C19486 VDD.t2269 VSS 0.03312f
C19487 VDD.t2267 VSS 0.032359f
C19488 VDD.t2869 VSS 0.053677f
C19489 VDD.n4152 VSS 0.078132f
C19490 VDD.n4153 VSS 0.011881f
C19491 VDD.n4154 VSS 0.011881f
C19492 VDD.n4155 VSS 0.013668f
C19493 VDD.n4157 VSS 0.011881f
C19494 VDD.n4158 VSS 0.011881f
C19495 VDD.t1681 VSS 0.014745f
C19496 VDD.n4159 VSS 0.013668f
C19497 VDD.n4160 VSS 0.013668f
C19498 VDD.n4161 VSS 0.03134f
C19499 VDD.t105 VSS 0.010137f
C19500 VDD.t3794 VSS 0.021516f
C19501 VDD.n4163 VSS 0.055166f
C19502 VDD.t106 VSS 0.010137f
C19503 VDD.n4164 VSS 0.030049f
C19504 VDD.t194 VSS 0.010137f
C19505 VDD.t3792 VSS 0.021516f
C19506 VDD.n4166 VSS 0.055166f
C19507 VDD.t195 VSS 0.010137f
C19508 VDD.n4167 VSS 0.030049f
C19509 VDD.n4168 VSS 0.02678f
C19510 VDD.t2561 VSS 0.014745f
C19511 VDD.t947 VSS 0.014745f
C19512 VDD.n4170 VSS 0.035938f
C19513 VDD.n4172 VSS 0.053216f
C19514 VDD.n4173 VSS 0.011881f
C19515 VDD.n4174 VSS 0.011881f
C19516 VDD.n4176 VSS 0.020244f
C19517 VDD.n4177 VSS 0.017065f
C19518 VDD.n4178 VSS 0.017111f
C19519 VDD.n4179 VSS 0.02392f
C19520 VDD.n4180 VSS 0.019581f
C19521 VDD.n4181 VSS 0.017065f
C19522 VDD.n4182 VSS 0.017774f
C19523 VDD.n4184 VSS 0.011881f
C19524 VDD.n4185 VSS 0.011881f
C19525 VDD.n4186 VSS 0.011881f
C19526 VDD.n4188 VSS 0.020244f
C19527 VDD.n4189 VSS 0.017088f
C19528 VDD.n4190 VSS 0.023848f
C19529 VDD.n4192 VSS 0.011881f
C19530 VDD.n4193 VSS 0.011881f
C19531 VDD.n4197 VSS 0.012061f
C19532 VDD.n4200 VSS 0.011881f
C19533 VDD.n4201 VSS 0.011881f
C19534 VDD.n4203 VSS 0.01576f
C19535 VDD.n4205 VSS 0.011881f
C19536 VDD.n4206 VSS 0.011881f
C19537 VDD.n4210 VSS 0.011917f
C19538 VDD.n4211 VSS 0.011881f
C19539 VDD.n4212 VSS 0.011881f
C19540 VDD.n4213 VSS 0.022712f
C19541 VDD.n4214 VSS 0.100348f
C19542 VDD.n4215 VSS 0.023051f
C19543 VDD.n4216 VSS 0.022101f
C19544 VDD.n4217 VSS 0.018814f
C19545 VDD.n4218 VSS 0.011881f
C19546 VDD.n4219 VSS 0.011881f
C19547 VDD.n4220 VSS 0.011881f
C19548 VDD.n4221 VSS 0.031187f
C19549 VDD.n4222 VSS 0.015933f
C19550 VDD.n4223 VSS 0.023316f
C19551 VDD.t136 VSS 0.010055f
C19552 VDD.n4224 VSS 0.017371f
C19553 VDD.n4225 VSS 0.011038f
C19554 VDD.n4226 VSS 0.011881f
C19555 VDD.n4227 VSS 0.011881f
C19556 VDD.n4228 VSS 0.011881f
C19557 VDD.n4230 VSS 0.018529f
C19558 VDD.n4232 VSS 0.01723f
C19559 VDD.n4233 VSS 0.011881f
C19560 VDD.n4234 VSS 0.011881f
C19561 VDD.n4235 VSS 0.011881f
C19562 VDD.n4237 VSS 0.025979f
C19563 VDD.n4239 VSS 0.011881f
C19564 VDD.n4240 VSS 0.011881f
C19565 VDD.n4241 VSS 0.011881f
C19566 VDD.n4243 VSS 0.014846f
C19567 VDD.n4244 VSS 0.017385f
C19568 VDD.n4245 VSS 0.010335f
C19569 VDD.n4246 VSS 0.011881f
C19570 VDD.n4247 VSS 0.011881f
C19571 VDD.n4248 VSS 0.011881f
C19572 VDD.n4250 VSS 0.011327f
C19573 VDD.n4251 VSS 0.016753f
C19574 VDD.n4252 VSS 0.010435f
C19575 VDD.n4253 VSS 0.011881f
C19576 VDD.n4254 VSS 0.011881f
C19577 VDD.n4255 VSS 0.011881f
C19578 VDD.n4257 VSS 0.025626f
C19579 VDD.n4259 VSS 0.011881f
C19580 VDD.n4260 VSS 0.011881f
C19581 VDD.n4261 VSS 0.011881f
C19582 VDD.n4263 VSS 0.010076f
C19583 VDD.n4267 VSS 0.011881f
C19584 VDD.n4268 VSS 0.011881f
C19585 VDD.n4269 VSS 0.011881f
C19586 VDD.n4270 VSS 0.010708f
C19587 VDD.n4271 VSS 0.011881f
C19588 VDD.n4275 VSS 0.011881f
C19589 VDD.n4277 VSS 0.011881f
C19590 VDD.n4279 VSS 0.014361f
C19591 VDD.n4280 VSS 0.010146f
C19592 VDD.t3787 VSS 0.041965f
C19593 VDD.n4282 VSS 0.03017f
C19594 VDD.n4283 VSS 0.011881f
C19595 VDD.t182 VSS 0.010055f
C19596 VDD.n4284 VSS 0.01771f
C19597 VDD.n4286 VSS 0.012758f
C19598 VDD.n4287 VSS 0.011881f
C19599 VDD.t809 VSS 0.014745f
C19600 VDD.n4288 VSS 0.020199f
C19601 VDD.n4289 VSS 0.011881f
C19602 VDD.n4290 VSS 0.013523f
C19603 VDD.t2576 VSS 0.013611f
C19604 VDD.n4292 VSS 0.013894f
C19605 VDD.n4293 VSS 0.015038f
C19606 VDD.n4295 VSS 0.011881f
C19607 VDD.n4296 VSS 0.011881f
C19608 VDD.n4297 VSS 0.011881f
C19609 VDD.n4299 VSS 0.017093f
C19610 VDD.t1188 VSS 0.012738f
C19611 VDD.n4301 VSS 0.013851f
C19612 VDD.n4302 VSS 0.011881f
C19613 VDD.n4303 VSS 0.011881f
C19614 VDD.n4304 VSS 0.011881f
C19615 VDD.n4306 VSS 0.018139f
C19616 VDD.n4308 VSS 0.014399f
C19617 VDD.n4310 VSS 0.011881f
C19618 VDD.n4311 VSS 0.011881f
C19619 VDD.n4312 VSS 0.011881f
C19620 VDD.n4313 VSS 0.02339f
C19621 VDD.n4314 VSS 0.037956f
C19622 VDD.t181 VSS 0.010055f
C19623 VDD.n4316 VSS 0.011917f
C19624 VDD.n4318 VSS 0.011881f
C19625 VDD.n4319 VSS 0.011881f
C19626 VDD.n4320 VSS 0.011881f
C19627 VDD.t1723 VSS 0.010846f
C19628 VDD.n4322 VSS 0.015964f
C19629 VDD.n4324 VSS 0.011881f
C19630 VDD.n4325 VSS 0.011881f
C19631 VDD.n4326 VSS 0.011881f
C19632 VDD.n4332 VSS 0.011881f
C19633 VDD.n4333 VSS 0.011881f
C19634 VDD.t889 VSS 0.015916f
C19635 VDD.n4335 VSS 0.024123f
C19636 VDD.t3203 VSS 0.014477f
C19637 VDD.n4336 VSS 0.017372f
C19638 VDD.n4337 VSS 0.011881f
C19639 VDD.n4338 VSS 0.011881f
C19640 VDD.n4339 VSS 0.011881f
C19641 VDD.n4340 VSS 0.036529f
C19642 VDD.n4341 VSS 0.082319f
C19643 VDD.t3180 VSS 0.051012f
C19644 VDD.t3202 VSS 0.037308f
C19645 VDD.t890 VSS 0.037308f
C19646 VDD.t888 VSS 0.113826f
C19647 VDD.t886 VSS 0.113826f
C19648 VDD.t3414 VSS 0.040734f
C19649 VDD.t658 VSS 0.041114f
C19650 VDD.t892 VSS 0.036546f
C19651 VDD.t2265 VSS 0.031597f
C19652 VDD.t1486 VSS 0.02779f
C19653 VDD.t2245 VSS 0.03312f
C19654 VDD.t1719 VSS 0.070428f
C19655 VDD.t1722 VSS 0.048348f
C19656 VDD.t3642 VSS 0.04987f
C19657 VDD.t656 VSS 0.064337f
C19658 VDD.t3359 VSS 0.041495f
C19659 VDD.t1584 VSS 0.036927f
C19660 VDD.t2275 VSS 0.073854f
C19661 VDD.t1720 VSS 0.085275f
C19662 VDD.t180 VSS 0.037688f
C19663 VDD.t2244 VSS 0.040734f
C19664 VDD.t1179 VSS 0.100502f
C19665 VDD.t1995 VSS 0.101644f
C19666 VDD.t1185 VSS 0.068144f
C19667 VDD.t1187 VSS 0.10469f
C19668 VDD.t2763 VSS 0.105451f
C19669 VDD.t2669 VSS 0.065098f
C19670 VDD.t1822 VSS 0.036546f
C19671 VDD.t808 VSS 0.036166f
C19672 VDD.t810 VSS 0.067382f
C19673 VDD.t2575 VSS 0.036166f
C19674 VDD.t2972 VSS 0.054058f
C19675 VDD.t642 VSS 0.067763f
C19676 VDD.t1429 VSS 0.090223f
C19677 VDD.t1835 VSS 0.054819f
C19678 VDD.t85 VSS 0.074996f
C19679 VDD.t1427 VSS 0.094792f
C19680 VDD.t641 VSS 0.070428f
C19681 VDD.t1443 VSS 0.064717f
C19682 VDD.t2802 VSS 0.049109f
C19683 VDD.t3756 VSS 0.041114f
C19684 VDD.t1829 VSS 0.031978f
C19685 VDD.t3754 VSS 0.031978f
C19686 VDD.t3484 VSS 0.072331f
C19687 VDD.t2953 VSS 0.081848f
C19688 VDD.t2804 VSS 0.07157f
C19689 VDD.t788 VSS 0.078422f
C19690 VDD.t2111 VSS 0.047206f
C19691 VDD.t2841 VSS 0.031978f
C19692 VDD.t2886 VSS 0.031978f
C19693 VDD.t3088 VSS 0.031978f
C19694 VDD.t3198 VSS 0.041114f
C19695 VDD.t2527 VSS 0.040353f
C19696 VDD.t795 VSS 0.056342f
C19697 VDD.t793 VSS 0.063956f
C19698 VDD.t791 VSS 0.063956f
C19699 VDD.t789 VSS 0.041495f
C19700 VDD.t2620 VSS 0.048728f
C19701 VDD.t1881 VSS 0.063575f
C19702 VDD.t1768 VSS 0.057865f
C19703 VDD.t409 VSS 0.057103f
C19704 VDD.t2529 VSS 0.051012f
C19705 VDD.t775 VSS 0.063956f
C19706 VDD.t2618 VSS 0.037308f
C19707 VDD.t82 VSS 0.070808f
C19708 VDD.n4342 VSS 0.136467f
C19709 VDD.n4343 VSS 0.044113f
C19710 VDD.n4344 VSS 0.01978f
C19711 VDD.n4345 VSS 0.019845f
C19712 VDD.n4346 VSS 0.019778f
C19713 VDD.n4348 VSS 0.018529f
C19714 VDD.n4350 VSS 0.011881f
C19715 VDD.n4351 VSS 0.011881f
C19716 VDD.n4352 VSS 0.011881f
C19717 VDD.n4354 VSS 0.010558f
C19718 VDD.n4355 VSS 0.015834f
C19719 VDD.n4357 VSS 0.012786f
C19720 VDD.n4358 VSS 0.013931f
C19721 VDD.n4359 VSS 0.01469f
C19722 VDD.n4361 VSS 0.011881f
C19723 VDD.n4362 VSS 0.011881f
C19724 VDD.n4363 VSS 0.011881f
C19725 VDD.n4365 VSS 0.013652f
C19726 VDD.n4368 VSS 0.011881f
C19727 VDD.n4369 VSS 0.011881f
C19728 VDD.n4370 VSS 0.011881f
C19729 VDD.n4374 VSS 0.017807f
C19730 VDD.n4375 VSS 0.010242f
C19731 VDD.n4376 VSS 0.011881f
C19732 VDD.n4377 VSS 0.011881f
C19733 VDD.n4378 VSS 0.011881f
C19734 VDD.n4380 VSS 0.011917f
C19735 VDD.t86 VSS 0.010055f
C19736 VDD.n4381 VSS 0.01771f
C19737 VDD.n4382 VSS 0.069744f
C19738 VDD.n4383 VSS 0.011881f
C19739 VDD.n4384 VSS 0.011881f
C19740 VDD.n4385 VSS 0.026102f
C19741 VDD.n4386 VSS 0.022882f
C19742 VDD.n4387 VSS 0.023127f
C19743 VDD.t87 VSS 0.010055f
C19744 VDD.n4388 VSS 0.01771f
C19745 VDD.n4389 VSS 0.022882f
C19746 VDD.n4390 VSS 0.011881f
C19747 VDD.n4391 VSS 0.011881f
C19748 VDD.n4392 VSS 0.01978f
C19749 VDD.n4393 VSS 0.024416f
C19750 VDD.n4394 VSS 0.026206f
C19751 VDD.n4395 VSS 0.017703f
C19752 VDD.n4396 VSS 0.012964f
C19753 VDD.n4397 VSS 0.010731f
C19754 VDD.n4399 VSS 0.014847f
C19755 VDD.n4402 VSS 0.011881f
C19756 VDD.n4403 VSS 0.011881f
C19757 VDD.n4404 VSS 0.011881f
C19758 VDD.n4407 VSS 0.015927f
C19759 VDD.n4410 VSS 0.011881f
C19760 VDD.n4411 VSS 0.023665f
C19761 VDD.n4413 VSS 0.022583f
C19762 VDD.t152 VSS 0.010055f
C19763 VDD.n4414 VSS 0.025888f
C19764 VDD.n4415 VSS 0.033189f
C19765 VDD.n4416 VSS 0.025594f
C19766 VDD.n4417 VSS 0.023665f
C19767 VDD.n4418 VSS 0.011881f
C19768 VDD.n4419 VSS 0.011881f
C19769 VDD.n4420 VSS 0.028983f
C19770 VDD.n4421 VSS 0.020659f
C19771 VDD.t153 VSS 0.010055f
C19772 VDD.n4423 VSS 0.011917f
C19773 VDD.n4424 VSS 0.011634f
C19774 VDD.n4426 VSS 0.011881f
C19775 VDD.n4427 VSS 0.011881f
C19776 VDD.n4430 VSS 0.020349f
C19777 VDD.n4431 VSS 0.014576f
C19778 VDD.n4433 VSS 0.011881f
C19779 VDD.n4434 VSS 0.011881f
C19780 VDD.n4435 VSS 0.011881f
C19781 VDD.t3236 VSS 0.014207f
C19782 VDD.n4438 VSS 0.011881f
C19783 VDD.n4440 VSS 0.01708f
C19784 VDD.n4441 VSS 0.021988f
C19785 VDD.n4442 VSS 0.011881f
C19786 VDD.t3798 VSS 0.075443f
C19787 VDD.n4443 VSS 0.126327f
C19788 VDD.t117 VSS 0.010055f
C19789 VDD.n4444 VSS 0.025888f
C19790 VDD.n4445 VSS 0.033189f
C19791 VDD.t412 VSS 0.010806f
C19792 VDD.n4446 VSS 0.02468f
C19793 VDD.n4447 VSS 0.011881f
C19794 VDD.t118 VSS 0.010055f
C19795 VDD.n4448 VSS 0.012625f
C19796 VDD.n4449 VSS 0.014066f
C19797 VDD.n4450 VSS 0.016065f
C19798 VDD.n4451 VSS 0.011881f
C19799 VDD.n4452 VSS 0.011401f
C19800 VDD.n4453 VSS 0.011881f
C19801 VDD.n4456 VSS 0.011881f
C19802 VDD.n4458 VSS 0.018262f
C19803 VDD.n4459 VSS 0.011881f
C19804 VDD.n4460 VSS 0.011881f
C19805 VDD.n4461 VSS 0.011881f
C19806 VDD.n4463 VSS 0.020571f
C19807 VDD.t733 VSS 0.01592f
C19808 VDD.n4465 VSS 0.018069f
C19809 VDD.n4466 VSS 0.011881f
C19810 VDD.n4467 VSS 0.011881f
C19811 VDD.n4468 VSS 0.011881f
C19812 VDD.n4470 VSS 0.013652f
C19813 VDD.n4473 VSS 0.011881f
C19814 VDD.n4474 VSS 0.011881f
C19815 VDD.n4477 VSS 0.011101f
C19816 VDD.n4479 VSS 0.011917f
C19817 VDD.n4480 VSS 0.011881f
C19818 VDD.n4481 VSS 0.011881f
C19819 VDD.n4482 VSS 0.020678f
C19820 VDD.n4483 VSS 0.031187f
C19821 VDD.n4484 VSS 0.025594f
C19822 VDD.n4485 VSS 0.023665f
C19823 VDD.n4486 VSS 0.023955f
C19824 VDD.n4487 VSS 0.023665f
C19825 VDD.t909 VSS 0.015916f
C19826 VDD.n4488 VSS 0.023368f
C19827 VDD.n4490 VSS 0.016753f
C19828 VDD.t907 VSS 0.014483f
C19829 VDD.n4491 VSS 0.019302f
C19830 VDD.n4492 VSS 0.011881f
C19831 VDD.n4493 VSS 0.011881f
C19832 VDD.n4495 VSS 0.015995f
C19833 VDD.t1214 VSS 0.01592f
C19834 VDD.t3238 VSS 0.014403f
C19835 VDD.n4497 VSS 0.031542f
C19836 VDD.n4498 VSS 0.011881f
C19837 VDD.n4499 VSS 0.011881f
C19838 VDD.n4500 VSS 0.011881f
C19839 VDD.n4501 VSS 0.044341f
C19840 VDD.n4502 VSS 0.158547f
C19841 VDD.t3237 VSS 0.091746f
C19842 VDD.t1213 VSS 0.031978f
C19843 VDD.t3235 VSS 0.032739f
C19844 VDD.t1215 VSS 0.036166f
C19845 VDD.t1217 VSS 0.065479f
C19846 VDD.t1211 VSS 0.039211f
C19847 VDD.t906 VSS 0.036546f
C19848 VDD.t2191 VSS 0.031978f
C19849 VDD.t908 VSS 0.083752f
C19850 VDD.t2157 VSS 0.113826f
C19851 VDD.t2970 VSS 0.073092f
C19852 VDD.t904 VSS 0.06053f
C19853 VDD.t116 VSS 0.031978f
C19854 VDD.t1716 VSS 0.045302f
C19855 VDD.t1093 VSS 0.070428f
C19856 VDD.t411 VSS 0.112684f
C19857 VDD.t2980 VSS 0.109639f
C19858 VDD.t2541 VSS 0.036927f
C19859 VDD.t413 VSS 0.041114f
C19860 VDD.t1783 VSS 0.053297f
C19861 VDD.t1094 VSS 0.031978f
C19862 VDD.t3239 VSS 0.037688f
C19863 VDD.t1715 VSS 0.0552f
C19864 VDD.t2632 VSS 0.103548f
C19865 VDD.t732 VSS 0.101264f
C19866 VDD.t734 VSS 0.03312f
C19867 VDD.t1091 VSS 0.032359f
C19868 VDD.t3126 VSS 0.032359f
C19869 VDD.t736 VSS 0.03312f
C19870 VDD.t738 VSS 0.069286f
C19871 VDD.t2240 VSS 0.090223f
C19872 VDD.t1592 VSS 0.085275f
C19873 VDD.t2467 VSS 0.041495f
C19874 VDD.t2019 VSS 0.048728f
C19875 VDD.t3753 VSS 0.092127f
C19876 VDD.t1672 VSS 0.081468f
C19877 VDD.t3257 VSS 0.035023f
C19878 VDD.t1220 VSS 0.02741f
C19879 VDD.t2153 VSS 0.037688f
C19880 VDD.t2470 VSS 0.036546f
C19881 VDD.t2009 VSS 0.053297f
C19882 VDD.t1191 VSS 0.070428f
C19883 VDD.t3367 VSS 0.072331f
C19884 VDD.t101 VSS 0.074996f
C19885 VDD.t1189 VSS 0.07728f
C19886 VDD.t2469 VSS 0.052155f
C19887 VDD.t1344 VSS 0.032739f
C19888 VDD.t1219 VSS 0.032739f
C19889 VDD.t1342 VSS 0.031978f
C19890 VDD.t1494 VSS 0.032739f
C19891 VDD.t1340 VSS 0.041114f
C19892 VDD.t3383 VSS 0.032739f
C19893 VDD.t1338 VSS 0.031978f
C19894 VDD.t1221 VSS 0.036546f
C19895 VDD.t2976 VSS 0.081848f
C19896 VDD.t1496 VSS 0.141997f
C19897 VDD.t2847 VSS 0.072331f
C19898 VDD.t2441 VSS 0.032739f
C19899 VDD.t2443 VSS 0.040734f
C19900 VDD.t1931 VSS 0.047967f
C19901 VDD.t2840 VSS 0.064337f
C19902 VDD.t2238 VSS 0.057103f
C19903 VDD.t2236 VSS 0.056342f
C19904 VDD.t323 VSS 0.051774f
C19905 VDD.t567 VSS 0.063956f
C19906 VDD.t1907 VSS 0.037308f
C19907 VDD.n4503 VSS 0.061001f
C19908 VDD.n4504 VSS 0.024103f
C19909 VDD.n4507 VSS 0.011881f
C19910 VDD.n4508 VSS 0.011881f
C19911 VDD.n4509 VSS 0.011881f
C19912 VDD.n4511 VSS 0.018401f
C19913 VDD.n4512 VSS 0.018401f
C19914 VDD.n4513 VSS 0.014361f
C19915 VDD.n4514 VSS 0.010695f
C19916 VDD.n4516 VSS 0.011881f
C19917 VDD.n4517 VSS 0.011881f
C19918 VDD.n4518 VSS 0.011881f
C19919 VDD.n4520 VSS 0.024603f
C19920 VDD.n4522 VSS 0.011881f
C19921 VDD.n4523 VSS 0.011881f
C19922 VDD.n4525 VSS 0.014618f
C19923 VDD.n4526 VSS 0.010631f
C19924 VDD.n4527 VSS 0.010663f
C19925 VDD.n4529 VSS 0.018412f
C19926 VDD.n4530 VSS 0.01978f
C19927 VDD.n4531 VSS 0.019845f
C19928 VDD.n4532 VSS 0.019778f
C19929 VDD.n4533 VSS 0.011881f
C19930 VDD.n4538 VSS 0.011881f
C19931 VDD.n4539 VSS 0.011881f
C19932 VDD.n4540 VSS 0.011881f
C19933 VDD.n4543 VSS 0.02343f
C19934 VDD.n4544 VSS 0.011881f
C19935 VDD.n4545 VSS 0.011881f
C19936 VDD.n4546 VSS 0.01978f
C19937 VDD.n4547 VSS 0.044113f
C19938 VDD.n4548 VSS 0.017356f
C19939 VDD.t1058 VSS 0.015709f
C19940 VDD.n4550 VSS 0.019343f
C19941 VDD.n4551 VSS 0.014801f
C19942 VDD.n4553 VSS 0.019778f
C19943 VDD.n4554 VSS 0.011881f
C19944 VDD.n4555 VSS 0.011881f
C19945 VDD.n4557 VSS 0.010227f
C19946 VDD.n4558 VSS 0.017052f
C19947 VDD.n4559 VSS 0.010242f
C19948 VDD.n4560 VSS 0.016701f
C19949 VDD.n4561 VSS 0.011881f
C19950 VDD.n4562 VSS 0.011881f
C19951 VDD.n4563 VSS 0.011881f
C19952 VDD.n4566 VSS 0.014912f
C19953 VDD.n4569 VSS 0.011101f
C19954 VDD.n4571 VSS 0.011881f
C19955 VDD.n4572 VSS 0.011881f
C19956 VDD.n4573 VSS 0.011881f
C19957 VDD.n4576 VSS 0.011267f
C19958 VDD.n4578 VSS 0.011881f
C19959 VDD.n4579 VSS 0.011881f
C19960 VDD.n4580 VSS 0.011881f
C19961 VDD.n4584 VSS 0.014404f
C19962 VDD.n4585 VSS 0.011881f
C19963 VDD.n4586 VSS 0.011881f
C19964 VDD.n4587 VSS 0.011881f
C19965 VDD.n4589 VSS 0.011798f
C19966 VDD.n4590 VSS 0.014361f
C19967 VDD.n4591 VSS 0.010626f
C19968 VDD.n4593 VSS 0.011881f
C19969 VDD.n4594 VSS 0.011881f
C19970 VDD.n4595 VSS 0.011881f
C19971 VDD.t1474 VSS 0.015994f
C19972 VDD.t2113 VSS 0.015761f
C19973 VDD.n4596 VSS 0.014865f
C19974 VDD.n4601 VSS 0.014892f
C19975 VDD.n4602 VSS 0.011881f
C19976 VDD.t1472 VSS 0.013927f
C19977 VDD.n4604 VSS 0.010242f
C19978 VDD.t2355 VSS 0.014477f
C19979 VDD.n4605 VSS 0.019845f
C19980 VDD.t2314 VSS 0.01592f
C19981 VDD.n4607 VSS 0.011881f
C19982 VDD.n4614 VSS 0.011812f
C19983 VDD.n4616 VSS 0.011881f
C19984 VDD.n4617 VSS 0.011881f
C19985 VDD.n4618 VSS 0.018262f
C19986 VDD.n4622 VSS 0.011881f
C19987 VDD.n4623 VSS 0.011881f
C19988 VDD.n4624 VSS 0.019778f
C19989 VDD.n4625 VSS 0.017543f
C19990 VDD.t99 VSS 0.010137f
C19991 VDD.t3770 VSS 0.021516f
C19992 VDD.n4627 VSS 0.055166f
C19993 VDD.t100 VSS 0.010137f
C19994 VDD.n4628 VSS 0.030049f
C19995 VDD.t2256 VSS 0.010831f
C19996 VDD.n4629 VSS 0.030933f
C19997 VDD.t2357 VSS 0.01447f
C19998 VDD.n4630 VSS 0.016038f
C19999 VDD.n4631 VSS 0.01978f
C20000 VDD.n4632 VSS 0.011881f
C20001 VDD.n4633 VSS 0.011881f
C20002 VDD.n4634 VSS 0.017052f
C20003 VDD.n4635 VSS 0.010227f
C20004 VDD.n4637 VSS 0.011863f
C20005 VDD.n4639 VSS 0.011881f
C20006 VDD.n4640 VSS 0.011881f
C20007 VDD.n4646 VSS 0.011881f
C20008 VDD.n4647 VSS 0.011881f
C20009 VDD.n4648 VSS 0.011881f
C20010 VDD.n4649 VSS 0.024652f
C20011 VDD.n4650 VSS 0.081558f
C20012 VDD.t2112 VSS 0.070047f
C20013 VDD.t1473 VSS 0.032739f
C20014 VDD.t2116 VSS 0.031978f
C20015 VDD.t1469 VSS 0.032739f
C20016 VDD.t2118 VSS 0.031978f
C20017 VDD.t1477 VSS 0.032739f
C20018 VDD.t2114 VSS 0.031978f
C20019 VDD.t1471 VSS 0.036546f
C20020 VDD.t2358 VSS 0.074235f
C20021 VDD.t1467 VSS 0.072712f
C20022 VDD.t2354 VSS 0.031978f
C20023 VDD.t3387 VSS 0.031978f
C20024 VDD.t2356 VSS 0.041114f
C20025 VDD.t1475 VSS 0.049109f
C20026 VDD.t2728 VSS 0.064717f
C20027 VDD.t2207 VSS 0.039972f
C20028 VDD.t98 VSS 0.037688f
C20029 VDD.t2255 VSS 0.091746f
C20030 VDD.t2313 VSS 0.074996f
C20031 VDD.t3401 VSS 0.032739f
C20032 VDD.t2315 VSS 0.036927f
C20033 VDD.t2257 VSS 0.032739f
C20034 VDD.t2311 VSS 0.047586f
C20035 VDD.t2309 VSS 0.03845f
C20036 VDD.t2210 VSS 0.036546f
C20037 VDD.t3499 VSS 0.037688f
C20038 VDD.t2727 VSS 0.041876f
C20039 VDD.t762 VSS 0.08261f
C20040 VDD.t1921 VSS 0.084132f
C20041 VDD.t2536 VSS 0.054058f
C20042 VDD.t2208 VSS 0.02741f
C20043 VDD.t1252 VSS 0.031978f
C20044 VDD.t3737 VSS 0.081468f
C20045 VDD.t3242 VSS 0.098599f
C20046 VDD.t1909 VSS 0.046444f
C20047 VDD.t94 VSS 0.041495f
C20048 VDD.t1547 VSS 0.087559f
C20049 VDD.t137 VSS 0.222704f
C20050 VDD.t1133 VSS 0.091746f
C20051 VDD.t419 VSS 0.031978f
C20052 VDD.t1131 VSS 0.032739f
C20053 VDD.t417 VSS 0.036166f
C20054 VDD.t2039 VSS 0.032739f
C20055 VDD.t415 VSS 0.03312f
C20056 VDD.t421 VSS 0.069286f
C20057 VDD.t2640 VSS 0.03883f
C20058 VDD.t573 VSS 0.034262f
C20059 VDD.t575 VSS 0.068144f
C20060 VDD.t2878 VSS 0.038069f
C20061 VDD.t843 VSS 0.033881f
C20062 VDD.t845 VSS 0.068144f
C20063 VDD.t3650 VSS 0.038069f
C20064 VDD.t3330 VSS 0.033881f
C20065 VDD.t3328 VSS 0.068144f
C20066 VDD.t1987 VSS 0.038069f
C20067 VDD.t1173 VSS 0.033881f
C20068 VDD.t1171 VSS 0.068144f
C20069 VDD.t2109 VSS 0.107735f
C20070 VDD.t1933 VSS 0.10507f
C20071 VDD.t2465 VSS 0.034262f
C20072 VDD.t203 VSS 0.105832f
C20073 VDD.t191 VSS 0.189584f
C20074 VDD.t1886 VSS 0.116491f
C20075 VDD.t1785 VSS 0.057103f
C20076 VDD.t3497 VSS 0.041114f
C20077 VDD.t637 VSS 0.031978f
C20078 VDD.t3495 VSS 0.070047f
C20079 VDD.n4651 VSS 0.120479f
C20080 VDD.n4652 VSS 0.04422f
C20081 VDD.n4653 VSS 0.011038f
C20082 VDD.n4654 VSS 0.011881f
C20083 VDD.n4655 VSS 0.011881f
C20084 VDD.n4656 VSS 0.015933f
C20085 VDD.n4657 VSS 0.02339f
C20086 VDD.n4658 VSS 0.037956f
C20087 VDD.t95 VSS 0.010055f
C20088 VDD.n4660 VSS 0.011917f
C20089 VDD.n4661 VSS 0.011881f
C20090 VDD.n4671 VSS 0.014404f
C20091 VDD.n4678 VSS 0.292366f
C20092 VDD.n4679 VSS 0.115767f
C20093 a_8912_37509.t13 VSS 0.177274f
C20094 a_8912_37509.n0 VSS 0.308192f
C20095 a_8912_37509.t32 VSS 0.890777f
C20096 a_8912_37509.n1 VSS 0.475921f
C20097 a_8912_37509.t34 VSS 0.890777f
C20098 a_8912_37509.t33 VSS 0.890777f
C20099 a_8912_37509.n2 VSS 1.34409f
C20100 a_8912_37509.t37 VSS 0.890777f
C20101 a_8912_37509.n3 VSS 0.548555f
C20102 a_8912_37509.n4 VSS 1.31827f
C20103 a_8912_37509.n5 VSS 0.502978f
C20104 a_8912_37509.t35 VSS 0.890777f
C20105 a_8912_37509.n6 VSS 1.31827f
C20106 a_8912_37509.n7 VSS 0.453882f
C20107 a_8912_37509.n8 VSS 0.459486f
C20108 a_8912_37509.n9 VSS 1.31827f
C20109 a_8912_37509.n10 VSS 0.481525f
C20110 a_8912_37509.t36 VSS 0.890777f
C20111 a_8912_37509.n11 VSS 1.31827f
C20112 a_8912_37509.n12 VSS 0.330231f
C20113 a_8912_37509.t14 VSS 0.784296f
C20114 a_8912_37509.t2 VSS 0.177274f
C20115 a_8912_37509.t11 VSS 0.177274f
C20116 a_8912_37509.n13 VSS 0.494639f
C20117 a_8912_37509.n14 VSS 2.08091f
C20118 a_8912_37509.t3 VSS 0.177274f
C20119 a_8912_37509.t0 VSS 0.177274f
C20120 a_8912_37509.n15 VSS 0.494639f
C20121 a_8912_37509.n16 VSS 1.04163f
C20122 a_8912_37509.t6 VSS 0.177274f
C20123 a_8912_37509.t7 VSS 0.177274f
C20124 a_8912_37509.n17 VSS 0.494639f
C20125 a_8912_37509.n18 VSS 1.04724f
C20126 a_8912_37509.t9 VSS 0.779123f
C20127 a_8912_37509.n19 VSS 1.13411f
C20128 a_8912_37509.t27 VSS 0.779123f
C20129 a_8912_37509.n20 VSS 1.12851f
C20130 a_8912_37509.t21 VSS 0.177274f
C20131 a_8912_37509.t17 VSS 0.177274f
C20132 a_8912_37509.n21 VSS 0.494639f
C20133 a_8912_37509.n22 VSS 1.04163f
C20134 a_8912_37509.t19 VSS 0.177274f
C20135 a_8912_37509.t22 VSS 0.177274f
C20136 a_8912_37509.n23 VSS 0.494639f
C20137 a_8912_37509.n24 VSS 1.04163f
C20138 a_8912_37509.t18 VSS 0.177274f
C20139 a_8912_37509.t26 VSS 0.177274f
C20140 a_8912_37509.n25 VSS 0.494639f
C20141 a_8912_37509.n26 VSS 1.04163f
C20142 a_8912_37509.t16 VSS 0.779123f
C20143 a_8912_37509.n27 VSS 1.59247f
C20144 a_8912_37509.n28 VSS 0.760578f
C20145 a_8912_37509.n29 VSS 1.31827f
C20146 a_8912_37509.n30 VSS 0.736298f
C20147 a_8912_37509.t5 VSS 0.76733f
C20148 a_8912_37509.n31 VSS 1.51956f
C20149 a_8912_37509.t31 VSS 0.772205f
C20150 a_8912_37509.t29 VSS 0.177274f
C20151 a_8912_37509.t28 VSS 0.177274f
C20152 a_8912_37509.n32 VSS 0.481849f
C20153 a_8912_37509.n33 VSS 1.95207f
C20154 a_8912_37509.t25 VSS 0.177274f
C20155 a_8912_37509.t24 VSS 0.177274f
C20156 a_8912_37509.n34 VSS 0.481849f
C20157 a_8912_37509.n35 VSS 0.977562f
C20158 a_8912_37509.t30 VSS 0.177274f
C20159 a_8912_37509.t20 VSS 0.177274f
C20160 a_8912_37509.n36 VSS 0.481849f
C20161 a_8912_37509.n37 VSS 0.983166f
C20162 a_8912_37509.t23 VSS 0.76733f
C20163 a_8912_37509.n38 VSS 1.06904f
C20164 a_8912_37509.t4 VSS 0.76733f
C20165 a_8912_37509.n39 VSS 1.06344f
C20166 a_8912_37509.t8 VSS 0.177274f
C20167 a_8912_37509.t12 VSS 0.177274f
C20168 a_8912_37509.n40 VSS 0.481849f
C20169 a_8912_37509.n41 VSS 0.977562f
C20170 a_8912_37509.t10 VSS 0.177274f
C20171 a_8912_37509.t1 VSS 0.177274f
C20172 a_8912_37509.n42 VSS 0.481849f
C20173 a_8912_37509.n43 VSS 0.983166f
C20174 a_8912_37509.n44 VSS 0.977562f
C20175 a_8912_37509.n45 VSS 0.481849f
C20176 a_8912_37509.t15 VSS 0.177274f
C20177 a_5088_37509.t8 VSS 0.140614f
C20178 a_5088_37509.t4 VSS 0.140614f
C20179 a_5088_37509.t1 VSS 0.140614f
C20180 a_5088_37509.n0 VSS 0.381086f
C20181 a_5088_37509.t2 VSS 0.140614f
C20182 a_5088_37509.t14 VSS 0.140614f
C20183 a_5088_37509.n1 VSS 0.376291f
C20184 a_5088_37509.n2 VSS 1.35312f
C20185 a_5088_37509.t11 VSS 0.140614f
C20186 a_5088_37509.t13 VSS 0.140614f
C20187 a_5088_37509.n3 VSS 0.376291f
C20188 a_5088_37509.n4 VSS 0.701585f
C20189 a_5088_37509.t6 VSS 0.140614f
C20190 a_5088_37509.t9 VSS 0.140614f
C20191 a_5088_37509.n5 VSS 0.376291f
C20192 a_5088_37509.n6 VSS 0.698353f
C20193 a_5088_37509.t19 VSS 0.194513f
C20194 a_5088_37509.t18 VSS 0.053336f
C20195 a_5088_37509.t16 VSS 0.053336f
C20196 a_5088_37509.n7 VSS 0.121722f
C20197 a_5088_37509.n8 VSS 0.755758f
C20198 a_5088_37509.t17 VSS 0.193609f
C20199 a_5088_37509.n9 VSS 1.98688f
C20200 a_5088_37509.n10 VSS 1.64996f
C20201 a_5088_37509.t7 VSS 0.140614f
C20202 a_5088_37509.t15 VSS 0.140614f
C20203 a_5088_37509.n11 VSS 0.360133f
C20204 a_5088_37509.n12 VSS 1.42395f
C20205 a_5088_37509.t12 VSS 0.140614f
C20206 a_5088_37509.t3 VSS 0.140614f
C20207 a_5088_37509.n13 VSS 0.360133f
C20208 a_5088_37509.n14 VSS 0.619605f
C20209 a_5088_37509.t10 VSS 0.140614f
C20210 a_5088_37509.t5 VSS 0.140614f
C20211 a_5088_37509.n15 VSS 0.360133f
C20212 a_5088_37509.n16 VSS 1.18972f
C20213 a_5088_37509.n17 VSS 0.364369f
C20214 a_5088_37509.t0 VSS 0.140614f
C20215 VDAC_P.t16 VSS 0.506361f
C20216 VDAC_P.t22 VSS 0.506152f
C20217 VDAC_P.n0 VSS 0.565956f
C20218 VDAC_P.t11 VSS 0.506152f
C20219 VDAC_P.n1 VSS 0.296568f
C20220 VDAC_P.t15 VSS 0.506152f
C20221 VDAC_P.n2 VSS 0.559117f
C20222 VDAC_P.t19 VSS 0.506361f
C20223 VDAC_P.t21 VSS 0.506152f
C20224 VDAC_P.n3 VSS 0.565956f
C20225 VDAC_P.t17 VSS 0.506152f
C20226 VDAC_P.n4 VSS 0.296568f
C20227 VDAC_P.t14 VSS 0.506152f
C20228 VDAC_P.n5 VSS 0.286437f
C20229 VDAC_P.n6 VSS 0.389891f
C20230 VDAC_P.t13 VSS 0.506324f
C20231 VDAC_P.t12 VSS 0.506152f
C20232 VDAC_P.n7 VSS 0.590358f
C20233 VDAC_P.t23 VSS 0.506152f
C20234 VDAC_P.n8 VSS 0.314549f
C20235 VDAC_P.t18 VSS 0.506152f
C20236 VDAC_P.n9 VSS -0.682165f
C20237 VDAC_P.t9 VSS 0.506152f
C20238 VDAC_P.n10 VSS -0.058656f
C20239 VDAC_P.t20 VSS 0.506152f
C20240 VDAC_P.n11 VSS 0.296568f
C20241 VDAC_P.t8 VSS 0.506152f
C20242 VDAC_P.n12 VSS 0.294714f
C20243 VDAC_P.t10 VSS 0.506154f
C20244 VDAC_P.n13 VSS 0.293364f
C20245 VDAC_P.n14 VSS 1.95614f
C20246 VDAC_P.t7 VSS 0.343978f
C20247 VDAC_P.t4 VSS 0.343978f
C20248 VDAC_P.n15 VSS 1.3174f
C20249 VDAC_P.t6 VSS 0.343978f
C20250 VDAC_P.t0 VSS 0.343978f
C20251 VDAC_P.n16 VSS 1.28659f
C20252 VDAC_P.n17 VSS 1.81217f
C20253 VDAC_P.t1 VSS 0.343978f
C20254 VDAC_P.t3 VSS 0.343978f
C20255 VDAC_P.n18 VSS 1.3174f
C20256 VDAC_P.t5 VSS 0.343978f
C20257 VDAC_P.t2 VSS 0.343978f
C20258 VDAC_P.n19 VSS 1.28659f
C20259 VDAC_P.n20 VSS 1.81477f
C20260 VDAC_P.n21 VSS 1.71275f
C20261 VDAC_P.n22 VSS 43.4479f
C20262 a_13259_45724.n0 VSS 0.017414f
C20263 a_13259_45724.t10 VSS 0.010342f
C20264 a_13259_45724.n1 VSS 0.068561f
C20265 a_13259_45724.n2 VSS 0.014887f
C20266 a_13259_45724.n3 VSS 0.533254f
C20267 a_13259_45724.t11 VSS 0.010237f
C20268 a_13259_45724.t18 VSS 0.022077f
C20269 a_13259_45724.n4 VSS 0.186314f
C20270 a_13259_45724.n5 VSS 0.016048f
C20271 a_13259_45724.t23 VSS 0.010757f
C20272 a_13259_45724.n6 VSS 0.02395f
C20273 a_13259_45724.n7 VSS 0.019305f
C20274 a_13259_45724.n8 VSS 0.188173f
C20275 a_13259_45724.t4 VSS 0.010465f
C20276 a_13259_45724.n9 VSS 0.022353f
C20277 a_13259_45724.t8 VSS 0.010465f
C20278 a_13259_45724.n10 VSS 0.015561f
C20279 a_13259_45724.n11 VSS 0.164122f
C20280 a_13259_45724.n12 VSS 0.101255f
C20281 a_13259_45724.n13 VSS 0.021024f
C20282 a_13259_45724.n14 VSS 0.209317f
C20283 a_13259_45724.n15 VSS 0.017473f
C20284 a_13259_45724.n16 VSS 0.183796f
C20285 a_13259_45724.n17 VSS 0.191922f
C20286 a_13259_45724.n18 VSS 0.148647f
C20287 a_13259_45724.n19 VSS 0.070694f
C20288 a_13259_45724.n20 VSS 0.012443f
.ends

