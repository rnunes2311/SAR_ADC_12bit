magic
tech sky130A
magscale 1 2
timestamp 1713020991
<< viali >>
rect 2053 7497 2087 7531
rect 6837 7497 6871 7531
rect 9137 7497 9171 7531
rect 10333 7497 10367 7531
rect 12081 7497 12115 7531
rect 15761 7497 15795 7531
rect 19073 7497 19107 7531
rect 26249 7497 26283 7531
rect 26709 7497 26743 7531
rect 27445 7497 27479 7531
rect 1409 7429 1443 7463
rect 3157 7429 3191 7463
rect 4905 7429 4939 7463
rect 14105 7429 14139 7463
rect 15577 7429 15611 7463
rect 22569 7429 22603 7463
rect 24593 7429 24627 7463
rect 1777 7361 1811 7395
rect 2237 7361 2271 7395
rect 2605 7361 2639 7395
rect 2697 7361 2731 7395
rect 3525 7361 3559 7395
rect 5273 7361 5307 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 6745 7361 6779 7395
rect 9045 7361 9079 7395
rect 10241 7361 10275 7395
rect 11529 7361 11563 7395
rect 11621 7361 11655 7395
rect 11989 7361 12023 7395
rect 14473 7361 14507 7395
rect 14841 7361 14875 7395
rect 15945 7361 15979 7395
rect 17325 7361 17359 7395
rect 18889 7361 18923 7395
rect 19441 7361 19475 7395
rect 19717 7361 19751 7395
rect 20637 7361 20671 7395
rect 26065 7361 26099 7395
rect 26433 7361 26467 7395
rect 26525 7361 26559 7395
rect 27169 7361 27203 7395
rect 27261 7361 27295 7395
rect 15025 7293 15059 7327
rect 19625 7293 19659 7327
rect 19993 7293 20027 7327
rect 17141 7225 17175 7259
rect 20269 7225 20303 7259
rect 22385 7225 22419 7259
rect 2421 7157 2455 7191
rect 2881 7157 2915 7191
rect 14657 7157 14691 7191
rect 15485 7157 15519 7191
rect 19533 7157 19567 7191
rect 19901 7157 19935 7191
rect 20453 7157 20487 7191
rect 20821 7157 20855 7191
rect 24501 7157 24535 7191
rect 25881 7157 25915 7191
rect 26985 7157 27019 7191
rect 1501 6953 1535 6987
rect 1869 6953 1903 6987
rect 3893 6953 3927 6987
rect 6653 6953 6687 6987
rect 8401 6953 8435 6987
rect 10149 6953 10183 6987
rect 11253 6953 11287 6987
rect 17601 6953 17635 6987
rect 18705 6953 18739 6987
rect 27445 6953 27479 6987
rect 5825 6885 5859 6919
rect 9597 6885 9631 6919
rect 20913 6885 20947 6919
rect 5181 6817 5215 6851
rect 9229 6817 9263 6851
rect 9321 6817 9355 6851
rect 11805 6817 11839 6851
rect 12449 6817 12483 6851
rect 17417 6817 17451 6851
rect 19257 6817 19291 6851
rect 19625 6817 19659 6851
rect 19717 6817 19751 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 23121 6817 23155 6851
rect 1685 6749 1719 6783
rect 2053 6749 2087 6783
rect 2421 6749 2455 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 6561 6749 6595 6783
rect 8493 6749 8527 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 10057 6749 10091 6783
rect 11621 6749 11655 6783
rect 12265 6749 12299 6783
rect 13829 6749 13863 6783
rect 15945 6749 15979 6783
rect 16037 6749 16071 6783
rect 17049 6749 17083 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 19901 6749 19935 6783
rect 20361 6749 20395 6783
rect 20821 6749 20855 6783
rect 22569 6749 22603 6783
rect 22661 6749 22695 6783
rect 22753 6749 22787 6783
rect 22937 6749 22971 6783
rect 23213 6749 23247 6783
rect 23397 6749 23431 6783
rect 26525 6749 26559 6783
rect 26893 6749 26927 6783
rect 27261 6749 27295 6783
rect 4445 6681 4479 6715
rect 4997 6681 5031 6715
rect 5549 6681 5583 6715
rect 11069 6681 11103 6715
rect 11713 6681 11747 6715
rect 13001 6681 13035 6715
rect 13645 6681 13679 6715
rect 15669 6681 15703 6715
rect 16405 6681 16439 6715
rect 18521 6681 18555 6715
rect 18737 6681 18771 6715
rect 20729 6681 20763 6715
rect 21189 6681 21223 6715
rect 22201 6681 22235 6715
rect 23305 6681 23339 6715
rect 2237 6613 2271 6647
rect 4537 6613 4571 6647
rect 4905 6613 4939 6647
rect 5457 6613 5491 6647
rect 6193 6613 6227 6647
rect 8953 6613 8987 6647
rect 10977 6613 11011 6647
rect 12081 6613 12115 6647
rect 12725 6613 12759 6647
rect 14197 6613 14231 6647
rect 17233 6613 17267 6647
rect 18889 6613 18923 6647
rect 20637 6613 20671 6647
rect 21097 6613 21131 6647
rect 22385 6613 22419 6647
rect 26709 6613 26743 6647
rect 27077 6613 27111 6647
rect 1501 6409 1535 6443
rect 5457 6409 5491 6443
rect 6469 6409 6503 6443
rect 6929 6409 6963 6443
rect 9689 6409 9723 6443
rect 11253 6409 11287 6443
rect 13277 6409 13311 6443
rect 13829 6409 13863 6443
rect 16129 6409 16163 6443
rect 19441 6409 19475 6443
rect 23857 6409 23891 6443
rect 27445 6409 27479 6443
rect 3893 6341 3927 6375
rect 16405 6341 16439 6375
rect 23305 6341 23339 6375
rect 1685 6273 1719 6307
rect 2053 6273 2087 6307
rect 5825 6273 5859 6307
rect 6837 6273 6871 6307
rect 9865 6273 9899 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 10517 6273 10551 6307
rect 11345 6273 11379 6307
rect 11529 6273 11563 6307
rect 13921 6273 13955 6307
rect 16865 6273 16899 6307
rect 17233 6273 17267 6307
rect 17693 6273 17727 6307
rect 18429 6273 18463 6307
rect 18546 6273 18580 6307
rect 19809 6273 19843 6307
rect 20269 6273 20303 6307
rect 20729 6273 20763 6307
rect 21097 6273 21131 6307
rect 21189 6273 21223 6307
rect 21373 6273 21407 6307
rect 21557 6273 21591 6307
rect 23581 6273 23615 6307
rect 26525 6273 26559 6307
rect 27261 6273 27295 6307
rect 3617 6205 3651 6239
rect 5365 6205 5399 6239
rect 5917 6205 5951 6239
rect 6009 6205 6043 6239
rect 7021 6205 7055 6239
rect 7573 6205 7607 6239
rect 7849 6205 7883 6239
rect 9597 6205 9631 6239
rect 10057 6205 10091 6239
rect 11805 6205 11839 6239
rect 13737 6205 13771 6239
rect 14381 6205 14415 6239
rect 14657 6205 14691 6239
rect 16221 6205 16255 6239
rect 17509 6205 17543 6239
rect 18705 6205 18739 6239
rect 19625 6205 19659 6239
rect 19717 6205 19751 6239
rect 19901 6205 19935 6239
rect 23673 6205 23707 6239
rect 24041 6205 24075 6239
rect 9965 6137 9999 6171
rect 16681 6137 16715 6171
rect 18153 6137 18187 6171
rect 21833 6137 21867 6171
rect 1869 6069 1903 6103
rect 10517 6069 10551 6103
rect 10793 6069 10827 6103
rect 14289 6069 14323 6103
rect 17049 6069 17083 6103
rect 19349 6069 19383 6103
rect 20177 6069 20211 6103
rect 20545 6069 20579 6103
rect 20821 6069 20855 6103
rect 21465 6069 21499 6103
rect 24133 6069 24167 6103
rect 26709 6069 26743 6103
rect 5641 5865 5675 5899
rect 8309 5865 8343 5899
rect 8953 5865 8987 5899
rect 11805 5865 11839 5899
rect 13093 5865 13127 5899
rect 15945 5865 15979 5899
rect 19073 5865 19107 5899
rect 19901 5865 19935 5899
rect 20913 5865 20947 5899
rect 21465 5865 21499 5899
rect 23673 5865 23707 5899
rect 27445 5865 27479 5899
rect 1501 5797 1535 5831
rect 12633 5797 12667 5831
rect 20545 5797 20579 5831
rect 21005 5797 21039 5831
rect 3893 5729 3927 5763
rect 5733 5729 5767 5763
rect 7481 5729 7515 5763
rect 8125 5729 8159 5763
rect 9505 5729 9539 5763
rect 9965 5729 9999 5763
rect 11713 5729 11747 5763
rect 12265 5729 12299 5763
rect 12449 5729 12483 5763
rect 12909 5729 12943 5763
rect 14381 5729 14415 5763
rect 16589 5729 16623 5763
rect 17417 5729 17451 5763
rect 17877 5729 17911 5763
rect 18153 5729 18187 5763
rect 18429 5729 18463 5763
rect 21373 5729 21407 5763
rect 22201 5729 22235 5763
rect 1685 5661 1719 5695
rect 2053 5661 2087 5695
rect 7757 5661 7791 5695
rect 7849 5661 7883 5695
rect 8493 5661 8527 5695
rect 8769 5661 8803 5695
rect 9321 5661 9355 5695
rect 13185 5661 13219 5695
rect 14105 5661 14139 5695
rect 17233 5661 17267 5695
rect 18291 5661 18325 5695
rect 19257 5661 19291 5695
rect 19405 5661 19439 5695
rect 19763 5661 19797 5695
rect 20269 5661 20303 5695
rect 20453 5661 20487 5695
rect 20637 5661 20671 5695
rect 20729 5661 20763 5695
rect 21189 5661 21223 5695
rect 21925 5661 21959 5695
rect 26893 5661 26927 5695
rect 27261 5661 27295 5695
rect 4169 5593 4203 5627
rect 6009 5593 6043 5627
rect 8217 5593 8251 5627
rect 9413 5593 9447 5627
rect 11437 5593 11471 5627
rect 13737 5593 13771 5627
rect 13921 5593 13955 5627
rect 19533 5593 19567 5627
rect 19625 5593 19659 5627
rect 20177 5593 20211 5627
rect 21465 5593 21499 5627
rect 1869 5525 1903 5559
rect 7573 5525 7607 5559
rect 8677 5525 8711 5559
rect 12173 5525 12207 5559
rect 15853 5525 15887 5559
rect 16313 5525 16347 5559
rect 16405 5525 16439 5559
rect 27077 5525 27111 5559
rect 1501 5321 1535 5355
rect 4813 5321 4847 5355
rect 5181 5321 5215 5355
rect 6377 5321 6411 5355
rect 9965 5321 9999 5355
rect 10149 5321 10183 5355
rect 11529 5321 11563 5355
rect 12541 5321 12575 5355
rect 14841 5321 14875 5355
rect 15209 5321 15243 5355
rect 19625 5321 19659 5355
rect 20361 5321 20395 5355
rect 22477 5321 22511 5355
rect 27445 5321 27479 5355
rect 8309 5253 8343 5287
rect 19441 5253 19475 5287
rect 19717 5253 19751 5287
rect 27077 5253 27111 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 2605 5185 2639 5219
rect 2881 5185 2915 5219
rect 4077 5185 4111 5219
rect 4537 5185 4571 5219
rect 6193 5185 6227 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 6837 5185 6871 5219
rect 8033 5185 8067 5219
rect 9873 5185 9907 5219
rect 10517 5185 10551 5219
rect 10977 5185 11011 5219
rect 11161 5185 11195 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 12725 5185 12759 5219
rect 13277 5185 13311 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 14381 5185 14415 5219
rect 14565 5185 14599 5219
rect 16221 5185 16255 5219
rect 16865 5185 16899 5219
rect 17233 5185 17267 5219
rect 17325 5185 17359 5219
rect 17509 5185 17543 5219
rect 17693 5185 17727 5219
rect 17969 5185 18003 5219
rect 18153 5185 18187 5219
rect 19901 5185 19935 5219
rect 19993 5185 20027 5219
rect 20177 5185 20211 5219
rect 20269 5185 20303 5219
rect 20821 5185 20855 5219
rect 22201 5185 22235 5219
rect 22397 5185 22431 5219
rect 22691 5185 22725 5219
rect 22845 5185 22879 5219
rect 23129 5175 23163 5209
rect 23397 5185 23431 5219
rect 23673 5185 23707 5219
rect 23857 5185 23891 5219
rect 26249 5185 26283 5219
rect 26801 5185 26835 5219
rect 26985 5185 27019 5219
rect 27261 5185 27295 5219
rect 3893 5117 3927 5151
rect 4353 5117 4387 5151
rect 4721 5117 4755 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 5917 5117 5951 5151
rect 10609 5117 10643 5151
rect 10793 5117 10827 5151
rect 11345 5117 11379 5151
rect 11989 5117 12023 5151
rect 12081 5117 12115 5151
rect 14749 5117 14783 5151
rect 15301 5117 15335 5151
rect 15393 5117 15427 5151
rect 15945 5117 15979 5151
rect 19073 5117 19107 5151
rect 5641 5049 5675 5083
rect 13645 5049 13679 5083
rect 15669 5049 15703 5083
rect 16957 5049 16991 5083
rect 20545 5049 20579 5083
rect 23765 5049 23799 5083
rect 1869 4981 1903 5015
rect 2237 4981 2271 5015
rect 2513 4981 2547 5015
rect 2789 4981 2823 5015
rect 4261 4981 4295 5015
rect 6101 4981 6135 5015
rect 9781 4981 9815 5015
rect 12909 4981 12943 5015
rect 15853 4981 15887 5015
rect 19441 4981 19475 5015
rect 22201 4981 22235 5015
rect 23029 4981 23063 5015
rect 26341 4981 26375 5015
rect 26617 4981 26651 5015
rect 5825 4777 5859 4811
rect 6101 4777 6135 4811
rect 9597 4777 9631 4811
rect 11989 4777 12023 4811
rect 12357 4777 12391 4811
rect 13553 4777 13587 4811
rect 14657 4777 14691 4811
rect 17141 4777 17175 4811
rect 21281 4777 21315 4811
rect 27445 4777 27479 4811
rect 1501 4709 1535 4743
rect 5917 4709 5951 4743
rect 19441 4709 19475 4743
rect 19809 4709 19843 4743
rect 22569 4709 22603 4743
rect 22753 4709 22787 4743
rect 5273 4641 5307 4675
rect 10241 4641 10275 4675
rect 12449 4641 12483 4675
rect 13369 4641 13403 4675
rect 16747 4641 16781 4675
rect 16957 4641 16991 4675
rect 21833 4641 21867 4675
rect 1685 4573 1719 4607
rect 2053 4573 2087 4607
rect 2237 4573 2271 4607
rect 2329 4573 2363 4607
rect 2605 4573 2639 4607
rect 6193 4573 6227 4607
rect 6469 4573 6503 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 7113 4573 7147 4607
rect 7277 4573 7311 4607
rect 9137 4573 9171 4607
rect 9505 4573 9539 4607
rect 12541 4573 12575 4607
rect 13001 4573 13035 4607
rect 14473 4573 14507 4607
rect 14749 4573 14783 4607
rect 16589 4573 16623 4607
rect 17417 4573 17451 4607
rect 17601 4573 17635 4607
rect 19533 4573 19567 4607
rect 19625 4573 19659 4607
rect 20269 4573 20303 4607
rect 20544 4573 20578 4607
rect 20637 4573 20671 4607
rect 20729 4573 20763 4607
rect 21097 4573 21131 4607
rect 22017 4573 22051 4607
rect 22109 4573 22143 4607
rect 23029 4573 23063 4607
rect 26341 4573 26375 4607
rect 26617 4573 26651 4607
rect 26893 4573 26927 4607
rect 27261 4573 27295 4607
rect 10517 4505 10551 4539
rect 17233 4505 17267 4539
rect 19257 4505 19291 4539
rect 22385 4505 22419 4539
rect 26433 4505 26467 4539
rect 1869 4437 1903 4471
rect 2513 4437 2547 4471
rect 5365 4437 5399 4471
rect 5457 4437 5491 4471
rect 6745 4437 6779 4471
rect 12173 4437 12207 4471
rect 13185 4437 13219 4471
rect 14197 4437 14231 4471
rect 17509 4437 17543 4471
rect 17785 4437 17819 4471
rect 19533 4437 19567 4471
rect 20913 4437 20947 4471
rect 21833 4437 21867 4471
rect 22293 4437 22327 4471
rect 26709 4437 26743 4471
rect 27077 4437 27111 4471
rect 4353 4233 4387 4267
rect 7665 4233 7699 4267
rect 9873 4233 9907 4267
rect 10977 4233 11011 4267
rect 11345 4233 11379 4267
rect 12081 4233 12115 4267
rect 17601 4233 17635 4267
rect 17693 4233 17727 4267
rect 19073 4233 19107 4267
rect 19717 4233 19751 4267
rect 9137 4165 9171 4199
rect 14907 4165 14941 4199
rect 16865 4165 16899 4199
rect 17325 4165 17359 4199
rect 19993 4165 20027 4199
rect 20453 4165 20487 4199
rect 22293 4165 22327 4199
rect 24041 4165 24075 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5457 4097 5491 4131
rect 5917 4097 5951 4131
rect 6193 4097 6227 4131
rect 6561 4097 6595 4131
rect 6929 4097 6963 4131
rect 7021 4097 7055 4131
rect 7849 4097 7883 4131
rect 8309 4097 8343 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 8953 4097 8987 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 9689 4097 9723 4131
rect 10057 4097 10091 4131
rect 11069 4097 11103 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 15485 4097 15519 4131
rect 15669 4097 15703 4131
rect 15761 4097 15795 4131
rect 15853 4097 15887 4131
rect 16681 4097 16715 4131
rect 16957 4097 16991 4131
rect 17049 4097 17083 4131
rect 17509 4097 17543 4131
rect 17877 4097 17911 4131
rect 18153 4097 18187 4131
rect 18981 4097 19015 4131
rect 19349 4097 19383 4131
rect 19625 4097 19659 4131
rect 19901 4097 19935 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 20637 4097 20671 4131
rect 20821 4097 20855 4131
rect 21097 4097 21131 4131
rect 21373 4097 21407 4131
rect 21557 4097 21591 4131
rect 22017 4097 22051 4131
rect 25973 4097 26007 4131
rect 26249 4097 26283 4131
rect 26525 4097 26559 4131
rect 26985 4097 27019 4131
rect 27261 4097 27295 4131
rect 4445 4029 4479 4063
rect 4629 4029 4663 4063
rect 7481 4029 7515 4063
rect 10793 4029 10827 4063
rect 11805 4029 11839 4063
rect 14381 4029 14415 4063
rect 14657 4029 14691 4063
rect 14749 4029 14783 4063
rect 15117 4029 15151 4063
rect 18061 4029 18095 4063
rect 18245 4029 18279 4063
rect 18337 4029 18371 4063
rect 26065 4029 26099 4063
rect 1501 3961 1535 3995
rect 2513 3961 2547 3995
rect 4905 3961 4939 3995
rect 5641 3961 5675 3995
rect 6837 3961 6871 3995
rect 8677 3961 8711 3995
rect 18521 3961 18555 3995
rect 21465 3961 21499 3995
rect 26341 3961 26375 3995
rect 27445 3961 27479 3995
rect 1869 3893 1903 3927
rect 2237 3893 2271 3927
rect 2789 3893 2823 3927
rect 3985 3893 4019 3927
rect 6009 3893 6043 3927
rect 8033 3893 8067 3927
rect 9505 3893 9539 3927
rect 10241 3893 10275 3927
rect 11897 3893 11931 3927
rect 12909 3893 12943 3927
rect 15301 3893 15335 3927
rect 16037 3893 16071 3927
rect 17233 3893 17267 3927
rect 18797 3893 18831 3927
rect 19257 3893 19291 3927
rect 26709 3893 26743 3927
rect 27077 3893 27111 3927
rect 6285 3689 6319 3723
rect 7008 3689 7042 3723
rect 13829 3689 13863 3723
rect 15025 3689 15059 3723
rect 15932 3689 15966 3723
rect 17877 3689 17911 3723
rect 27445 3689 27479 3723
rect 1501 3621 1535 3655
rect 4169 3553 4203 3587
rect 4445 3553 4479 3587
rect 6653 3553 6687 3587
rect 6745 3553 6779 3587
rect 9137 3553 9171 3587
rect 9413 3553 9447 3587
rect 11161 3553 11195 3587
rect 14473 3553 14507 3587
rect 15669 3553 15703 3587
rect 17693 3553 17727 3587
rect 18521 3553 18555 3587
rect 21833 3553 21867 3587
rect 22201 3553 22235 3587
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2329 3485 2363 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 11529 3485 11563 3519
rect 14289 3485 14323 3519
rect 14841 3485 14875 3519
rect 15209 3485 15243 3519
rect 15301 3485 15335 3519
rect 18061 3485 18095 3519
rect 19257 3485 19291 3519
rect 21373 3485 21407 3519
rect 21649 3485 21683 3519
rect 21925 3485 21959 3519
rect 23949 3485 23983 3519
rect 24501 3485 24535 3519
rect 26065 3485 26099 3519
rect 26341 3485 26375 3519
rect 26617 3485 26651 3519
rect 26893 3485 26927 3519
rect 27261 3485 27295 3519
rect 8769 3417 8803 3451
rect 11805 3417 11839 3451
rect 13553 3417 13587 3451
rect 13737 3417 13771 3451
rect 18705 3417 18739 3451
rect 19533 3417 19567 3451
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 14105 3349 14139 3383
rect 18613 3349 18647 3383
rect 19073 3349 19107 3383
rect 21005 3349 21039 3383
rect 21465 3349 21499 3383
rect 24593 3349 24627 3383
rect 26157 3349 26191 3383
rect 26433 3349 26467 3383
rect 26709 3349 26743 3383
rect 27077 3349 27111 3383
rect 1501 3145 1535 3179
rect 5825 3145 5859 3179
rect 7481 3145 7515 3179
rect 10793 3145 10827 3179
rect 13277 3145 13311 3179
rect 13461 3145 13495 3179
rect 13921 3145 13955 3179
rect 18889 3145 18923 3179
rect 23305 3145 23339 3179
rect 25605 3145 25639 3179
rect 27445 3145 27479 3179
rect 7849 3077 7883 3111
rect 11897 3077 11931 3111
rect 16957 3077 16991 3111
rect 18705 3077 18739 3111
rect 19901 3077 19935 3111
rect 21649 3077 21683 3111
rect 23949 3077 23983 3111
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 2697 3009 2731 3043
rect 2973 3009 3007 3043
rect 3617 3009 3651 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 9689 3009 9723 3043
rect 9873 3009 9907 3043
rect 10977 3009 11011 3043
rect 11069 3009 11103 3043
rect 11161 3009 11195 3043
rect 11345 3009 11379 3043
rect 11805 3009 11839 3043
rect 11989 3009 12023 3043
rect 12173 3009 12207 3043
rect 12265 3009 12299 3043
rect 12461 3009 12495 3043
rect 13185 3009 13219 3043
rect 13369 3009 13403 3043
rect 13829 3009 13863 3043
rect 14473 3009 14507 3043
rect 16681 3009 16715 3043
rect 19073 3009 19107 3043
rect 19165 3009 19199 3043
rect 19349 3009 19383 3043
rect 19533 3009 19567 3043
rect 19625 3009 19659 3043
rect 22845 3009 22879 3043
rect 23673 3009 23707 3043
rect 24225 3009 24259 3043
rect 24501 3009 24535 3043
rect 25513 3009 25547 3043
rect 26065 3009 26099 3043
rect 26433 3009 26467 3043
rect 26525 3009 26559 3043
rect 26985 3009 27019 3043
rect 27261 3009 27295 3043
rect 5641 2941 5675 2975
rect 6009 2941 6043 2975
rect 9597 2941 9631 2975
rect 12357 2941 12391 2975
rect 14105 2941 14139 2975
rect 14749 2941 14783 2975
rect 16497 2941 16531 2975
rect 22385 2941 22419 2975
rect 22569 2941 22603 2975
rect 23213 2941 23247 2975
rect 23765 2941 23799 2975
rect 24041 2941 24075 2975
rect 24409 2941 24443 2975
rect 27077 2941 27111 2975
rect 11621 2873 11655 2907
rect 22477 2873 22511 2907
rect 1869 2805 1903 2839
rect 2237 2805 2271 2839
rect 2605 2805 2639 2839
rect 2881 2805 2915 2839
rect 3880 2805 3914 2839
rect 5365 2805 5399 2839
rect 6193 2805 6227 2839
rect 6377 2805 6411 2839
rect 9873 2805 9907 2839
rect 19533 2805 19567 2839
rect 24593 2805 24627 2839
rect 25881 2805 25915 2839
rect 26249 2805 26283 2839
rect 26709 2805 26743 2839
rect 3249 2601 3283 2635
rect 4905 2601 4939 2635
rect 5641 2601 5675 2635
rect 6929 2601 6963 2635
rect 8493 2601 8527 2635
rect 9045 2601 9079 2635
rect 10885 2601 10919 2635
rect 12909 2601 12943 2635
rect 14841 2601 14875 2635
rect 15853 2601 15887 2635
rect 16681 2601 16715 2635
rect 18245 2601 18279 2635
rect 20085 2601 20119 2635
rect 21925 2601 21959 2635
rect 24041 2601 24075 2635
rect 25513 2601 25547 2635
rect 2421 2533 2455 2567
rect 2789 2533 2823 2567
rect 7941 2533 7975 2567
rect 23673 2533 23707 2567
rect 4905 2465 4939 2499
rect 17141 2465 17175 2499
rect 20821 2465 20855 2499
rect 23029 2465 23063 2499
rect 23397 2465 23431 2499
rect 2237 2397 2271 2431
rect 2605 2397 2639 2431
rect 2973 2397 3007 2431
rect 3065 2397 3099 2431
rect 3801 2397 3835 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 5365 2397 5399 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 6377 2397 6411 2431
rect 7113 2397 7147 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8125 2397 8159 2431
rect 8677 2397 8711 2431
rect 9229 2397 9263 2431
rect 9965 2397 9999 2431
rect 11069 2397 11103 2431
rect 12081 2397 12115 2431
rect 12725 2397 12759 2431
rect 13645 2397 13679 2431
rect 14289 2397 14323 2431
rect 14473 2397 14507 2431
rect 14657 2397 14691 2431
rect 15117 2397 15151 2431
rect 15301 2397 15335 2431
rect 15491 2397 15525 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 17049 2397 17083 2431
rect 17233 2397 17267 2431
rect 17325 2397 17359 2431
rect 18429 2397 18463 2431
rect 19533 2397 19567 2431
rect 20269 2397 20303 2431
rect 20729 2397 20763 2431
rect 20913 2397 20947 2431
rect 21005 2397 21039 2431
rect 22109 2397 22143 2431
rect 22661 2397 22695 2431
rect 22845 2397 22879 2431
rect 23213 2397 23247 2431
rect 23489 2397 23523 2431
rect 23857 2397 23891 2431
rect 24685 2397 24719 2431
rect 25329 2397 25363 2431
rect 25605 2397 25639 2431
rect 26157 2397 26191 2431
rect 26525 2397 26559 2431
rect 27169 2397 27203 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 5457 2329 5491 2363
rect 7297 2329 7331 2363
rect 14565 2329 14599 2363
rect 15209 2329 15243 2363
rect 22753 2329 22787 2363
rect 27537 2329 27571 2363
rect 2053 2261 2087 2295
rect 3985 2261 4019 2295
rect 4445 2261 4479 2295
rect 5089 2261 5123 2295
rect 6561 2261 6595 2295
rect 8309 2261 8343 2295
rect 10149 2261 10183 2295
rect 11897 2261 11931 2295
rect 13829 2261 13863 2295
rect 15669 2261 15703 2295
rect 17509 2261 17543 2295
rect 19349 2261 19383 2295
rect 21189 2261 21223 2295
rect 24869 2261 24903 2295
rect 25789 2261 25823 2295
rect 26341 2261 26375 2295
rect 26709 2261 26743 2295
<< metal1 >>
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 24302 8004 24308 8016
rect 10376 7976 24308 8004
rect 10376 7964 10382 7976
rect 24302 7964 24308 7976
rect 24360 7964 24366 8016
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 17310 7936 17316 7948
rect 1728 7908 17316 7936
rect 1728 7896 1734 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 26878 7868 26884 7880
rect 8812 7840 26884 7868
rect 8812 7828 8818 7840
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 23842 7800 23848 7812
rect 2746 7772 23848 7800
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 2746 7732 2774 7772
rect 23842 7760 23848 7772
rect 23900 7760 23906 7812
rect 2280 7704 2774 7732
rect 2280 7692 2286 7704
rect 1104 7642 27876 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 27876 7642
rect 1104 7568 27876 7590
rect 1026 7488 1032 7540
rect 1084 7528 1090 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1084 7500 2053 7528
rect 1084 7488 1090 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 5994 7488 6000 7540
rect 6052 7488 6058 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6604 7500 6837 7528
rect 6604 7488 6610 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8352 7500 9137 7528
rect 8352 7488 8358 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10100 7500 10333 7528
rect 10100 7488 10106 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11848 7500 12081 7528
rect 11848 7488 11854 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 12406 7500 15240 7528
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 1397 7463 1455 7469
rect 1397 7460 1409 7463
rect 1360 7432 1409 7460
rect 1360 7420 1366 7432
rect 1397 7429 1409 7432
rect 1443 7429 1455 7463
rect 1397 7423 1455 7429
rect 1780 7432 3096 7460
rect 1780 7401 1808 7432
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 2590 7352 2596 7404
rect 2648 7352 2654 7404
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 2700 7324 2728 7355
rect 1176 7296 2728 7324
rect 1176 7284 1182 7296
rect 3068 7256 3096 7432
rect 3142 7420 3148 7472
rect 3200 7420 3206 7472
rect 4706 7420 4712 7472
rect 4764 7460 4770 7472
rect 4893 7463 4951 7469
rect 4893 7460 4905 7463
rect 4764 7432 4905 7460
rect 4764 7420 4770 7432
rect 4893 7429 4905 7432
rect 4939 7429 4951 7463
rect 6012 7460 6040 7488
rect 12406 7460 12434 7500
rect 6012 7432 12434 7460
rect 4893 7423 4951 7429
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 14093 7463 14151 7469
rect 14093 7460 14105 7463
rect 13596 7432 14105 7460
rect 13596 7420 13602 7432
rect 14093 7429 14105 7432
rect 14139 7429 14151 7463
rect 14093 7423 14151 7429
rect 14292 7432 14872 7460
rect 14292 7404 14320 7432
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5307 7364 5549 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 9030 7352 9036 7404
rect 9088 7352 9094 7404
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11655 7364 11989 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 14844 7401 14872 7432
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 6972 7296 15025 7324
rect 6972 7284 6978 7296
rect 15013 7293 15025 7296
rect 15059 7324 15071 7327
rect 15102 7324 15108 7336
rect 15059 7296 15108 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15212 7324 15240 7500
rect 15286 7488 15292 7540
rect 15344 7488 15350 7540
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7497 15807 7531
rect 15749 7491 15807 7497
rect 15304 7392 15332 7488
rect 15565 7463 15623 7469
rect 15565 7429 15577 7463
rect 15611 7460 15623 7463
rect 15764 7460 15792 7491
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 19061 7531 19119 7537
rect 19061 7497 19073 7531
rect 19107 7528 19119 7531
rect 22738 7528 22744 7540
rect 19107 7500 22744 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 26237 7531 26295 7537
rect 26237 7528 26249 7531
rect 22848 7500 26249 7528
rect 15611 7432 15792 7460
rect 15611 7429 15623 7432
rect 15565 7423 15623 7429
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 15304 7364 15945 7392
rect 15933 7361 15945 7364
rect 15979 7361 15991 7395
rect 17052 7392 17080 7488
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17052 7364 17325 7392
rect 15933 7355 15991 7361
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 18800 7392 18828 7488
rect 18984 7432 20484 7460
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18800 7364 18889 7392
rect 17313 7355 17371 7361
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 18984 7324 19012 7432
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19536 7364 19717 7392
rect 15212 7296 19012 7324
rect 8294 7256 8300 7268
rect 3068 7228 8300 7256
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 17129 7259 17187 7265
rect 17129 7256 17141 7259
rect 14424 7228 17141 7256
rect 14424 7216 14430 7228
rect 17129 7225 17141 7228
rect 17175 7225 17187 7259
rect 19536 7256 19564 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 19659 7296 19993 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 19981 7293 19993 7296
rect 20027 7324 20039 7327
rect 20070 7324 20076 7336
rect 20027 7296 20076 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 20456 7324 20484 7432
rect 20530 7420 20536 7472
rect 20588 7420 20594 7472
rect 22278 7420 22284 7472
rect 22336 7460 22342 7472
rect 22557 7463 22615 7469
rect 22557 7460 22569 7463
rect 22336 7432 22569 7460
rect 22336 7420 22342 7432
rect 22557 7429 22569 7432
rect 22603 7429 22615 7463
rect 22557 7423 22615 7429
rect 20548 7392 20576 7420
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 20548 7364 20637 7392
rect 20625 7361 20637 7364
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 22848 7324 22876 7500
rect 26237 7497 26249 7500
rect 26283 7497 26295 7531
rect 26237 7491 26295 7497
rect 26694 7488 26700 7540
rect 26752 7488 26758 7540
rect 27430 7488 27436 7540
rect 27488 7488 27494 7540
rect 27522 7488 27528 7540
rect 27580 7488 27586 7540
rect 24026 7420 24032 7472
rect 24084 7460 24090 7472
rect 24581 7463 24639 7469
rect 24581 7460 24593 7463
rect 24084 7432 24593 7460
rect 24084 7420 24090 7432
rect 24581 7429 24593 7432
rect 24627 7429 24639 7463
rect 24581 7423 24639 7429
rect 25774 7420 25780 7472
rect 25832 7460 25838 7472
rect 27540 7460 27568 7488
rect 25832 7432 26096 7460
rect 25832 7420 25838 7432
rect 26068 7401 26096 7432
rect 27172 7432 27568 7460
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 27172 7401 27200 7432
rect 26513 7395 26571 7401
rect 26513 7361 26525 7395
rect 26559 7361 26571 7395
rect 26513 7355 26571 7361
rect 27157 7395 27215 7401
rect 27157 7361 27169 7395
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 20456 7296 22876 7324
rect 23014 7284 23020 7336
rect 23072 7324 23078 7336
rect 26528 7324 26556 7355
rect 23072 7296 26556 7324
rect 23072 7284 23078 7296
rect 17129 7219 17187 7225
rect 18708 7228 19564 7256
rect 20257 7259 20315 7265
rect 18708 7200 18736 7228
rect 20257 7225 20269 7259
rect 20303 7225 20315 7259
rect 20257 7219 20315 7225
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 5810 7188 5816 7200
rect 2915 7160 5816 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 14642 7148 14648 7200
rect 14700 7148 14706 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15436 7160 15485 7188
rect 15436 7148 15442 7160
rect 15473 7157 15485 7160
rect 15519 7188 15531 7191
rect 16390 7188 16396 7200
rect 15519 7160 16396 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 18690 7148 18696 7200
rect 18748 7148 18754 7200
rect 19518 7148 19524 7200
rect 19576 7148 19582 7200
rect 19886 7148 19892 7200
rect 19944 7148 19950 7200
rect 19978 7148 19984 7200
rect 20036 7188 20042 7200
rect 20272 7188 20300 7219
rect 21634 7216 21640 7268
rect 21692 7256 21698 7268
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 21692 7228 22385 7256
rect 21692 7216 21698 7228
rect 22373 7225 22385 7228
rect 22419 7225 22431 7259
rect 22373 7219 22431 7225
rect 23952 7228 25912 7256
rect 20346 7188 20352 7200
rect 20036 7160 20352 7188
rect 20036 7148 20042 7160
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20438 7148 20444 7200
rect 20496 7148 20502 7200
rect 20809 7191 20867 7197
rect 20809 7157 20821 7191
rect 20855 7188 20867 7191
rect 20898 7188 20904 7200
rect 20855 7160 20904 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 20990 7148 20996 7200
rect 21048 7188 21054 7200
rect 23952 7188 23980 7228
rect 21048 7160 23980 7188
rect 21048 7148 21054 7160
rect 24486 7148 24492 7200
rect 24544 7148 24550 7200
rect 25884 7197 25912 7228
rect 26326 7216 26332 7268
rect 26384 7256 26390 7268
rect 27264 7256 27292 7355
rect 26384 7228 27292 7256
rect 26384 7216 26390 7228
rect 25869 7191 25927 7197
rect 25869 7157 25881 7191
rect 25915 7157 25927 7191
rect 25869 7151 25927 7157
rect 26970 7148 26976 7200
rect 27028 7148 27034 7200
rect 1104 7098 27876 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 27876 7098
rect 1104 7024 27876 7046
rect 1486 6944 1492 6996
rect 1544 6944 1550 6996
rect 1854 6944 1860 6996
rect 1912 6944 1918 6996
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3568 6956 3893 6984
rect 3568 6944 3574 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 5442 6984 5448 6996
rect 4212 6956 5448 6984
rect 4212 6944 4218 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6641 6987 6699 6993
rect 6641 6953 6653 6987
rect 6687 6984 6699 6987
rect 6730 6984 6736 6996
rect 6687 6956 6736 6984
rect 6687 6953 6699 6956
rect 6641 6947 6699 6953
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 9030 6984 9036 6996
rect 8435 6956 9036 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6984 10195 6987
rect 10226 6984 10232 6996
rect 10183 6956 10232 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 11514 6984 11520 6996
rect 11287 6956 11520 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 17589 6987 17647 6993
rect 14516 6956 16896 6984
rect 14516 6944 14522 6956
rect 5810 6876 5816 6928
rect 5868 6876 5874 6928
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 9232 6888 9597 6916
rect 4706 6848 4712 6860
rect 3988 6820 4712 6848
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 3988 6789 4016 6820
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5534 6848 5540 6860
rect 5215 6820 5540 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5644 6820 6224 6848
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 5644 6780 5672 6820
rect 6196 6792 6224 6820
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8662 6848 8668 6860
rect 8352 6820 8668 6848
rect 8352 6808 8358 6820
rect 8662 6808 8668 6820
rect 8720 6848 8726 6860
rect 9232 6857 9260 6888
rect 9585 6885 9597 6888
rect 9631 6885 9643 6919
rect 11054 6916 11060 6928
rect 9585 6879 9643 6885
rect 10612 6888 11060 6916
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 8720 6820 9229 6848
rect 8720 6808 8726 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9950 6848 9956 6860
rect 9355 6820 9956 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9950 6808 9956 6820
rect 10008 6848 10014 6860
rect 10502 6848 10508 6860
rect 10008 6820 10508 6848
rect 10008 6808 10014 6820
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 4295 6752 5672 6780
rect 5721 6783 5779 6789
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 4433 6715 4491 6721
rect 4433 6681 4445 6715
rect 4479 6712 4491 6715
rect 4985 6715 5043 6721
rect 4985 6712 4997 6715
rect 4479 6684 4997 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 4985 6681 4997 6684
rect 5031 6681 5043 6715
rect 4985 6675 5043 6681
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6681 5595 6715
rect 5736 6712 5764 6743
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9858 6780 9864 6792
rect 9815 6752 9864 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 6270 6712 6276 6724
rect 5736 6684 6276 6712
rect 5537 6675 5595 6681
rect 1118 6604 1124 6656
rect 1176 6644 1182 6656
rect 2225 6647 2283 6653
rect 2225 6644 2237 6647
rect 1176 6616 2237 6644
rect 1176 6604 1182 6616
rect 2225 6613 2237 6616
rect 2271 6613 2283 6647
rect 2225 6607 2283 6613
rect 4522 6604 4528 6656
rect 4580 6604 4586 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5350 6644 5356 6656
rect 4939 6616 5356 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5350 6604 5356 6616
rect 5408 6644 5414 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5408 6616 5457 6644
rect 5408 6604 5414 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5552 6644 5580 6675
rect 6270 6672 6276 6684
rect 6328 6712 6334 6724
rect 9600 6712 9628 6743
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10612 6780 10640 6888
rect 11054 6876 11060 6888
rect 11112 6916 11118 6928
rect 16868 6916 16896 6956
rect 17589 6953 17601 6987
rect 17635 6984 17647 6987
rect 18138 6984 18144 6996
rect 17635 6956 18144 6984
rect 17635 6953 17647 6956
rect 17589 6947 17647 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 20622 6984 20628 6996
rect 18748 6956 20628 6984
rect 18748 6944 18754 6956
rect 20622 6944 20628 6956
rect 20680 6984 20686 6996
rect 21450 6984 21456 6996
rect 20680 6956 21456 6984
rect 20680 6944 20686 6956
rect 21450 6944 21456 6956
rect 21508 6984 21514 6996
rect 24486 6984 24492 6996
rect 21508 6956 24492 6984
rect 21508 6944 21514 6956
rect 24486 6944 24492 6956
rect 24544 6944 24550 6996
rect 26970 6944 26976 6996
rect 27028 6944 27034 6996
rect 27430 6944 27436 6996
rect 27488 6944 27494 6996
rect 11112 6888 11928 6916
rect 11112 6876 11118 6888
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 10744 6820 11805 6848
rect 10744 6808 10750 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11900 6848 11928 6888
rect 12360 6888 12664 6916
rect 16868 6888 19288 6916
rect 12360 6848 12388 6888
rect 11900 6820 12388 6848
rect 11793 6811 11851 6817
rect 10284 6752 10640 6780
rect 10284 6740 10290 6752
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11020 6752 11621 6780
rect 11020 6740 11026 6752
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12360 6780 12388 6820
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12636 6848 12664 6888
rect 14090 6848 14096 6860
rect 12483 6820 12572 6848
rect 12636 6820 14096 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12299 6752 12388 6780
rect 12544 6780 12572 6820
rect 14090 6808 14096 6820
rect 14148 6848 14154 6860
rect 14274 6848 14280 6860
rect 14148 6820 14280 6848
rect 14148 6808 14154 6820
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 15010 6848 15016 6860
rect 14332 6820 15016 6848
rect 14332 6808 14338 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15620 6820 16068 6848
rect 15620 6808 15626 6820
rect 16040 6792 16068 6820
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 19260 6857 19288 6888
rect 19886 6876 19892 6928
rect 19944 6916 19950 6928
rect 19944 6888 20024 6916
rect 19944 6876 19950 6888
rect 19996 6857 20024 6888
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 20901 6919 20959 6925
rect 20901 6916 20913 6919
rect 20128 6888 20913 6916
rect 20128 6876 20134 6888
rect 20901 6885 20913 6888
rect 20947 6916 20959 6919
rect 26988 6916 27016 6944
rect 20947 6888 27016 6916
rect 20947 6885 20959 6888
rect 20901 6879 20959 6885
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16172 6820 17417 6848
rect 16172 6808 16178 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6817 19303 6851
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 19245 6811 19303 6817
rect 19352 6820 19625 6848
rect 13170 6780 13176 6792
rect 12544 6752 13176 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6780 13875 6783
rect 14366 6780 14372 6792
rect 13863 6752 14372 6780
rect 13863 6749 13875 6752
rect 13817 6743 13875 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 9876 6712 9904 6740
rect 10870 6712 10876 6724
rect 6328 6684 9674 6712
rect 9876 6684 10876 6712
rect 6328 6672 6334 6684
rect 5718 6644 5724 6656
rect 5552 6616 5724 6644
rect 5445 6607 5503 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6181 6647 6239 6653
rect 6181 6613 6193 6647
rect 6227 6644 6239 6647
rect 6362 6644 6368 6656
rect 6227 6616 6368 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8628 6616 8953 6644
rect 8628 6604 8634 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 9646 6644 9674 6684
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 11146 6712 11152 6724
rect 11103 6684 11152 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 11701 6715 11759 6721
rect 11701 6681 11713 6715
rect 11747 6712 11759 6715
rect 11747 6684 12848 6712
rect 11747 6681 11759 6684
rect 11701 6675 11759 6681
rect 9766 6644 9772 6656
rect 9646 6616 9772 6644
rect 8941 6607 8999 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10965 6647 11023 6653
rect 10965 6644 10977 6647
rect 10192 6616 10977 6644
rect 10192 6604 10198 6616
rect 10965 6613 10977 6616
rect 11011 6644 11023 6647
rect 11422 6644 11428 6656
rect 11011 6616 11428 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 12066 6604 12072 6656
rect 12124 6604 12130 6656
rect 12710 6604 12716 6656
rect 12768 6604 12774 6656
rect 12820 6644 12848 6684
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13446 6712 13452 6724
rect 13044 6684 13452 6712
rect 13044 6672 13050 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 13633 6715 13691 6721
rect 13633 6681 13645 6715
rect 13679 6712 13691 6715
rect 13722 6712 13728 6724
rect 13679 6684 13728 6712
rect 13679 6681 13691 6684
rect 13633 6675 13691 6681
rect 13722 6672 13728 6684
rect 13780 6672 13786 6724
rect 15562 6712 15568 6724
rect 15226 6684 15568 6712
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 15654 6672 15660 6724
rect 15712 6672 15718 6724
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 15948 6712 15976 6743
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16080 6752 16620 6780
rect 16080 6740 16086 6752
rect 15804 6684 15976 6712
rect 15804 6672 15810 6684
rect 16390 6672 16396 6724
rect 16448 6672 16454 6724
rect 16592 6712 16620 6752
rect 17034 6740 17040 6792
rect 17092 6740 17098 6792
rect 19058 6780 19064 6792
rect 17144 6752 19064 6780
rect 17144 6712 17172 6752
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 16592 6684 17172 6712
rect 18506 6672 18512 6724
rect 18564 6672 18570 6724
rect 18725 6715 18783 6721
rect 18725 6681 18737 6715
rect 18771 6712 18783 6715
rect 19242 6712 19248 6724
rect 18771 6684 19248 6712
rect 18771 6681 18783 6684
rect 18725 6675 18783 6681
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 12820 6616 14197 6644
rect 14185 6613 14197 6616
rect 14231 6644 14243 6647
rect 16482 6644 16488 6656
rect 14231 6616 16488 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17310 6644 17316 6656
rect 17267 6616 17316 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 18874 6604 18880 6656
rect 18932 6604 18938 6656
rect 19352 6644 19380 6820
rect 19613 6817 19625 6820
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 19705 6851 19763 6857
rect 19705 6817 19717 6851
rect 19751 6848 19763 6851
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 19751 6820 19993 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 19981 6817 19993 6820
rect 20027 6817 20039 6851
rect 19981 6811 20039 6817
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20990 6848 20996 6860
rect 20824 6820 20996 6848
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 19536 6712 19564 6743
rect 19794 6740 19800 6792
rect 19852 6780 19858 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19852 6752 19901 6780
rect 19852 6740 19858 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 20128 6752 20361 6780
rect 20128 6740 20134 6752
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 20824 6789 20852 6820
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21634 6848 21640 6860
rect 21140 6820 21640 6848
rect 21140 6808 21146 6820
rect 21634 6808 21640 6820
rect 21692 6808 21698 6860
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6848 23167 6851
rect 23290 6848 23296 6860
rect 23155 6820 23296 6848
rect 23155 6817 23167 6820
rect 23109 6811 23167 6817
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 20809 6783 20867 6789
rect 20809 6780 20821 6783
rect 20588 6752 20821 6780
rect 20588 6740 20594 6752
rect 20809 6749 20821 6752
rect 20855 6749 20867 6783
rect 22462 6780 22468 6792
rect 20809 6743 20867 6749
rect 21008 6752 22468 6780
rect 20717 6715 20775 6721
rect 20717 6712 20729 6715
rect 19536 6684 20729 6712
rect 20717 6681 20729 6684
rect 20763 6681 20775 6715
rect 21008 6712 21036 6752
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6749 22615 6783
rect 22557 6743 22615 6749
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 20717 6675 20775 6681
rect 20824 6684 21036 6712
rect 20824 6656 20852 6684
rect 21174 6672 21180 6724
rect 21232 6672 21238 6724
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 22572 6712 22600 6743
rect 22244 6684 22600 6712
rect 22244 6672 22250 6684
rect 22664 6656 22692 6743
rect 22738 6740 22744 6792
rect 22796 6740 22802 6792
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 22848 6752 22937 6780
rect 22848 6712 22876 6752
rect 22925 6749 22937 6752
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23198 6740 23204 6792
rect 23256 6740 23262 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 26510 6740 26516 6792
rect 26568 6740 26574 6792
rect 26786 6740 26792 6792
rect 26844 6780 26850 6792
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26844 6752 26893 6780
rect 26844 6740 26850 6752
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 26881 6743 26939 6749
rect 26970 6740 26976 6792
rect 27028 6780 27034 6792
rect 27249 6783 27307 6789
rect 27249 6780 27261 6783
rect 27028 6752 27261 6780
rect 27028 6740 27034 6752
rect 27249 6749 27261 6752
rect 27295 6749 27307 6783
rect 27249 6743 27307 6749
rect 23293 6715 23351 6721
rect 23293 6712 23305 6715
rect 22848 6684 23305 6712
rect 22848 6656 22876 6684
rect 23293 6681 23305 6684
rect 23339 6681 23351 6715
rect 23293 6675 23351 6681
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 19352 6616 20637 6644
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 20806 6604 20812 6656
rect 20864 6604 20870 6656
rect 21082 6604 21088 6656
rect 21140 6604 21146 6656
rect 22370 6604 22376 6656
rect 22428 6604 22434 6656
rect 22646 6604 22652 6656
rect 22704 6604 22710 6656
rect 22830 6604 22836 6656
rect 22888 6604 22894 6656
rect 26694 6604 26700 6656
rect 26752 6604 26758 6656
rect 27062 6604 27068 6656
rect 27120 6604 27126 6656
rect 1104 6554 27876 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 27876 6554
rect 1104 6480 27876 6502
rect 950 6400 956 6452
rect 1008 6440 1014 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 1008 6412 1501 6440
rect 1008 6400 1014 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 4522 6440 4528 6452
rect 1489 6403 1547 6409
rect 3896 6412 4528 6440
rect 3896 6381 3924 6412
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 4764 6412 5457 6440
rect 4764 6400 4770 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 6457 6443 6515 6449
rect 6457 6409 6469 6443
rect 6503 6440 6515 6443
rect 6546 6440 6552 6452
rect 6503 6412 6552 6440
rect 6503 6409 6515 6412
rect 6457 6403 6515 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6914 6400 6920 6452
rect 6972 6400 6978 6452
rect 7024 6412 9168 6440
rect 3881 6375 3939 6381
rect 3881 6341 3893 6375
rect 3927 6341 3939 6375
rect 3881 6335 3939 6341
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 6730 6372 6736 6384
rect 5408 6344 6736 6372
rect 5408 6332 5414 6344
rect 6730 6332 6736 6344
rect 6788 6372 6794 6384
rect 7024 6372 7052 6412
rect 9140 6384 9168 6412
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9456 6412 9689 6440
rect 9456 6400 9462 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 10244 6412 10824 6440
rect 7742 6372 7748 6384
rect 6788 6344 7052 6372
rect 7576 6344 7748 6372
rect 6788 6332 6794 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1946 6304 1952 6316
rect 1719 6276 1952 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 5442 6304 5448 6316
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 3878 6236 3884 6248
rect 3651 6208 3884 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 1034 6128 1040 6180
rect 1092 6168 1098 6180
rect 5000 6168 5028 6290
rect 5368 6276 5448 6304
rect 5368 6245 5396 6276
rect 5442 6264 5448 6276
rect 5500 6304 5506 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5500 6276 5825 6304
rect 5500 6264 5506 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6144 6276 6837 6304
rect 6144 6264 6150 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 7576 6304 7604 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 10244 6372 10272 6412
rect 9180 6344 10272 6372
rect 10336 6344 10640 6372
rect 9180 6332 9186 6344
rect 6825 6267 6883 6273
rect 7024 6276 7604 6304
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 5902 6196 5908 6248
rect 5960 6196 5966 6248
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 6638 6236 6644 6248
rect 6043 6208 6644 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 6638 6196 6644 6208
rect 6696 6236 6702 6248
rect 7024 6245 7052 6276
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9214 6304 9220 6316
rect 8996 6276 9220 6304
rect 8996 6264 9002 6276
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9858 6313 9864 6316
rect 9853 6304 9864 6313
rect 9819 6276 9864 6304
rect 9853 6267 9864 6276
rect 9858 6264 9864 6267
rect 9916 6264 9922 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10336 6313 10364 6344
rect 10612 6316 10640 6344
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10410 6264 10416 6316
rect 10468 6264 10474 6316
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10796 6304 10824 6412
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 11241 6443 11299 6449
rect 11241 6440 11253 6443
rect 10928 6412 11253 6440
rect 10928 6400 10934 6412
rect 11241 6409 11253 6412
rect 11287 6440 11299 6443
rect 12434 6440 12440 6452
rect 11287 6412 12440 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 12768 6412 12940 6440
rect 12768 6400 12774 6412
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 11480 6344 11560 6372
rect 11480 6332 11486 6344
rect 10796 6276 11192 6304
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6696 6208 7021 6236
rect 6696 6196 6702 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 5442 6168 5448 6180
rect 1092 6140 1900 6168
rect 5000 6140 5448 6168
rect 1092 6128 1098 6140
rect 1872 6109 1900 6140
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 7576 6112 7604 6199
rect 7834 6196 7840 6248
rect 7892 6196 7898 6248
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 9631 6208 9665 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 9600 6168 9628 6199
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 10045 6239 10103 6245
rect 10045 6236 10057 6239
rect 9824 6208 10057 6236
rect 9824 6196 9830 6208
rect 10045 6205 10057 6208
rect 10091 6236 10103 6239
rect 10091 6208 11100 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 9364 6140 9965 6168
rect 9364 6128 9370 6140
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 10134 6128 10140 6180
rect 10192 6128 10198 6180
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 7006 6100 7012 6112
rect 2096 6072 7012 6100
rect 2096 6060 2102 6072
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8018 6100 8024 6112
rect 7616 6072 8024 6100
rect 7616 6060 7622 6072
rect 8018 6060 8024 6072
rect 8076 6100 8082 6112
rect 10152 6100 10180 6128
rect 8076 6072 10180 6100
rect 8076 6060 8082 6072
rect 10502 6060 10508 6112
rect 10560 6060 10566 6112
rect 10778 6060 10784 6112
rect 10836 6060 10842 6112
rect 11072 6100 11100 6208
rect 11164 6168 11192 6276
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11532 6313 11560 6344
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 11296 6276 11345 6304
rect 11296 6264 11302 6276
rect 11333 6273 11345 6276
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 11514 6168 11520 6180
rect 11164 6140 11520 6168
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 11882 6100 11888 6112
rect 11072 6072 11888 6100
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12912 6100 12940 6412
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 13228 6412 13277 6440
rect 13228 6400 13234 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6440 13875 6443
rect 14642 6440 14648 6452
rect 13863 6412 14648 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 16114 6440 16120 6452
rect 15028 6412 16120 6440
rect 15028 6372 15056 6412
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16408 6412 19380 6440
rect 16022 6372 16028 6384
rect 14016 6344 15056 6372
rect 15870 6344 16028 6372
rect 14016 6316 14044 6344
rect 16022 6332 16028 6344
rect 16080 6332 16086 6384
rect 16408 6381 16436 6412
rect 16393 6375 16451 6381
rect 16393 6341 16405 6375
rect 16439 6341 16451 6375
rect 19352 6372 19380 6412
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 20588 6412 21128 6440
rect 20588 6400 20594 6412
rect 20806 6372 20812 6384
rect 19352 6344 20812 6372
rect 16393 6335 16451 6341
rect 20806 6332 20812 6344
rect 20864 6332 20870 6384
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13596 6276 13921 6304
rect 13596 6264 13602 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 13998 6264 14004 6316
rect 14056 6264 14062 6316
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 14274 6236 14280 6248
rect 13771 6208 14280 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 14415 6208 14504 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 14476 6112 14504 6208
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 15010 6196 15016 6248
rect 15068 6236 15074 6248
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 15068 6208 16221 6236
rect 15068 6196 15074 6208
rect 16209 6205 16221 6208
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 16868 6236 16896 6267
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 17000 6276 17233 6304
rect 17000 6264 17006 6276
rect 17221 6273 17233 6276
rect 17267 6304 17279 6307
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 17267 6276 17693 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 18414 6264 18420 6316
rect 18472 6264 18478 6316
rect 18534 6307 18592 6313
rect 18534 6304 18546 6307
rect 18524 6273 18546 6304
rect 18580 6273 18592 6307
rect 18524 6267 18592 6273
rect 17034 6236 17040 6248
rect 16868 6208 17040 6236
rect 16669 6171 16727 6177
rect 16669 6168 16681 6171
rect 15672 6140 16681 6168
rect 12032 6072 12940 6100
rect 14277 6103 14335 6109
rect 12032 6060 12038 6072
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14366 6100 14372 6112
rect 14323 6072 14372 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 14458 6060 14464 6112
rect 14516 6060 14522 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 15672 6100 15700 6140
rect 16669 6137 16681 6140
rect 16715 6137 16727 6171
rect 16669 6131 16727 6137
rect 15436 6072 15700 6100
rect 15436 6060 15442 6072
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16868 6100 16896 6208
rect 17034 6196 17040 6208
rect 17092 6236 17098 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 17092 6208 17509 6236
rect 17092 6196 17098 6208
rect 17497 6205 17509 6208
rect 17543 6205 17555 6239
rect 18524 6236 18552 6267
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 19484 6276 19809 6304
rect 19484 6264 19490 6276
rect 19797 6273 19809 6276
rect 19843 6304 19855 6307
rect 19978 6304 19984 6316
rect 19843 6276 19984 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20622 6304 20628 6316
rect 20303 6276 20628 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 21100 6313 21128 6412
rect 21450 6400 21456 6452
rect 21508 6400 21514 6452
rect 21634 6400 21640 6452
rect 21692 6400 21698 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22428 6412 23526 6440
rect 22428 6400 22434 6412
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21223 6276 21373 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21361 6273 21373 6276
rect 21407 6304 21419 6307
rect 21468 6304 21496 6400
rect 21407 6276 21496 6304
rect 21545 6307 21603 6313
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 21545 6273 21557 6307
rect 21591 6304 21603 6307
rect 21652 6304 21680 6400
rect 22738 6332 22744 6384
rect 22796 6332 22802 6384
rect 23290 6332 23296 6384
rect 23348 6332 23354 6384
rect 23498 6372 23526 6412
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 23900 6412 26464 6440
rect 23900 6400 23906 6412
rect 26436 6384 26464 6412
rect 27430 6400 27436 6452
rect 27488 6400 27494 6452
rect 23498 6344 23612 6372
rect 23584 6313 23612 6344
rect 26418 6332 26424 6384
rect 26476 6332 26482 6384
rect 21591 6276 21680 6304
rect 23569 6307 23627 6313
rect 21591 6273 21603 6276
rect 21545 6267 21603 6273
rect 23569 6273 23581 6307
rect 23615 6273 23627 6307
rect 23569 6267 23627 6273
rect 17497 6199 17555 6205
rect 17604 6208 18552 6236
rect 17218 6128 17224 6180
rect 17276 6168 17282 6180
rect 17604 6168 17632 6208
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19116 6208 19625 6236
rect 19116 6196 19122 6208
rect 19613 6205 19625 6208
rect 19659 6205 19671 6239
rect 19613 6199 19671 6205
rect 19702 6196 19708 6248
rect 19760 6196 19766 6248
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 20732 6236 20760 6267
rect 24302 6264 24308 6316
rect 24360 6304 24366 6316
rect 26513 6307 26571 6313
rect 26513 6304 26525 6307
rect 24360 6276 26525 6304
rect 24360 6264 24366 6276
rect 26513 6273 26525 6276
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 27249 6307 27307 6313
rect 27249 6273 27261 6307
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 20732 6208 21128 6236
rect 17276 6140 17632 6168
rect 18141 6171 18199 6177
rect 17276 6128 17282 6140
rect 18141 6137 18153 6171
rect 18187 6137 18199 6171
rect 19518 6168 19524 6180
rect 18141 6131 18199 6137
rect 19076 6140 19524 6168
rect 16264 6072 16896 6100
rect 16264 6060 16270 6072
rect 17034 6060 17040 6112
rect 17092 6060 17098 6112
rect 18156 6100 18184 6131
rect 18414 6100 18420 6112
rect 18156 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6100 18478 6112
rect 19076 6100 19104 6140
rect 19518 6128 19524 6140
rect 19576 6168 19582 6180
rect 20254 6168 20260 6180
rect 19576 6140 20260 6168
rect 19576 6128 19582 6140
rect 20254 6128 20260 6140
rect 20312 6168 20318 6180
rect 21100 6168 21128 6208
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 21784 6208 23520 6236
rect 21784 6196 21790 6208
rect 21266 6168 21272 6180
rect 20312 6140 20852 6168
rect 21100 6140 21272 6168
rect 20312 6128 20318 6140
rect 18472 6072 19104 6100
rect 18472 6060 18478 6072
rect 19334 6060 19340 6112
rect 19392 6060 19398 6112
rect 20165 6103 20223 6109
rect 20165 6069 20177 6103
rect 20211 6100 20223 6103
rect 20346 6100 20352 6112
rect 20211 6072 20352 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 20824 6109 20852 6140
rect 21266 6128 21272 6140
rect 21324 6168 21330 6180
rect 21821 6171 21879 6177
rect 21821 6168 21833 6171
rect 21324 6140 21833 6168
rect 21324 6128 21330 6140
rect 21821 6137 21833 6140
rect 21867 6137 21879 6171
rect 23492 6168 23520 6208
rect 23658 6196 23664 6248
rect 23716 6196 23722 6248
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23992 6208 24041 6236
rect 23992 6196 23998 6208
rect 24029 6205 24041 6208
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 27264 6168 27292 6267
rect 23492 6140 27292 6168
rect 21821 6131 21879 6137
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 20496 6072 20545 6100
rect 20496 6060 20502 6072
rect 20533 6069 20545 6072
rect 20579 6069 20591 6103
rect 20533 6063 20591 6069
rect 20809 6103 20867 6109
rect 20809 6069 20821 6103
rect 20855 6100 20867 6103
rect 20990 6100 20996 6112
rect 20855 6072 20996 6100
rect 20855 6069 20867 6072
rect 20809 6063 20867 6069
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 21450 6060 21456 6112
rect 21508 6060 21514 6112
rect 21836 6100 21864 6131
rect 22554 6100 22560 6112
rect 21836 6072 22560 6100
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 22738 6060 22744 6112
rect 22796 6100 22802 6112
rect 23290 6100 23296 6112
rect 22796 6072 23296 6100
rect 22796 6060 22802 6072
rect 23290 6060 23296 6072
rect 23348 6060 23354 6112
rect 24118 6060 24124 6112
rect 24176 6060 24182 6112
rect 26694 6060 26700 6112
rect 26752 6060 26758 6112
rect 1104 6010 27876 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 27876 6010
rect 1104 5936 27876 5958
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 6086 5896 6092 5908
rect 5675 5868 6092 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 6546 5896 6552 5908
rect 6236 5868 6552 5896
rect 6236 5856 6242 5868
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7558 5896 7564 5908
rect 7024 5868 7564 5896
rect 950 5788 956 5840
rect 1008 5828 1014 5840
rect 1489 5831 1547 5837
rect 1489 5828 1501 5831
rect 1008 5800 1501 5828
rect 1008 5788 1014 5800
rect 1489 5797 1501 5800
rect 1535 5797 1547 5831
rect 1489 5791 1547 5797
rect 3878 5720 3884 5772
rect 3936 5760 3942 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 3936 5732 5733 5760
rect 3936 5720 3942 5732
rect 5721 5729 5733 5732
rect 5767 5760 5779 5763
rect 6454 5760 6460 5772
rect 5767 5732 6460 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6454 5720 6460 5732
rect 6512 5760 6518 5772
rect 7024 5760 7052 5868
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 7892 5868 8309 5896
rect 7892 5856 7898 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8536 5868 8953 5896
rect 8536 5856 8542 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 10686 5896 10692 5908
rect 8941 5859 8999 5865
rect 9646 5868 10692 5896
rect 8846 5828 8852 5840
rect 6512 5732 7052 5760
rect 7116 5800 8852 5828
rect 6512 5720 6518 5732
rect 7116 5704 7144 5800
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7926 5760 7932 5772
rect 7515 5732 7932 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7926 5720 7932 5732
rect 7984 5760 7990 5772
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7984 5732 8125 5760
rect 7984 5720 7990 5732
rect 8113 5729 8125 5732
rect 8159 5760 8171 5763
rect 8159 5732 9352 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 7098 5652 7104 5704
rect 7156 5652 7162 5704
rect 7742 5652 7748 5704
rect 7800 5652 7806 5704
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5691 8539 5695
rect 8662 5692 8668 5704
rect 8588 5691 8668 5692
rect 8527 5664 8668 5691
rect 8527 5663 8616 5664
rect 8527 5661 8539 5663
rect 8481 5655 8539 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9324 5701 9352 5732
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9646 5760 9674 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11790 5856 11796 5908
rect 11848 5856 11854 5908
rect 12066 5856 12072 5908
rect 12124 5856 12130 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13814 5896 13820 5908
rect 13127 5868 13820 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13814 5856 13820 5868
rect 13872 5896 13878 5908
rect 13872 5868 15424 5896
rect 13872 5856 13878 5868
rect 9548 5732 9674 5760
rect 9953 5763 10011 5769
rect 9548 5720 9554 5732
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10962 5760 10968 5772
rect 9999 5732 10968 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11698 5720 11704 5772
rect 11756 5720 11762 5772
rect 12084 5760 12112 5856
rect 12621 5831 12679 5837
rect 12621 5797 12633 5831
rect 12667 5797 12679 5831
rect 15396 5828 15424 5868
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15712 5868 15945 5896
rect 15712 5856 15718 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 18598 5896 18604 5908
rect 15933 5859 15991 5865
rect 17880 5868 18604 5896
rect 15396 5800 17448 5828
rect 12621 5791 12679 5797
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 12084 5732 12265 5760
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 12253 5723 12311 5729
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 12636 5760 12664 5791
rect 12483 5732 12664 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12894 5720 12900 5772
rect 12952 5720 12958 5772
rect 13906 5760 13912 5772
rect 13188 5732 13912 5760
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 4154 5584 4160 5636
rect 4212 5584 4218 5636
rect 5442 5624 5448 5636
rect 5382 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5624 5506 5636
rect 5902 5624 5908 5636
rect 5500 5596 5908 5624
rect 5500 5584 5506 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 5994 5584 6000 5636
rect 6052 5584 6058 5636
rect 7300 5596 7604 5624
rect 1854 5516 1860 5568
rect 1912 5516 1918 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 6178 5556 6184 5568
rect 4856 5528 6184 5556
rect 4856 5516 4862 5528
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7300 5556 7328 5596
rect 7576 5565 7604 5596
rect 8202 5584 8208 5636
rect 8260 5584 8266 5636
rect 8772 5624 8800 5655
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 12912 5692 12940 5720
rect 13188 5701 13216 5732
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 15562 5720 15568 5772
rect 15620 5720 15626 5772
rect 17420 5769 17448 5800
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 17405 5763 17463 5769
rect 16623 5732 17356 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 11940 5664 12940 5692
rect 13173 5695 13231 5701
rect 11940 5652 11946 5664
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13998 5692 14004 5704
rect 13173 5655 13231 5661
rect 13648 5664 14004 5692
rect 9030 5624 9036 5636
rect 8772 5596 9036 5624
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 9401 5627 9459 5633
rect 9401 5593 9413 5627
rect 9447 5624 9459 5627
rect 9447 5596 10180 5624
rect 9447 5593 9459 5596
rect 9401 5587 9459 5593
rect 6880 5528 7328 5556
rect 7561 5559 7619 5565
rect 6880 5516 6886 5528
rect 7561 5525 7573 5559
rect 7607 5525 7619 5559
rect 7561 5519 7619 5525
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 10152 5556 10180 5596
rect 10778 5584 10784 5636
rect 10836 5584 10842 5636
rect 11422 5584 11428 5636
rect 11480 5584 11486 5636
rect 13648 5624 13676 5664
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 15580 5692 15608 5720
rect 15502 5664 15608 5692
rect 14093 5655 14151 5661
rect 11532 5596 13676 5624
rect 11532 5556 11560 5596
rect 13722 5584 13728 5636
rect 13780 5584 13786 5636
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 14108 5624 14136 5655
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 15712 5664 17233 5692
rect 15712 5652 15718 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17328 5692 17356 5732
rect 17405 5729 17417 5763
rect 17451 5729 17463 5763
rect 17770 5760 17776 5772
rect 17405 5723 17463 5729
rect 17604 5732 17776 5760
rect 17604 5692 17632 5732
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 17880 5769 17908 5868
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 18874 5856 18880 5908
rect 18932 5856 18938 5908
rect 18966 5856 18972 5908
rect 19024 5896 19030 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 19024 5868 19073 5896
rect 19024 5856 19030 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 19889 5899 19947 5905
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 20070 5896 20076 5908
rect 19935 5868 20076 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 20901 5899 20959 5905
rect 20680 5868 20852 5896
rect 20680 5856 20686 5868
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18141 5763 18199 5769
rect 18141 5760 18153 5763
rect 18012 5732 18153 5760
rect 18012 5720 18018 5732
rect 18141 5729 18153 5732
rect 18187 5729 18199 5763
rect 18141 5723 18199 5729
rect 18414 5720 18420 5772
rect 18472 5720 18478 5772
rect 18892 5760 18920 5856
rect 19150 5788 19156 5840
rect 19208 5828 19214 5840
rect 19978 5828 19984 5840
rect 19208 5800 19984 5828
rect 19208 5788 19214 5800
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20533 5831 20591 5837
rect 20533 5797 20545 5831
rect 20579 5828 20591 5831
rect 20714 5828 20720 5840
rect 20579 5800 20720 5828
rect 20579 5797 20591 5800
rect 20533 5791 20591 5797
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 20346 5760 20352 5772
rect 18892 5732 19288 5760
rect 18322 5701 18328 5704
rect 17328 5664 17632 5692
rect 18279 5695 18328 5701
rect 17221 5655 17279 5661
rect 18279 5661 18291 5695
rect 18325 5661 18328 5695
rect 18279 5655 18328 5661
rect 18322 5652 18328 5655
rect 18380 5652 18386 5704
rect 19260 5701 19288 5732
rect 19408 5732 20352 5760
rect 19408 5701 19436 5732
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19393 5695 19451 5701
rect 19393 5661 19405 5695
rect 19439 5661 19451 5695
rect 19393 5655 19451 5661
rect 19751 5695 19809 5701
rect 19751 5661 19763 5695
rect 19797 5692 19809 5695
rect 19978 5692 19984 5704
rect 19797 5664 19984 5692
rect 19797 5661 19809 5664
rect 19751 5655 19809 5661
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 20254 5652 20260 5704
rect 20312 5652 20318 5704
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 20824 5692 20852 5868
rect 20901 5865 20913 5899
rect 20947 5896 20959 5899
rect 21082 5896 21088 5908
rect 20947 5868 21088 5896
rect 20947 5865 20959 5868
rect 20901 5859 20959 5865
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 21174 5856 21180 5908
rect 21232 5856 21238 5908
rect 21450 5856 21456 5908
rect 21508 5856 21514 5908
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 23661 5899 23719 5905
rect 23661 5896 23673 5899
rect 23440 5868 23673 5896
rect 23440 5856 23446 5868
rect 23661 5865 23673 5868
rect 23707 5865 23719 5899
rect 23661 5859 23719 5865
rect 27430 5856 27436 5908
rect 27488 5856 27494 5908
rect 20993 5831 21051 5837
rect 20993 5797 21005 5831
rect 21039 5828 21051 5831
rect 21192 5828 21220 5856
rect 21039 5800 21220 5828
rect 21039 5797 21051 5800
rect 20993 5791 21051 5797
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5760 21419 5763
rect 21542 5760 21548 5772
rect 21407 5732 21548 5760
rect 21407 5729 21419 5732
rect 21361 5723 21419 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5760 22247 5763
rect 22830 5760 22836 5772
rect 22235 5732 22836 5760
rect 22235 5729 22247 5732
rect 22189 5723 22247 5729
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 20763 5664 20852 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 14458 5624 14464 5636
rect 13955 5596 14464 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 14458 5584 14464 5596
rect 14516 5584 14522 5636
rect 16850 5624 16856 5636
rect 15856 5596 16856 5624
rect 10152 5528 11560 5556
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11664 5528 12173 5556
rect 11664 5516 11670 5528
rect 12161 5525 12173 5528
rect 12207 5556 12219 5559
rect 13538 5556 13544 5568
rect 12207 5528 13544 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 13538 5516 13544 5528
rect 13596 5556 13602 5568
rect 14366 5556 14372 5568
rect 13596 5528 14372 5556
rect 13596 5516 13602 5528
rect 14366 5516 14372 5528
rect 14424 5556 14430 5568
rect 15102 5556 15108 5568
rect 14424 5528 15108 5556
rect 14424 5516 14430 5528
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15856 5565 15884 5596
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 18966 5584 18972 5636
rect 19024 5624 19030 5636
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 19024 5596 19533 5624
rect 19024 5584 19030 5596
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19613 5627 19671 5633
rect 19613 5593 19625 5627
rect 19659 5624 19671 5627
rect 20165 5627 20223 5633
rect 20165 5624 20177 5627
rect 19659 5596 20177 5624
rect 19659 5593 19671 5596
rect 19613 5587 19671 5593
rect 20165 5593 20177 5596
rect 20211 5624 20223 5627
rect 20211 5596 20392 5624
rect 20211 5593 20223 5596
rect 20165 5587 20223 5593
rect 15841 5559 15899 5565
rect 15841 5556 15853 5559
rect 15252 5528 15853 5556
rect 15252 5516 15258 5528
rect 15841 5525 15853 5528
rect 15887 5525 15899 5559
rect 15841 5519 15899 5525
rect 16298 5516 16304 5568
rect 16356 5516 16362 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16482 5556 16488 5568
rect 16439 5528 16488 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16482 5516 16488 5528
rect 16540 5556 16546 5568
rect 20254 5556 20260 5568
rect 16540 5528 20260 5556
rect 16540 5516 16546 5528
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20364 5556 20392 5596
rect 20640 5556 20668 5655
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21048 5664 21189 5692
rect 21048 5652 21054 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21177 5655 21235 5661
rect 21376 5664 21925 5692
rect 21192 5624 21220 5655
rect 21376 5624 21404 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 23290 5652 23296 5704
rect 23348 5652 23354 5704
rect 26878 5652 26884 5704
rect 26936 5652 26942 5704
rect 27246 5652 27252 5704
rect 27304 5652 27310 5704
rect 21192 5596 21404 5624
rect 21450 5584 21456 5636
rect 21508 5584 21514 5636
rect 20364 5528 20668 5556
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 23198 5556 23204 5568
rect 20772 5528 23204 5556
rect 20772 5516 20778 5528
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 27062 5516 27068 5568
rect 27120 5516 27126 5568
rect 1104 5466 27876 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 27876 5466
rect 1104 5392 27876 5414
rect 950 5312 956 5364
rect 1008 5352 1014 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 1008 5324 1501 5352
rect 1008 5312 1014 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 1489 5315 1547 5321
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4212 5324 4813 5352
rect 4212 5312 4218 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 4948 5324 5181 5352
rect 4948 5312 4954 5324
rect 5169 5321 5181 5324
rect 5215 5352 5227 5355
rect 5350 5352 5356 5364
rect 5215 5324 5356 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5994 5312 6000 5364
rect 6052 5352 6058 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6052 5324 6377 5352
rect 6052 5312 6058 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 7576 5324 9628 5352
rect 1964 5284 1992 5312
rect 7576 5284 7604 5324
rect 1964 5256 7604 5284
rect 8297 5287 8355 5293
rect 8297 5253 8309 5287
rect 8343 5284 8355 5287
rect 8570 5284 8576 5296
rect 8343 5256 8576 5284
rect 8343 5253 8355 5256
rect 8297 5247 8355 5253
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 8938 5244 8944 5296
rect 8996 5244 9002 5296
rect 9600 5284 9628 5324
rect 9950 5312 9956 5364
rect 10008 5312 10014 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 10100 5324 10149 5352
rect 10100 5312 10106 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 10137 5315 10195 5321
rect 10980 5324 11376 5352
rect 10870 5284 10876 5296
rect 9600 5256 10876 5284
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 10980 5228 11008 5324
rect 11348 5284 11376 5324
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 11480 5324 11529 5352
rect 11480 5312 11486 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 12400 5324 12541 5352
rect 12400 5312 12406 5324
rect 12529 5321 12541 5324
rect 12575 5352 12587 5355
rect 13722 5352 13728 5364
rect 12575 5324 13728 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13814 5312 13820 5364
rect 13872 5312 13878 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14700 5324 14841 5352
rect 14700 5312 14706 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 15160 5324 15209 5352
rect 15160 5312 15166 5324
rect 15197 5321 15209 5324
rect 15243 5352 15255 5355
rect 16298 5352 16304 5364
rect 15243 5324 16304 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16448 5324 17908 5352
rect 16448 5312 16454 5324
rect 11348 5256 12388 5284
rect 12360 5228 12388 5256
rect 13170 5244 13176 5296
rect 13228 5244 13234 5296
rect 13832 5284 13860 5312
rect 17880 5284 17908 5324
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 19613 5355 19671 5361
rect 18012 5324 19564 5352
rect 18012 5312 18018 5324
rect 19058 5284 19064 5296
rect 13648 5256 13860 5284
rect 14384 5256 17724 5284
rect 17880 5256 19064 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1854 5216 1860 5228
rect 1719 5188 1860 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2222 5216 2228 5228
rect 2087 5188 2228 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2332 5080 2360 5179
rect 2590 5176 2596 5228
rect 2648 5176 2654 5228
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3786 5216 3792 5228
rect 2915 5188 3792 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4111 5188 4537 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4525 5185 4537 5188
rect 4571 5216 4583 5219
rect 4798 5216 4804 5228
rect 4571 5188 4804 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 6181 5219 6239 5225
rect 5368 5188 6132 5216
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3292 5120 3893 5148
rect 3292 5108 3298 5120
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4755 5120 5273 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 4356 5080 4384 5111
rect 5368 5080 5396 5188
rect 6104 5160 6132 5188
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6227 5188 6561 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5491 5120 5672 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5644 5089 5672 5120
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 5905 5151 5963 5157
rect 5905 5148 5917 5151
rect 5868 5120 5917 5148
rect 5868 5108 5874 5120
rect 5905 5117 5917 5120
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 6086 5108 6092 5160
rect 6144 5108 6150 5160
rect 6564 5148 6592 5179
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9646 5188 9873 5216
rect 7760 5148 7788 5176
rect 6564 5120 7788 5148
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9306 5148 9312 5160
rect 8720 5120 9312 5148
rect 8720 5108 8726 5120
rect 9306 5108 9312 5120
rect 9364 5148 9370 5160
rect 9646 5148 9674 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 10502 5176 10508 5228
rect 10560 5176 10566 5228
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10744 5188 10824 5216
rect 10744 5176 10750 5188
rect 9364 5120 9674 5148
rect 9364 5108 9370 5120
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10520 5148 10548 5176
rect 9824 5120 10548 5148
rect 9824 5108 9830 5120
rect 10594 5108 10600 5160
rect 10652 5108 10658 5160
rect 10796 5157 10824 5188
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11112 5188 11161 5216
rect 11112 5176 11118 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11480 5188 11897 5216
rect 11480 5176 11486 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12492 5188 12725 5216
rect 12492 5176 12498 5188
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 13188 5216 13216 5244
rect 13648 5228 13676 5256
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13188 5188 13277 5216
rect 12713 5179 12771 5185
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14384 5225 14412 5256
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 14056 5188 14381 5216
rect 14056 5176 14062 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 15838 5216 15844 5228
rect 14660 5188 15844 5216
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11379 5120 11989 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 14660 5148 14688 5188
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 16206 5176 16212 5228
rect 16264 5176 16270 5228
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 17218 5216 17224 5228
rect 16960 5188 17224 5216
rect 12176 5120 14688 5148
rect 14737 5151 14795 5157
rect 2332 5052 2728 5080
rect 4356 5052 5396 5080
rect 5629 5083 5687 5089
rect 2700 5024 2728 5052
rect 5629 5049 5641 5083
rect 5675 5049 5687 5083
rect 10686 5080 10692 5092
rect 5629 5043 5687 5049
rect 5828 5052 7236 5080
rect 1034 4972 1040 5024
rect 1092 5012 1098 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1092 4984 1869 5012
rect 1092 4972 1098 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 2222 4972 2228 5024
rect 2280 4972 2286 5024
rect 2498 4972 2504 5024
rect 2556 4972 2562 5024
rect 2682 4972 2688 5024
rect 2740 4972 2746 5024
rect 2774 4972 2780 5024
rect 2832 4972 2838 5024
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 5718 5012 5724 5024
rect 4295 4984 5724 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 5718 4972 5724 4984
rect 5776 5012 5782 5024
rect 5828 5012 5856 5052
rect 5776 4984 5856 5012
rect 5776 4972 5782 4984
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 6052 4984 6101 5012
rect 6052 4972 6058 4984
rect 6089 4981 6101 4984
rect 6135 5012 6147 5015
rect 6270 5012 6276 5024
rect 6135 4984 6276 5012
rect 6135 4981 6147 4984
rect 6089 4975 6147 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7208 5012 7236 5052
rect 9324 5052 10692 5080
rect 9324 5012 9352 5052
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 7208 4984 9352 5012
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 9769 4975 9827 4981
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 12176 5012 12204 5120
rect 13648 5089 13676 5120
rect 14737 5117 14749 5151
rect 14783 5148 14795 5151
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14783 5120 15301 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 15378 5108 15384 5160
rect 15436 5108 15442 5160
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16960 5148 16988 5188
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 15979 5120 16988 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 17126 5108 17132 5160
rect 17184 5148 17190 5160
rect 17328 5148 17356 5179
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17696 5225 17724 5256
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 19426 5244 19432 5296
rect 19484 5244 19490 5296
rect 19536 5284 19564 5324
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19886 5352 19892 5364
rect 19659 5324 19892 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20349 5355 20407 5361
rect 20349 5321 20361 5355
rect 20395 5352 20407 5355
rect 20806 5352 20812 5364
rect 20395 5324 20812 5352
rect 20395 5321 20407 5324
rect 20349 5315 20407 5321
rect 20806 5312 20812 5324
rect 20864 5352 20870 5364
rect 21450 5352 21456 5364
rect 20864 5324 21456 5352
rect 20864 5312 20870 5324
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 21836 5324 22416 5352
rect 19705 5287 19763 5293
rect 19705 5284 19717 5287
rect 19536 5256 19717 5284
rect 19705 5253 19717 5256
rect 19751 5253 19763 5287
rect 19705 5247 19763 5253
rect 19812 5256 21772 5284
rect 17681 5219 17739 5225
rect 17681 5185 17693 5219
rect 17727 5185 17739 5219
rect 17681 5179 17739 5185
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17828 5188 17969 5216
rect 17828 5176 17834 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18782 5216 18788 5228
rect 18196 5188 18788 5216
rect 18196 5176 18202 5188
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 18874 5176 18880 5228
rect 18932 5216 18938 5228
rect 19812 5216 19840 5256
rect 21744 5228 21772 5256
rect 18932 5188 19840 5216
rect 18932 5176 18938 5188
rect 19886 5176 19892 5228
rect 19944 5176 19950 5228
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5216 20039 5219
rect 20070 5216 20076 5228
rect 20027 5188 20076 5216
rect 20027 5185 20039 5188
rect 19981 5179 20039 5185
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20438 5216 20444 5228
rect 20303 5188 20444 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 17184 5120 17356 5148
rect 19061 5151 19119 5157
rect 17184 5108 17190 5120
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 19702 5148 19708 5160
rect 19107 5120 19708 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 19794 5108 19800 5160
rect 19852 5148 19858 5160
rect 20180 5148 20208 5179
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 20898 5216 20904 5228
rect 20855 5188 20904 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 20898 5176 20904 5188
rect 20956 5216 20962 5228
rect 21634 5216 21640 5228
rect 20956 5188 21640 5216
rect 20956 5176 20962 5188
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 21726 5176 21732 5228
rect 21784 5176 21790 5228
rect 19852 5120 20300 5148
rect 19852 5108 19858 5120
rect 20272 5092 20300 5120
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 21836 5148 21864 5324
rect 22388 5284 22416 5324
rect 22462 5312 22468 5364
rect 22520 5312 22526 5364
rect 27430 5312 27436 5364
rect 27488 5312 27494 5364
rect 23934 5284 23940 5296
rect 22388 5256 23940 5284
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22278 5216 22284 5228
rect 22235 5188 22284 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22385 5219 22443 5225
rect 22385 5185 22397 5219
rect 22431 5216 22443 5219
rect 22554 5216 22560 5228
rect 22431 5188 22560 5216
rect 22431 5185 22443 5188
rect 22385 5179 22443 5185
rect 22554 5176 22560 5188
rect 22612 5216 22618 5228
rect 23400 5225 23428 5256
rect 23934 5244 23940 5256
rect 23992 5244 23998 5296
rect 27065 5287 27123 5293
rect 27065 5284 27077 5287
rect 26804 5256 27077 5284
rect 22679 5219 22737 5225
rect 22679 5216 22691 5219
rect 22612 5188 22691 5216
rect 22612 5176 22618 5188
rect 22679 5185 22691 5188
rect 22725 5185 22737 5219
rect 22679 5179 22737 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23385 5219 23443 5225
rect 22879 5188 22968 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 20404 5120 21864 5148
rect 22296 5148 22324 5176
rect 22940 5148 22968 5188
rect 23117 5209 23175 5215
rect 23117 5175 23129 5209
rect 23163 5206 23175 5209
rect 23163 5178 23244 5206
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 23163 5175 23175 5178
rect 23117 5169 23175 5175
rect 22296 5120 22968 5148
rect 23216 5148 23244 5178
rect 23658 5176 23664 5228
rect 23716 5176 23722 5228
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5216 23903 5219
rect 24118 5216 24124 5228
rect 23891 5188 24124 5216
rect 23891 5185 23903 5188
rect 23845 5179 23903 5185
rect 24118 5176 24124 5188
rect 24176 5176 24182 5228
rect 26234 5176 26240 5228
rect 26292 5176 26298 5228
rect 26804 5225 26832 5256
rect 27065 5253 27077 5256
rect 27111 5253 27123 5287
rect 27065 5247 27123 5253
rect 26789 5219 26847 5225
rect 26789 5185 26801 5219
rect 26835 5185 26847 5219
rect 26789 5179 26847 5185
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5185 27031 5219
rect 26973 5179 27031 5185
rect 23216 5120 23428 5148
rect 20404 5108 20410 5120
rect 23400 5092 23428 5120
rect 13633 5083 13691 5089
rect 13633 5049 13645 5083
rect 13679 5049 13691 5083
rect 13633 5043 13691 5049
rect 14274 5040 14280 5092
rect 14332 5080 14338 5092
rect 15657 5083 15715 5089
rect 15657 5080 15669 5083
rect 14332 5052 15669 5080
rect 14332 5040 14338 5052
rect 15657 5049 15669 5052
rect 15703 5049 15715 5083
rect 15657 5043 15715 5049
rect 16945 5083 17003 5089
rect 16945 5049 16957 5083
rect 16991 5080 17003 5083
rect 17310 5080 17316 5092
rect 16991 5052 17316 5080
rect 16991 5049 17003 5052
rect 16945 5043 17003 5049
rect 17310 5040 17316 5052
rect 17368 5080 17374 5092
rect 19978 5080 19984 5092
rect 17368 5052 19984 5080
rect 17368 5040 17374 5052
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 20254 5040 20260 5092
rect 20312 5040 20318 5092
rect 20533 5083 20591 5089
rect 20533 5049 20545 5083
rect 20579 5080 20591 5083
rect 20714 5080 20720 5092
rect 20579 5052 20720 5080
rect 20579 5049 20591 5052
rect 20533 5043 20591 5049
rect 20714 5040 20720 5052
rect 20772 5080 20778 5092
rect 22830 5080 22836 5092
rect 20772 5052 22836 5080
rect 20772 5040 20778 5052
rect 22830 5040 22836 5052
rect 22888 5040 22894 5092
rect 23382 5040 23388 5092
rect 23440 5040 23446 5092
rect 23566 5040 23572 5092
rect 23624 5080 23630 5092
rect 23753 5083 23811 5089
rect 23753 5080 23765 5083
rect 23624 5052 23765 5080
rect 23624 5040 23630 5052
rect 23753 5049 23765 5052
rect 23799 5080 23811 5083
rect 26234 5080 26240 5092
rect 23799 5052 26240 5080
rect 23799 5049 23811 5052
rect 23753 5043 23811 5049
rect 26234 5040 26240 5052
rect 26292 5040 26298 5092
rect 26418 5040 26424 5092
rect 26476 5080 26482 5092
rect 26988 5080 27016 5179
rect 27246 5176 27252 5228
rect 27304 5176 27310 5228
rect 26476 5052 27016 5080
rect 26476 5040 26482 5052
rect 10192 4984 12204 5012
rect 10192 4972 10198 4984
rect 12894 4972 12900 5024
rect 12952 4972 12958 5024
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 14700 4984 15853 5012
rect 14700 4972 14706 4984
rect 15841 4981 15853 4984
rect 15887 5012 15899 5015
rect 17034 5012 17040 5024
rect 15887 4984 17040 5012
rect 15887 4981 15899 4984
rect 15841 4975 15899 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 19392 4984 19441 5012
rect 19392 4972 19398 4984
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 19429 4975 19487 4981
rect 20622 4972 20628 5024
rect 20680 5012 20686 5024
rect 22189 5015 22247 5021
rect 22189 5012 22201 5015
rect 20680 4984 22201 5012
rect 20680 4972 20686 4984
rect 22189 4981 22201 4984
rect 22235 5012 22247 5015
rect 22646 5012 22652 5024
rect 22235 4984 22652 5012
rect 22235 4981 22247 4984
rect 22189 4975 22247 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 22738 4972 22744 5024
rect 22796 5012 22802 5024
rect 23017 5015 23075 5021
rect 23017 5012 23029 5015
rect 22796 4984 23029 5012
rect 22796 4972 22802 4984
rect 23017 4981 23029 4984
rect 23063 4981 23075 5015
rect 23017 4975 23075 4981
rect 26326 4972 26332 5024
rect 26384 4972 26390 5024
rect 26602 4972 26608 5024
rect 26660 4972 26666 5024
rect 1104 4922 27876 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 27876 4922
rect 1104 4848 27876 4870
rect 2222 4768 2228 4820
rect 2280 4768 2286 4820
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 4614 4808 4620 4820
rect 2372 4780 4620 4808
rect 2372 4768 2378 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5684 4780 5825 4808
rect 5684 4768 5690 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 6052 4780 6101 4808
rect 6052 4768 6058 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 9490 4808 9496 4820
rect 7892 4780 9496 4808
rect 7892 4768 7898 4780
rect 9490 4768 9496 4780
rect 9548 4808 9554 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 9548 4780 9597 4808
rect 9548 4768 9554 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11790 4808 11796 4820
rect 11296 4780 11796 4808
rect 11296 4768 11302 4780
rect 11790 4768 11796 4780
rect 11848 4808 11854 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11848 4780 11989 4808
rect 11848 4768 11854 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 11977 4771 12035 4777
rect 12342 4768 12348 4820
rect 12400 4768 12406 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13722 4808 13728 4820
rect 13587 4780 13728 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13722 4768 13728 4780
rect 13780 4808 13786 4820
rect 13780 4780 14320 4808
rect 13780 4768 13786 4780
rect 950 4700 956 4752
rect 1008 4740 1014 4752
rect 1489 4743 1547 4749
rect 1489 4740 1501 4743
rect 1008 4712 1501 4740
rect 1008 4700 1014 4712
rect 1489 4709 1501 4712
rect 1535 4709 1547 4743
rect 1489 4703 1547 4709
rect 2240 4672 2268 4768
rect 5552 4740 5580 4768
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 5552 4712 5917 4740
rect 5905 4709 5917 4712
rect 5951 4709 5963 4743
rect 5905 4703 5963 4709
rect 6104 4712 7144 4740
rect 1688 4644 2268 4672
rect 1688 4613 1716 4644
rect 5258 4632 5264 4684
rect 5316 4632 5322 4684
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 2087 4576 2237 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 6104 4604 6132 4712
rect 7116 4672 7144 4712
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 9030 4740 9036 4752
rect 7432 4712 9036 4740
rect 7432 4700 7438 4712
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 14292 4740 14320 4780
rect 14642 4768 14648 4820
rect 14700 4768 14706 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 17586 4768 17592 4820
rect 17644 4808 17650 4820
rect 20714 4808 20720 4820
rect 17644 4780 20720 4808
rect 17644 4768 17650 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21269 4811 21327 4817
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 21542 4808 21548 4820
rect 21315 4780 21548 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 22336 4780 22784 4808
rect 22336 4768 22342 4780
rect 15378 4740 15384 4752
rect 14292 4712 15384 4740
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 18874 4740 18880 4752
rect 15764 4712 18880 4740
rect 10134 4672 10140 4684
rect 6748 4644 7052 4672
rect 7116 4644 10140 4672
rect 6748 4616 6776 4644
rect 2639 4576 6132 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4606 6515 4607
rect 6503 4604 6684 4606
rect 6730 4604 6736 4616
rect 6503 4578 6736 4604
rect 6503 4573 6515 4578
rect 6656 4576 6736 4578
rect 6457 4567 6515 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7024 4613 7052 4644
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10229 4675 10287 4681
rect 10229 4641 10241 4675
rect 10275 4672 10287 4675
rect 11698 4672 11704 4684
rect 10275 4644 11704 4672
rect 10275 4641 10287 4644
rect 10229 4635 10287 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 12434 4632 12440 4684
rect 12492 4632 12498 4684
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 13228 4644 13369 4672
rect 13228 4632 13234 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 13357 4635 13415 4641
rect 13630 4632 13636 4684
rect 13688 4632 13694 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15764 4672 15792 4712
rect 18874 4700 18880 4712
rect 18932 4700 18938 4752
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 19518 4740 19524 4752
rect 19475 4712 19524 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 19518 4700 19524 4712
rect 19576 4740 19582 4752
rect 19797 4743 19855 4749
rect 19797 4740 19809 4743
rect 19576 4712 19809 4740
rect 19576 4700 19582 4712
rect 19797 4709 19809 4712
rect 19843 4709 19855 4743
rect 19797 4703 19855 4709
rect 20346 4700 20352 4752
rect 20404 4740 20410 4752
rect 20404 4712 21864 4740
rect 20404 4700 20410 4712
rect 16758 4681 16764 4684
rect 15252 4644 15792 4672
rect 16735 4675 16764 4681
rect 15252 4632 15258 4644
rect 16735 4641 16747 4675
rect 16735 4635 16764 4641
rect 16758 4632 16764 4635
rect 16816 4632 16822 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 16945 4675 17003 4681
rect 16945 4672 16957 4675
rect 16908 4644 16957 4672
rect 16908 4632 16914 4644
rect 16945 4641 16957 4644
rect 16991 4641 17003 4675
rect 16945 4635 17003 4641
rect 18506 4632 18512 4684
rect 18564 4632 18570 4684
rect 19150 4632 19156 4684
rect 19208 4632 19214 4684
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 19300 4644 19656 4672
rect 19300 4632 19306 4644
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 6932 4536 6960 4567
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7282 4613 7288 4616
rect 7265 4607 7288 4613
rect 7265 4573 7277 4607
rect 7265 4567 7288 4573
rect 7282 4564 7288 4567
rect 7340 4564 7346 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4604 9183 4607
rect 9214 4604 9220 4616
rect 9171 4576 9220 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9456 4576 9505 4604
rect 9456 4564 9462 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12894 4604 12900 4616
rect 12575 4576 12900 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13648 4604 13676 4632
rect 13044 4576 13676 4604
rect 13044 4564 13050 4576
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13964 4576 14473 4604
rect 13964 4564 13970 4576
rect 14461 4573 14473 4576
rect 14507 4604 14519 4607
rect 14642 4604 14648 4616
rect 14507 4576 14648 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 16574 4604 16580 4616
rect 14783 4576 16580 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 18524 4604 18552 4632
rect 17635 4576 18552 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 6196 4508 6776 4536
rect 6932 4508 7236 4536
rect 1034 4428 1040 4480
rect 1092 4468 1098 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1092 4440 1869 4468
rect 1092 4428 1098 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 1857 4431 1915 4437
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2280 4440 2513 4468
rect 2280 4428 2286 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5316 4440 5365 4468
rect 5316 4428 5322 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 5442 4428 5448 4480
rect 5500 4428 5506 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 6196 4468 6224 4508
rect 6748 4477 6776 4508
rect 7208 4480 7236 4508
rect 10502 4496 10508 4548
rect 10560 4496 10566 4548
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 10836 4508 10994 4536
rect 12084 4508 14780 4536
rect 10836 4496 10842 4508
rect 5592 4440 6224 4468
rect 6733 4471 6791 4477
rect 5592 4428 5598 4440
rect 6733 4437 6745 4471
rect 6779 4437 6791 4471
rect 6733 4431 6791 4437
rect 7190 4428 7196 4480
rect 7248 4428 7254 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 12084 4468 12112 4508
rect 7340 4440 12112 4468
rect 7340 4428 7346 4440
rect 12158 4428 12164 4480
rect 12216 4428 12222 4480
rect 13170 4428 13176 4480
rect 13228 4428 13234 4480
rect 14182 4428 14188 4480
rect 14240 4428 14246 4480
rect 14752 4468 14780 4508
rect 15102 4496 15108 4548
rect 15160 4536 15166 4548
rect 17221 4539 17279 4545
rect 17221 4536 17233 4539
rect 15160 4508 17233 4536
rect 15160 4496 15166 4508
rect 17221 4505 17233 4508
rect 17267 4536 17279 4539
rect 18322 4536 18328 4548
rect 17267 4508 18328 4536
rect 17267 4505 17279 4508
rect 17221 4499 17279 4505
rect 18322 4496 18328 4508
rect 18380 4496 18386 4548
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 14752 4440 17509 4468
rect 17497 4437 17509 4440
rect 17543 4468 17555 4471
rect 17586 4468 17592 4480
rect 17543 4440 17592 4468
rect 17543 4437 17555 4440
rect 17497 4431 17555 4437
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 18230 4468 18236 4480
rect 17819 4440 18236 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18432 4468 18460 4576
rect 18506 4496 18512 4548
rect 18564 4536 18570 4548
rect 19168 4536 19196 4632
rect 19628 4613 19656 4644
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 21836 4681 21864 4712
rect 22554 4700 22560 4752
rect 22612 4700 22618 4752
rect 22756 4749 22784 4780
rect 27430 4768 27436 4820
rect 27488 4768 27494 4820
rect 22741 4743 22799 4749
rect 22741 4709 22753 4743
rect 22787 4740 22799 4743
rect 23106 4740 23112 4752
rect 22787 4712 23112 4740
rect 22787 4709 22799 4712
rect 22741 4703 22799 4709
rect 23106 4700 23112 4712
rect 23164 4740 23170 4752
rect 24026 4740 24032 4752
rect 23164 4712 24032 4740
rect 23164 4700 23170 4712
rect 24026 4700 24032 4712
rect 24084 4700 24090 4752
rect 21821 4675 21879 4681
rect 20128 4644 20575 4672
rect 20128 4632 20134 4644
rect 20547 4616 20575 4644
rect 20640 4644 21312 4672
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 19659 4576 20269 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20530 4604 20536 4616
rect 20491 4576 20536 4604
rect 20257 4567 20315 4573
rect 19245 4539 19303 4545
rect 19245 4536 19257 4539
rect 18564 4508 19257 4536
rect 18564 4496 18570 4508
rect 19245 4505 19257 4508
rect 19291 4505 19303 4539
rect 19536 4536 19564 4567
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 20640 4613 20668 4644
rect 21284 4616 21312 4644
rect 21821 4641 21833 4675
rect 21867 4641 21879 4675
rect 21821 4635 21879 4641
rect 21928 4644 26372 4672
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 20717 4607 20775 4613
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 20898 4604 20904 4616
rect 20763 4576 20904 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 20990 4564 20996 4616
rect 21048 4604 21054 4616
rect 21085 4607 21143 4613
rect 21085 4604 21097 4607
rect 21048 4576 21097 4604
rect 21048 4564 21054 4576
rect 21085 4573 21097 4576
rect 21131 4573 21143 4607
rect 21085 4567 21143 4573
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 20806 4536 20812 4548
rect 19536 4508 20812 4536
rect 19245 4499 19303 4505
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 21928 4536 21956 4644
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4604 22155 4607
rect 22738 4604 22744 4616
rect 22143 4576 22744 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 20916 4508 21956 4536
rect 22020 4536 22048 4567
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 26344 4613 26372 4644
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 26329 4607 26387 4613
rect 26329 4573 26341 4607
rect 26375 4573 26387 4607
rect 26329 4567 26387 4573
rect 22373 4539 22431 4545
rect 22020 4508 22324 4536
rect 19334 4468 19340 4480
rect 18432 4440 19340 4468
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19518 4428 19524 4480
rect 19576 4428 19582 4480
rect 20254 4428 20260 4480
rect 20312 4468 20318 4480
rect 20622 4468 20628 4480
rect 20312 4440 20628 4468
rect 20312 4428 20318 4440
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 20916 4477 20944 4508
rect 20901 4471 20959 4477
rect 20901 4468 20913 4471
rect 20772 4440 20913 4468
rect 20772 4428 20778 4440
rect 20901 4437 20913 4440
rect 20947 4437 20959 4471
rect 20901 4431 20959 4437
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22186 4468 22192 4480
rect 21867 4440 22192 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 22296 4477 22324 4508
rect 22373 4505 22385 4539
rect 22419 4536 22431 4539
rect 22462 4536 22468 4548
rect 22419 4508 22468 4536
rect 22419 4505 22431 4508
rect 22373 4499 22431 4505
rect 22462 4496 22468 4508
rect 22520 4496 22526 4548
rect 22646 4496 22652 4548
rect 22704 4536 22710 4548
rect 23032 4536 23060 4567
rect 26602 4564 26608 4616
rect 26660 4564 26666 4616
rect 26881 4607 26939 4613
rect 26881 4573 26893 4607
rect 26927 4573 26939 4607
rect 26881 4567 26939 4573
rect 22704 4508 23060 4536
rect 26421 4539 26479 4545
rect 22704 4496 22710 4508
rect 26421 4505 26433 4539
rect 26467 4536 26479 4539
rect 26896 4536 26924 4567
rect 27246 4564 27252 4616
rect 27304 4564 27310 4616
rect 26467 4508 26924 4536
rect 26467 4505 26479 4508
rect 26421 4499 26479 4505
rect 22281 4471 22339 4477
rect 22281 4437 22293 4471
rect 22327 4468 22339 4471
rect 23198 4468 23204 4480
rect 22327 4440 23204 4468
rect 22327 4437 22339 4440
rect 22281 4431 22339 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 26697 4471 26755 4477
rect 26697 4437 26709 4471
rect 26743 4468 26755 4471
rect 26786 4468 26792 4480
rect 26743 4440 26792 4468
rect 26743 4437 26755 4440
rect 26697 4431 26755 4437
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 27062 4428 27068 4480
rect 27120 4428 27126 4480
rect 1104 4378 27876 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 27876 4378
rect 1104 4304 27876 4326
rect 2774 4264 2780 4276
rect 2240 4236 2780 4264
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2240 4128 2268 4236
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 4341 4267 4399 4273
rect 4341 4233 4353 4267
rect 4387 4264 4399 4267
rect 4798 4264 4804 4276
rect 4387 4236 4804 4264
rect 4387 4233 4399 4236
rect 4341 4227 4399 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5442 4264 5448 4276
rect 5184 4236 5448 4264
rect 5184 4140 5212 4236
rect 5442 4224 5448 4236
rect 5500 4264 5506 4276
rect 5626 4264 5632 4276
rect 5500 4236 5632 4264
rect 5500 4224 5506 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 6730 4264 6736 4276
rect 5920 4236 6736 4264
rect 5920 4196 5948 4236
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7650 4264 7656 4276
rect 7064 4236 7656 4264
rect 7064 4224 7070 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 7760 4236 9873 4264
rect 5368 4168 5948 4196
rect 2087 4100 2268 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1688 4060 1716 4091
rect 2314 4088 2320 4140
rect 2372 4088 2378 4140
rect 2498 4088 2504 4140
rect 2556 4088 2562 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2516 4060 2544 4088
rect 1688 4032 2544 4060
rect 1486 3952 1492 4004
rect 1544 3952 1550 4004
rect 2130 3952 2136 4004
rect 2188 3992 2194 4004
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 2188 3964 2513 3992
rect 2188 3952 2194 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2608 3992 2636 4091
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 5368 4137 5396 4168
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 5920 4137 5948 4168
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 7760 4196 7788 4236
rect 9861 4233 9873 4236
rect 9907 4264 9919 4267
rect 10318 4264 10324 4276
rect 9907 4236 10324 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 11238 4264 11244 4276
rect 11011 4236 11244 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 11333 4267 11391 4273
rect 11333 4233 11345 4267
rect 11379 4264 11391 4267
rect 11974 4264 11980 4276
rect 11379 4236 11980 4264
rect 11379 4233 11391 4236
rect 11333 4227 11391 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12066 4224 12072 4276
rect 12124 4224 12130 4276
rect 15102 4264 15108 4276
rect 13096 4236 15108 4264
rect 6052 4168 7788 4196
rect 6052 4156 6058 4168
rect 9030 4156 9036 4208
rect 9088 4196 9094 4208
rect 9125 4199 9183 4205
rect 9125 4196 9137 4199
rect 9088 4168 9137 4196
rect 9088 4156 9094 4168
rect 9125 4165 9137 4168
rect 9171 4165 9183 4199
rect 13096 4196 13124 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 16574 4264 16580 4276
rect 15488 4236 16580 4264
rect 9125 4159 9183 4165
rect 9600 4168 13124 4196
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 4663 4032 5672 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 4448 3992 4476 4023
rect 4798 3992 4804 4004
rect 2608 3964 4384 3992
rect 4448 3964 4804 3992
rect 2501 3955 2559 3961
rect 1034 3884 1040 3936
rect 1092 3924 1098 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1092 3896 1869 3924
rect 1092 3884 1098 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2004 3896 2237 3924
rect 2004 3884 2010 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4356 3924 4384 3964
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 4890 3952 4896 4004
rect 4948 3952 4954 4004
rect 5644 4001 5672 4032
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6196 4060 6224 4091
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6328 4100 6561 4128
rect 6328 4088 6334 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7098 4128 7104 4140
rect 7055 4100 7104 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 6932 4060 6960 4091
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 7926 4128 7932 4140
rect 7883 4100 7932 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 7926 4088 7932 4100
rect 7984 4128 7990 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 7984 4100 8309 4128
rect 7984 4088 7990 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 8846 4128 8852 4140
rect 8803 4100 8852 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 7190 4060 7196 4072
rect 5868 4032 7196 4060
rect 5868 4020 5874 4032
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7742 4060 7748 4072
rect 7515 4032 7748 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7742 4020 7748 4032
rect 7800 4060 7806 4072
rect 8680 4060 8708 4091
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 8987 4100 9076 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9048 4060 9076 4100
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 7800 4032 9076 4060
rect 9232 4060 9260 4088
rect 9600 4060 9628 4168
rect 13722 4156 13728 4208
rect 13780 4156 13786 4208
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 14918 4205 14924 4208
rect 14895 4199 14924 4205
rect 14424 4168 14688 4196
rect 14424 4156 14430 4168
rect 9674 4088 9680 4140
rect 9732 4088 9738 4140
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 11054 4128 11060 4140
rect 10045 4091 10103 4097
rect 10152 4100 11060 4128
rect 9232 4032 9628 4060
rect 7800 4020 7806 4032
rect 5629 3995 5687 4001
rect 5629 3961 5641 3995
rect 5675 3961 5687 3995
rect 5629 3955 5687 3961
rect 5902 3952 5908 4004
rect 5960 3952 5966 4004
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 6822 3992 6828 4004
rect 6144 3964 6828 3992
rect 6144 3952 6150 3964
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 8662 3952 8668 4004
rect 8720 3952 8726 4004
rect 9048 3992 9076 4032
rect 10152 3992 10180 4100
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11422 4128 11428 4140
rect 11195 4100 11428 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 12986 4128 12992 4140
rect 11563 4100 12992 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 11532 4060 11560 4091
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 14660 4128 14688 4168
rect 14895 4165 14907 4199
rect 14895 4159 14924 4165
rect 14918 4156 14924 4159
rect 14976 4156 14982 4208
rect 15488 4137 15516 4236
rect 16574 4224 16580 4236
rect 16632 4264 16638 4276
rect 17218 4264 17224 4276
rect 16632 4236 17224 4264
rect 16632 4224 16638 4236
rect 17218 4224 17224 4236
rect 17276 4264 17282 4276
rect 17586 4264 17592 4276
rect 17276 4236 17592 4264
rect 17276 4224 17282 4236
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 17681 4267 17739 4273
rect 17681 4233 17693 4267
rect 17727 4264 17739 4267
rect 18138 4264 18144 4276
rect 17727 4236 18144 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 18138 4224 18144 4236
rect 18196 4224 18202 4276
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18932 4236 19073 4264
rect 18932 4224 18938 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 19242 4224 19248 4276
rect 19300 4224 19306 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19392 4236 19656 4264
rect 19392 4224 19398 4236
rect 16482 4196 16488 4208
rect 15672 4168 16488 4196
rect 15672 4137 15700 4168
rect 16482 4156 16488 4168
rect 16540 4196 16546 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 16540 4168 16865 4196
rect 16540 4156 16546 4168
rect 16853 4165 16865 4168
rect 16899 4165 16911 4199
rect 17313 4199 17371 4205
rect 17313 4196 17325 4199
rect 16853 4159 16911 4165
rect 16960 4168 17325 4196
rect 16960 4140 16988 4168
rect 17313 4165 17325 4168
rect 17359 4165 17371 4199
rect 17313 4159 17371 4165
rect 17420 4168 18276 4196
rect 15473 4131 15531 4137
rect 14660 4100 15424 4128
rect 10827 4032 11560 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 11072 4004 11100 4032
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12066 4060 12072 4072
rect 11848 4032 12072 4060
rect 11848 4020 11854 4032
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 13872 4032 14381 4060
rect 13872 4020 13878 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 14642 4020 14648 4072
rect 14700 4020 14706 4072
rect 14734 4020 14740 4072
rect 14792 4020 14798 4072
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14884 4032 15117 4060
rect 14884 4020 14890 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15396 4060 15424 4100
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 15930 4128 15936 4140
rect 15887 4100 15936 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 15672 4060 15700 4091
rect 15396 4032 15700 4060
rect 15105 4023 15163 4029
rect 9048 3964 10180 3992
rect 11054 3952 11060 4004
rect 11112 3952 11118 4004
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 15654 3992 15660 4004
rect 11480 3964 13032 3992
rect 11480 3952 11486 3964
rect 5810 3924 5816 3936
rect 4356 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 5920 3924 5948 3952
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5920 3896 6009 3924
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8846 3924 8852 3936
rect 8067 3896 8852 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 9490 3884 9496 3936
rect 9548 3884 9554 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 10410 3924 10416 3936
rect 10275 3896 10416 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10410 3884 10416 3896
rect 10468 3924 10474 3936
rect 10870 3924 10876 3936
rect 10468 3896 10876 3924
rect 10468 3884 10474 3896
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12710 3924 12716 3936
rect 11931 3896 12716 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12860 3896 12909 3924
rect 12860 3884 12866 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 13004 3924 13032 3964
rect 14568 3964 15660 3992
rect 14568 3924 14596 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15764 3992 15792 4091
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16206 4060 16212 4072
rect 15935 4032 16212 4060
rect 15935 3992 15963 4032
rect 16206 4020 16212 4032
rect 16264 4060 16270 4072
rect 16684 4060 16712 4091
rect 16942 4088 16948 4140
rect 17000 4088 17006 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17420 4128 17448 4168
rect 17083 4100 17448 4128
rect 17497 4131 17555 4137
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17678 4128 17684 4140
rect 17543 4100 17684 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17512 4060 17540 4091
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 17911 4100 18153 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18141 4097 18153 4100
rect 18187 4097 18199 4131
rect 18248 4128 18276 4168
rect 18969 4131 19027 4137
rect 18248 4100 18920 4128
rect 18141 4091 18199 4097
rect 16264 4032 17540 4060
rect 18049 4063 18107 4069
rect 16264 4020 16270 4032
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 15764 3964 15963 3992
rect 17034 3952 17040 4004
rect 17092 3992 17098 4004
rect 18064 3992 18092 4023
rect 18230 4020 18236 4072
rect 18288 4020 18294 4072
rect 18322 4020 18328 4072
rect 18380 4020 18386 4072
rect 18892 4060 18920 4100
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19260 4128 19288 4224
rect 19628 4196 19656 4236
rect 19702 4224 19708 4276
rect 19760 4224 19766 4276
rect 19886 4224 19892 4276
rect 19944 4264 19950 4276
rect 20254 4264 20260 4276
rect 19944 4236 20260 4264
rect 19944 4224 19950 4236
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 21266 4224 21272 4276
rect 21324 4224 21330 4276
rect 22370 4264 22376 4276
rect 22020 4236 22376 4264
rect 19904 4196 19932 4224
rect 19981 4199 20039 4205
rect 19981 4196 19993 4199
rect 19628 4168 19993 4196
rect 19015 4100 19288 4128
rect 19337 4131 19395 4137
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 19518 4128 19524 4140
rect 19383 4100 19524 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 19518 4088 19524 4100
rect 19576 4088 19582 4140
rect 19628 4137 19656 4168
rect 19981 4165 19993 4168
rect 20027 4165 20039 4199
rect 20438 4196 20444 4208
rect 19981 4159 20039 4165
rect 20088 4168 20444 4196
rect 20088 4140 20116 4168
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 21284 4196 21312 4224
rect 20824 4168 21312 4196
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4097 19671 4131
rect 19886 4128 19892 4140
rect 19613 4091 19671 4097
rect 19812 4100 19892 4128
rect 19812 4060 19840 4100
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20303 4100 20484 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 18892 4032 19840 4060
rect 20346 4020 20352 4072
rect 20404 4020 20410 4072
rect 17092 3964 18092 3992
rect 17092 3952 17098 3964
rect 13004 3896 14596 3924
rect 12897 3887 12955 3893
rect 15286 3884 15292 3936
rect 15344 3884 15350 3936
rect 16022 3884 16028 3936
rect 16080 3884 16086 3936
rect 17218 3884 17224 3936
rect 17276 3884 17282 3936
rect 18064 3924 18092 3964
rect 18509 3995 18567 4001
rect 18509 3961 18521 3995
rect 18555 3992 18567 3995
rect 20364 3992 20392 4020
rect 18555 3964 20392 3992
rect 20456 3992 20484 4100
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 20824 4137 20852 4168
rect 20625 4131 20683 4137
rect 20625 4128 20637 4131
rect 20588 4100 20637 4128
rect 20588 4088 20594 4100
rect 20625 4097 20637 4100
rect 20671 4097 20683 4131
rect 20625 4091 20683 4097
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 20640 4060 20668 4091
rect 20990 4088 20996 4140
rect 21048 4128 21054 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 21048 4100 21097 4128
rect 21048 4088 21054 4100
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 21358 4088 21364 4140
rect 21416 4088 21422 4140
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 21726 4128 21732 4140
rect 21600 4100 21732 4128
rect 21600 4088 21606 4100
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 22020 4137 22048 4236
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 22186 4156 22192 4208
rect 22244 4196 22250 4208
rect 22281 4199 22339 4205
rect 22281 4196 22293 4199
rect 22244 4168 22293 4196
rect 22244 4156 22250 4168
rect 22281 4165 22293 4168
rect 22327 4165 22339 4199
rect 22281 4159 22339 4165
rect 24026 4156 24032 4208
rect 24084 4156 24090 4208
rect 26344 4168 27292 4196
rect 26344 4140 26372 4168
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21928 4100 22017 4128
rect 21266 4060 21272 4072
rect 20640 4032 21272 4060
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 21928 4060 21956 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 23348 4114 23414 4128
rect 23348 4100 23428 4114
rect 23348 4088 23354 4100
rect 23014 4060 23020 4072
rect 21876 4032 21956 4060
rect 22112 4032 23020 4060
rect 21876 4020 21882 4032
rect 20898 3992 20904 4004
rect 20456 3964 20904 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 18785 3927 18843 3933
rect 18785 3924 18797 3927
rect 18064 3896 18797 3924
rect 18785 3893 18797 3896
rect 18831 3924 18843 3927
rect 19245 3927 19303 3933
rect 19245 3924 19257 3927
rect 18831 3896 19257 3924
rect 18831 3893 18843 3896
rect 18785 3887 18843 3893
rect 19245 3893 19257 3896
rect 19291 3893 19303 3927
rect 19245 3887 19303 3893
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 20456 3924 20484 3964
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 21450 3952 21456 4004
rect 21508 3992 21514 4004
rect 22112 3992 22140 4032
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23400 4060 23428 4100
rect 25958 4088 25964 4140
rect 26016 4088 26022 4140
rect 26234 4088 26240 4140
rect 26292 4088 26298 4140
rect 26326 4088 26332 4140
rect 26384 4088 26390 4140
rect 26513 4131 26571 4137
rect 26513 4097 26525 4131
rect 26559 4097 26571 4131
rect 26513 4091 26571 4097
rect 26053 4063 26111 4069
rect 23400 4032 23888 4060
rect 23860 4004 23888 4032
rect 26053 4029 26065 4063
rect 26099 4060 26111 4063
rect 26528 4060 26556 4091
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 27264 4137 27292 4168
rect 27249 4131 27307 4137
rect 27249 4097 27261 4131
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 26099 4032 26556 4060
rect 26099 4029 26111 4032
rect 26053 4023 26111 4029
rect 21508 3964 22140 3992
rect 21508 3952 21514 3964
rect 23842 3952 23848 4004
rect 23900 3952 23906 4004
rect 26329 3995 26387 4001
rect 26329 3961 26341 3995
rect 26375 3992 26387 3995
rect 26878 3992 26884 4004
rect 26375 3964 26884 3992
rect 26375 3961 26387 3964
rect 26329 3955 26387 3961
rect 26878 3952 26884 3964
rect 26936 3952 26942 4004
rect 27430 3952 27436 4004
rect 27488 3952 27494 4004
rect 19576 3896 20484 3924
rect 20916 3924 20944 3952
rect 21358 3924 21364 3936
rect 20916 3896 21364 3924
rect 19576 3884 19582 3896
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 26694 3884 26700 3936
rect 26752 3884 26758 3936
rect 27062 3884 27068 3936
rect 27120 3884 27126 3936
rect 1104 3834 27876 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 27876 3834
rect 1104 3760 27876 3782
rect 2774 3720 2780 3732
rect 2746 3680 2780 3720
rect 2832 3680 2838 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 4856 3692 6285 3720
rect 4856 3680 4862 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6273 3683 6331 3689
rect 6454 3680 6460 3732
rect 6512 3680 6518 3732
rect 7006 3729 7012 3732
rect 6996 3723 7012 3729
rect 6996 3689 7008 3723
rect 6996 3683 7012 3689
rect 7006 3680 7012 3683
rect 7064 3680 7070 3732
rect 9140 3692 11560 3720
rect 950 3612 956 3664
rect 1008 3652 1014 3664
rect 1489 3655 1547 3661
rect 1489 3652 1501 3655
rect 1008 3624 1501 3652
rect 1008 3612 1014 3624
rect 1489 3621 1501 3624
rect 1535 3621 1547 3655
rect 1489 3615 1547 3621
rect 2746 3584 2774 3680
rect 5534 3652 5540 3664
rect 5460 3624 5540 3652
rect 1688 3556 2774 3584
rect 1688 3525 1716 3556
rect 4154 3544 4160 3596
rect 4212 3544 4218 3596
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 5460 3584 5488 3624
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 6472 3652 6500 3680
rect 6472 3624 6776 3652
rect 4479 3556 5488 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 6748 3593 6776 3624
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 5684 3556 6653 3584
rect 5684 3544 5690 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 7558 3584 7564 3596
rect 6779 3556 7564 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 9140 3593 9168 3692
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3584 9459 3587
rect 9490 3584 9496 3596
rect 9447 3556 9496 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 11146 3544 11152 3596
rect 11204 3544 11210 3596
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1854 3476 1860 3528
rect 1912 3476 1918 3528
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2222 3516 2228 3528
rect 2087 3488 2228 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5718 3516 5724 3528
rect 5592 3488 5724 3516
rect 5592 3476 5598 3488
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6178 3476 6184 3528
rect 6236 3476 6242 3528
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3516 6515 3519
rect 6546 3516 6552 3528
rect 6503 3488 6552 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 10778 3516 10784 3528
rect 10534 3488 10784 3516
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 11532 3525 11560 3692
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13780 3692 13829 3720
rect 13780 3680 13786 3692
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14700 3692 15025 3720
rect 14700 3680 14706 3692
rect 15013 3689 15025 3692
rect 15059 3720 15071 3723
rect 15194 3720 15200 3732
rect 15059 3692 15200 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15920 3723 15978 3729
rect 15920 3689 15932 3723
rect 15966 3720 15978 3723
rect 16022 3720 16028 3732
rect 15966 3692 16028 3720
rect 15966 3689 15978 3692
rect 15920 3683 15978 3689
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 16540 3692 17877 3720
rect 16540 3680 16546 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 19518 3720 19524 3732
rect 17865 3683 17923 3689
rect 19352 3692 19524 3720
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 14608 3624 15700 3652
rect 14608 3612 14614 3624
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 12860 3556 14473 3584
rect 12860 3544 12866 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3485 11575 3519
rect 13630 3516 13636 3528
rect 11517 3479 11575 3485
rect 13188 3488 13636 3516
rect 1872 3448 1900 3476
rect 5736 3448 5764 3476
rect 8757 3451 8815 3457
rect 1872 3420 2774 3448
rect 5736 3420 7498 3448
rect 1034 3340 1040 3392
rect 1092 3380 1098 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1092 3352 1869 3380
rect 1092 3340 1098 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 2746 3380 2774 3420
rect 8757 3417 8769 3451
rect 8803 3417 8815 3451
rect 11422 3448 11428 3460
rect 8757 3411 8815 3417
rect 10704 3420 11428 3448
rect 5718 3380 5724 3392
rect 2746 3352 5724 3380
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7190 3380 7196 3392
rect 6880 3352 7196 3380
rect 6880 3340 6886 3352
rect 7190 3340 7196 3352
rect 7248 3380 7254 3392
rect 7374 3380 7380 3392
rect 7248 3352 7380 3380
rect 7248 3340 7254 3352
rect 7374 3340 7380 3352
rect 7432 3380 7438 3392
rect 8772 3380 8800 3411
rect 10704 3380 10732 3420
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 11532 3448 11560 3479
rect 11698 3448 11704 3460
rect 11532 3420 11704 3448
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11790 3408 11796 3460
rect 11848 3408 11854 3460
rect 11900 3420 12282 3448
rect 7432 3352 10732 3380
rect 7432 3340 7438 3352
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11900 3380 11928 3420
rect 10836 3352 11928 3380
rect 12176 3380 12204 3420
rect 13188 3380 13216 3488
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14148 3488 14289 3516
rect 14148 3476 14154 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14476 3516 14504 3547
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15672 3593 15700 3624
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 19352 3652 19380 3692
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 22554 3720 22560 3732
rect 19944 3692 22560 3720
rect 19944 3680 19950 3692
rect 17092 3624 19380 3652
rect 17092 3612 17098 3624
rect 15657 3587 15715 3593
rect 14792 3556 15240 3584
rect 14792 3544 14798 3556
rect 15212 3528 15240 3556
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 16666 3584 16672 3596
rect 15703 3556 16672 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17586 3584 17592 3596
rect 17000 3556 17592 3584
rect 17000 3544 17006 3556
rect 17586 3544 17592 3556
rect 17644 3584 17650 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 17644 3556 17693 3584
rect 17644 3544 17650 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 18874 3584 18880 3596
rect 18555 3556 18880 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 20070 3584 20076 3596
rect 19168 3556 20076 3584
rect 14826 3516 14832 3528
rect 14476 3488 14832 3516
rect 14277 3479 14335 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15194 3476 15200 3528
rect 15252 3476 15258 3528
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 15562 3476 15568 3528
rect 15620 3476 15626 3528
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3516 18107 3519
rect 19168 3516 19196 3556
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 20312 3556 21404 3584
rect 20312 3544 20318 3556
rect 21376 3525 21404 3556
rect 18095 3488 19196 3516
rect 19245 3519 19303 3525
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 21361 3519 21419 3525
rect 21361 3485 21373 3519
rect 21407 3516 21419 3519
rect 21450 3516 21456 3528
rect 21407 3488 21456 3516
rect 21407 3485 21419 3488
rect 21361 3479 21419 3485
rect 13262 3408 13268 3460
rect 13320 3448 13326 3460
rect 13538 3448 13544 3460
rect 13320 3420 13544 3448
rect 13320 3408 13326 3420
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 13725 3451 13783 3457
rect 13725 3417 13737 3451
rect 13771 3417 13783 3451
rect 13725 3411 13783 3417
rect 12176 3352 13216 3380
rect 10836 3340 10842 3352
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 13740 3380 13768 3411
rect 13504 3352 13768 3380
rect 13504 3340 13510 3352
rect 14090 3340 14096 3392
rect 14148 3340 14154 3392
rect 15304 3380 15332 3476
rect 15580 3448 15608 3476
rect 15580 3420 16422 3448
rect 18506 3408 18512 3460
rect 18564 3408 18570 3460
rect 18690 3408 18696 3460
rect 18748 3448 18754 3460
rect 18966 3448 18972 3460
rect 18748 3420 18972 3448
rect 18748 3408 18754 3420
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 19260 3448 19288 3479
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21652 3525 21680 3692
rect 22554 3680 22560 3692
rect 22612 3720 22618 3732
rect 22612 3692 24532 3720
rect 22612 3680 22618 3692
rect 21821 3587 21879 3593
rect 21821 3553 21833 3587
rect 21867 3584 21879 3587
rect 22189 3587 22247 3593
rect 22189 3584 22201 3587
rect 21867 3556 22201 3584
rect 21867 3553 21879 3556
rect 21821 3547 21879 3553
rect 22189 3553 22201 3556
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 21913 3519 21971 3525
rect 21913 3485 21925 3519
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 19426 3448 19432 3460
rect 19260 3420 19432 3448
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 19521 3451 19579 3457
rect 19521 3417 19533 3451
rect 19567 3417 19579 3451
rect 19521 3411 19579 3417
rect 16666 3380 16672 3392
rect 15304 3352 16672 3380
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 16850 3340 16856 3392
rect 16908 3380 16914 3392
rect 18524 3380 18552 3408
rect 16908 3352 18552 3380
rect 16908 3340 16914 3352
rect 18598 3340 18604 3392
rect 18656 3340 18662 3392
rect 19061 3383 19119 3389
rect 19061 3349 19073 3383
rect 19107 3380 19119 3383
rect 19536 3380 19564 3411
rect 19794 3408 19800 3460
rect 19852 3448 19858 3460
rect 19978 3448 19984 3460
rect 19852 3420 19984 3448
rect 19852 3408 19858 3420
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 21818 3448 21824 3460
rect 20916 3420 21824 3448
rect 19107 3352 19564 3380
rect 19107 3349 19119 3352
rect 19061 3343 19119 3349
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 20916 3380 20944 3420
rect 21818 3408 21824 3420
rect 21876 3448 21882 3460
rect 21928 3448 21956 3479
rect 23658 3476 23664 3528
rect 23716 3516 23722 3528
rect 24504 3525 24532 3692
rect 27062 3680 27068 3732
rect 27120 3680 27126 3732
rect 27430 3680 27436 3732
rect 27488 3680 27494 3732
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23716 3488 23949 3516
rect 23716 3476 23722 3488
rect 23937 3485 23949 3488
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 24489 3519 24547 3525
rect 24489 3485 24501 3519
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 24854 3476 24860 3528
rect 24912 3516 24918 3528
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 24912 3488 26065 3516
rect 24912 3476 24918 3488
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26053 3479 26111 3485
rect 26326 3476 26332 3528
rect 26384 3476 26390 3528
rect 26602 3476 26608 3528
rect 26660 3476 26666 3528
rect 26786 3476 26792 3528
rect 26844 3476 26850 3528
rect 26881 3519 26939 3525
rect 26881 3485 26893 3519
rect 26927 3516 26939 3519
rect 27080 3516 27108 3680
rect 26927 3488 27108 3516
rect 27249 3519 27307 3525
rect 26927 3485 26939 3488
rect 26881 3479 26939 3485
rect 27249 3485 27261 3519
rect 27295 3485 27307 3519
rect 27249 3479 27307 3485
rect 21876 3420 21956 3448
rect 21876 3408 21882 3420
rect 22646 3408 22652 3460
rect 22704 3408 22710 3460
rect 19668 3352 20944 3380
rect 19668 3340 19674 3352
rect 20990 3340 20996 3392
rect 21048 3340 21054 3392
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 21453 3383 21511 3389
rect 21453 3380 21465 3383
rect 21324 3352 21465 3380
rect 21324 3340 21330 3352
rect 21453 3349 21465 3352
rect 21499 3380 21511 3383
rect 21910 3380 21916 3392
rect 21499 3352 21916 3380
rect 21499 3349 21511 3352
rect 21453 3343 21511 3349
rect 21910 3340 21916 3352
rect 21968 3340 21974 3392
rect 22370 3340 22376 3392
rect 22428 3380 22434 3392
rect 23676 3380 23704 3476
rect 26804 3448 26832 3476
rect 27264 3448 27292 3479
rect 26804 3420 27292 3448
rect 22428 3352 23704 3380
rect 22428 3340 22434 3352
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 24581 3383 24639 3389
rect 24581 3380 24593 3383
rect 23808 3352 24593 3380
rect 23808 3340 23814 3352
rect 24581 3349 24593 3352
rect 24627 3349 24639 3383
rect 24581 3343 24639 3349
rect 26142 3340 26148 3392
rect 26200 3340 26206 3392
rect 26418 3340 26424 3392
rect 26476 3340 26482 3392
rect 26694 3340 26700 3392
rect 26752 3340 26758 3392
rect 27062 3340 27068 3392
rect 27120 3340 27126 3392
rect 1104 3290 27876 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 27876 3290
rect 1104 3216 27876 3238
rect 950 3136 956 3188
rect 1008 3176 1014 3188
rect 1489 3179 1547 3185
rect 1489 3176 1501 3179
rect 1008 3148 1501 3176
rect 1008 3136 1014 3148
rect 1489 3145 1501 3148
rect 1535 3145 1547 3179
rect 1489 3139 1547 3145
rect 1946 3136 1952 3188
rect 2004 3136 2010 3188
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2700 3148 5212 3176
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1964 3040 1992 3136
rect 1719 3012 1992 3040
rect 2041 3043 2099 3049
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2148 3040 2176 3136
rect 2087 3012 2176 3040
rect 2240 3040 2268 3136
rect 2700 3049 2728 3148
rect 4154 3108 4160 3120
rect 3620 3080 4160 3108
rect 3620 3049 3648 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 5184 3108 5212 3148
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 5813 3179 5871 3185
rect 5813 3176 5825 3179
rect 5776 3148 5825 3176
rect 5776 3136 5782 3148
rect 5813 3145 5825 3148
rect 5859 3145 5871 3179
rect 5813 3139 5871 3145
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 7469 3179 7527 3185
rect 5960 3148 6592 3176
rect 5960 3136 5966 3148
rect 6086 3108 6092 3120
rect 5184 3080 6092 3108
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2240 3012 2421 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 2976 2904 3004 3003
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 5534 3040 5540 3052
rect 5014 3012 5540 3040
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 6270 3040 6276 3052
rect 6012 3012 6276 3040
rect 4908 2972 4936 3000
rect 3712 2944 4936 2972
rect 5629 2975 5687 2981
rect 3712 2904 3740 2944
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 5902 2972 5908 2984
rect 5675 2944 5908 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6012 2981 6040 3012
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6564 3049 6592 3148
rect 7469 3145 7481 3179
rect 7515 3145 7527 3179
rect 7469 3139 7527 3145
rect 7484 3108 7512 3139
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 7984 3148 9904 3176
rect 7984 3136 7990 3148
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7116 3080 7420 3108
rect 7484 3080 7849 3108
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6822 3040 6828 3052
rect 6595 3012 6828 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7116 3049 7144 3080
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6932 2972 6960 3003
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 7392 3040 7420 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 9306 3068 9312 3120
rect 9364 3108 9370 3120
rect 9364 3080 9812 3108
rect 9364 3068 9370 3080
rect 7466 3040 7472 3052
rect 7392 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9272 3012 9689 3040
rect 9272 3000 9278 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 7300 2972 7328 3000
rect 6788 2944 6960 2972
rect 7208 2944 7328 2972
rect 6788 2932 6794 2944
rect 7208 2916 7236 2944
rect 9582 2932 9588 2984
rect 9640 2932 9646 2984
rect 9784 2972 9812 3080
rect 9876 3049 9904 3148
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 10560 3148 10793 3176
rect 10560 3136 10566 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 13265 3179 13323 3185
rect 10781 3139 10839 3145
rect 10888 3148 12388 3176
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10888 3040 10916 3148
rect 11514 3108 11520 3120
rect 10980 3080 11520 3108
rect 10980 3049 11008 3080
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 11882 3068 11888 3120
rect 11940 3068 11946 3120
rect 9907 3012 10916 3040
rect 10965 3043 11023 3049
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 10980 2972 11008 3003
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11164 2972 11192 3003
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 11296 3012 11345 3040
rect 11296 3000 11302 3012
rect 11333 3009 11345 3012
rect 11379 3009 11391 3043
rect 11532 3040 11560 3068
rect 11793 3043 11851 3049
rect 11532 3038 11652 3040
rect 11793 3038 11805 3043
rect 11532 3012 11805 3038
rect 11624 3010 11805 3012
rect 11333 3003 11391 3009
rect 11793 3009 11805 3010
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 11977 3043 12035 3049
rect 12161 3046 12219 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12084 3043 12219 3046
rect 12084 3018 12173 3043
rect 11992 2972 12020 3003
rect 9784 2944 11008 2972
rect 11072 2944 12020 2972
rect 12084 2972 12112 3018
rect 12161 3009 12173 3018
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 12360 3040 12388 3148
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 13354 3176 13360 3188
rect 13311 3148 13360 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 13814 3176 13820 3188
rect 13495 3148 13820 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 13909 3179 13967 3185
rect 13909 3145 13921 3179
rect 13955 3176 13967 3179
rect 14090 3176 14096 3188
rect 13955 3148 14096 3176
rect 13955 3145 13967 3148
rect 13909 3139 13967 3145
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14274 3136 14280 3188
rect 14332 3136 14338 3188
rect 14550 3136 14556 3188
rect 14608 3136 14614 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15620 3148 17356 3176
rect 15620 3136 15626 3148
rect 12449 3043 12507 3049
rect 12449 3040 12461 3043
rect 12360 3012 12461 3040
rect 12449 3009 12461 3012
rect 12495 3040 12507 3043
rect 13173 3043 13231 3049
rect 12495 3012 13124 3040
rect 12495 3009 12507 3012
rect 12449 3003 12507 3009
rect 12084 2944 12204 2972
rect 2976 2876 3740 2904
rect 6196 2876 7144 2904
rect 1034 2796 1040 2848
rect 1092 2836 1098 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 1092 2808 1869 2836
rect 1092 2796 1098 2808
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 1857 2799 1915 2805
rect 2222 2796 2228 2848
rect 2280 2796 2286 2848
rect 2590 2796 2596 2848
rect 2648 2796 2654 2848
rect 2866 2796 2872 2848
rect 2924 2796 2930 2848
rect 3868 2839 3926 2845
rect 3868 2805 3880 2839
rect 3914 2836 3926 2839
rect 3970 2836 3976 2848
rect 3914 2808 3976 2836
rect 3914 2805 3926 2808
rect 3868 2799 3926 2805
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5258 2836 5264 2848
rect 4948 2808 5264 2836
rect 4948 2796 4954 2808
rect 5258 2796 5264 2808
rect 5316 2836 5322 2848
rect 6196 2845 6224 2876
rect 7116 2848 7144 2876
rect 7190 2864 7196 2916
rect 7248 2864 7254 2916
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 11072 2904 11100 2944
rect 9088 2876 11100 2904
rect 11609 2907 11667 2913
rect 9088 2864 9094 2876
rect 11609 2873 11621 2907
rect 11655 2904 11667 2907
rect 11698 2904 11704 2916
rect 11655 2876 11704 2904
rect 11655 2873 11667 2876
rect 11609 2867 11667 2873
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 5316 2808 5365 2836
rect 5316 2796 5322 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2805 6239 2839
rect 6181 2799 6239 2805
rect 6362 2796 6368 2848
rect 6420 2796 6426 2848
rect 7098 2796 7104 2848
rect 7156 2796 7162 2848
rect 9858 2796 9864 2848
rect 9916 2796 9922 2848
rect 11992 2836 12020 2944
rect 12176 2904 12204 2944
rect 12342 2932 12348 2984
rect 12400 2932 12406 2984
rect 12986 2932 12992 2984
rect 13044 2932 13050 2984
rect 13096 2972 13124 3012
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13262 3040 13268 3052
rect 13219 3012 13268 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3040 13415 3043
rect 13817 3043 13875 3049
rect 13403 3012 13768 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 13372 2972 13400 3003
rect 13096 2944 13400 2972
rect 13004 2904 13032 2932
rect 12176 2876 13032 2904
rect 13170 2836 13176 2848
rect 11992 2808 13176 2836
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13740 2836 13768 3012
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 14292 3040 14320 3136
rect 14568 3108 14596 3136
rect 14476 3080 14596 3108
rect 14476 3049 14504 3080
rect 13863 3012 14320 3040
rect 14461 3043 14519 3049
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 15856 3026 15884 3148
rect 16850 3108 16856 3120
rect 16684 3080 16856 3108
rect 16684 3049 16712 3080
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 16945 3111 17003 3117
rect 16945 3077 16957 3111
rect 16991 3108 17003 3111
rect 17218 3108 17224 3120
rect 16991 3080 17224 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 17328 3108 17356 3148
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 17736 3148 18276 3176
rect 17736 3136 17742 3148
rect 18248 3108 18276 3148
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 18656 3148 18889 3176
rect 18656 3136 18662 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 19702 3136 19708 3188
rect 19760 3176 19766 3188
rect 22646 3176 22652 3188
rect 19760 3148 19932 3176
rect 19760 3136 19766 3148
rect 18693 3111 18751 3117
rect 18693 3108 18705 3111
rect 17328 3080 17434 3108
rect 18248 3080 18705 3108
rect 18693 3077 18705 3080
rect 18739 3108 18751 3111
rect 18739 3080 19380 3108
rect 18739 3077 18751 3080
rect 18693 3071 18751 3077
rect 16669 3043 16727 3049
rect 14461 3003 14519 3009
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 19058 3000 19064 3052
rect 19116 3000 19122 3052
rect 19150 3000 19156 3052
rect 19208 3000 19214 3052
rect 19352 3049 19380 3080
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19904 3117 19932 3148
rect 20272 3148 22652 3176
rect 19889 3111 19947 3117
rect 19484 3080 19656 3108
rect 19484 3068 19490 3080
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19518 3000 19524 3052
rect 19576 3000 19582 3052
rect 19628 3049 19656 3080
rect 19889 3077 19901 3111
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 19978 3068 19984 3120
rect 20036 3108 20042 3120
rect 20272 3108 20300 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23106 3136 23112 3188
rect 23164 3136 23170 3188
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 23256 3148 23305 3176
rect 23256 3136 23262 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 25593 3179 25651 3185
rect 25593 3176 25605 3179
rect 23293 3139 23351 3145
rect 23400 3148 25605 3176
rect 20036 3080 20378 3108
rect 20036 3068 20042 3080
rect 21358 3068 21364 3120
rect 21416 3108 21422 3120
rect 21637 3111 21695 3117
rect 21637 3108 21649 3111
rect 21416 3080 21649 3108
rect 21416 3068 21422 3080
rect 21637 3077 21649 3080
rect 21683 3077 21695 3111
rect 21637 3071 21695 3077
rect 21910 3068 21916 3120
rect 21968 3108 21974 3120
rect 23124 3108 23152 3136
rect 23400 3108 23428 3148
rect 25593 3145 25605 3148
rect 25639 3145 25651 3179
rect 25593 3139 25651 3145
rect 26418 3136 26424 3188
rect 26476 3136 26482 3188
rect 26694 3136 26700 3188
rect 26752 3136 26758 3188
rect 26878 3136 26884 3188
rect 26936 3136 26942 3188
rect 27430 3136 27436 3188
rect 27488 3136 27494 3188
rect 21968 3080 23152 3108
rect 23216 3080 23428 3108
rect 23937 3111 23995 3117
rect 21968 3068 21974 3080
rect 22848 3049 22876 3080
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14182 2972 14188 2984
rect 14139 2944 14188 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14734 2932 14740 2984
rect 14792 2932 14798 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 15252 2944 16497 2972
rect 15252 2932 15258 2944
rect 16485 2941 16497 2944
rect 16531 2972 16543 2975
rect 18138 2972 18144 2984
rect 16531 2944 18144 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 21450 2932 21456 2984
rect 21508 2972 21514 2984
rect 22370 2972 22376 2984
rect 21508 2944 22376 2972
rect 21508 2932 21514 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2972 22615 2975
rect 22922 2972 22928 2984
rect 22603 2944 22928 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 23216 2981 23244 3080
rect 23937 3077 23949 3111
rect 23983 3108 23995 3111
rect 25406 3108 25412 3120
rect 23983 3080 25412 3108
rect 23983 3077 23995 3080
rect 23937 3071 23995 3077
rect 25406 3068 25412 3080
rect 25464 3068 25470 3120
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 23661 3043 23719 3049
rect 23661 3040 23673 3043
rect 23348 3012 23673 3040
rect 23348 3000 23354 3012
rect 23661 3009 23673 3012
rect 23707 3009 23719 3043
rect 23661 3003 23719 3009
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23900 3012 24225 3040
rect 23900 3000 23906 3012
rect 24213 3009 24225 3012
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 24486 3000 24492 3052
rect 24544 3000 24550 3052
rect 25498 3000 25504 3052
rect 25556 3000 25562 3052
rect 26436 3049 26464 3136
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3040 26571 3043
rect 26712 3040 26740 3136
rect 26896 3108 26924 3136
rect 26896 3080 27292 3108
rect 26559 3012 26740 3040
rect 26559 3009 26571 3012
rect 26513 3003 26571 3009
rect 23201 2975 23259 2981
rect 23201 2941 23213 2975
rect 23247 2941 23259 2975
rect 23750 2972 23756 2984
rect 23201 2935 23259 2941
rect 23308 2944 23756 2972
rect 19306 2876 19748 2904
rect 15378 2836 15384 2848
rect 13740 2808 15384 2836
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 15930 2836 15936 2848
rect 15528 2808 15936 2836
rect 15528 2796 15534 2808
rect 15930 2796 15936 2808
rect 15988 2836 15994 2848
rect 19306 2836 19334 2876
rect 15988 2808 19334 2836
rect 15988 2796 15994 2808
rect 19518 2796 19524 2848
rect 19576 2796 19582 2848
rect 19720 2836 19748 2876
rect 22462 2864 22468 2916
rect 22520 2864 22526 2916
rect 23308 2836 23336 2944
rect 23750 2932 23756 2944
rect 23808 2932 23814 2984
rect 23934 2932 23940 2984
rect 23992 2972 23998 2984
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23992 2944 24041 2972
rect 23992 2932 23998 2944
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2972 24455 2975
rect 26068 2972 26096 3003
rect 26970 3000 26976 3052
rect 27028 3000 27034 3052
rect 27264 3049 27292 3080
rect 27249 3043 27307 3049
rect 27249 3009 27261 3043
rect 27295 3009 27307 3043
rect 27249 3003 27307 3009
rect 27065 2975 27123 2981
rect 27065 2972 27077 2975
rect 24443 2944 26004 2972
rect 26068 2944 27077 2972
rect 24443 2941 24455 2944
rect 24397 2935 24455 2941
rect 25976 2904 26004 2944
rect 27065 2941 27077 2944
rect 27111 2941 27123 2975
rect 27065 2935 27123 2941
rect 26602 2904 26608 2916
rect 25976 2876 26608 2904
rect 26602 2864 26608 2876
rect 26660 2864 26666 2916
rect 19720 2808 23336 2836
rect 24578 2796 24584 2848
rect 24636 2796 24642 2848
rect 25866 2796 25872 2848
rect 25924 2796 25930 2848
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26237 2839 26295 2845
rect 26237 2836 26249 2839
rect 26108 2808 26249 2836
rect 26108 2796 26114 2808
rect 26237 2805 26249 2808
rect 26283 2805 26295 2839
rect 26237 2799 26295 2805
rect 26694 2796 26700 2848
rect 26752 2796 26758 2848
rect 1104 2746 27876 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 27876 2746
rect 1104 2672 27876 2694
rect 3234 2592 3240 2644
rect 3292 2592 3298 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5442 2632 5448 2644
rect 4939 2604 5448 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5442 2592 5448 2604
rect 5500 2632 5506 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5500 2604 5641 2632
rect 5500 2592 5506 2604
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 6730 2632 6736 2644
rect 5629 2595 5687 2601
rect 5736 2604 6736 2632
rect 1210 2524 1216 2576
rect 1268 2564 1274 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 1268 2536 2421 2564
rect 1268 2524 1274 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2533 2835 2567
rect 5736 2564 5764 2604
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7006 2632 7012 2644
rect 6963 2604 7012 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 7156 2604 8493 2632
rect 7156 2592 7162 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8904 2604 9045 2632
rect 8904 2592 8910 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 10870 2592 10876 2644
rect 10928 2592 10934 2644
rect 12894 2592 12900 2644
rect 12952 2592 12958 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 14366 2632 14372 2644
rect 13228 2604 14372 2632
rect 13228 2592 13234 2604
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14792 2604 14841 2632
rect 14792 2592 14798 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15470 2632 15476 2644
rect 14976 2604 15476 2632
rect 14976 2592 14982 2604
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 15620 2604 15853 2632
rect 15620 2592 15626 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 16666 2592 16672 2644
rect 16724 2592 16730 2644
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 17184 2604 18245 2632
rect 17184 2592 17190 2604
rect 18233 2601 18245 2604
rect 18279 2601 18291 2635
rect 18233 2595 18291 2601
rect 18782 2592 18788 2644
rect 18840 2632 18846 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 18840 2604 20085 2632
rect 18840 2592 18846 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 21910 2592 21916 2644
rect 21968 2592 21974 2644
rect 22664 2604 23796 2632
rect 7929 2567 7987 2573
rect 2777 2527 2835 2533
rect 5368 2536 5764 2564
rect 6288 2536 7861 2564
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 2792 2496 2820 2527
rect 1360 2468 2820 2496
rect 1360 2456 1366 2468
rect 4890 2456 4896 2508
rect 4948 2456 4954 2508
rect 2222 2388 2228 2440
rect 2280 2388 2286 2440
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 1036 2320 1042 2372
rect 1094 2360 1100 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 1094 2332 1409 2360
rect 1094 2320 1100 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1762 2320 1768 2372
rect 1820 2320 1826 2372
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 3068 2360 3096 2391
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 5368 2437 5396 2536
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5500 2468 5856 2496
rect 5500 2456 5506 2468
rect 5828 2437 5856 2468
rect 6288 2440 6316 2536
rect 7208 2468 7696 2496
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3476 2400 3801 2428
rect 3476 2388 3482 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5307 2400 5365 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 2556 2332 3096 2360
rect 4632 2360 4660 2391
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 4632 2332 5457 2360
rect 2556 2320 2562 2332
rect 5445 2329 5457 2332
rect 5491 2329 5503 2363
rect 5552 2360 5580 2391
rect 6270 2388 6276 2440
rect 6328 2388 6334 2440
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7208 2437 7236 2468
rect 7668 2440 7696 2468
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 7650 2388 7656 2440
rect 7708 2428 7714 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7708 2400 7757 2428
rect 7708 2388 7714 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7833 2428 7861 2536
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 7975 2536 8156 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 7926 2428 7932 2440
rect 7833 2400 7932 2428
rect 7745 2391 7803 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8128 2437 8156 2536
rect 11882 2524 11888 2576
rect 11940 2564 11946 2576
rect 15102 2564 15108 2576
rect 11940 2536 15108 2564
rect 11940 2524 11946 2536
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8260 2468 14228 2496
rect 8260 2456 8266 2468
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 6288 2360 6316 2388
rect 5552 2332 6316 2360
rect 7285 2363 7343 2369
rect 5445 2323 5503 2329
rect 7285 2329 7297 2363
rect 7331 2360 7343 2363
rect 7576 2360 7604 2388
rect 8680 2360 8708 2391
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8996 2400 9229 2428
rect 8996 2388 9002 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 10836 2400 11069 2428
rect 10836 2388 10842 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12342 2428 12348 2440
rect 12115 2400 12348 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12710 2388 12716 2440
rect 12768 2388 12774 2440
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13320 2400 13645 2428
rect 13320 2388 13326 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 7331 2332 7604 2360
rect 7944 2332 8708 2360
rect 7331 2329 7343 2332
rect 7285 2323 7343 2329
rect 1578 2252 1584 2304
rect 1636 2292 1642 2304
rect 2041 2295 2099 2301
rect 2041 2292 2053 2295
rect 1636 2264 2053 2292
rect 1636 2252 1642 2264
rect 2041 2261 2053 2264
rect 2087 2261 2099 2295
rect 2041 2255 2099 2261
rect 3970 2252 3976 2304
rect 4028 2252 4034 2304
rect 4430 2252 4436 2304
rect 4488 2252 4494 2304
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 5077 2295 5135 2301
rect 5077 2292 5089 2295
rect 4672 2264 5089 2292
rect 4672 2252 4678 2264
rect 5077 2261 5089 2264
rect 5123 2261 5135 2295
rect 5077 2255 5135 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6236 2264 6561 2292
rect 6236 2252 6242 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7944 2292 7972 2332
rect 14200 2304 14228 2468
rect 14292 2437 14320 2536
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 16942 2564 16948 2576
rect 15344 2536 16948 2564
rect 15344 2524 15350 2536
rect 16942 2524 16948 2536
rect 17000 2564 17006 2576
rect 21358 2564 21364 2576
rect 17000 2536 17080 2564
rect 17000 2524 17006 2536
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 14608 2468 16068 2496
rect 14608 2456 14614 2468
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14424 2400 14473 2428
rect 14424 2388 14430 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 14918 2428 14924 2440
rect 14691 2400 14924 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15378 2428 15384 2440
rect 15335 2400 15384 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 16040 2437 16068 2468
rect 15479 2431 15537 2437
rect 15479 2397 15491 2431
rect 15525 2397 15537 2431
rect 15479 2391 15537 2397
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 14553 2363 14611 2369
rect 14553 2329 14565 2363
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 15488 2360 15516 2391
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 17052 2437 17080 2536
rect 20732 2536 21364 2564
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2496 17187 2499
rect 17175 2468 17356 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17328 2437 17356 2468
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 15243 2332 15516 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 7156 2264 7972 2292
rect 7156 2252 7162 2264
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8076 2264 8309 2292
rect 8076 2252 8082 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 10137 2295 10195 2301
rect 10137 2292 10149 2295
rect 9916 2264 10149 2292
rect 9916 2252 9922 2264
rect 10137 2261 10149 2264
rect 10183 2261 10195 2295
rect 10137 2255 10195 2261
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 13596 2264 13829 2292
rect 13596 2252 13602 2264
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 13817 2255 13875 2261
rect 14178 2252 14184 2304
rect 14236 2252 14242 2304
rect 14568 2292 14596 2323
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 17236 2360 17264 2391
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18196 2400 18429 2428
rect 18196 2388 18202 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20732 2437 20760 2536
rect 21358 2524 21364 2536
rect 21416 2524 21422 2576
rect 22664 2564 22692 2604
rect 21468 2536 22692 2564
rect 20809 2499 20867 2505
rect 20809 2465 20821 2499
rect 20855 2496 20867 2499
rect 20855 2468 21036 2496
rect 20855 2465 20867 2468
rect 20809 2459 20867 2465
rect 21008 2437 21036 2468
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 19794 2360 19800 2372
rect 15620 2332 19800 2360
rect 15620 2320 15626 2332
rect 19794 2320 19800 2332
rect 19852 2360 19858 2372
rect 20916 2360 20944 2391
rect 21468 2360 21496 2536
rect 22664 2496 22692 2536
rect 22738 2524 22744 2576
rect 22796 2564 22802 2576
rect 23661 2567 23719 2573
rect 23661 2564 23673 2567
rect 22796 2536 23673 2564
rect 22796 2524 22802 2536
rect 23661 2533 23673 2536
rect 23707 2533 23719 2567
rect 23768 2564 23796 2604
rect 24026 2592 24032 2644
rect 24084 2592 24090 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 24486 2564 24492 2576
rect 23768 2536 24492 2564
rect 23661 2527 23719 2533
rect 24486 2524 24492 2536
rect 24544 2524 24550 2576
rect 22664 2468 22876 2496
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21876 2400 22109 2428
rect 21876 2388 21882 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 22848 2437 22876 2468
rect 23014 2456 23020 2508
rect 23072 2456 23078 2508
rect 23385 2499 23443 2505
rect 23385 2465 23397 2499
rect 23431 2496 23443 2499
rect 23431 2468 26556 2496
rect 23431 2465 23443 2468
rect 23385 2459 23443 2465
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22428 2400 22661 2428
rect 22428 2388 22434 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22922 2388 22928 2440
rect 22980 2428 22986 2440
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 22980 2400 23213 2428
rect 22980 2388 22986 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 19852 2332 21496 2360
rect 22741 2363 22799 2369
rect 19852 2320 19858 2332
rect 22741 2329 22753 2363
rect 22787 2360 22799 2363
rect 23492 2360 23520 2391
rect 23842 2388 23848 2440
rect 23900 2388 23906 2440
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 25317 2431 25375 2437
rect 25317 2397 25329 2431
rect 25363 2397 25375 2431
rect 25317 2391 25375 2397
rect 22787 2332 23520 2360
rect 25332 2360 25360 2391
rect 25590 2388 25596 2440
rect 25648 2388 25654 2440
rect 26142 2388 26148 2440
rect 26200 2388 26206 2440
rect 26528 2437 26556 2468
rect 26513 2431 26571 2437
rect 26513 2397 26525 2431
rect 26559 2397 26571 2431
rect 26513 2391 26571 2397
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26660 2400 27169 2428
rect 26660 2388 26666 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 26418 2360 26424 2372
rect 25332 2332 26424 2360
rect 22787 2329 22799 2332
rect 22741 2323 22799 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 27525 2363 27583 2369
rect 27525 2329 27537 2363
rect 27571 2360 27583 2363
rect 27821 2360 27827 2372
rect 27571 2332 27827 2360
rect 27571 2329 27583 2332
rect 27525 2323 27583 2329
rect 27821 2320 27827 2332
rect 27879 2320 27885 2372
rect 15286 2292 15292 2304
rect 14568 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15436 2264 15669 2292
rect 15436 2252 15442 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17497 2295 17555 2301
rect 17497 2292 17509 2295
rect 17276 2264 17509 2292
rect 17276 2252 17282 2264
rect 17497 2261 17509 2264
rect 17543 2261 17555 2295
rect 17497 2255 17555 2261
rect 19058 2252 19064 2304
rect 19116 2292 19122 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 19116 2264 19349 2292
rect 19116 2252 19122 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 20898 2252 20904 2304
rect 20956 2292 20962 2304
rect 21177 2295 21235 2301
rect 21177 2292 21189 2295
rect 20956 2264 21189 2292
rect 20956 2252 20962 2264
rect 21177 2261 21189 2264
rect 21223 2261 21235 2295
rect 21177 2255 21235 2261
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 22922 2292 22928 2304
rect 21692 2264 22928 2292
rect 21692 2252 21698 2264
rect 22922 2252 22928 2264
rect 22980 2292 22986 2304
rect 23934 2292 23940 2304
rect 22980 2264 23940 2292
rect 22980 2252 22986 2264
rect 23934 2252 23940 2264
rect 23992 2252 23998 2304
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 24857 2295 24915 2301
rect 24857 2292 24869 2295
rect 24636 2264 24869 2292
rect 24636 2252 24642 2264
rect 24857 2261 24869 2264
rect 24903 2261 24915 2295
rect 24857 2255 24915 2261
rect 25498 2252 25504 2304
rect 25556 2292 25562 2304
rect 25777 2295 25835 2301
rect 25777 2292 25789 2295
rect 25556 2264 25789 2292
rect 25556 2252 25562 2264
rect 25777 2261 25789 2264
rect 25823 2261 25835 2295
rect 25777 2255 25835 2261
rect 26326 2252 26332 2304
rect 26384 2252 26390 2304
rect 26697 2295 26755 2301
rect 26697 2261 26709 2295
rect 26743 2292 26755 2295
rect 27062 2292 27068 2304
rect 26743 2264 27068 2292
rect 26743 2261 26755 2264
rect 26697 2255 26755 2261
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 1104 2202 27876 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 27876 2202
rect 1104 2128 27876 2150
rect 2682 2048 2688 2100
rect 2740 2088 2746 2100
rect 2740 2060 12434 2088
rect 2740 2048 2746 2060
rect 2314 1912 2320 1964
rect 2372 1952 2378 1964
rect 8386 1952 8392 1964
rect 2372 1924 8392 1952
rect 2372 1912 2378 1924
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 12406 1952 12434 2060
rect 14178 2048 14184 2100
rect 14236 2088 14242 2100
rect 27194 2088 27200 2100
rect 14236 2060 27200 2088
rect 14236 2048 14242 2060
rect 27194 2048 27200 2060
rect 27252 2048 27258 2100
rect 17386 1980 17392 2032
rect 17444 2020 17450 2032
rect 24854 2020 24860 2032
rect 17444 1992 24860 2020
rect 17444 1980 17450 1992
rect 24854 1980 24860 1992
rect 24912 1980 24918 2032
rect 23406 1952 23412 1964
rect 12406 1924 23412 1952
rect 23406 1912 23412 1924
rect 23464 1912 23470 1964
rect 4798 1844 4804 1896
rect 4856 1884 4862 1896
rect 27286 1884 27292 1896
rect 4856 1856 27292 1884
rect 4856 1844 4862 1856
rect 27286 1844 27292 1856
rect 27344 1844 27350 1896
rect 3786 1776 3792 1828
rect 3844 1816 3850 1828
rect 17034 1816 17040 1828
rect 3844 1788 17040 1816
rect 3844 1776 3850 1788
rect 17034 1776 17040 1788
rect 17092 1776 17098 1828
rect 17386 1776 17392 1828
rect 17444 1776 17450 1828
rect 5626 1708 5632 1760
rect 5684 1748 5690 1760
rect 17404 1748 17432 1776
rect 5684 1720 17432 1748
rect 5684 1708 5690 1720
<< via1 >>
rect 10324 7964 10376 8016
rect 24308 7964 24360 8016
rect 1676 7896 1728 7948
rect 17316 7896 17368 7948
rect 8760 7828 8812 7880
rect 26884 7828 26936 7880
rect 2228 7692 2280 7744
rect 23848 7760 23900 7812
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1032 7488 1084 7540
rect 6000 7488 6052 7540
rect 6552 7488 6604 7540
rect 8300 7488 8352 7540
rect 10048 7488 10100 7540
rect 11796 7488 11848 7540
rect 1308 7420 1360 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 1124 7284 1176 7336
rect 3148 7463 3200 7472
rect 3148 7429 3157 7463
rect 3157 7429 3191 7463
rect 3191 7429 3200 7463
rect 3148 7420 3200 7429
rect 4712 7420 4764 7472
rect 13544 7420 13596 7472
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 14280 7352 14332 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 6920 7284 6972 7336
rect 15108 7284 15160 7336
rect 15292 7488 15344 7540
rect 17040 7488 17092 7540
rect 18788 7488 18840 7540
rect 22744 7488 22796 7540
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 8300 7216 8352 7268
rect 14372 7216 14424 7268
rect 20076 7284 20128 7336
rect 20536 7420 20588 7472
rect 22284 7420 22336 7472
rect 26700 7531 26752 7540
rect 26700 7497 26709 7531
rect 26709 7497 26743 7531
rect 26743 7497 26752 7531
rect 26700 7488 26752 7497
rect 27436 7531 27488 7540
rect 27436 7497 27445 7531
rect 27445 7497 27479 7531
rect 27479 7497 27488 7531
rect 27436 7488 27488 7497
rect 27528 7488 27580 7540
rect 24032 7420 24084 7472
rect 25780 7420 25832 7472
rect 26424 7395 26476 7404
rect 26424 7361 26433 7395
rect 26433 7361 26467 7395
rect 26467 7361 26476 7395
rect 26424 7352 26476 7361
rect 23020 7284 23072 7336
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 5816 7148 5868 7200
rect 14648 7191 14700 7200
rect 14648 7157 14657 7191
rect 14657 7157 14691 7191
rect 14691 7157 14700 7191
rect 14648 7148 14700 7157
rect 15384 7148 15436 7200
rect 16396 7148 16448 7200
rect 18696 7148 18748 7200
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 19892 7191 19944 7200
rect 19892 7157 19901 7191
rect 19901 7157 19935 7191
rect 19935 7157 19944 7191
rect 19892 7148 19944 7157
rect 19984 7148 20036 7200
rect 21640 7216 21692 7268
rect 20352 7148 20404 7200
rect 20444 7191 20496 7200
rect 20444 7157 20453 7191
rect 20453 7157 20487 7191
rect 20487 7157 20496 7191
rect 20444 7148 20496 7157
rect 20904 7148 20956 7200
rect 20996 7148 21048 7200
rect 24492 7191 24544 7200
rect 24492 7157 24501 7191
rect 24501 7157 24535 7191
rect 24535 7157 24544 7191
rect 24492 7148 24544 7157
rect 26332 7216 26384 7268
rect 26976 7191 27028 7200
rect 26976 7157 26985 7191
rect 26985 7157 27019 7191
rect 27019 7157 27028 7191
rect 26976 7148 27028 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1860 6987 1912 6996
rect 1860 6953 1869 6987
rect 1869 6953 1903 6987
rect 1903 6953 1912 6987
rect 1860 6944 1912 6953
rect 3516 6944 3568 6996
rect 4160 6944 4212 6996
rect 5448 6944 5500 6996
rect 6736 6944 6788 6996
rect 9036 6944 9088 6996
rect 10232 6944 10284 6996
rect 11520 6944 11572 6996
rect 14464 6944 14516 6996
rect 5816 6919 5868 6928
rect 5816 6885 5825 6919
rect 5825 6885 5859 6919
rect 5859 6885 5868 6919
rect 5816 6876 5868 6885
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 4712 6808 4764 6860
rect 5540 6808 5592 6860
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 8300 6808 8352 6860
rect 8668 6808 8720 6860
rect 9956 6808 10008 6860
rect 10508 6808 10560 6860
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6184 6740 6236 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 1124 6604 1176 6656
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 5356 6604 5408 6656
rect 6276 6672 6328 6724
rect 9864 6740 9916 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10232 6740 10284 6792
rect 11060 6876 11112 6928
rect 18144 6944 18196 6996
rect 18696 6987 18748 6996
rect 18696 6953 18705 6987
rect 18705 6953 18739 6987
rect 18739 6953 18748 6987
rect 18696 6944 18748 6953
rect 20628 6944 20680 6996
rect 21456 6944 21508 6996
rect 24492 6944 24544 6996
rect 26976 6944 27028 6996
rect 27436 6987 27488 6996
rect 27436 6953 27445 6987
rect 27445 6953 27479 6987
rect 27479 6953 27488 6987
rect 27436 6944 27488 6953
rect 10692 6808 10744 6860
rect 10968 6740 11020 6792
rect 14096 6808 14148 6860
rect 14280 6808 14332 6860
rect 15016 6808 15068 6860
rect 15568 6808 15620 6860
rect 16120 6808 16172 6860
rect 19892 6876 19944 6928
rect 20076 6876 20128 6928
rect 13176 6740 13228 6792
rect 14372 6740 14424 6792
rect 5724 6604 5776 6656
rect 6368 6604 6420 6656
rect 8576 6604 8628 6656
rect 10876 6672 10928 6724
rect 11152 6672 11204 6724
rect 9772 6604 9824 6656
rect 10140 6604 10192 6656
rect 11428 6604 11480 6656
rect 12072 6647 12124 6656
rect 12072 6613 12081 6647
rect 12081 6613 12115 6647
rect 12115 6613 12124 6647
rect 12072 6604 12124 6613
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 12992 6715 13044 6724
rect 12992 6681 13001 6715
rect 13001 6681 13035 6715
rect 13035 6681 13044 6715
rect 12992 6672 13044 6681
rect 13452 6672 13504 6724
rect 13728 6672 13780 6724
rect 15568 6672 15620 6724
rect 15660 6715 15712 6724
rect 15660 6681 15669 6715
rect 15669 6681 15703 6715
rect 15703 6681 15712 6715
rect 15660 6672 15712 6681
rect 15752 6672 15804 6724
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 16396 6715 16448 6724
rect 16396 6681 16405 6715
rect 16405 6681 16439 6715
rect 16439 6681 16448 6715
rect 16396 6672 16448 6681
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 19064 6740 19116 6792
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 19248 6672 19300 6724
rect 16488 6604 16540 6656
rect 17316 6604 17368 6656
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19800 6740 19852 6792
rect 20076 6740 20128 6792
rect 20536 6740 20588 6792
rect 20996 6808 21048 6860
rect 21088 6808 21140 6860
rect 21640 6808 21692 6860
rect 23296 6808 23348 6860
rect 22468 6740 22520 6792
rect 21180 6715 21232 6724
rect 21180 6681 21189 6715
rect 21189 6681 21223 6715
rect 21223 6681 21232 6715
rect 21180 6672 21232 6681
rect 22192 6715 22244 6724
rect 22192 6681 22201 6715
rect 22201 6681 22235 6715
rect 22235 6681 22244 6715
rect 22192 6672 22244 6681
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 23204 6783 23256 6792
rect 23204 6749 23213 6783
rect 23213 6749 23247 6783
rect 23247 6749 23256 6783
rect 23204 6740 23256 6749
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 26792 6740 26844 6792
rect 26976 6740 27028 6792
rect 20812 6604 20864 6656
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 22376 6647 22428 6656
rect 22376 6613 22385 6647
rect 22385 6613 22419 6647
rect 22419 6613 22428 6647
rect 22376 6604 22428 6613
rect 22652 6604 22704 6656
rect 22836 6604 22888 6656
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 27068 6647 27120 6656
rect 27068 6613 27077 6647
rect 27077 6613 27111 6647
rect 27111 6613 27120 6647
rect 27068 6604 27120 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 956 6400 1008 6452
rect 4528 6400 4580 6452
rect 4712 6400 4764 6452
rect 6552 6400 6604 6452
rect 6920 6443 6972 6452
rect 6920 6409 6929 6443
rect 6929 6409 6963 6443
rect 6963 6409 6972 6443
rect 6920 6400 6972 6409
rect 5356 6332 5408 6384
rect 6736 6332 6788 6384
rect 9404 6400 9456 6452
rect 1952 6264 2004 6316
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 3884 6196 3936 6248
rect 1040 6128 1092 6180
rect 5448 6264 5500 6316
rect 6092 6264 6144 6316
rect 7748 6332 7800 6384
rect 9128 6332 9180 6384
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6644 6196 6696 6248
rect 8944 6264 8996 6316
rect 9220 6264 9272 6316
rect 9864 6307 9916 6316
rect 9864 6273 9865 6307
rect 9865 6273 9899 6307
rect 9899 6273 9916 6307
rect 9864 6264 9916 6273
rect 10232 6264 10284 6316
rect 10416 6307 10468 6316
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 10600 6264 10652 6316
rect 10876 6400 10928 6452
rect 12440 6400 12492 6452
rect 12716 6400 12768 6452
rect 11428 6332 11480 6384
rect 5448 6128 5500 6180
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 9312 6128 9364 6180
rect 9772 6196 9824 6248
rect 10140 6128 10192 6180
rect 2044 6060 2096 6112
rect 7012 6060 7064 6112
rect 7564 6060 7616 6112
rect 8024 6060 8076 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 11244 6264 11296 6316
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 11520 6128 11572 6180
rect 11888 6060 11940 6112
rect 11980 6060 12032 6112
rect 13176 6400 13228 6452
rect 14648 6400 14700 6452
rect 16120 6443 16172 6452
rect 16120 6409 16129 6443
rect 16129 6409 16163 6443
rect 16163 6409 16172 6443
rect 16120 6400 16172 6409
rect 16028 6332 16080 6384
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20536 6400 20588 6452
rect 20812 6332 20864 6384
rect 13544 6264 13596 6316
rect 14004 6264 14056 6316
rect 14280 6196 14332 6248
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15016 6196 15068 6248
rect 16948 6264 17000 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 14372 6060 14424 6112
rect 14464 6060 14516 6112
rect 15384 6060 15436 6112
rect 16212 6060 16264 6112
rect 17040 6196 17092 6248
rect 19432 6264 19484 6316
rect 19984 6264 20036 6316
rect 20628 6264 20680 6316
rect 21456 6400 21508 6452
rect 21640 6400 21692 6452
rect 22376 6400 22428 6452
rect 22744 6332 22796 6384
rect 23296 6375 23348 6384
rect 23296 6341 23305 6375
rect 23305 6341 23339 6375
rect 23339 6341 23348 6375
rect 23296 6332 23348 6341
rect 23848 6443 23900 6452
rect 23848 6409 23857 6443
rect 23857 6409 23891 6443
rect 23891 6409 23900 6443
rect 23848 6400 23900 6409
rect 27436 6443 27488 6452
rect 27436 6409 27445 6443
rect 27445 6409 27479 6443
rect 27479 6409 27488 6443
rect 27436 6400 27488 6409
rect 26424 6332 26476 6384
rect 17224 6128 17276 6180
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 19064 6196 19116 6248
rect 19708 6239 19760 6248
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 24308 6264 24360 6316
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18420 6060 18472 6112
rect 19524 6128 19576 6180
rect 20260 6128 20312 6180
rect 21732 6196 21784 6248
rect 19340 6103 19392 6112
rect 19340 6069 19349 6103
rect 19349 6069 19383 6103
rect 19383 6069 19392 6103
rect 19340 6060 19392 6069
rect 20352 6060 20404 6112
rect 20444 6060 20496 6112
rect 21272 6128 21324 6180
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 23940 6196 23992 6248
rect 20996 6060 21048 6112
rect 21456 6103 21508 6112
rect 21456 6069 21465 6103
rect 21465 6069 21499 6103
rect 21499 6069 21508 6103
rect 21456 6060 21508 6069
rect 22560 6060 22612 6112
rect 22744 6060 22796 6112
rect 23296 6060 23348 6112
rect 24124 6103 24176 6112
rect 24124 6069 24133 6103
rect 24133 6069 24167 6103
rect 24167 6069 24176 6103
rect 24124 6060 24176 6069
rect 26700 6103 26752 6112
rect 26700 6069 26709 6103
rect 26709 6069 26743 6103
rect 26743 6069 26752 6103
rect 26700 6060 26752 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 6092 5856 6144 5908
rect 6184 5856 6236 5908
rect 6552 5856 6604 5908
rect 956 5788 1008 5840
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 6460 5720 6512 5772
rect 7564 5856 7616 5908
rect 7840 5856 7892 5908
rect 8484 5856 8536 5908
rect 8852 5788 8904 5840
rect 7932 5720 7984 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 7104 5652 7156 5704
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8668 5652 8720 5704
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 10692 5856 10744 5908
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 12072 5856 12124 5908
rect 13820 5856 13872 5908
rect 9496 5720 9548 5729
rect 10968 5720 11020 5772
rect 11704 5763 11756 5772
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 15660 5856 15712 5908
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 5448 5584 5500 5636
rect 5908 5584 5960 5636
rect 6000 5627 6052 5636
rect 6000 5593 6009 5627
rect 6009 5593 6043 5627
rect 6043 5593 6052 5627
rect 6000 5584 6052 5593
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 4804 5516 4856 5568
rect 6184 5516 6236 5568
rect 6828 5516 6880 5568
rect 8208 5627 8260 5636
rect 8208 5593 8217 5627
rect 8217 5593 8251 5627
rect 8251 5593 8260 5627
rect 8208 5584 8260 5593
rect 11888 5652 11940 5704
rect 13912 5720 13964 5772
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 15568 5720 15620 5772
rect 9036 5584 9088 5636
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 10784 5584 10836 5636
rect 11428 5627 11480 5636
rect 11428 5593 11437 5627
rect 11437 5593 11471 5627
rect 11471 5593 11480 5627
rect 11428 5584 11480 5593
rect 14004 5652 14056 5704
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 15660 5652 15712 5704
rect 17776 5720 17828 5772
rect 18604 5856 18656 5908
rect 18880 5856 18932 5908
rect 18972 5856 19024 5908
rect 20076 5856 20128 5908
rect 20628 5856 20680 5908
rect 17960 5720 18012 5772
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 19156 5788 19208 5840
rect 19984 5788 20036 5840
rect 20720 5788 20772 5840
rect 18328 5652 18380 5704
rect 20352 5720 20404 5772
rect 19984 5652 20036 5704
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 21088 5856 21140 5908
rect 21180 5856 21232 5908
rect 21456 5899 21508 5908
rect 21456 5865 21465 5899
rect 21465 5865 21499 5899
rect 21499 5865 21508 5899
rect 21456 5856 21508 5865
rect 23388 5856 23440 5908
rect 27436 5899 27488 5908
rect 27436 5865 27445 5899
rect 27445 5865 27479 5899
rect 27479 5865 27488 5899
rect 27436 5856 27488 5865
rect 21548 5720 21600 5772
rect 22836 5720 22888 5772
rect 14464 5584 14516 5636
rect 11612 5516 11664 5568
rect 13544 5516 13596 5568
rect 14372 5516 14424 5568
rect 15108 5516 15160 5568
rect 15200 5516 15252 5568
rect 16856 5584 16908 5636
rect 18972 5584 19024 5636
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 16488 5516 16540 5568
rect 20260 5516 20312 5568
rect 20996 5652 21048 5704
rect 23296 5652 23348 5704
rect 26884 5695 26936 5704
rect 26884 5661 26893 5695
rect 26893 5661 26927 5695
rect 26927 5661 26936 5695
rect 26884 5652 26936 5661
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 21456 5627 21508 5636
rect 21456 5593 21465 5627
rect 21465 5593 21499 5627
rect 21499 5593 21508 5627
rect 21456 5584 21508 5593
rect 20720 5516 20772 5568
rect 23204 5516 23256 5568
rect 27068 5559 27120 5568
rect 27068 5525 27077 5559
rect 27077 5525 27111 5559
rect 27111 5525 27120 5559
rect 27068 5516 27120 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 956 5312 1008 5364
rect 1952 5312 2004 5364
rect 4160 5312 4212 5364
rect 4896 5312 4948 5364
rect 5356 5312 5408 5364
rect 6000 5312 6052 5364
rect 8576 5244 8628 5296
rect 8944 5244 8996 5296
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10048 5312 10100 5364
rect 10876 5244 10928 5296
rect 11428 5312 11480 5364
rect 12348 5312 12400 5364
rect 13728 5312 13780 5364
rect 13820 5312 13872 5364
rect 14648 5312 14700 5364
rect 15108 5312 15160 5364
rect 16304 5312 16356 5364
rect 16396 5312 16448 5364
rect 13176 5244 13228 5296
rect 17960 5312 18012 5364
rect 1860 5176 1912 5228
rect 2228 5176 2280 5228
rect 2596 5219 2648 5228
rect 2596 5185 2605 5219
rect 2605 5185 2639 5219
rect 2639 5185 2648 5219
rect 2596 5176 2648 5185
rect 3792 5176 3844 5228
rect 4804 5176 4856 5228
rect 3240 5108 3292 5160
rect 5816 5108 5868 5160
rect 6092 5108 6144 5160
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 7748 5176 7800 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8668 5108 8720 5160
rect 9312 5108 9364 5160
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10692 5176 10744 5228
rect 9772 5108 9824 5160
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11060 5176 11112 5228
rect 11428 5176 11480 5228
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 12440 5176 12492 5228
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 14004 5176 14056 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 15844 5176 15896 5228
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17224 5219 17276 5228
rect 1040 4972 1092 5024
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 2688 4972 2740 5024
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 5724 4972 5776 5024
rect 6000 4972 6052 5024
rect 6276 4972 6328 5024
rect 10692 5040 10744 5092
rect 9680 4972 9732 5024
rect 10140 4972 10192 5024
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17132 5108 17184 5160
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 19064 5244 19116 5296
rect 19432 5287 19484 5296
rect 19432 5253 19441 5287
rect 19441 5253 19475 5287
rect 19475 5253 19484 5287
rect 19432 5244 19484 5253
rect 19892 5312 19944 5364
rect 20812 5312 20864 5364
rect 21456 5312 21508 5364
rect 17776 5176 17828 5228
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 18788 5176 18840 5228
rect 18880 5176 18932 5228
rect 19892 5219 19944 5228
rect 19892 5185 19901 5219
rect 19901 5185 19935 5219
rect 19935 5185 19944 5219
rect 19892 5176 19944 5185
rect 20076 5176 20128 5228
rect 19708 5108 19760 5160
rect 19800 5108 19852 5160
rect 20444 5176 20496 5228
rect 20904 5176 20956 5228
rect 21640 5176 21692 5228
rect 21732 5176 21784 5228
rect 20352 5108 20404 5160
rect 22468 5355 22520 5364
rect 22468 5321 22477 5355
rect 22477 5321 22511 5355
rect 22511 5321 22520 5355
rect 22468 5312 22520 5321
rect 27436 5355 27488 5364
rect 27436 5321 27445 5355
rect 27445 5321 27479 5355
rect 27479 5321 27488 5355
rect 27436 5312 27488 5321
rect 22284 5176 22336 5228
rect 22560 5176 22612 5228
rect 23940 5244 23992 5296
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 24124 5176 24176 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 14280 5040 14332 5092
rect 17316 5040 17368 5092
rect 19984 5040 20036 5092
rect 20260 5040 20312 5092
rect 20720 5040 20772 5092
rect 22836 5040 22888 5092
rect 23388 5040 23440 5092
rect 23572 5040 23624 5092
rect 26240 5040 26292 5092
rect 26424 5040 26476 5092
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 14648 4972 14700 5024
rect 17040 4972 17092 5024
rect 19340 4972 19392 5024
rect 20628 4972 20680 5024
rect 22652 4972 22704 5024
rect 22744 4972 22796 5024
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2228 4768 2280 4820
rect 2320 4768 2372 4820
rect 4620 4768 4672 4820
rect 5540 4768 5592 4820
rect 5632 4768 5684 4820
rect 6000 4768 6052 4820
rect 7840 4768 7892 4820
rect 9496 4768 9548 4820
rect 11244 4768 11296 4820
rect 11796 4768 11848 4820
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 13728 4768 13780 4820
rect 956 4700 1008 4752
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 7380 4700 7432 4752
rect 9036 4700 9088 4752
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 17132 4811 17184 4820
rect 17132 4777 17141 4811
rect 17141 4777 17175 4811
rect 17175 4777 17184 4811
rect 17132 4768 17184 4777
rect 17592 4768 17644 4820
rect 20720 4768 20772 4820
rect 21548 4768 21600 4820
rect 22284 4768 22336 4820
rect 15384 4700 15436 4752
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6736 4564 6788 4616
rect 10140 4632 10192 4684
rect 11704 4632 11756 4684
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 13176 4632 13228 4684
rect 13636 4632 13688 4684
rect 15200 4632 15252 4684
rect 18880 4700 18932 4752
rect 19524 4700 19576 4752
rect 20352 4700 20404 4752
rect 16764 4675 16816 4684
rect 16764 4641 16781 4675
rect 16781 4641 16816 4675
rect 16764 4632 16816 4641
rect 16856 4632 16908 4684
rect 18512 4632 18564 4684
rect 19156 4632 19208 4684
rect 19248 4632 19300 4684
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 7288 4607 7340 4616
rect 7288 4573 7311 4607
rect 7311 4573 7340 4607
rect 7288 4564 7340 4573
rect 9220 4564 9272 4616
rect 9404 4564 9456 4616
rect 12900 4564 12952 4616
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 13912 4564 13964 4616
rect 14648 4564 14700 4616
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 1040 4428 1092 4480
rect 2228 4428 2280 4480
rect 5264 4428 5316 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 5540 4428 5592 4480
rect 10508 4539 10560 4548
rect 10508 4505 10517 4539
rect 10517 4505 10551 4539
rect 10551 4505 10560 4539
rect 10508 4496 10560 4505
rect 10784 4496 10836 4548
rect 7196 4428 7248 4480
rect 7288 4428 7340 4480
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 15108 4496 15160 4548
rect 18328 4496 18380 4548
rect 17592 4428 17644 4480
rect 18236 4428 18288 4480
rect 18512 4496 18564 4548
rect 20076 4632 20128 4684
rect 22560 4743 22612 4752
rect 22560 4709 22569 4743
rect 22569 4709 22603 4743
rect 22603 4709 22612 4743
rect 22560 4700 22612 4709
rect 27436 4811 27488 4820
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 23112 4700 23164 4752
rect 24032 4700 24084 4752
rect 20536 4607 20588 4616
rect 20536 4573 20544 4607
rect 20544 4573 20578 4607
rect 20578 4573 20588 4607
rect 20536 4564 20588 4573
rect 20904 4564 20956 4616
rect 20996 4564 21048 4616
rect 21272 4564 21324 4616
rect 20812 4496 20864 4548
rect 22744 4564 22796 4616
rect 19340 4428 19392 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 20260 4428 20312 4480
rect 20628 4428 20680 4480
rect 20720 4428 20772 4480
rect 22192 4428 22244 4480
rect 22468 4496 22520 4548
rect 22652 4496 22704 4548
rect 26608 4607 26660 4616
rect 26608 4573 26617 4607
rect 26617 4573 26651 4607
rect 26651 4573 26660 4607
rect 26608 4564 26660 4573
rect 27252 4607 27304 4616
rect 27252 4573 27261 4607
rect 27261 4573 27295 4607
rect 27295 4573 27304 4607
rect 27252 4564 27304 4573
rect 23204 4428 23256 4480
rect 26792 4428 26844 4480
rect 27068 4471 27120 4480
rect 27068 4437 27077 4471
rect 27077 4437 27111 4471
rect 27111 4437 27120 4471
rect 27068 4428 27120 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2780 4224 2832 4276
rect 4804 4224 4856 4276
rect 5448 4224 5500 4276
rect 5632 4224 5684 4276
rect 6736 4224 6788 4276
rect 7012 4224 7064 4276
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2504 4088 2556 4140
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 2136 3952 2188 4004
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6000 4156 6052 4208
rect 10324 4224 10376 4276
rect 11244 4224 11296 4276
rect 11980 4224 12032 4276
rect 12072 4267 12124 4276
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 9036 4156 9088 4208
rect 15108 4224 15160 4276
rect 1040 3884 1092 3936
rect 1952 3884 2004 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 4804 3952 4856 4004
rect 4896 3995 4948 4004
rect 4896 3961 4905 3995
rect 4905 3961 4939 3995
rect 4939 3961 4948 3995
rect 4896 3952 4948 3961
rect 5816 4020 5868 4072
rect 6276 4088 6328 4140
rect 7104 4088 7156 4140
rect 7932 4088 7984 4140
rect 7196 4020 7248 4072
rect 7748 4020 7800 4072
rect 8852 4088 8904 4140
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 13728 4156 13780 4208
rect 14372 4156 14424 4208
rect 14924 4199 14976 4208
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 9956 4088 10008 4140
rect 11060 4131 11112 4140
rect 5908 3952 5960 4004
rect 6092 3952 6144 4004
rect 6828 3995 6880 4004
rect 6828 3961 6837 3995
rect 6837 3961 6871 3995
rect 6871 3961 6880 3995
rect 6828 3952 6880 3961
rect 8668 3995 8720 4004
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 11428 4088 11480 4140
rect 12992 4088 13044 4140
rect 14924 4165 14941 4199
rect 14941 4165 14976 4199
rect 14924 4156 14976 4165
rect 16580 4224 16632 4276
rect 17224 4224 17276 4276
rect 17592 4267 17644 4276
rect 17592 4233 17601 4267
rect 17601 4233 17635 4267
rect 17635 4233 17644 4267
rect 17592 4224 17644 4233
rect 18144 4224 18196 4276
rect 18880 4224 18932 4276
rect 19248 4224 19300 4276
rect 19340 4224 19392 4276
rect 16488 4156 16540 4208
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 12072 4020 12124 4072
rect 13820 4020 13872 4072
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 14740 4020 14792 4029
rect 14832 4020 14884 4072
rect 11060 3952 11112 4004
rect 11428 3952 11480 4004
rect 5816 3884 5868 3936
rect 8852 3884 8904 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 10416 3884 10468 3936
rect 10876 3884 10928 3936
rect 12716 3884 12768 3936
rect 12808 3884 12860 3936
rect 15660 3952 15712 4004
rect 15936 4088 15988 4140
rect 16212 4020 16264 4072
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 17684 4088 17736 4140
rect 17040 3952 17092 4004
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 19892 4224 19944 4276
rect 20260 4224 20312 4276
rect 21272 4224 21324 4276
rect 19524 4088 19576 4140
rect 20444 4199 20496 4208
rect 20444 4165 20453 4199
rect 20453 4165 20487 4199
rect 20487 4165 20496 4199
rect 20444 4156 20496 4165
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20352 4020 20404 4072
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16028 3884 16080 3893
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 20536 4088 20588 4140
rect 20996 4088 21048 4140
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 21732 4088 21784 4140
rect 22376 4224 22428 4276
rect 22192 4156 22244 4208
rect 24032 4199 24084 4208
rect 24032 4165 24041 4199
rect 24041 4165 24075 4199
rect 24075 4165 24084 4199
rect 24032 4156 24084 4165
rect 21272 4020 21324 4072
rect 21824 4020 21876 4072
rect 23296 4088 23348 4140
rect 19524 3884 19576 3936
rect 20904 3952 20956 4004
rect 21456 3995 21508 4004
rect 21456 3961 21465 3995
rect 21465 3961 21499 3995
rect 21499 3961 21508 3995
rect 23020 4020 23072 4072
rect 25964 4131 26016 4140
rect 25964 4097 25973 4131
rect 25973 4097 26007 4131
rect 26007 4097 26016 4131
rect 25964 4088 26016 4097
rect 26240 4131 26292 4140
rect 26240 4097 26249 4131
rect 26249 4097 26283 4131
rect 26283 4097 26292 4131
rect 26240 4088 26292 4097
rect 26332 4088 26384 4140
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 21456 3952 21508 3961
rect 23848 3952 23900 4004
rect 26884 3952 26936 4004
rect 27436 3995 27488 4004
rect 27436 3961 27445 3995
rect 27445 3961 27479 3995
rect 27479 3961 27488 3995
rect 27436 3952 27488 3961
rect 21364 3884 21416 3936
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 27068 3927 27120 3936
rect 27068 3893 27077 3927
rect 27077 3893 27111 3927
rect 27111 3893 27120 3927
rect 27068 3884 27120 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2780 3680 2832 3732
rect 4804 3680 4856 3732
rect 6460 3680 6512 3732
rect 7012 3723 7064 3732
rect 7012 3689 7042 3723
rect 7042 3689 7064 3723
rect 7012 3680 7064 3689
rect 956 3612 1008 3664
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 5540 3612 5592 3664
rect 5632 3544 5684 3596
rect 7564 3544 7616 3596
rect 9496 3544 9548 3596
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 1860 3476 1912 3528
rect 2228 3476 2280 3528
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 5540 3476 5592 3528
rect 5724 3476 5776 3528
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 6552 3476 6604 3528
rect 10784 3476 10836 3528
rect 13728 3680 13780 3732
rect 14648 3680 14700 3732
rect 15200 3680 15252 3732
rect 16028 3680 16080 3732
rect 16488 3680 16540 3732
rect 14556 3612 14608 3664
rect 12808 3544 12860 3596
rect 1040 3340 1092 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 5724 3340 5776 3392
rect 6828 3340 6880 3392
rect 7196 3340 7248 3392
rect 7380 3340 7432 3392
rect 11428 3408 11480 3460
rect 11704 3408 11756 3460
rect 11796 3451 11848 3460
rect 11796 3417 11805 3451
rect 11805 3417 11839 3451
rect 11839 3417 11848 3451
rect 11796 3408 11848 3417
rect 10784 3340 10836 3392
rect 13636 3476 13688 3528
rect 14096 3476 14148 3528
rect 14740 3544 14792 3596
rect 17040 3612 17092 3664
rect 19524 3680 19576 3732
rect 19892 3680 19944 3732
rect 16672 3544 16724 3596
rect 16948 3544 17000 3596
rect 17592 3544 17644 3596
rect 18880 3544 18932 3596
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15568 3476 15620 3528
rect 20076 3544 20128 3596
rect 20260 3544 20312 3596
rect 13268 3408 13320 3460
rect 13544 3451 13596 3460
rect 13544 3417 13553 3451
rect 13553 3417 13587 3451
rect 13587 3417 13596 3451
rect 13544 3408 13596 3417
rect 13452 3340 13504 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 18512 3408 18564 3460
rect 18696 3451 18748 3460
rect 18696 3417 18705 3451
rect 18705 3417 18739 3451
rect 18739 3417 18748 3451
rect 18696 3408 18748 3417
rect 18972 3408 19024 3460
rect 21456 3476 21508 3528
rect 22560 3680 22612 3732
rect 19432 3408 19484 3460
rect 16672 3340 16724 3392
rect 16856 3340 16908 3392
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 19800 3408 19852 3460
rect 19984 3408 20036 3460
rect 19616 3340 19668 3392
rect 21824 3408 21876 3460
rect 23664 3476 23716 3528
rect 27068 3680 27120 3732
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 24860 3476 24912 3528
rect 26332 3519 26384 3528
rect 26332 3485 26341 3519
rect 26341 3485 26375 3519
rect 26375 3485 26384 3519
rect 26332 3476 26384 3485
rect 26608 3519 26660 3528
rect 26608 3485 26617 3519
rect 26617 3485 26651 3519
rect 26651 3485 26660 3519
rect 26608 3476 26660 3485
rect 26792 3476 26844 3528
rect 22652 3408 22704 3460
rect 20996 3383 21048 3392
rect 20996 3349 21005 3383
rect 21005 3349 21039 3383
rect 21039 3349 21048 3383
rect 20996 3340 21048 3349
rect 21272 3340 21324 3392
rect 21916 3340 21968 3392
rect 22376 3340 22428 3392
rect 23756 3340 23808 3392
rect 26148 3383 26200 3392
rect 26148 3349 26157 3383
rect 26157 3349 26191 3383
rect 26191 3349 26200 3383
rect 26148 3340 26200 3349
rect 26424 3383 26476 3392
rect 26424 3349 26433 3383
rect 26433 3349 26467 3383
rect 26467 3349 26476 3383
rect 26424 3340 26476 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 27068 3383 27120 3392
rect 27068 3349 27077 3383
rect 27077 3349 27111 3383
rect 27111 3349 27120 3383
rect 27068 3340 27120 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 956 3136 1008 3188
rect 1952 3136 2004 3188
rect 2136 3136 2188 3188
rect 2228 3136 2280 3188
rect 4160 3068 4212 3120
rect 5724 3136 5776 3188
rect 5908 3136 5960 3188
rect 6092 3068 6144 3120
rect 4896 3000 4948 3052
rect 5540 3000 5592 3052
rect 5908 2932 5960 2984
rect 6276 3000 6328 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7932 3136 7984 3188
rect 6828 3000 6880 3052
rect 6736 2932 6788 2984
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 9312 3068 9364 3120
rect 7472 3000 7524 3052
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8944 3000 8996 3052
rect 9220 3000 9272 3052
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 10508 3136 10560 3188
rect 11520 3068 11572 3120
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11244 3000 11296 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 13360 3136 13412 3188
rect 13820 3136 13872 3188
rect 14096 3136 14148 3188
rect 14280 3136 14332 3188
rect 14556 3136 14608 3188
rect 15568 3136 15620 3188
rect 1040 2796 1092 2848
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 3976 2796 4028 2848
rect 4896 2796 4948 2848
rect 5264 2796 5316 2848
rect 7196 2864 7248 2916
rect 9036 2864 9088 2916
rect 11704 2864 11756 2916
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 7104 2796 7156 2848
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 12348 2975 12400 2984
rect 12348 2941 12357 2975
rect 12357 2941 12391 2975
rect 12391 2941 12400 2975
rect 12348 2932 12400 2941
rect 12992 2932 13044 2984
rect 13268 3000 13320 3052
rect 13176 2796 13228 2848
rect 16856 3068 16908 3120
rect 17224 3068 17276 3120
rect 17684 3136 17736 3188
rect 18604 3136 18656 3188
rect 19708 3136 19760 3188
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19156 3043 19208 3052
rect 19156 3009 19165 3043
rect 19165 3009 19199 3043
rect 19199 3009 19208 3043
rect 19156 3000 19208 3009
rect 19432 3068 19484 3120
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 19984 3068 20036 3120
rect 22652 3136 22704 3188
rect 23112 3136 23164 3188
rect 23204 3136 23256 3188
rect 21364 3068 21416 3120
rect 21916 3068 21968 3120
rect 26424 3136 26476 3188
rect 26700 3136 26752 3188
rect 26884 3136 26936 3188
rect 27436 3179 27488 3188
rect 27436 3145 27445 3179
rect 27445 3145 27479 3179
rect 27479 3145 27488 3179
rect 27436 3136 27488 3145
rect 14188 2932 14240 2984
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 15200 2932 15252 2984
rect 18144 2932 18196 2984
rect 21456 2932 21508 2984
rect 22376 2975 22428 2984
rect 22376 2941 22385 2975
rect 22385 2941 22419 2975
rect 22419 2941 22428 2975
rect 22376 2932 22428 2941
rect 22928 2932 22980 2984
rect 25412 3068 25464 3120
rect 23296 3000 23348 3052
rect 23848 3000 23900 3052
rect 24492 3043 24544 3052
rect 24492 3009 24501 3043
rect 24501 3009 24535 3043
rect 24535 3009 24544 3043
rect 24492 3000 24544 3009
rect 25504 3043 25556 3052
rect 25504 3009 25513 3043
rect 25513 3009 25547 3043
rect 25547 3009 25556 3043
rect 25504 3000 25556 3009
rect 23756 2975 23808 2984
rect 15384 2796 15436 2848
rect 15476 2796 15528 2848
rect 15936 2796 15988 2848
rect 19524 2839 19576 2848
rect 19524 2805 19533 2839
rect 19533 2805 19567 2839
rect 19567 2805 19576 2839
rect 19524 2796 19576 2805
rect 22468 2907 22520 2916
rect 22468 2873 22477 2907
rect 22477 2873 22511 2907
rect 22511 2873 22520 2907
rect 22468 2864 22520 2873
rect 23756 2941 23765 2975
rect 23765 2941 23799 2975
rect 23799 2941 23808 2975
rect 23756 2932 23808 2941
rect 23940 2932 23992 2984
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 26608 2864 26660 2916
rect 24584 2839 24636 2848
rect 24584 2805 24593 2839
rect 24593 2805 24627 2839
rect 24627 2805 24636 2839
rect 24584 2796 24636 2805
rect 25872 2839 25924 2848
rect 25872 2805 25881 2839
rect 25881 2805 25915 2839
rect 25915 2805 25924 2839
rect 25872 2796 25924 2805
rect 26056 2796 26108 2848
rect 26700 2839 26752 2848
rect 26700 2805 26709 2839
rect 26709 2805 26743 2839
rect 26743 2805 26752 2839
rect 26700 2796 26752 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 5448 2592 5500 2644
rect 1216 2524 1268 2576
rect 6736 2592 6788 2644
rect 7012 2592 7064 2644
rect 7104 2592 7156 2644
rect 8852 2592 8904 2644
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13176 2592 13228 2644
rect 14372 2592 14424 2644
rect 14740 2592 14792 2644
rect 14924 2592 14976 2644
rect 15476 2592 15528 2644
rect 15568 2592 15620 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 17132 2592 17184 2644
rect 18788 2592 18840 2644
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 1308 2456 1360 2508
rect 4896 2499 4948 2508
rect 4896 2465 4905 2499
rect 4905 2465 4939 2499
rect 4939 2465 4948 2499
rect 4896 2456 4948 2465
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 1042 2320 1094 2372
rect 1768 2363 1820 2372
rect 1768 2329 1777 2363
rect 1777 2329 1811 2363
rect 1811 2329 1820 2363
rect 1768 2320 1820 2329
rect 2504 2320 2556 2372
rect 3424 2388 3476 2440
rect 5448 2456 5500 2508
rect 6276 2388 6328 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7564 2388 7616 2440
rect 7656 2388 7708 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 11888 2524 11940 2576
rect 8208 2456 8260 2508
rect 8944 2388 8996 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10784 2388 10836 2440
rect 12348 2388 12400 2440
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 13268 2388 13320 2440
rect 1584 2252 1636 2304
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 4620 2252 4672 2304
rect 6184 2252 6236 2304
rect 7104 2252 7156 2304
rect 15108 2524 15160 2576
rect 15292 2524 15344 2576
rect 16948 2524 17000 2576
rect 14556 2456 14608 2508
rect 14372 2388 14424 2440
rect 14924 2388 14976 2440
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15384 2388 15436 2440
rect 16304 2388 16356 2440
rect 8024 2252 8076 2304
rect 9864 2252 9916 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 13544 2252 13596 2304
rect 14184 2252 14236 2304
rect 15568 2320 15620 2372
rect 18144 2388 18196 2440
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 19984 2388 20036 2440
rect 21364 2524 21416 2576
rect 19800 2320 19852 2372
rect 22744 2524 22796 2576
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 24492 2524 24544 2576
rect 21824 2388 21876 2440
rect 22376 2388 22428 2440
rect 23020 2499 23072 2508
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 22928 2388 22980 2440
rect 23848 2431 23900 2440
rect 23848 2397 23857 2431
rect 23857 2397 23891 2431
rect 23891 2397 23900 2431
rect 23848 2388 23900 2397
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 26148 2431 26200 2440
rect 26148 2397 26157 2431
rect 26157 2397 26191 2431
rect 26191 2397 26200 2431
rect 26148 2388 26200 2397
rect 26608 2388 26660 2440
rect 26424 2320 26476 2372
rect 27827 2320 27879 2372
rect 15292 2252 15344 2304
rect 15384 2252 15436 2304
rect 17224 2252 17276 2304
rect 19064 2252 19116 2304
rect 20904 2252 20956 2304
rect 21640 2252 21692 2304
rect 22928 2252 22980 2304
rect 23940 2252 23992 2304
rect 24584 2252 24636 2304
rect 25504 2252 25556 2304
rect 26332 2295 26384 2304
rect 26332 2261 26341 2295
rect 26341 2261 26375 2295
rect 26375 2261 26384 2295
rect 26332 2252 26384 2261
rect 27068 2252 27120 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 2688 2048 2740 2100
rect 2320 1912 2372 1964
rect 8392 1912 8444 1964
rect 14184 2048 14236 2100
rect 27200 2048 27252 2100
rect 17392 1980 17444 2032
rect 24860 1980 24912 2032
rect 23412 1912 23464 1964
rect 4804 1844 4856 1896
rect 27292 1844 27344 1896
rect 3792 1776 3844 1828
rect 17040 1776 17092 1828
rect 17392 1776 17444 1828
rect 5632 1708 5684 1760
<< metal2 >>
rect 10324 8016 10376 8022
rect 1122 7984 1178 7993
rect 1122 7919 1178 7928
rect 1030 7712 1086 7721
rect 1030 7647 1086 7656
rect 1044 7546 1072 7647
rect 1032 7540 1084 7546
rect 1032 7482 1084 7488
rect 1136 7342 1164 7919
rect 1306 7580 1362 7980
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1320 7478 1348 7580
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1490 7168 1546 7177
rect 1490 7103 1546 7112
rect 1504 7002 1532 7103
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1688 6798 1716 7890
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 1858 7440 1914 7449
rect 2240 7410 2268 7686
rect 3146 7580 3202 7980
rect 4709 7580 4765 7980
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 3160 7478 3188 7580
rect 4724 7478 4752 7580
rect 4874 7579 5182 7588
rect 6550 7580 6606 7980
rect 8298 7580 8354 7980
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 6564 7546 6592 7580
rect 8312 7546 8340 7580
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 1858 7375 1914 7384
rect 2228 7404 2280 7410
rect 1872 7002 1900 7375
rect 2228 7346 2280 7352
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 2424 6905 2452 7142
rect 2608 6914 2636 7346
rect 3528 7002 3556 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 2410 6896 2466 6905
rect 2608 6886 2728 6914
rect 2410 6831 2466 6840
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 1124 6656 1176 6662
rect 954 6624 1010 6633
rect 1124 6598 1176 6604
rect 954 6559 1010 6568
rect 968 6458 996 6559
rect 956 6452 1008 6458
rect 956 6394 1008 6400
rect 1136 6361 1164 6598
rect 2056 6440 2084 6734
rect 2056 6412 2176 6440
rect 1122 6352 1178 6361
rect 2042 6352 2098 6361
rect 1122 6287 1178 6296
rect 1952 6316 2004 6322
rect 2042 6287 2044 6296
rect 1952 6258 2004 6264
rect 2096 6287 2098 6296
rect 2044 6258 2096 6264
rect 1040 6180 1092 6186
rect 1040 6122 1092 6128
rect 1052 6089 1080 6122
rect 1038 6080 1094 6089
rect 1038 6015 1094 6024
rect 956 5840 1008 5846
rect 954 5808 956 5817
rect 1008 5808 1010 5817
rect 954 5743 1010 5752
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 1688 5710 1716 5743
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1860 5568 1912 5574
rect 1858 5536 1860 5545
rect 1912 5536 1914 5545
rect 1858 5471 1914 5480
rect 1964 5370 1992 6258
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5710 2084 6054
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 956 5364 1008 5370
rect 956 5306 1008 5312
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 968 5273 996 5306
rect 954 5264 1010 5273
rect 954 5199 1010 5208
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1040 5024 1092 5030
rect 1038 4992 1040 5001
rect 1092 4992 1094 5001
rect 1038 4927 1094 4936
rect 956 4752 1008 4758
rect 954 4720 956 4729
rect 1008 4720 1010 4729
rect 954 4655 1010 4664
rect 1040 4480 1092 4486
rect 1038 4448 1040 4457
rect 1092 4448 1094 4457
rect 1038 4383 1094 4392
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1504 4010 1532 4111
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1040 3936 1092 3942
rect 1038 3904 1040 3913
rect 1092 3904 1094 3913
rect 1038 3839 1094 3848
rect 956 3664 1008 3670
rect 954 3632 956 3641
rect 1008 3632 1010 3641
rect 954 3567 1010 3576
rect 1872 3534 1900 5170
rect 2148 4593 2176 6412
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2240 5114 2268 5170
rect 2240 5086 2360 5114
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4826 2268 4966
rect 2332 4826 2360 5086
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2318 4720 2374 4729
rect 2318 4655 2374 4664
rect 2332 4622 2360 4655
rect 2320 4616 2372 4622
rect 2134 4584 2190 4593
rect 2320 4558 2372 4564
rect 2134 4519 2190 4528
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1040 3392 1092 3398
rect 1038 3360 1040 3369
rect 1092 3360 1094 3369
rect 1038 3295 1094 3304
rect 1964 3194 1992 3878
rect 2148 3194 2176 3946
rect 2240 3534 2268 4422
rect 2424 4185 2452 6734
rect 2594 5264 2650 5273
rect 2594 5199 2596 5208
rect 2648 5199 2650 5208
rect 2596 5170 2648 5176
rect 2594 5128 2650 5137
rect 2700 5114 2728 6886
rect 4172 6798 4200 6938
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6458 4568 6598
rect 4724 6458 4752 6802
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5368 6390 5396 6598
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5778 3924 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4172 5370 4200 5578
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4816 5234 4844 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5368 5370 5396 6326
rect 5460 6322 5488 6938
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5642 5488 6122
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 2650 5086 2728 5114
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 2594 5063 2650 5072
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2410 4176 2466 4185
rect 2320 4140 2372 4146
rect 2516 4146 2544 4966
rect 2410 4111 2466 4120
rect 2504 4140 2556 4146
rect 2320 4082 2372 4088
rect 2504 4082 2556 4088
rect 2332 4049 2360 4082
rect 2318 4040 2374 4049
rect 2318 3975 2374 3984
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3194 2268 3334
rect 956 3188 1008 3194
rect 956 3130 1008 3136
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 968 3097 996 3130
rect 954 3088 1010 3097
rect 954 3023 1010 3032
rect 1040 2848 1092 2854
rect 1038 2816 1040 2825
rect 2228 2848 2280 2854
rect 1092 2816 1094 2825
rect 2228 2790 2280 2796
rect 1038 2751 1094 2760
rect 2240 2689 2268 2790
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 1216 2576 1268 2582
rect 1216 2518 1268 2524
rect 2226 2544 2282 2553
rect 1042 2372 1094 2378
rect 1042 2314 1094 2320
rect 1054 1760 1082 2314
rect 1228 2281 1256 2518
rect 1308 2508 1360 2514
rect 2226 2479 2282 2488
rect 1308 2450 1360 2456
rect 1214 2272 1270 2281
rect 1214 2207 1270 2216
rect 1320 2009 1348 2450
rect 2240 2446 2268 2479
rect 2228 2440 2280 2446
rect 1766 2408 1822 2417
rect 2228 2382 2280 2388
rect 1766 2343 1768 2352
rect 1820 2343 1822 2352
rect 1768 2314 1820 2320
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1596 1760 1624 2246
rect 2332 1970 2360 3470
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 2446 2636 2790
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 2516 1760 2544 2314
rect 2700 2106 2728 4966
rect 2792 4282 2820 4966
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3738 2820 3878
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2884 2961 2912 4082
rect 3252 3505 3280 5102
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2428 2912 2790
rect 3252 2650 3280 3431
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2964 2440 3016 2446
rect 2884 2400 2964 2428
rect 2964 2382 3016 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 3436 1760 3464 2382
rect 3804 1834 3832 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3988 2854 4016 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4250 3632 4306 3641
rect 4160 3596 4212 3602
rect 4212 3576 4250 3584
rect 4212 3567 4306 3576
rect 4212 3556 4292 3567
rect 4160 3538 4212 3544
rect 4172 3126 4200 3538
rect 4160 3120 4212 3126
rect 4632 3097 4660 4762
rect 4908 4570 4936 5306
rect 5262 4992 5318 5001
rect 5262 4927 5318 4936
rect 5276 4690 5304 4927
rect 5460 4706 5488 5578
rect 5552 4826 5580 6802
rect 5644 4826 5672 7346
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6934 5856 7142
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 6012 6798 6040 7482
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 7002 6776 7346
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 5030 5764 6598
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5908 6248 5960 6254
rect 5906 6216 5908 6225
rect 5960 6216 5962 6225
rect 5906 6151 5962 6160
rect 6104 5914 6132 6258
rect 6196 5914 6224 6734
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 5906 5672 5962 5681
rect 5906 5607 5908 5616
rect 5960 5607 5962 5616
rect 6000 5636 6052 5642
rect 5908 5578 5960 5584
rect 6000 5578 6052 5584
rect 6012 5370 6040 5578
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6104 5166 6132 5850
rect 6196 5574 6224 5850
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5264 4684 5316 4690
rect 5460 4678 5764 4706
rect 5264 4626 5316 4632
rect 4816 4542 4936 4570
rect 4816 4282 4844 4542
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4816 3738 4844 3946
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4908 3584 4936 3946
rect 4816 3556 4936 3584
rect 5184 3584 5212 4082
rect 5276 3777 5304 4422
rect 5460 4282 5488 4422
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5184 3556 5304 3584
rect 4160 3062 4212 3068
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 4816 3040 4844 3556
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4896 3052 4948 3058
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2310 4660 3023
rect 4816 3012 4896 3040
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 3988 2009 4016 2246
rect 4448 2190 4476 2246
rect 4356 2162 4476 2190
rect 3974 2000 4030 2009
rect 3974 1935 4030 1944
rect 3792 1828 3844 1834
rect 3792 1770 3844 1776
rect 4356 1760 4384 2162
rect 4816 1902 4844 3012
rect 4896 2994 4948 3000
rect 5276 2854 5304 3556
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 4908 2514 4936 2790
rect 5460 2650 5488 4082
rect 5552 3670 5580 4422
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5644 3602 5672 4218
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5736 3534 5764 4678
rect 5828 4078 5856 5102
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4826 6040 4966
rect 6000 4820 6052 4826
rect 5920 4780 6000 4808
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5920 4010 5948 4780
rect 6000 4762 6052 4768
rect 6104 4706 6132 5102
rect 6288 5030 6316 6666
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6104 4678 6316 4706
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 4457 6224 4558
rect 6182 4448 6238 4457
rect 6182 4383 6238 4392
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5816 3936 5868 3942
rect 6012 3890 6040 4150
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5868 3884 6040 3890
rect 5816 3878 6040 3884
rect 5828 3862 6040 3878
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5552 3058 5580 3470
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3194 5764 3334
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5736 2774 5764 3130
rect 5920 2990 5948 3130
rect 6104 3126 6132 3946
rect 6196 3534 6224 4383
rect 6288 4146 6316 4678
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6288 3058 6316 4082
rect 6380 3058 6408 6598
rect 6564 6458 6592 6734
rect 6932 6458 6960 7278
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6866 8340 7210
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6550 5944 6606 5953
rect 6550 5879 6552 5888
rect 6604 5879 6606 5888
rect 6552 5850 6604 5856
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6472 3738 6500 5714
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6472 3641 6500 3674
rect 6458 3632 6514 3641
rect 6458 3567 6514 3576
rect 6564 3534 6592 5850
rect 6656 5234 6684 6190
rect 6748 5234 6776 6326
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5234 6868 5510
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6656 5001 6684 5170
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4282 6776 4558
rect 7024 4282 7052 6054
rect 7576 5914 7604 6054
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7760 5794 7788 6326
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5914 7880 6190
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7760 5766 7880 5794
rect 7852 5710 7880 5766
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7104 5704 7156 5710
rect 7102 5672 7104 5681
rect 7748 5704 7800 5710
rect 7156 5672 7158 5681
rect 7748 5646 7800 5652
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7102 5607 7158 5616
rect 7760 5234 7788 5646
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7380 4752 7432 4758
rect 7116 4712 7380 4740
rect 7116 4622 7144 4712
rect 7432 4712 7512 4740
rect 7380 4694 7432 4700
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4486 7328 4558
rect 7196 4480 7248 4486
rect 7288 4480 7340 4486
rect 7196 4422 7248 4428
rect 7286 4448 7288 4457
rect 7340 4448 7342 4457
rect 7208 4298 7236 4422
rect 7286 4383 7342 4392
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 7012 4276 7064 4282
rect 7208 4270 7328 4298
rect 7012 4218 7064 4224
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6748 3233 6776 4218
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6840 3890 6868 3946
rect 6918 3904 6974 3913
rect 6840 3862 6918 3890
rect 6918 3839 6974 3848
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6734 3224 6790 3233
rect 6734 3159 6790 3168
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5908 2984 5960 2990
rect 6380 2938 6408 2994
rect 6748 2990 6776 3159
rect 6840 3058 6868 3334
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 5908 2926 5960 2932
rect 5644 2746 5764 2774
rect 6288 2910 6408 2938
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 4874 2204 5182 2213
rect 5460 2206 5488 2450
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 2178 5488 2206
rect 4804 1896 4856 1902
rect 4804 1838 4856 1844
rect 5276 1760 5304 2178
rect 5644 1766 5672 2746
rect 6288 2446 6316 2910
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6380 2446 6408 2790
rect 6748 2650 6776 2926
rect 7024 2650 7052 3674
rect 7116 2854 7144 4082
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3398 7236 4014
rect 7300 3641 7328 4270
rect 7286 3632 7342 3641
rect 7286 3567 7342 3576
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3058 7236 3334
rect 7300 3058 7328 3567
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2650 7144 2790
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7104 2440 7156 2446
rect 7208 2428 7236 2858
rect 7392 2774 7420 3334
rect 7484 3058 7512 4712
rect 7654 4312 7710 4321
rect 7654 4247 7656 4256
rect 7708 4247 7710 4256
rect 7656 4218 7708 4224
rect 7760 4078 7788 5170
rect 7852 4826 7880 5646
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7944 4146 7972 5714
rect 8036 5234 8064 6054
rect 8298 5944 8354 5953
rect 8220 5902 8298 5930
rect 8220 5642 8248 5902
rect 8496 5914 8524 6734
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8298 5879 8354 5888
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8588 5302 8616 6598
rect 8680 5710 8708 6802
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8680 5166 8708 5510
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7748 4072 7800 4078
rect 8772 4026 8800 7822
rect 10046 7580 10102 7980
rect 24308 8016 24360 8022
rect 10324 7958 10376 7964
rect 10060 7546 10088 7580
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9048 7002 9076 7346
rect 10244 7002 10272 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9140 6390 9168 6734
rect 9416 6458 9444 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8852 5840 8904 5846
rect 8956 5828 8984 6258
rect 9232 6089 9260 6258
rect 9784 6254 9812 6598
rect 9876 6322 9904 6734
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9218 6080 9274 6089
rect 9218 6015 9274 6024
rect 8904 5800 8984 5828
rect 8852 5782 8904 5788
rect 8956 5302 8984 5800
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 7748 4014 7800 4020
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7576 3058 7604 3538
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7484 2836 7512 2994
rect 7484 2808 7604 2836
rect 7392 2746 7512 2774
rect 7484 2446 7512 2746
rect 7576 2446 7604 2808
rect 7156 2400 7236 2428
rect 7472 2440 7524 2446
rect 7104 2382 7156 2388
rect 7472 2382 7524 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7656 2440 7708 2446
rect 7760 2428 7788 4014
rect 8680 4010 8800 4026
rect 8668 4004 8800 4010
rect 8720 3998 8800 4004
rect 8668 3946 8720 3952
rect 8206 3904 8262 3913
rect 8206 3839 8262 3848
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7944 2446 7972 3130
rect 8220 2514 8248 3839
rect 8680 2774 8708 3946
rect 8864 3942 8892 4082
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8404 2746 8708 2774
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 7708 2400 7788 2428
rect 7932 2440 7984 2446
rect 7656 2382 7708 2388
rect 7932 2382 7984 2388
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 5632 1760 5684 1766
rect 6196 1760 6224 2246
rect 7116 1760 7144 2246
rect 8036 1760 8064 2246
rect 8404 1970 8432 2746
rect 8864 2650 8892 3878
rect 8956 3058 8984 5238
rect 9048 4758 9076 5578
rect 9324 5166 9352 6122
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 9048 4214 9076 4694
rect 9220 4616 9272 4622
rect 9324 4604 9352 5102
rect 9508 4826 9536 5714
rect 9968 5370 9996 6802
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10060 5370 10088 6734
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6186 10180 6598
rect 10244 6322 10272 6734
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10244 5953 10272 6258
rect 10230 5944 10286 5953
rect 10230 5879 10286 5888
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 5024 9732 5030
rect 9784 5012 9812 5102
rect 9732 4984 9812 5012
rect 9680 4966 9732 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9272 4576 9352 4604
rect 9404 4616 9456 4622
rect 9220 4558 9272 4564
rect 9404 4558 9456 4564
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9048 2922 9076 4150
rect 9232 4146 9260 4558
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9312 4140 9364 4146
rect 9416 4128 9444 4558
rect 9586 4312 9642 4321
rect 9586 4247 9642 4256
rect 9364 4100 9444 4128
rect 9312 4082 9364 4088
rect 9232 3058 9260 4082
rect 9324 3641 9352 4082
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9310 3632 9366 3641
rect 9508 3602 9536 3878
rect 9310 3567 9366 3576
rect 9496 3596 9548 3602
rect 9324 3126 9352 3567
rect 9496 3538 9548 3544
rect 9600 3233 9628 4247
rect 9692 4146 9720 4966
rect 9968 4146 9996 5306
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4690 10180 4966
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10336 4282 10364 7958
rect 11794 7580 11850 7980
rect 13542 7580 13598 7980
rect 15290 7580 15346 7980
rect 17038 7580 17094 7980
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 11808 7546 11836 7580
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 13556 7478 13584 7580
rect 15304 7546 15332 7580
rect 17052 7546 17080 7580
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 11532 7002 11560 7346
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 12990 6896 13046 6905
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10520 6322 10548 6802
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10428 3942 10456 6258
rect 10508 6112 10560 6118
rect 10612 6100 10640 6258
rect 10560 6072 10640 6100
rect 10508 6054 10560 6060
rect 10520 5234 10548 6054
rect 10704 5914 10732 6802
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 6458 10916 6666
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5234 10732 5850
rect 10796 5817 10824 6054
rect 10782 5808 10838 5817
rect 10980 5778 11008 6734
rect 10782 5743 10838 5752
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 9586 3224 9642 3233
rect 10520 3194 10548 4490
rect 10612 3233 10640 5102
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 5001 10732 5034
rect 10690 4992 10746 5001
rect 10690 4927 10746 4936
rect 10796 4554 10824 5578
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10888 4865 10916 5238
rect 10980 5234 11008 5714
rect 11072 5234 11100 6870
rect 14292 6866 14320 7346
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 12990 6831 13046 6840
rect 14096 6860 14148 6866
rect 11150 6760 11206 6769
rect 11150 6695 11152 6704
rect 11204 6695 11206 6704
rect 11702 6760 11758 6769
rect 13004 6730 13032 6831
rect 14096 6802 14148 6808
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13726 6760 13782 6769
rect 11702 6695 11758 6704
rect 12992 6724 13044 6730
rect 11152 6666 11204 6672
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11440 6390 11468 6598
rect 11428 6384 11480 6390
rect 11334 6352 11390 6361
rect 11244 6316 11296 6322
rect 11428 6326 11480 6332
rect 11334 6287 11390 6296
rect 11244 6258 11296 6264
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10874 4856 10930 4865
rect 11256 4826 11284 6258
rect 10874 4791 10930 4800
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 3534 10824 4490
rect 11256 4282 11284 4762
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11060 4140 11112 4146
rect 11112 4100 11192 4128
rect 11060 4082 11112 4088
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3398 10824 3470
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10598 3224 10654 3233
rect 9586 3159 9642 3168
rect 10508 3188 10560 3194
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9600 2990 9628 3159
rect 10598 3159 10654 3168
rect 10508 3130 10560 3136
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8944 2440 8996 2446
rect 9876 2428 9904 2790
rect 10888 2650 10916 3878
rect 11072 3058 11100 3946
rect 11164 3602 11192 4100
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11256 3058 11284 4218
rect 11348 3913 11376 6287
rect 11520 6180 11572 6186
rect 11572 6140 11652 6168
rect 11520 6122 11572 6128
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11440 5370 11468 5578
rect 11624 5574 11652 6140
rect 11716 5778 11744 6695
rect 12992 6666 13044 6672
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5914 11836 6190
rect 11888 6112 11940 6118
rect 11980 6112 12032 6118
rect 11888 6054 11940 6060
rect 11978 6080 11980 6089
rect 12032 6080 12034 6089
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11440 5001 11468 5170
rect 11426 4992 11482 5001
rect 11426 4927 11482 4936
rect 11716 4690 11744 5714
rect 11900 5710 11928 6054
rect 11978 6015 12034 6024
rect 12084 5914 12112 6598
rect 12728 6458 12756 6598
rect 13188 6458 13216 6734
rect 13452 6724 13504 6730
rect 13726 6695 13728 6704
rect 13452 6666 13504 6672
rect 13780 6695 13782 6704
rect 13728 6666 13780 6672
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 12268 5370 12388 5386
rect 12268 5364 12400 5370
rect 12268 5358 12348 5364
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11440 4010 11468 4082
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11334 3904 11390 3913
rect 11334 3839 11390 3848
rect 11440 3466 11468 3946
rect 11716 3466 11744 4626
rect 11808 4078 11836 4762
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 11992 4282 12020 4383
rect 12084 4282 12112 5102
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 3210 11836 3402
rect 11716 3182 11836 3210
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11532 2825 11560 3062
rect 11716 2922 11744 3182
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11900 2582 11928 3062
rect 12084 3040 12112 4014
rect 12176 3913 12204 4422
rect 12268 4049 12296 5358
rect 12348 5306 12400 5312
rect 12452 5234 12480 6394
rect 13188 6225 13216 6394
rect 13174 6216 13230 6225
rect 13174 6151 13230 6160
rect 12898 5808 12954 5817
rect 12728 5752 12898 5760
rect 12728 5732 12900 5752
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12360 4826 12388 5170
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12452 4690 12480 5170
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12254 4040 12310 4049
rect 12254 3975 12310 3984
rect 12728 3942 12756 5732
rect 12952 5743 12954 5752
rect 12900 5714 12952 5720
rect 13188 5302 13216 6151
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4622 12940 4966
rect 13188 4690 13216 5238
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12716 3936 12768 3942
rect 12162 3904 12218 3913
rect 12716 3878 12768 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12162 3839 12218 3848
rect 12820 3641 12848 3878
rect 12806 3632 12862 3641
rect 12806 3567 12808 3576
rect 12860 3567 12862 3576
rect 12808 3538 12860 3544
rect 12256 3052 12308 3058
rect 12084 3012 12256 3040
rect 12256 2994 12308 3000
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 12360 2446 12388 2926
rect 12912 2650 12940 4558
rect 13004 4146 13032 4558
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4185 13216 4422
rect 13174 4176 13230 4185
rect 12992 4140 13044 4146
rect 13174 4111 13230 4120
rect 12992 4082 13044 4088
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13280 3176 13308 3402
rect 13464 3398 13492 6666
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5574 13584 6258
rect 13740 5642 13768 6666
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13726 5536 13782 5545
rect 13726 5471 13782 5480
rect 13740 5370 13768 5471
rect 13832 5370 13860 5850
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13648 4690 13676 5170
rect 13740 4826 13768 5170
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13636 4684 13688 4690
rect 13556 4644 13636 4672
rect 13556 3466 13584 4644
rect 13636 4626 13688 4632
rect 13924 4622 13952 5714
rect 14016 5710 14044 6258
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14016 5234 14044 5646
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 14002 4176 14058 4185
rect 13740 3738 13768 4150
rect 14002 4111 14058 4120
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13740 3618 13768 3674
rect 13648 3590 13768 3618
rect 13648 3534 13676 3590
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13832 3194 13860 4014
rect 14016 3913 14044 4111
rect 14002 3904 14058 3913
rect 14002 3839 14058 3848
rect 14108 3534 14136 6802
rect 14384 6798 14412 7210
rect 14476 7002 14504 7346
rect 15108 7336 15160 7342
rect 15160 7284 15240 7290
rect 15108 7278 15240 7284
rect 15120 7262 15240 7278
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14660 6458 14688 7142
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15028 6254 15056 6802
rect 14280 6248 14332 6254
rect 14648 6248 14700 6254
rect 14280 6190 14332 6196
rect 14462 6216 14518 6225
rect 14292 5098 14320 6190
rect 14648 6190 14700 6196
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 14462 6151 14518 6160
rect 14476 6118 14504 6151
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14384 5778 14412 6054
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14476 5642 14504 6054
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3194 14136 3334
rect 13004 3148 13308 3176
rect 13004 2990 13032 3148
rect 13280 3058 13308 3148
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13188 2650 13216 2790
rect 13372 2774 13400 3130
rect 14200 2990 14228 4422
rect 14384 4298 14412 5510
rect 14292 4270 14412 4298
rect 14292 3194 14320 4270
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13280 2746 13400 2774
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13280 2446 13308 2746
rect 14384 2650 14412 4150
rect 14476 4060 14504 5578
rect 14554 5400 14610 5409
rect 14660 5370 14688 6190
rect 15014 5672 15070 5681
rect 15014 5607 15070 5616
rect 14554 5335 14610 5344
rect 14648 5364 14700 5370
rect 14568 5234 14596 5335
rect 14648 5306 14700 5312
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4826 14688 4966
rect 14922 4856 14978 4865
rect 14648 4820 14700 4826
rect 14922 4791 14978 4800
rect 14648 4762 14700 4768
rect 14648 4616 14700 4622
rect 14700 4576 14780 4604
rect 14648 4558 14700 4564
rect 14752 4078 14780 4576
rect 14936 4214 14964 4791
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14648 4072 14700 4078
rect 14476 4032 14648 4060
rect 14568 3670 14596 4032
rect 14648 4014 14700 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14568 3194 14596 3606
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14660 2961 14688 3674
rect 14752 3602 14780 4014
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14844 3534 14872 4014
rect 14936 3777 14964 4150
rect 14922 3768 14978 3777
rect 14922 3703 14978 3712
rect 15028 3641 15056 5607
rect 15212 5574 15240 7262
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 15396 6905 15424 7142
rect 15382 6896 15438 6905
rect 15842 6896 15898 6905
rect 15382 6831 15438 6840
rect 15568 6860 15620 6866
rect 15842 6831 15898 6840
rect 16120 6860 16172 6866
rect 15568 6802 15620 6808
rect 15580 6730 15608 6802
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15120 5370 15148 5510
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15396 5166 15424 6054
rect 15580 5778 15608 6666
rect 15672 5914 15700 6666
rect 15764 6225 15792 6666
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15120 4282 15148 4490
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15212 3738 15240 4626
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15014 3632 15070 3641
rect 15014 3567 15070 3576
rect 15304 3534 15332 3878
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15212 2990 15240 3470
rect 15396 3074 15424 4694
rect 15580 3534 15608 5714
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 4010 15700 5646
rect 15856 5234 15884 6831
rect 16120 6802 16172 6808
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6390 16068 6734
rect 16132 6458 16160 6802
rect 16408 6730 16436 7142
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5234 16252 6054
rect 16408 5953 16436 6666
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16394 5944 16450 5953
rect 16394 5879 16450 5888
rect 16500 5574 16528 6598
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16316 5370 16344 5510
rect 16394 5400 16450 5409
rect 16304 5364 16356 5370
rect 16394 5335 16396 5344
rect 16304 5306 16356 5312
rect 16448 5335 16450 5344
rect 16396 5306 16448 5312
rect 16868 5234 16896 5578
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3194 15608 3470
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15396 3046 15608 3074
rect 14740 2984 14792 2990
rect 14646 2952 14702 2961
rect 15200 2984 15252 2990
rect 14740 2926 14792 2932
rect 15120 2944 15200 2972
rect 14646 2887 14702 2896
rect 14752 2650 14780 2926
rect 14922 2816 14978 2825
rect 14922 2751 14978 2760
rect 14936 2650 14964 2751
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14384 2446 14412 2586
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 9956 2440 10008 2446
rect 9876 2400 9956 2428
rect 8944 2382 8996 2388
rect 9956 2382 10008 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 12348 2440 12400 2446
rect 12716 2440 12768 2446
rect 12348 2382 12400 2388
rect 12636 2400 12716 2428
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8956 1760 8984 2382
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9876 1760 9904 2246
rect 10796 1760 10824 2382
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 2190 11928 2246
rect 11716 2162 11928 2190
rect 11716 1760 11744 2162
rect 12636 1760 12664 2400
rect 12716 2382 12768 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14184 2304 14236 2310
rect 14184 2246 14236 2252
rect 13556 1760 13584 2246
rect 14196 2106 14224 2246
rect 14568 2186 14596 2450
rect 14936 2446 14964 2586
rect 15120 2582 15148 2944
rect 15200 2926 15252 2932
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15120 2446 15148 2518
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15304 2310 15332 2518
rect 15396 2446 15424 2790
rect 15488 2650 15516 2790
rect 15580 2650 15608 3046
rect 15948 2854 15976 4082
rect 16224 4078 16252 5170
rect 16762 4992 16818 5001
rect 16762 4927 16818 4936
rect 16776 4690 16804 4927
rect 16868 4690 16896 5170
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 4282 16620 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 3738 16068 3878
rect 16500 3738 16528 4150
rect 16960 4146 16988 6258
rect 17052 6254 17080 6734
rect 17328 6662 17356 7890
rect 18786 7580 18842 7980
rect 20534 7580 20590 7980
rect 22282 7580 22338 7980
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 18800 7546 18828 7580
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 20548 7478 20576 7580
rect 22296 7478 22324 7580
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19444 7290 19472 7346
rect 20076 7336 20128 7342
rect 19444 7262 20024 7290
rect 20076 7278 20128 7284
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 18708 7002 18736 7142
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5030 17080 6054
rect 17236 5234 17264 6122
rect 17328 5409 17356 6598
rect 17604 5868 18000 5896
rect 17314 5400 17370 5409
rect 17314 5335 17370 5344
rect 17498 5264 17554 5273
rect 17224 5228 17276 5234
rect 17498 5199 17500 5208
rect 17224 5170 17276 5176
rect 17552 5199 17554 5208
rect 17500 5170 17552 5176
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 3754 16988 4082
rect 17052 4010 17080 4966
rect 17144 4826 17172 5102
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16488 3732 16540 3738
rect 16960 3726 17080 3754
rect 16488 3674 16540 3680
rect 17052 3670 17080 3726
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16672 3596 16724 3602
rect 16948 3596 17000 3602
rect 16724 3556 16896 3584
rect 16672 3538 16724 3544
rect 16868 3398 16896 3556
rect 16948 3538 17000 3544
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 16684 2650 16712 3334
rect 16868 3126 16896 3334
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16960 2582 16988 3538
rect 17144 2650 17172 4762
rect 17236 4282 17264 5170
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17236 3126 17264 3878
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 15384 2440 15436 2446
rect 16304 2440 16356 2446
rect 15436 2388 15608 2394
rect 15384 2382 15608 2388
rect 17328 2394 17356 5034
rect 17604 4826 17632 5868
rect 17972 5778 18000 5868
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17788 5658 17816 5714
rect 17788 5630 18000 5658
rect 17972 5370 18000 5630
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18156 5234 18184 6938
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18420 6316 18472 6322
rect 18248 6276 18420 6304
rect 17776 5228 17828 5234
rect 17696 5188 17776 5216
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4321 17448 4558
rect 17604 4486 17632 4762
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17406 4312 17462 4321
rect 17406 4247 17462 4256
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17604 3602 17632 4218
rect 17696 4146 17724 5188
rect 17776 5170 17828 5176
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18248 4570 18276 6276
rect 18420 6258 18472 6264
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18432 5778 18460 6054
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18156 4542 18276 4570
rect 18340 4554 18368 5646
rect 18524 4690 18552 6666
rect 18708 6254 18736 6938
rect 19536 6882 19564 7142
rect 19352 6854 19564 6882
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18604 5908 18656 5914
rect 18708 5896 18736 6190
rect 18892 5914 18920 6598
rect 19076 6497 19104 6734
rect 19248 6724 19300 6730
rect 19352 6712 19380 6854
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19300 6684 19380 6712
rect 19248 6666 19300 6672
rect 19062 6488 19118 6497
rect 19444 6458 19472 6734
rect 19062 6423 19118 6432
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19076 6066 19104 6190
rect 18984 6038 19104 6066
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 18984 5914 19012 6038
rect 18656 5868 18736 5896
rect 18880 5908 18932 5914
rect 18604 5850 18656 5856
rect 18880 5850 18932 5856
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4548 18380 4554
rect 18156 4282 18184 4542
rect 18328 4490 18380 4496
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18326 4448 18382 4457
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17696 3194 17724 4082
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 18156 2990 18184 4218
rect 18248 4078 18276 4422
rect 18326 4383 18382 4392
rect 18340 4078 18368 4383
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18524 3466 18552 4490
rect 18694 3496 18750 3505
rect 18512 3460 18564 3466
rect 18694 3431 18696 3440
rect 18512 3402 18564 3408
rect 18748 3431 18750 3440
rect 18696 3402 18748 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3194 18644 3334
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18800 2650 18828 5170
rect 18892 4758 18920 5170
rect 18880 4752 18932 4758
rect 18880 4694 18932 4700
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18892 3602 18920 4218
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18984 3466 19012 5578
rect 19168 5522 19196 5782
rect 19076 5494 19196 5522
rect 19076 5302 19104 5494
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 19076 3058 19104 5238
rect 19246 5128 19302 5137
rect 19168 5086 19246 5114
rect 19168 4690 19196 5086
rect 19246 5063 19302 5072
rect 19352 5030 19380 6054
rect 19444 5302 19472 6258
rect 19536 6186 19564 6854
rect 19720 6254 19748 7262
rect 19996 7206 20024 7262
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19904 6934 19932 7142
rect 20088 6934 20116 7278
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 19892 6928 19944 6934
rect 20076 6928 20128 6934
rect 19892 6870 19944 6876
rect 19996 6876 20076 6882
rect 19996 6870 20128 6876
rect 19996 6854 20116 6870
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19522 5944 19578 5953
rect 19578 5888 19656 5896
rect 19522 5879 19656 5888
rect 19536 5868 19656 5879
rect 19522 5808 19578 5817
rect 19522 5743 19578 5752
rect 19536 5545 19564 5743
rect 19522 5536 19578 5545
rect 19522 5471 19578 5480
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19536 4758 19564 5471
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4282 19288 4626
rect 19340 4480 19392 4486
rect 19524 4480 19576 4486
rect 19340 4422 19392 4428
rect 19444 4440 19524 4468
rect 19352 4282 19380 4422
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19444 3618 19472 4440
rect 19524 4422 19576 4428
rect 19628 4434 19656 5868
rect 19720 5166 19748 6190
rect 19812 5166 19840 6734
rect 19996 6322 20024 6854
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20364 6746 20392 7142
rect 20456 6866 20484 7142
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20536 6792 20588 6798
rect 20364 6740 20536 6746
rect 20364 6734 20588 6740
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19904 5370 19932 6190
rect 20088 5914 20116 6734
rect 20364 6718 20576 6734
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5840 20036 5846
rect 20166 5808 20222 5817
rect 20036 5788 20166 5794
rect 19984 5782 20166 5788
rect 19996 5766 20166 5782
rect 20166 5743 20222 5752
rect 20272 5710 20300 6122
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20364 5778 20392 6054
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20456 5710 20484 6054
rect 19984 5704 20036 5710
rect 20260 5704 20312 5710
rect 20036 5664 20208 5692
rect 19984 5646 20036 5652
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19628 4406 19840 4434
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3942 19564 4082
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19536 3738 19564 3878
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19352 3590 19472 3618
rect 19154 3224 19210 3233
rect 19154 3159 19210 3168
rect 19168 3058 19196 3159
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 19352 2553 19380 3590
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 3346 19472 3402
rect 19616 3392 19668 3398
rect 19444 3340 19616 3346
rect 19444 3334 19668 3340
rect 19444 3318 19656 3334
rect 19444 3126 19472 3318
rect 19720 3194 19748 4218
rect 19812 3466 19840 4406
rect 19904 4282 19932 5170
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19996 4865 20024 5034
rect 19982 4856 20038 4865
rect 19982 4791 20038 4800
rect 20088 4690 20116 5170
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19904 3738 19932 4082
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20088 3602 20116 4082
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19996 3126 20024 3402
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19524 3052 19576 3058
rect 19576 3012 19840 3040
rect 19524 2994 19576 3000
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19338 2544 19394 2553
rect 19338 2479 19394 2488
rect 19536 2446 19564 2790
rect 16304 2382 16356 2388
rect 15396 2378 15608 2382
rect 15396 2372 15620 2378
rect 15396 2366 15568 2372
rect 15568 2314 15620 2320
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 14476 2158 14596 2186
rect 14184 2100 14236 2106
rect 14184 2042 14236 2048
rect 14476 1760 14504 2158
rect 15396 1760 15424 2246
rect 16316 1760 16344 2382
rect 17052 2366 17356 2394
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 17052 1834 17080 2366
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17040 1828 17092 1834
rect 17040 1770 17092 1776
rect 17236 1760 17264 2246
rect 17392 2032 17444 2038
rect 17392 1974 17444 1980
rect 17404 1834 17432 1974
rect 17392 1828 17444 1834
rect 17392 1770 17444 1776
rect 18156 1760 18184 2382
rect 19812 2378 19840 3012
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19800 2372 19852 2378
rect 19800 2314 19852 2320
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 1760 19104 2246
rect 19996 1760 20024 2382
rect 20180 2009 20208 5664
rect 20260 5646 20312 5652
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20260 5568 20312 5574
rect 20312 5528 20392 5556
rect 20260 5510 20312 5516
rect 20364 5166 20392 5528
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20272 4486 20300 5034
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20272 3602 20300 4218
rect 20364 4078 20392 4694
rect 20456 4214 20484 5170
rect 20548 4622 20576 6394
rect 20640 6322 20668 6938
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6390 20852 6598
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5914 20668 6258
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20720 5840 20772 5846
rect 20718 5808 20720 5817
rect 20772 5808 20774 5817
rect 20718 5743 20774 5752
rect 20732 5574 20760 5743
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20548 4146 20576 4558
rect 20640 4486 20668 4966
rect 20732 4826 20760 5034
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20718 4584 20774 4593
rect 20824 4554 20852 5306
rect 20916 5234 20944 7142
rect 21008 6866 21036 7142
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21100 6746 21128 6802
rect 21008 6718 21128 6746
rect 21180 6724 21232 6730
rect 21008 6118 21036 6718
rect 21180 6666 21232 6672
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21100 5914 21128 6598
rect 21192 5914 21220 6666
rect 21468 6458 21496 6938
rect 21652 6866 21680 7210
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21652 6458 21680 6802
rect 22756 6798 22784 7482
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22468 6792 22520 6798
rect 22190 6760 22246 6769
rect 22468 6734 22520 6740
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22190 6695 22192 6704
rect 22244 6695 22246 6704
rect 22192 6666 22244 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22388 6458 22416 6598
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21272 6180 21324 6186
rect 21272 6122 21324 6128
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20902 5128 20958 5137
rect 21008 5114 21036 5646
rect 20958 5086 21036 5114
rect 20902 5063 20958 5072
rect 21284 4622 21312 6122
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21468 5914 21496 6054
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21468 5370 21496 5578
rect 21560 5545 21588 5714
rect 21546 5536 21602 5545
rect 21546 5471 21602 5480
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21744 5234 21772 6190
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21454 4720 21510 4729
rect 21454 4655 21510 4664
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20718 4519 20774 4528
rect 20812 4548 20864 4554
rect 20732 4486 20760 4519
rect 20812 4490 20864 4496
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20916 4010 20944 4558
rect 21008 4146 21036 4558
rect 21284 4282 21312 4558
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 21008 3398 21036 4082
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21284 3398 21312 4014
rect 21376 3942 21404 4082
rect 21468 4010 21496 4655
rect 21560 4146 21588 4762
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21008 3233 21036 3334
rect 20994 3224 21050 3233
rect 20994 3159 21050 3168
rect 21376 3126 21404 3878
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21376 2582 21404 3062
rect 21468 2990 21496 3470
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 21652 2310 21680 5170
rect 22296 4826 22324 5170
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22204 4214 22232 4422
rect 22388 4282 22416 6394
rect 22480 5370 22508 6734
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22480 4554 22508 5306
rect 22572 5234 22600 6054
rect 22664 5250 22692 6598
rect 22742 6488 22798 6497
rect 22742 6423 22798 6432
rect 22756 6390 22784 6423
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22756 6118 22784 6326
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22848 5778 22876 6598
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22664 5222 22968 5250
rect 22572 4842 22600 5170
rect 22664 5030 22692 5222
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22572 4814 22692 4842
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21744 2774 21772 4082
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21836 3466 21864 4014
rect 22572 3738 22600 4694
rect 22664 4554 22692 4814
rect 22756 4622 22784 4966
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 21928 3126 21956 3334
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 22388 2990 22416 3334
rect 22664 3194 22692 3402
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 21744 2746 21956 2774
rect 21928 2650 21956 2746
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 22388 2446 22416 2926
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22376 2440 22428 2446
rect 22480 2417 22508 2858
rect 22848 2836 22876 5034
rect 22940 2990 22968 5222
rect 23032 4078 23060 7278
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23216 5574 23244 6734
rect 23308 6390 23336 6802
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23308 5710 23336 6054
rect 23400 5914 23428 6734
rect 23860 6458 23888 7754
rect 24030 7580 24086 7980
rect 26422 7984 26478 7993
rect 24308 7958 24360 7964
rect 24044 7478 24072 7580
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 24320 6322 24348 7958
rect 25778 7580 25834 7980
rect 26422 7919 26478 7928
rect 25792 7478 25820 7580
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 26436 7410 26464 7919
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26712 7449 26740 7482
rect 26698 7440 26754 7449
rect 26424 7404 26476 7410
rect 26698 7375 26754 7384
rect 26424 7346 26476 7352
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24504 7002 24532 7142
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23124 3194 23152 4694
rect 23216 4486 23244 5510
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23216 3194 23244 4422
rect 23308 4146 23336 5646
rect 23400 5098 23428 5850
rect 23676 5234 23704 6190
rect 23952 5302 23980 6190
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 23940 5296 23992 5302
rect 23940 5238 23992 5244
rect 24136 5234 24164 6054
rect 26238 5400 26294 5409
rect 26238 5335 26294 5344
rect 26252 5234 26280 5335
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23296 3052 23348 3058
rect 23032 3012 23296 3040
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 23032 2836 23060 3012
rect 23296 2994 23348 3000
rect 22848 2808 23060 2836
rect 22744 2576 22796 2582
rect 22744 2518 22796 2524
rect 22376 2382 22428 2388
rect 22466 2408 22522 2417
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 20916 1760 20944 2246
rect 21836 1760 21864 2382
rect 22466 2343 22522 2352
rect 22756 1760 22784 2518
rect 23032 2514 23060 2808
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22940 2310 22968 2382
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 23584 2194 23612 5034
rect 23676 3534 23704 5170
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 24044 4214 24072 4694
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 2990 23796 3334
rect 23860 3058 23888 3946
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 23848 2440 23900 2446
rect 23426 2166 23612 2194
rect 23676 2400 23848 2428
rect 23426 1970 23454 2166
rect 23412 1964 23464 1970
rect 23412 1906 23464 1912
rect 23676 1760 23704 2400
rect 23848 2382 23900 2388
rect 23952 2310 23980 2926
rect 24136 2774 24164 5170
rect 26344 5114 26372 7210
rect 26514 6896 26570 6905
rect 26514 6831 26570 6840
rect 26528 6798 26556 6831
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26424 6384 26476 6390
rect 26712 6361 26740 6598
rect 26424 6326 26476 6332
rect 26698 6352 26754 6361
rect 26252 5098 26372 5114
rect 26436 5098 26464 6326
rect 26698 6287 26754 6296
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 26712 5817 26740 6054
rect 26698 5808 26754 5817
rect 26698 5743 26754 5752
rect 26240 5092 26372 5098
rect 26292 5086 26372 5092
rect 26424 5092 26476 5098
rect 26240 5034 26292 5040
rect 26424 5034 26476 5040
rect 26332 5024 26384 5030
rect 26608 5024 26660 5030
rect 26332 4966 26384 4972
rect 26514 4992 26570 5001
rect 26344 4146 26372 4966
rect 26608 4966 26660 4972
rect 26514 4927 26570 4936
rect 26528 4604 26556 4927
rect 26620 4729 26648 4966
rect 26804 4865 26832 6734
rect 26896 5710 26924 7822
rect 27434 7712 27490 7721
rect 27434 7647 27490 7656
rect 27448 7546 27476 7647
rect 27526 7580 27582 7980
rect 27540 7546 27568 7580
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 27434 7168 27490 7177
rect 26988 7002 27016 7142
rect 27434 7103 27490 7112
rect 27448 7002 27476 7103
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27066 6896 27122 6905
rect 27066 6831 27122 6840
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 26988 5273 27016 6734
rect 27080 6662 27108 6831
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 27434 6624 27490 6633
rect 27434 6559 27490 6568
rect 27448 6458 27476 6559
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27434 6080 27490 6089
rect 27434 6015 27490 6024
rect 27448 5914 27476 6015
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27252 5704 27304 5710
rect 27250 5672 27252 5681
rect 27304 5672 27306 5681
rect 27250 5607 27306 5616
rect 27068 5568 27120 5574
rect 27066 5536 27068 5545
rect 27120 5536 27122 5545
rect 27066 5471 27122 5480
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27448 5273 27476 5306
rect 26974 5264 27030 5273
rect 27434 5264 27490 5273
rect 27252 5228 27304 5234
rect 26974 5199 27030 5208
rect 27172 5188 27252 5216
rect 26790 4856 26846 4865
rect 26790 4791 26846 4800
rect 26606 4720 26662 4729
rect 26606 4655 26662 4664
rect 26608 4616 26660 4622
rect 26528 4576 26608 4604
rect 26608 4558 26660 4564
rect 26792 4480 26844 4486
rect 27068 4480 27120 4486
rect 26792 4422 26844 4428
rect 27066 4448 27068 4457
rect 27120 4448 27122 4457
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 25976 3777 26004 4082
rect 26252 4049 26280 4082
rect 26238 4040 26294 4049
rect 26238 3975 26294 3984
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26712 3777 26740 3878
rect 25962 3768 26018 3777
rect 25962 3703 26018 3712
rect 26698 3768 26754 3777
rect 26698 3703 26754 3712
rect 26606 3632 26662 3641
rect 26606 3567 26662 3576
rect 26620 3534 26648 3567
rect 26804 3534 26832 4422
rect 27066 4383 27122 4392
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24044 2746 24164 2774
rect 24044 2650 24072 2746
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24504 2582 24532 2994
rect 24584 2848 24636 2854
rect 24636 2796 24716 2802
rect 24584 2790 24716 2796
rect 24596 2774 24716 2790
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24688 2446 24716 2774
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24596 1760 24624 2246
rect 24872 2038 24900 3470
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25424 2428 25452 3062
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25516 2650 25544 2994
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 25596 2440 25648 2446
rect 25424 2400 25596 2428
rect 25596 2382 25648 2388
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 25516 1760 25544 2246
rect 25884 2009 25912 2790
rect 26068 2553 26096 2790
rect 26054 2544 26110 2553
rect 26054 2479 26110 2488
rect 26160 2446 26188 3334
rect 26344 2689 26372 3470
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 26436 3194 26464 3334
rect 26712 3194 26740 3334
rect 26896 3194 26924 3946
rect 26988 3913 27016 4082
rect 27068 3936 27120 3942
rect 26974 3904 27030 3913
rect 27068 3878 27120 3884
rect 26974 3839 27030 3848
rect 27080 3738 27108 3878
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 27068 3392 27120 3398
rect 27066 3360 27068 3369
rect 27120 3360 27122 3369
rect 27066 3295 27122 3304
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26700 3188 26752 3194
rect 26700 3130 26752 3136
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 26974 3088 27030 3097
rect 26974 3023 26976 3032
rect 27028 3023 27030 3032
rect 26976 2994 27028 3000
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26330 2680 26386 2689
rect 26330 2615 26386 2624
rect 26620 2446 26648 2858
rect 26700 2848 26752 2854
rect 26698 2816 26700 2825
rect 26752 2816 26754 2825
rect 26698 2751 26754 2760
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 26332 2304 26384 2310
rect 26330 2272 26332 2281
rect 26384 2272 26386 2281
rect 26330 2207 26386 2216
rect 25870 2000 25926 2009
rect 25870 1935 25926 1944
rect 26436 1760 26464 2314
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27080 1760 27108 2246
rect 27172 2214 27200 5188
rect 27434 5199 27490 5208
rect 27252 5170 27304 5176
rect 27434 4992 27490 5001
rect 27434 4927 27490 4936
rect 27448 4826 27476 4927
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27172 2186 27234 2214
rect 27206 2106 27234 2186
rect 27264 2187 27292 4558
rect 27434 4176 27490 4185
rect 27434 4111 27490 4120
rect 27448 4010 27476 4111
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27434 3904 27490 3913
rect 27434 3839 27490 3848
rect 27448 3738 27476 3839
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27448 3097 27476 3130
rect 27434 3088 27490 3097
rect 27434 3023 27490 3032
rect 27827 2372 27879 2378
rect 27827 2314 27879 2320
rect 27264 2159 27332 2187
rect 27200 2100 27252 2106
rect 27200 2042 27252 2048
rect 27304 1902 27332 2159
rect 27292 1896 27344 1902
rect 27292 1838 27344 1844
rect 27839 1760 27867 2314
rect 1040 1360 1096 1760
rect 1582 1360 1638 1760
rect 2502 1360 2558 1760
rect 3422 1360 3478 1760
rect 4342 1360 4398 1760
rect 5262 1360 5318 1760
rect 5632 1702 5684 1708
rect 6182 1360 6238 1760
rect 7102 1360 7158 1760
rect 8022 1360 8078 1760
rect 8942 1360 8998 1760
rect 9862 1360 9918 1760
rect 10782 1360 10838 1760
rect 11702 1360 11758 1760
rect 12622 1360 12678 1760
rect 13542 1360 13598 1760
rect 14462 1360 14518 1760
rect 15382 1360 15438 1760
rect 16302 1360 16358 1760
rect 17222 1360 17278 1760
rect 18142 1360 18198 1760
rect 19062 1360 19118 1760
rect 19982 1360 20038 1760
rect 20902 1360 20958 1760
rect 21822 1360 21878 1760
rect 22742 1360 22798 1760
rect 23662 1360 23718 1760
rect 24582 1360 24638 1760
rect 25502 1360 25558 1760
rect 26422 1360 26478 1760
rect 27066 1360 27122 1760
rect 27825 1360 27881 1760
<< via2 >>
rect 1122 7928 1178 7984
rect 1030 7656 1086 7712
rect 1490 7112 1546 7168
rect 1858 7384 1914 7440
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2410 6840 2466 6896
rect 954 6568 1010 6624
rect 1122 6296 1178 6352
rect 2042 6316 2098 6352
rect 2042 6296 2044 6316
rect 2044 6296 2096 6316
rect 2096 6296 2098 6316
rect 1038 6024 1094 6080
rect 954 5788 956 5808
rect 956 5788 1008 5808
rect 1008 5788 1010 5808
rect 954 5752 1010 5788
rect 1674 5752 1730 5808
rect 1858 5516 1860 5536
rect 1860 5516 1912 5536
rect 1912 5516 1914 5536
rect 1858 5480 1914 5516
rect 954 5208 1010 5264
rect 1038 4972 1040 4992
rect 1040 4972 1092 4992
rect 1092 4972 1094 4992
rect 1038 4936 1094 4972
rect 954 4700 956 4720
rect 956 4700 1008 4720
rect 1008 4700 1010 4720
rect 954 4664 1010 4700
rect 1038 4428 1040 4448
rect 1040 4428 1092 4448
rect 1092 4428 1094 4448
rect 1038 4392 1094 4428
rect 1490 4120 1546 4176
rect 1038 3884 1040 3904
rect 1040 3884 1092 3904
rect 1092 3884 1094 3904
rect 1038 3848 1094 3884
rect 954 3612 956 3632
rect 956 3612 1008 3632
rect 1008 3612 1010 3632
rect 954 3576 1010 3612
rect 2318 4664 2374 4720
rect 2134 4528 2190 4584
rect 1038 3340 1040 3360
rect 1040 3340 1092 3360
rect 1092 3340 1094 3360
rect 1038 3304 1094 3340
rect 2594 5228 2650 5264
rect 2594 5208 2596 5228
rect 2596 5208 2648 5228
rect 2648 5208 2650 5228
rect 2594 5072 2650 5128
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 2410 4120 2466 4176
rect 2318 3984 2374 4040
rect 954 3032 1010 3088
rect 1038 2796 1040 2816
rect 1040 2796 1092 2816
rect 1092 2796 1094 2816
rect 1038 2760 1094 2796
rect 2226 2624 2282 2680
rect 2226 2488 2282 2544
rect 1214 2216 1270 2272
rect 1766 2372 1822 2408
rect 1766 2352 1768 2372
rect 1768 2352 1820 2372
rect 1820 2352 1822 2372
rect 1306 1944 1362 2000
rect 3238 3440 3294 3496
rect 2870 2896 2926 2952
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3576 4306 3632
rect 5262 4936 5318 4992
rect 5906 6196 5908 6216
rect 5908 6196 5960 6216
rect 5960 6196 5962 6216
rect 5906 6160 5962 6196
rect 5906 5636 5962 5672
rect 5906 5616 5908 5636
rect 5908 5616 5960 5636
rect 5960 5616 5962 5636
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 5262 3712 5318 3768
rect 4618 3032 4674 3088
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3974 1944 4030 2000
rect 6182 4392 6238 4448
rect 6550 5908 6606 5944
rect 6550 5888 6552 5908
rect 6552 5888 6604 5908
rect 6604 5888 6606 5908
rect 6458 3576 6514 3632
rect 6642 4936 6698 4992
rect 7102 5652 7104 5672
rect 7104 5652 7156 5672
rect 7156 5652 7158 5672
rect 7102 5616 7158 5652
rect 7286 4428 7288 4448
rect 7288 4428 7340 4448
rect 7340 4428 7342 4448
rect 7286 4392 7342 4428
rect 6918 3848 6974 3904
rect 6734 3168 6790 3224
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 7286 3576 7342 3632
rect 7654 4276 7710 4312
rect 7654 4256 7656 4276
rect 7656 4256 7708 4276
rect 7708 4256 7710 4276
rect 8298 5888 8354 5944
rect 9218 6024 9274 6080
rect 8206 3848 8262 3904
rect 10230 5888 10286 5944
rect 9586 4256 9642 4312
rect 9310 3576 9366 3632
rect 10782 5752 10838 5808
rect 9586 3168 9642 3224
rect 10690 4936 10746 4992
rect 12990 6840 13046 6896
rect 11150 6724 11206 6760
rect 11150 6704 11152 6724
rect 11152 6704 11204 6724
rect 11204 6704 11206 6724
rect 11702 6704 11758 6760
rect 11334 6296 11390 6352
rect 10874 4800 10930 4856
rect 10598 3168 10654 3224
rect 11978 6060 11980 6080
rect 11980 6060 12032 6080
rect 12032 6060 12034 6080
rect 11426 4936 11482 4992
rect 11978 6024 12034 6060
rect 13726 6724 13782 6760
rect 13726 6704 13728 6724
rect 13728 6704 13780 6724
rect 13780 6704 13782 6724
rect 11334 3848 11390 3904
rect 11978 4392 12034 4448
rect 11518 2760 11574 2816
rect 13174 6160 13230 6216
rect 12898 5772 12954 5808
rect 12898 5752 12900 5772
rect 12900 5752 12952 5772
rect 12952 5752 12954 5772
rect 12254 3984 12310 4040
rect 12162 3848 12218 3904
rect 12806 3596 12862 3632
rect 12806 3576 12808 3596
rect 12808 3576 12860 3596
rect 12860 3576 12862 3596
rect 13174 4120 13230 4176
rect 13726 5480 13782 5536
rect 14002 4120 14058 4176
rect 14002 3848 14058 3904
rect 14462 6160 14518 6216
rect 14554 5344 14610 5400
rect 15014 5616 15070 5672
rect 14922 4800 14978 4856
rect 14922 3712 14978 3768
rect 15382 6840 15438 6896
rect 15842 6840 15898 6896
rect 15750 6160 15806 6216
rect 15014 3576 15070 3632
rect 16394 5888 16450 5944
rect 16394 5364 16450 5400
rect 16394 5344 16396 5364
rect 16396 5344 16448 5364
rect 16448 5344 16450 5364
rect 14646 2896 14702 2952
rect 14922 2760 14978 2816
rect 16762 4936 16818 4992
rect 17314 5344 17370 5400
rect 17498 5228 17554 5264
rect 17498 5208 17500 5228
rect 17500 5208 17552 5228
rect 17552 5208 17554 5228
rect 17406 4256 17462 4312
rect 19062 6432 19118 6488
rect 18326 4392 18382 4448
rect 18694 3460 18750 3496
rect 18694 3440 18696 3460
rect 18696 3440 18748 3460
rect 18748 3440 18750 3460
rect 19246 5072 19302 5128
rect 19522 5888 19578 5944
rect 19522 5752 19578 5808
rect 19522 5480 19578 5536
rect 20166 5752 20222 5808
rect 19154 3168 19210 3224
rect 19982 4800 20038 4856
rect 19338 2488 19394 2544
rect 20718 5788 20720 5808
rect 20720 5788 20772 5808
rect 20772 5788 20774 5808
rect 20718 5752 20774 5788
rect 20718 4528 20774 4584
rect 22190 6724 22246 6760
rect 22190 6704 22192 6724
rect 22192 6704 22244 6724
rect 22244 6704 22246 6724
rect 20902 5072 20958 5128
rect 21546 5480 21602 5536
rect 21454 4664 21510 4720
rect 20994 3168 21050 3224
rect 22742 6432 22798 6488
rect 26422 7928 26478 7984
rect 26698 7384 26754 7440
rect 26238 5344 26294 5400
rect 20166 1944 20222 2000
rect 22466 2352 22522 2408
rect 26514 6840 26570 6896
rect 26698 6296 26754 6352
rect 26698 5752 26754 5808
rect 26514 4936 26570 4992
rect 27434 7656 27490 7712
rect 27434 7112 27490 7168
rect 27066 6840 27122 6896
rect 27434 6568 27490 6624
rect 27434 6024 27490 6080
rect 27250 5652 27252 5672
rect 27252 5652 27304 5672
rect 27304 5652 27306 5672
rect 27250 5616 27306 5652
rect 27066 5516 27068 5536
rect 27068 5516 27120 5536
rect 27120 5516 27122 5536
rect 27066 5480 27122 5516
rect 26974 5208 27030 5264
rect 26790 4800 26846 4856
rect 26606 4664 26662 4720
rect 27066 4428 27068 4448
rect 27068 4428 27120 4448
rect 27120 4428 27122 4448
rect 26238 3984 26294 4040
rect 25962 3712 26018 3768
rect 26698 3712 26754 3768
rect 26606 3576 26662 3632
rect 27066 4392 27122 4428
rect 26054 2488 26110 2544
rect 26974 3848 27030 3904
rect 27066 3340 27068 3360
rect 27068 3340 27120 3360
rect 27120 3340 27122 3360
rect 27066 3304 27122 3340
rect 26974 3052 27030 3088
rect 26974 3032 26976 3052
rect 26976 3032 27028 3052
rect 27028 3032 27030 3052
rect 26330 2624 26386 2680
rect 26698 2796 26700 2816
rect 26700 2796 26752 2816
rect 26752 2796 26754 2816
rect 26698 2760 26754 2796
rect 26330 2252 26332 2272
rect 26332 2252 26384 2272
rect 26384 2252 26386 2272
rect 26330 2216 26386 2252
rect 25870 1944 25926 2000
rect 27434 5208 27490 5264
rect 27434 4936 27490 4992
rect 27434 4120 27490 4176
rect 27434 3848 27490 3904
rect 27434 3032 27490 3088
<< metal3 >>
rect 480 7986 880 8016
rect 1117 7986 1183 7989
rect 480 7984 1183 7986
rect 480 7928 1122 7984
rect 1178 7928 1183 7984
rect 480 7926 1183 7928
rect 480 7896 880 7926
rect 1117 7923 1183 7926
rect 26417 7986 26483 7989
rect 28077 7986 28477 8016
rect 26417 7984 28477 7986
rect 26417 7928 26422 7984
rect 26478 7928 28477 7984
rect 26417 7926 28477 7928
rect 26417 7923 26483 7926
rect 28077 7896 28477 7926
rect 480 7714 880 7744
rect 1025 7714 1091 7717
rect 480 7712 1091 7714
rect 480 7656 1030 7712
rect 1086 7656 1091 7712
rect 480 7654 1091 7656
rect 480 7624 880 7654
rect 1025 7651 1091 7654
rect 27429 7714 27495 7717
rect 28077 7714 28477 7744
rect 27429 7712 28477 7714
rect 27429 7656 27434 7712
rect 27490 7656 28477 7712
rect 27429 7654 28477 7656
rect 27429 7651 27495 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 28077 7624 28477 7654
rect 4870 7583 5186 7584
rect 480 7442 880 7472
rect 1853 7442 1919 7445
rect 480 7440 1919 7442
rect 480 7384 1858 7440
rect 1914 7384 1919 7440
rect 480 7382 1919 7384
rect 480 7352 880 7382
rect 1853 7379 1919 7382
rect 26693 7442 26759 7445
rect 28077 7442 28477 7472
rect 26693 7440 28477 7442
rect 26693 7384 26698 7440
rect 26754 7384 28477 7440
rect 26693 7382 28477 7384
rect 26693 7379 26759 7382
rect 28077 7352 28477 7382
rect 480 7170 880 7200
rect 1485 7170 1551 7173
rect 480 7168 1551 7170
rect 480 7112 1490 7168
rect 1546 7112 1551 7168
rect 480 7110 1551 7112
rect 480 7080 880 7110
rect 1485 7107 1551 7110
rect 27429 7170 27495 7173
rect 28077 7170 28477 7200
rect 27429 7168 28477 7170
rect 27429 7112 27434 7168
rect 27490 7112 28477 7168
rect 27429 7110 28477 7112
rect 27429 7107 27495 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 28077 7080 28477 7110
rect 4210 7039 4526 7040
rect 480 6898 880 6928
rect 2405 6898 2471 6901
rect 480 6896 2471 6898
rect 480 6840 2410 6896
rect 2466 6840 2471 6896
rect 480 6838 2471 6840
rect 480 6808 880 6838
rect 2405 6835 2471 6838
rect 12985 6898 13051 6901
rect 15377 6898 15443 6901
rect 12985 6896 15443 6898
rect 12985 6840 12990 6896
rect 13046 6840 15382 6896
rect 15438 6840 15443 6896
rect 12985 6838 15443 6840
rect 12985 6835 13051 6838
rect 15377 6835 15443 6838
rect 15837 6898 15903 6901
rect 26509 6898 26575 6901
rect 15837 6896 26575 6898
rect 15837 6840 15842 6896
rect 15898 6840 26514 6896
rect 26570 6840 26575 6896
rect 15837 6838 26575 6840
rect 15837 6835 15903 6838
rect 26509 6835 26575 6838
rect 27061 6898 27127 6901
rect 28077 6898 28477 6928
rect 27061 6896 28477 6898
rect 27061 6840 27066 6896
rect 27122 6840 28477 6896
rect 27061 6838 28477 6840
rect 27061 6835 27127 6838
rect 28077 6808 28477 6838
rect 11145 6762 11211 6765
rect 11697 6762 11763 6765
rect 13721 6762 13787 6765
rect 22185 6762 22251 6765
rect 11145 6760 22251 6762
rect 11145 6704 11150 6760
rect 11206 6704 11702 6760
rect 11758 6704 13726 6760
rect 13782 6704 22190 6760
rect 22246 6704 22251 6760
rect 11145 6702 22251 6704
rect 11145 6699 11211 6702
rect 11697 6699 11763 6702
rect 13721 6699 13787 6702
rect 22185 6699 22251 6702
rect 480 6626 880 6656
rect 949 6626 1015 6629
rect 480 6624 1015 6626
rect 480 6568 954 6624
rect 1010 6568 1015 6624
rect 480 6566 1015 6568
rect 480 6536 880 6566
rect 949 6563 1015 6566
rect 27429 6626 27495 6629
rect 28077 6626 28477 6656
rect 27429 6624 28477 6626
rect 27429 6568 27434 6624
rect 27490 6568 28477 6624
rect 27429 6566 28477 6568
rect 27429 6563 27495 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 28077 6536 28477 6566
rect 4870 6495 5186 6496
rect 19057 6490 19123 6493
rect 22737 6490 22803 6493
rect 19057 6488 22803 6490
rect 19057 6432 19062 6488
rect 19118 6432 22742 6488
rect 22798 6432 22803 6488
rect 19057 6430 22803 6432
rect 19057 6427 19123 6430
rect 22737 6427 22803 6430
rect 480 6354 880 6384
rect 1117 6354 1183 6357
rect 480 6352 1183 6354
rect 480 6296 1122 6352
rect 1178 6296 1183 6352
rect 480 6294 1183 6296
rect 480 6264 880 6294
rect 1117 6291 1183 6294
rect 2037 6354 2103 6357
rect 11329 6354 11395 6357
rect 2037 6352 11395 6354
rect 2037 6296 2042 6352
rect 2098 6296 11334 6352
rect 11390 6296 11395 6352
rect 2037 6294 11395 6296
rect 2037 6291 2103 6294
rect 11329 6291 11395 6294
rect 26693 6354 26759 6357
rect 28077 6354 28477 6384
rect 26693 6352 28477 6354
rect 26693 6296 26698 6352
rect 26754 6296 28477 6352
rect 26693 6294 28477 6296
rect 26693 6291 26759 6294
rect 28077 6264 28477 6294
rect 5901 6218 5967 6221
rect 13169 6218 13235 6221
rect 5901 6216 13235 6218
rect 5901 6160 5906 6216
rect 5962 6160 13174 6216
rect 13230 6160 13235 6216
rect 5901 6158 13235 6160
rect 5901 6155 5967 6158
rect 13169 6155 13235 6158
rect 14457 6218 14523 6221
rect 15745 6218 15811 6221
rect 14457 6216 15811 6218
rect 14457 6160 14462 6216
rect 14518 6160 15750 6216
rect 15806 6160 15811 6216
rect 14457 6158 15811 6160
rect 14457 6155 14523 6158
rect 15745 6155 15811 6158
rect 480 6082 880 6112
rect 1033 6082 1099 6085
rect 480 6080 1099 6082
rect 480 6024 1038 6080
rect 1094 6024 1099 6080
rect 480 6022 1099 6024
rect 480 5992 880 6022
rect 1033 6019 1099 6022
rect 9213 6082 9279 6085
rect 11973 6082 12039 6085
rect 9213 6080 12039 6082
rect 9213 6024 9218 6080
rect 9274 6024 11978 6080
rect 12034 6024 12039 6080
rect 9213 6022 12039 6024
rect 9213 6019 9279 6022
rect 11973 6019 12039 6022
rect 27429 6082 27495 6085
rect 28077 6082 28477 6112
rect 27429 6080 28477 6082
rect 27429 6024 27434 6080
rect 27490 6024 28477 6080
rect 27429 6022 28477 6024
rect 27429 6019 27495 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 28077 5992 28477 6022
rect 4210 5951 4526 5952
rect 6545 5946 6611 5949
rect 8293 5946 8359 5949
rect 10225 5946 10291 5949
rect 6545 5944 10291 5946
rect 6545 5888 6550 5944
rect 6606 5888 8298 5944
rect 8354 5888 10230 5944
rect 10286 5888 10291 5944
rect 6545 5886 10291 5888
rect 6545 5883 6611 5886
rect 8293 5883 8359 5886
rect 10225 5883 10291 5886
rect 16389 5946 16455 5949
rect 19517 5946 19583 5949
rect 16389 5944 19583 5946
rect 16389 5888 16394 5944
rect 16450 5888 19522 5944
rect 19578 5888 19583 5944
rect 16389 5886 19583 5888
rect 16389 5883 16455 5886
rect 19517 5883 19583 5886
rect 480 5810 880 5840
rect 949 5810 1015 5813
rect 480 5808 1015 5810
rect 480 5752 954 5808
rect 1010 5752 1015 5808
rect 480 5750 1015 5752
rect 480 5720 880 5750
rect 949 5747 1015 5750
rect 1669 5810 1735 5813
rect 10777 5810 10843 5813
rect 12893 5810 12959 5813
rect 19517 5810 19583 5813
rect 1669 5808 12450 5810
rect 1669 5752 1674 5808
rect 1730 5752 10782 5808
rect 10838 5752 12450 5808
rect 1669 5750 12450 5752
rect 1669 5747 1735 5750
rect 10777 5747 10843 5750
rect 5901 5674 5967 5677
rect 7097 5674 7163 5677
rect 5901 5672 7163 5674
rect 5901 5616 5906 5672
rect 5962 5616 7102 5672
rect 7158 5616 7163 5672
rect 5901 5614 7163 5616
rect 12390 5674 12450 5750
rect 12893 5808 19583 5810
rect 12893 5752 12898 5808
rect 12954 5752 19522 5808
rect 19578 5752 19583 5808
rect 12893 5750 19583 5752
rect 12893 5747 12959 5750
rect 19517 5747 19583 5750
rect 20161 5810 20227 5813
rect 20713 5810 20779 5813
rect 20161 5808 20779 5810
rect 20161 5752 20166 5808
rect 20222 5752 20718 5808
rect 20774 5752 20779 5808
rect 20161 5750 20779 5752
rect 20161 5747 20227 5750
rect 20713 5747 20779 5750
rect 26693 5810 26759 5813
rect 28077 5810 28477 5840
rect 26693 5808 28477 5810
rect 26693 5752 26698 5808
rect 26754 5752 28477 5808
rect 26693 5750 28477 5752
rect 26693 5747 26759 5750
rect 28077 5720 28477 5750
rect 15009 5674 15075 5677
rect 27245 5674 27311 5677
rect 12390 5672 15075 5674
rect 12390 5616 15014 5672
rect 15070 5616 15075 5672
rect 12390 5614 15075 5616
rect 5901 5611 5967 5614
rect 7097 5611 7163 5614
rect 15009 5611 15075 5614
rect 15150 5672 27311 5674
rect 15150 5616 27250 5672
rect 27306 5616 27311 5672
rect 15150 5614 27311 5616
rect 480 5538 880 5568
rect 1853 5538 1919 5541
rect 480 5536 1919 5538
rect 480 5480 1858 5536
rect 1914 5480 1919 5536
rect 480 5478 1919 5480
rect 480 5448 880 5478
rect 1853 5475 1919 5478
rect 13721 5538 13787 5541
rect 15150 5538 15210 5614
rect 27245 5611 27311 5614
rect 13721 5536 15210 5538
rect 13721 5480 13726 5536
rect 13782 5480 15210 5536
rect 13721 5478 15210 5480
rect 19517 5538 19583 5541
rect 21541 5538 21607 5541
rect 19517 5536 21607 5538
rect 19517 5480 19522 5536
rect 19578 5480 21546 5536
rect 21602 5480 21607 5536
rect 19517 5478 21607 5480
rect 13721 5475 13787 5478
rect 19517 5475 19583 5478
rect 21541 5475 21607 5478
rect 27061 5538 27127 5541
rect 28077 5538 28477 5568
rect 27061 5536 28477 5538
rect 27061 5480 27066 5536
rect 27122 5480 28477 5536
rect 27061 5478 28477 5480
rect 27061 5475 27127 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 28077 5448 28477 5478
rect 4870 5407 5186 5408
rect 14549 5402 14615 5405
rect 16389 5402 16455 5405
rect 14549 5400 16455 5402
rect 14549 5344 14554 5400
rect 14610 5344 16394 5400
rect 16450 5344 16455 5400
rect 14549 5342 16455 5344
rect 14549 5339 14615 5342
rect 16389 5339 16455 5342
rect 17309 5402 17375 5405
rect 26233 5402 26299 5405
rect 17309 5400 26299 5402
rect 17309 5344 17314 5400
rect 17370 5344 26238 5400
rect 26294 5344 26299 5400
rect 17309 5342 26299 5344
rect 17309 5339 17375 5342
rect 26233 5339 26299 5342
rect 480 5266 880 5296
rect 949 5266 1015 5269
rect 480 5264 1015 5266
rect 480 5208 954 5264
rect 1010 5208 1015 5264
rect 480 5206 1015 5208
rect 480 5176 880 5206
rect 949 5203 1015 5206
rect 2589 5266 2655 5269
rect 17493 5266 17559 5269
rect 26969 5266 27035 5269
rect 2589 5264 27035 5266
rect 2589 5208 2594 5264
rect 2650 5208 17498 5264
rect 17554 5208 26974 5264
rect 27030 5208 27035 5264
rect 2589 5206 27035 5208
rect 2589 5203 2655 5206
rect 17493 5203 17559 5206
rect 26969 5203 27035 5206
rect 27429 5266 27495 5269
rect 28077 5266 28477 5296
rect 27429 5264 28477 5266
rect 27429 5208 27434 5264
rect 27490 5208 28477 5264
rect 27429 5206 28477 5208
rect 27429 5203 27495 5206
rect 28077 5176 28477 5206
rect 2589 5130 2655 5133
rect 19241 5130 19307 5133
rect 20897 5130 20963 5133
rect 2589 5128 12450 5130
rect 2589 5072 2594 5128
rect 2650 5072 12450 5128
rect 2589 5070 12450 5072
rect 2589 5067 2655 5070
rect 480 4994 880 5024
rect 1033 4994 1099 4997
rect 480 4992 1099 4994
rect 480 4936 1038 4992
rect 1094 4936 1099 4992
rect 480 4934 1099 4936
rect 480 4904 880 4934
rect 1033 4931 1099 4934
rect 5257 4994 5323 4997
rect 6637 4994 6703 4997
rect 5257 4992 6703 4994
rect 5257 4936 5262 4992
rect 5318 4936 6642 4992
rect 6698 4936 6703 4992
rect 5257 4934 6703 4936
rect 5257 4931 5323 4934
rect 6637 4931 6703 4934
rect 10685 4994 10751 4997
rect 11421 4994 11487 4997
rect 10685 4992 11487 4994
rect 10685 4936 10690 4992
rect 10746 4936 11426 4992
rect 11482 4936 11487 4992
rect 10685 4934 11487 4936
rect 12390 4994 12450 5070
rect 19241 5128 20963 5130
rect 19241 5072 19246 5128
rect 19302 5072 20902 5128
rect 20958 5072 20963 5128
rect 19241 5070 20963 5072
rect 19241 5067 19307 5070
rect 20897 5067 20963 5070
rect 16757 4994 16823 4997
rect 26509 4994 26575 4997
rect 12390 4992 26575 4994
rect 12390 4936 16762 4992
rect 16818 4936 26514 4992
rect 26570 4936 26575 4992
rect 12390 4934 26575 4936
rect 10685 4931 10751 4934
rect 11421 4931 11487 4934
rect 16757 4931 16823 4934
rect 26509 4931 26575 4934
rect 27429 4994 27495 4997
rect 28077 4994 28477 5024
rect 27429 4992 28477 4994
rect 27429 4936 27434 4992
rect 27490 4936 28477 4992
rect 27429 4934 28477 4936
rect 27429 4931 27495 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 28077 4904 28477 4934
rect 4210 4863 4526 4864
rect 10869 4858 10935 4861
rect 14917 4858 14983 4861
rect 10869 4856 14983 4858
rect 10869 4800 10874 4856
rect 10930 4800 14922 4856
rect 14978 4800 14983 4856
rect 10869 4798 14983 4800
rect 10869 4795 10935 4798
rect 14917 4795 14983 4798
rect 19977 4858 20043 4861
rect 26785 4858 26851 4861
rect 19977 4856 26851 4858
rect 19977 4800 19982 4856
rect 20038 4800 26790 4856
rect 26846 4800 26851 4856
rect 19977 4798 26851 4800
rect 19977 4795 20043 4798
rect 26785 4795 26851 4798
rect 480 4722 880 4752
rect 949 4722 1015 4725
rect 480 4720 1015 4722
rect 480 4664 954 4720
rect 1010 4664 1015 4720
rect 480 4662 1015 4664
rect 480 4632 880 4662
rect 949 4659 1015 4662
rect 2313 4722 2379 4725
rect 21449 4722 21515 4725
rect 2313 4720 21515 4722
rect 2313 4664 2318 4720
rect 2374 4664 21454 4720
rect 21510 4664 21515 4720
rect 2313 4662 21515 4664
rect 2313 4659 2379 4662
rect 21449 4659 21515 4662
rect 26601 4722 26667 4725
rect 28077 4722 28477 4752
rect 26601 4720 28477 4722
rect 26601 4664 26606 4720
rect 26662 4664 28477 4720
rect 26601 4662 28477 4664
rect 26601 4659 26667 4662
rect 28077 4632 28477 4662
rect 2129 4586 2195 4589
rect 20713 4586 20779 4589
rect 2129 4584 20779 4586
rect 2129 4528 2134 4584
rect 2190 4528 20718 4584
rect 20774 4528 20779 4584
rect 2129 4526 20779 4528
rect 2129 4523 2195 4526
rect 20713 4523 20779 4526
rect 480 4450 880 4480
rect 1033 4450 1099 4453
rect 480 4448 1099 4450
rect 480 4392 1038 4448
rect 1094 4392 1099 4448
rect 480 4390 1099 4392
rect 480 4360 880 4390
rect 1033 4387 1099 4390
rect 6177 4450 6243 4453
rect 7281 4450 7347 4453
rect 6177 4448 7347 4450
rect 6177 4392 6182 4448
rect 6238 4392 7286 4448
rect 7342 4392 7347 4448
rect 6177 4390 7347 4392
rect 6177 4387 6243 4390
rect 7281 4387 7347 4390
rect 11973 4450 12039 4453
rect 18321 4450 18387 4453
rect 11973 4448 18387 4450
rect 11973 4392 11978 4448
rect 12034 4392 18326 4448
rect 18382 4392 18387 4448
rect 11973 4390 18387 4392
rect 11973 4387 12039 4390
rect 18321 4387 18387 4390
rect 27061 4450 27127 4453
rect 28077 4450 28477 4480
rect 27061 4448 28477 4450
rect 27061 4392 27066 4448
rect 27122 4392 28477 4448
rect 27061 4390 28477 4392
rect 27061 4387 27127 4390
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 28077 4360 28477 4390
rect 4870 4319 5186 4320
rect 7649 4314 7715 4317
rect 8150 4314 8156 4316
rect 7649 4312 8156 4314
rect 7649 4256 7654 4312
rect 7710 4256 8156 4312
rect 7649 4254 8156 4256
rect 7649 4251 7715 4254
rect 8150 4252 8156 4254
rect 8220 4252 8226 4316
rect 9581 4314 9647 4317
rect 17401 4314 17467 4317
rect 9581 4312 17467 4314
rect 9581 4256 9586 4312
rect 9642 4256 17406 4312
rect 17462 4256 17467 4312
rect 9581 4254 17467 4256
rect 9581 4251 9647 4254
rect 17401 4251 17467 4254
rect 480 4178 880 4208
rect 1485 4178 1551 4181
rect 480 4176 1551 4178
rect 480 4120 1490 4176
rect 1546 4120 1551 4176
rect 480 4118 1551 4120
rect 480 4088 880 4118
rect 1485 4115 1551 4118
rect 2405 4178 2471 4181
rect 13169 4178 13235 4181
rect 13997 4178 14063 4181
rect 2405 4176 14063 4178
rect 2405 4120 2410 4176
rect 2466 4120 13174 4176
rect 13230 4120 14002 4176
rect 14058 4120 14063 4176
rect 2405 4118 14063 4120
rect 2405 4115 2471 4118
rect 13169 4115 13235 4118
rect 13997 4115 14063 4118
rect 27429 4178 27495 4181
rect 28077 4178 28477 4208
rect 27429 4176 28477 4178
rect 27429 4120 27434 4176
rect 27490 4120 28477 4176
rect 27429 4118 28477 4120
rect 27429 4115 27495 4118
rect 28077 4088 28477 4118
rect 2313 4042 2379 4045
rect 12249 4042 12315 4045
rect 26233 4042 26299 4045
rect 2313 4040 12315 4042
rect 2313 3984 2318 4040
rect 2374 3984 12254 4040
rect 12310 3984 12315 4040
rect 2313 3982 12315 3984
rect 2313 3979 2379 3982
rect 12249 3979 12315 3982
rect 12390 4040 26299 4042
rect 12390 3984 26238 4040
rect 26294 3984 26299 4040
rect 12390 3982 26299 3984
rect 480 3906 880 3936
rect 1033 3906 1099 3909
rect 480 3904 1099 3906
rect 480 3848 1038 3904
rect 1094 3848 1099 3904
rect 480 3846 1099 3848
rect 480 3816 880 3846
rect 1033 3843 1099 3846
rect 6913 3906 6979 3909
rect 8201 3906 8267 3909
rect 6913 3904 8267 3906
rect 6913 3848 6918 3904
rect 6974 3848 8206 3904
rect 8262 3848 8267 3904
rect 6913 3846 8267 3848
rect 6913 3843 6979 3846
rect 8201 3843 8267 3846
rect 11329 3906 11395 3909
rect 12157 3906 12223 3909
rect 12390 3906 12450 3982
rect 26233 3979 26299 3982
rect 11329 3904 12450 3906
rect 11329 3848 11334 3904
rect 11390 3848 12162 3904
rect 12218 3848 12450 3904
rect 11329 3846 12450 3848
rect 13997 3906 14063 3909
rect 26969 3906 27035 3909
rect 13997 3904 27035 3906
rect 13997 3848 14002 3904
rect 14058 3848 26974 3904
rect 27030 3848 27035 3904
rect 13997 3846 27035 3848
rect 11329 3843 11395 3846
rect 12157 3843 12223 3846
rect 13997 3843 14063 3846
rect 26969 3843 27035 3846
rect 27429 3906 27495 3909
rect 28077 3906 28477 3936
rect 27429 3904 28477 3906
rect 27429 3848 27434 3904
rect 27490 3848 28477 3904
rect 27429 3846 28477 3848
rect 27429 3843 27495 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 28077 3816 28477 3846
rect 4210 3775 4526 3776
rect 5257 3770 5323 3773
rect 14917 3770 14983 3773
rect 25957 3770 26023 3773
rect 5257 3768 12450 3770
rect 5257 3712 5262 3768
rect 5318 3712 12450 3768
rect 5257 3710 12450 3712
rect 5257 3707 5323 3710
rect 480 3634 880 3664
rect 949 3634 1015 3637
rect 480 3632 1015 3634
rect 480 3576 954 3632
rect 1010 3576 1015 3632
rect 480 3574 1015 3576
rect 480 3544 880 3574
rect 949 3571 1015 3574
rect 4245 3634 4311 3637
rect 6453 3634 6519 3637
rect 4245 3632 6519 3634
rect 4245 3576 4250 3632
rect 4306 3576 6458 3632
rect 6514 3576 6519 3632
rect 4245 3574 6519 3576
rect 4245 3571 4311 3574
rect 6453 3571 6519 3574
rect 7281 3634 7347 3637
rect 9305 3634 9371 3637
rect 7281 3632 9371 3634
rect 7281 3576 7286 3632
rect 7342 3576 9310 3632
rect 9366 3576 9371 3632
rect 7281 3574 9371 3576
rect 12390 3634 12450 3710
rect 14917 3768 26023 3770
rect 14917 3712 14922 3768
rect 14978 3712 25962 3768
rect 26018 3712 26023 3768
rect 14917 3710 26023 3712
rect 14917 3707 14983 3710
rect 25957 3707 26023 3710
rect 26693 3770 26759 3773
rect 26693 3768 27722 3770
rect 26693 3712 26698 3768
rect 26754 3712 27722 3768
rect 26693 3710 27722 3712
rect 26693 3707 26759 3710
rect 12801 3634 12867 3637
rect 12390 3632 12867 3634
rect 12390 3576 12806 3632
rect 12862 3576 12867 3632
rect 12390 3574 12867 3576
rect 7281 3571 7347 3574
rect 9305 3571 9371 3574
rect 12801 3571 12867 3574
rect 15009 3634 15075 3637
rect 26601 3634 26667 3637
rect 15009 3632 26667 3634
rect 15009 3576 15014 3632
rect 15070 3576 26606 3632
rect 26662 3576 26667 3632
rect 15009 3574 26667 3576
rect 27662 3634 27722 3710
rect 28077 3634 28477 3664
rect 27662 3574 28477 3634
rect 15009 3571 15075 3574
rect 26601 3571 26667 3574
rect 28077 3544 28477 3574
rect 3233 3498 3299 3501
rect 18689 3498 18755 3501
rect 3233 3496 18755 3498
rect 3233 3440 3238 3496
rect 3294 3440 18694 3496
rect 18750 3440 18755 3496
rect 3233 3438 18755 3440
rect 3233 3435 3299 3438
rect 18689 3435 18755 3438
rect 480 3362 880 3392
rect 1033 3362 1099 3365
rect 480 3360 1099 3362
rect 480 3304 1038 3360
rect 1094 3304 1099 3360
rect 480 3302 1099 3304
rect 480 3272 880 3302
rect 1033 3299 1099 3302
rect 27061 3362 27127 3365
rect 28077 3362 28477 3392
rect 27061 3360 28477 3362
rect 27061 3304 27066 3360
rect 27122 3304 28477 3360
rect 27061 3302 28477 3304
rect 27061 3299 27127 3302
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 28077 3272 28477 3302
rect 4870 3231 5186 3232
rect 6729 3226 6795 3229
rect 9581 3226 9647 3229
rect 6729 3224 9647 3226
rect 6729 3168 6734 3224
rect 6790 3168 9586 3224
rect 9642 3168 9647 3224
rect 6729 3166 9647 3168
rect 6729 3163 6795 3166
rect 9581 3163 9647 3166
rect 10593 3226 10659 3229
rect 19149 3226 19215 3229
rect 20989 3226 21055 3229
rect 10593 3224 21055 3226
rect 10593 3168 10598 3224
rect 10654 3168 19154 3224
rect 19210 3168 20994 3224
rect 21050 3168 21055 3224
rect 10593 3166 21055 3168
rect 10593 3163 10659 3166
rect 19149 3163 19215 3166
rect 20989 3163 21055 3166
rect 480 3090 880 3120
rect 949 3090 1015 3093
rect 480 3088 1015 3090
rect 480 3032 954 3088
rect 1010 3032 1015 3088
rect 480 3030 1015 3032
rect 480 3000 880 3030
rect 949 3027 1015 3030
rect 4613 3090 4679 3093
rect 26969 3090 27035 3093
rect 4613 3088 27035 3090
rect 4613 3032 4618 3088
rect 4674 3032 26974 3088
rect 27030 3032 27035 3088
rect 4613 3030 27035 3032
rect 4613 3027 4679 3030
rect 26969 3027 27035 3030
rect 27429 3090 27495 3093
rect 28077 3090 28477 3120
rect 27429 3088 28477 3090
rect 27429 3032 27434 3088
rect 27490 3032 28477 3088
rect 27429 3030 28477 3032
rect 27429 3027 27495 3030
rect 28077 3000 28477 3030
rect 2865 2954 2931 2957
rect 14641 2954 14707 2957
rect 2865 2952 14707 2954
rect 2865 2896 2870 2952
rect 2926 2896 14646 2952
rect 14702 2896 14707 2952
rect 2865 2894 14707 2896
rect 2865 2891 2931 2894
rect 14641 2891 14707 2894
rect 480 2818 880 2848
rect 1033 2818 1099 2821
rect 480 2816 1099 2818
rect 480 2760 1038 2816
rect 1094 2760 1099 2816
rect 480 2758 1099 2760
rect 480 2728 880 2758
rect 1033 2755 1099 2758
rect 11513 2818 11579 2821
rect 14917 2818 14983 2821
rect 11513 2816 14983 2818
rect 11513 2760 11518 2816
rect 11574 2760 14922 2816
rect 14978 2760 14983 2816
rect 11513 2758 14983 2760
rect 11513 2755 11579 2758
rect 14917 2755 14983 2758
rect 26693 2818 26759 2821
rect 28077 2818 28477 2848
rect 26693 2816 28477 2818
rect 26693 2760 26698 2816
rect 26754 2760 28477 2816
rect 26693 2758 28477 2760
rect 26693 2755 26759 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 28077 2728 28477 2758
rect 4210 2687 4526 2688
rect 2221 2682 2287 2685
rect 1166 2680 2287 2682
rect 1166 2624 2226 2680
rect 2282 2624 2287 2680
rect 1166 2622 2287 2624
rect 480 2546 880 2576
rect 1166 2546 1226 2622
rect 2221 2619 2287 2622
rect 8150 2620 8156 2684
rect 8220 2682 8226 2684
rect 26325 2682 26391 2685
rect 8220 2680 26391 2682
rect 8220 2624 26330 2680
rect 26386 2624 26391 2680
rect 8220 2622 26391 2624
rect 8220 2620 8226 2622
rect 26325 2619 26391 2622
rect 480 2486 1226 2546
rect 2221 2546 2287 2549
rect 19333 2546 19399 2549
rect 2221 2544 19399 2546
rect 2221 2488 2226 2544
rect 2282 2488 19338 2544
rect 19394 2488 19399 2544
rect 2221 2486 19399 2488
rect 480 2456 880 2486
rect 2221 2483 2287 2486
rect 19333 2483 19399 2486
rect 26049 2546 26115 2549
rect 28077 2546 28477 2576
rect 26049 2544 28477 2546
rect 26049 2488 26054 2544
rect 26110 2488 28477 2544
rect 26049 2486 28477 2488
rect 26049 2483 26115 2486
rect 28077 2456 28477 2486
rect 1761 2410 1827 2413
rect 22461 2410 22527 2413
rect 1761 2408 22527 2410
rect 1761 2352 1766 2408
rect 1822 2352 22466 2408
rect 22522 2352 22527 2408
rect 1761 2350 22527 2352
rect 1761 2347 1827 2350
rect 22461 2347 22527 2350
rect 480 2274 880 2304
rect 1209 2274 1275 2277
rect 480 2272 1275 2274
rect 480 2216 1214 2272
rect 1270 2216 1275 2272
rect 480 2214 1275 2216
rect 480 2184 880 2214
rect 1209 2211 1275 2214
rect 26325 2274 26391 2277
rect 28077 2274 28477 2304
rect 26325 2272 28477 2274
rect 26325 2216 26330 2272
rect 26386 2216 28477 2272
rect 26325 2214 28477 2216
rect 26325 2211 26391 2214
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 28077 2184 28477 2214
rect 4870 2143 5186 2144
rect 480 2002 880 2032
rect 1301 2002 1367 2005
rect 480 2000 1367 2002
rect 480 1944 1306 2000
rect 1362 1944 1367 2000
rect 480 1942 1367 1944
rect 480 1912 880 1942
rect 1301 1939 1367 1942
rect 3969 2002 4035 2005
rect 20161 2002 20227 2005
rect 3969 2000 20227 2002
rect 3969 1944 3974 2000
rect 4030 1944 20166 2000
rect 20222 1944 20227 2000
rect 3969 1942 20227 1944
rect 3969 1939 4035 1942
rect 20161 1939 20227 1942
rect 25865 2002 25931 2005
rect 28077 2002 28477 2032
rect 25865 2000 28477 2002
rect 25865 1944 25870 2000
rect 25926 1944 28477 2000
rect 25865 1942 28477 1944
rect 25865 1939 25931 1942
rect 28077 1912 28477 1942
<< via3 >>
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 8156 4252 8220 4316
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 8156 2620 8220 2684
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 7104 4528 7664
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 7648 5188 7664
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 8155 4316 8221 4317
rect 8155 4252 8156 4316
rect 8220 4252 8221 4316
rect 8155 4251 8221 4252
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 8158 2685 8218 4251
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1710522493
transform 1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1710522493
transform -1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1710522493
transform -1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1710522493
transform -1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1710522493
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 22908 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _096_
timestamp 1710522493
transform 1 0 22172 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 21620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 17480 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _099_
timestamp 1710522493
transform 1 0 17204 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19044 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19412 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 23092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _103_
timestamp 1710522493
transform -1 0 20700 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 21344 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 20976 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _106_
timestamp 1710522493
transform -1 0 20884 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _108_
timestamp 1710522493
transform -1 0 21528 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 21252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 18492 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _112_
timestamp 1710522493
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 23184 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 17296 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _117_
timestamp 1710522493
transform 1 0 17204 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _118_
timestamp 1710522493
transform 1 0 10764 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _119_
timestamp 1710522493
transform -1 0 18584 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 22172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1710522493
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1710522493
transform -1 0 5888 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1710522493
transform -1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 1710522493
transform 1 0 6440 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1710522493
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1710522493
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1710522493
transform -1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1710522493
transform 1 0 10120 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1710522493
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1710522493
transform 1 0 11224 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp 1710522493
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5704 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1710522493
transform 1 0 24472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _136_
timestamp 1710522493
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 1710522493
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _138_
timestamp 1710522493
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 1710522493
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 1710522493
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _141_
timestamp 1710522493
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1710522493
transform -1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _143_
timestamp 1710522493
transform -1 0 17296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _144_
timestamp 1710522493
transform -1 0 19596 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _145_
timestamp 1710522493
transform -1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1710522493
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 23000 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _148_
timestamp 1710522493
transform 1 0 24012 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 5336 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1710522493
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _151_
timestamp 1710522493
transform 1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1710522493
transform 1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _153_
timestamp 1710522493
transform 1 0 7452 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1710522493
transform 1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1710522493
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _157_
timestamp 1710522493
transform -1 0 12604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1710522493
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _159_
timestamp 1710522493
transform 1 0 12972 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1710522493
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _161_
timestamp 1710522493
transform 1 0 14720 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1710522493
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _163_
timestamp 1710522493
transform 1 0 16560 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1710522493
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _165_
timestamp 1710522493
transform 1 0 17020 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1710522493
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _167_
timestamp 1710522493
transform 1 0 20700 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1710522493
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _169_
timestamp 1710522493
transform 1 0 23644 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1710522493
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 5612 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1710522493
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _173_
timestamp 1710522493
transform -1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1710522493
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _175_
timestamp 1710522493
transform -1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1710522493
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _177_
timestamp 1710522493
transform 1 0 9660 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1710522493
transform -1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _179_
timestamp 1710522493
transform 1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1710522493
transform -1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _181_
timestamp 1710522493
transform -1 0 13892 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1710522493
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _183_
timestamp 1710522493
transform -1 0 15456 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1710522493
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _185_
timestamp 1710522493
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1710522493
transform -1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _187_
timestamp 1710522493
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1710522493
transform -1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _189_
timestamp 1710522493
transform -1 0 21712 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1710522493
transform -1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _191_
timestamp 1710522493
transform -1 0 24012 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1710522493
transform -1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _193_
timestamp 1710522493
transform -1 0 20884 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _194_
timestamp 1710522493
transform 1 0 23276 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 22356 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1710522493
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _197_
timestamp 1710522493
transform 1 0 3864 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 13248 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _199_
timestamp 1710522493
transform -1 0 12512 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 1710522493
transform 1 0 11776 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _201_
timestamp 1710522493
transform -1 0 6256 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1710522493
transform 1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1710522493
transform 1 0 4784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _204_
timestamp 1710522493
transform -1 0 6532 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1710522493
transform 1 0 4048 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1710522493
transform 1 0 4508 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _207_
timestamp 1710522493
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _208_
timestamp 1710522493
transform 1 0 10948 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1710522493
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 7360 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _211_
timestamp 1710522493
transform 1 0 6900 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _212_
timestamp 1710522493
transform -1 0 7544 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _213_
timestamp 1710522493
transform 1 0 8924 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _214_
timestamp 1710522493
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _215_
timestamp 1710522493
transform -1 0 11408 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _216_
timestamp 1710522493
transform -1 0 12236 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _217_
timestamp 1710522493
transform 1 0 14260 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _218_
timestamp 1710522493
transform 1 0 15456 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _219_
timestamp 1710522493
transform 1 0 16652 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _220_
timestamp 1710522493
transform -1 0 20332 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _221_
timestamp 1710522493
transform -1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 7544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _223_
timestamp 1710522493
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _225_
timestamp 1710522493
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _226_
timestamp 1710522493
transform -1 0 6256 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1710522493
transform -1 0 6716 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1710522493
transform 1 0 3956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 19688 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1710522493
transform 1 0 15916 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _231_
timestamp 1710522493
transform -1 0 19688 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp 1710522493
transform -1 0 19320 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1710522493
transform -1 0 19136 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _234_
timestamp 1710522493
transform -1 0 17296 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _235_
timestamp 1710522493
transform 1 0 14352 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1710522493
transform 1 0 14812 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _237_
timestamp 1710522493
transform -1 0 16284 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp 1710522493
transform -1 0 15088 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1710522493
transform -1 0 14352 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _240_
timestamp 1710522493
transform -1 0 14812 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _241_
timestamp 1710522493
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1710522493
transform 1 0 13432 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 1710522493
transform 1 0 3864 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 1710522493
transform 1 0 3588 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 1710522493
transform 1 0 21896 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 1710522493
transform -1 0 23644 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 21988 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 1710522493
transform -1 0 11776 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _250_
timestamp 1710522493
transform 1 0 4140 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _251_
timestamp 1710522493
transform 1 0 7544 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _252_
timestamp 1710522493
transform 1 0 6716 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _253_
timestamp 1710522493
transform 1 0 9108 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _254_
timestamp 1710522493
transform 1 0 7544 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 1710522493
transform 1 0 10212 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _256_
timestamp 1710522493
transform 1 0 11500 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _257_
timestamp 1710522493
transform 1 0 14444 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _258_
timestamp 1710522493
transform 1 0 15640 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _259_
timestamp 1710522493
transform 1 0 16652 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _260_
timestamp 1710522493
transform 1 0 19596 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _261_
timestamp 1710522493
transform 1 0 21896 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _262_
timestamp 1710522493
transform 1 0 5704 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _263_
timestamp 1710522493
transform 1 0 8004 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _264_
timestamp 1710522493
transform 1 0 3588 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1710522493
transform -1 0 16008 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1710522493
transform 1 0 19228 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _267_
timestamp 1710522493
transform 1 0 14352 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _268_
timestamp 1710522493
transform 1 0 14076 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 1710522493
transform -1 0 14720 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 1710522493
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout98 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 1710522493
transform -1 0 16560 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 1710522493
transform -1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 1710522493
transform -1 0 13156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp 1710522493
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 1710522493
transform -1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 1710522493
transform -1 0 15732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 1710522493
transform -1 0 11224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 1710522493
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout107
timestamp 1710522493
transform -1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 1710522493
transform -1 0 13984 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_52
timestamp 1710522493
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_70
timestamp 1710522493
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1710522493
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1710522493
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_89 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_95
timestamp 1710522493
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_100
timestamp 1710522493
transform 1 0 10304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1710522493
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1710522493
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_120
timestamp 1710522493
transform 1 0 12144 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_129
timestamp 1710522493
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_135
timestamp 1710522493
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1710522493
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_150
timestamp 1710522493
transform 1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_155
timestamp 1710522493
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_163
timestamp 1710522493
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1710522493
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_172
timestamp 1710522493
transform 1 0 16928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_180
timestamp 1710522493
transform 1 0 17664 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp 1710522493
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1710522493
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_201
timestamp 1710522493
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1710522493
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_209
timestamp 1710522493
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_220
timestamp 1710522493
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_225
timestamp 1710522493
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_229
timestamp 1710522493
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_233
timestamp 1710522493
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_237
timestamp 1710522493
transform 1 0 22908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1710522493
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1710522493
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_260
timestamp 1710522493
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_270
timestamp 1710522493
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_281
timestamp 1710522493
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_21
timestamp 1710522493
transform 1 0 3036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_47
timestamp 1710522493
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_60
timestamp 1710522493
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_96 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 9936 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_104
timestamp 1710522493
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1710522493
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_124
timestamp 1710522493
transform 1 0 12512 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_130
timestamp 1710522493
transform 1 0 13064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_143
timestamp 1710522493
transform 1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_192
timestamp 1710522493
transform 1 0 18768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_225
timestamp 1710522493
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_257
timestamp 1710522493
transform 1 0 24748 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1710522493
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1710522493
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1710522493
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_110
timestamp 1710522493
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_146
timestamp 1710522493
transform 1 0 14536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_156
timestamp 1710522493
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_185
timestamp 1710522493
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_217
timestamp 1710522493
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1710522493
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_259
timestamp 1710522493
transform 1 0 24932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_20
timestamp 1710522493
transform 1 0 2944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_28
timestamp 1710522493
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_66
timestamp 1710522493
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_92
timestamp 1710522493
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_100
timestamp 1710522493
transform 1 0 10304 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_104
timestamp 1710522493
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_120
timestamp 1710522493
transform 1 0 12144 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_155
timestamp 1710522493
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_163
timestamp 1710522493
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1710522493
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_190
timestamp 1710522493
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_209
timestamp 1710522493
transform 1 0 20332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1710522493
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_250
timestamp 1710522493
transform 1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_262
timestamp 1710522493
transform 1 0 25208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_17
timestamp 1710522493
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1710522493
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1710522493
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_41
timestamp 1710522493
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_59
timestamp 1710522493
transform 1 0 6532 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_68
timestamp 1710522493
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1710522493
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_94
timestamp 1710522493
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_98
timestamp 1710522493
transform 1 0 10120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_125
timestamp 1710522493
transform 1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1710522493
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1710522493
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_149
timestamp 1710522493
transform 1 0 14812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_161
timestamp 1710522493
transform 1 0 15916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_167
timestamp 1710522493
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_182
timestamp 1710522493
transform 1 0 17848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1710522493
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_205
timestamp 1710522493
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_220
timestamp 1710522493
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_224
timestamp 1710522493
transform 1 0 21712 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_239
timestamp 1710522493
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1710522493
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1710522493
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_265
timestamp 1710522493
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_273
timestamp 1710522493
transform 1 0 26220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_20
timestamp 1710522493
transform 1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_28
timestamp 1710522493
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_64
timestamp 1710522493
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_72
timestamp 1710522493
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_129
timestamp 1710522493
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_139
timestamp 1710522493
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_143
timestamp 1710522493
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1710522493
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_187
timestamp 1710522493
transform 1 0 18308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_215
timestamp 1710522493
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1710522493
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1710522493
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1710522493
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1710522493
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_11
timestamp 1710522493
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_23
timestamp 1710522493
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1710522493
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1710522493
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_94
timestamp 1710522493
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_132
timestamp 1710522493
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_170
timestamp 1710522493
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_174
timestamp 1710522493
transform 1 0 17112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_205
timestamp 1710522493
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_222
timestamp 1710522493
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_246
timestamp 1710522493
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1710522493
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1710522493
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_277
timestamp 1710522493
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_11
timestamp 1710522493
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_23
timestamp 1710522493
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1710522493
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_67
timestamp 1710522493
transform 1 0 7268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_107
timestamp 1710522493
transform 1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_133
timestamp 1710522493
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_176
timestamp 1710522493
transform 1 0 17296 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_209
timestamp 1710522493
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1710522493
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_252
timestamp 1710522493
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_264
timestamp 1710522493
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_281
timestamp 1710522493
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1710522493
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1710522493
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_62
timestamp 1710522493
transform 1 0 6808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_74
timestamp 1710522493
transform 1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1710522493
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_95
timestamp 1710522493
transform 1 0 9844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_100
timestamp 1710522493
transform 1 0 10304 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_124
timestamp 1710522493
transform 1 0 12512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_131
timestamp 1710522493
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_135
timestamp 1710522493
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1710522493
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_168
timestamp 1710522493
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_172
timestamp 1710522493
transform 1 0 16928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_180
timestamp 1710522493
transform 1 0 17664 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_188
timestamp 1710522493
transform 1 0 18400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1710522493
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_219
timestamp 1710522493
transform 1 0 21252 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_227
timestamp 1710522493
transform 1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1710522493
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1710522493
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1710522493
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_265
timestamp 1710522493
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_273
timestamp 1710522493
transform 1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_20
timestamp 1710522493
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 1710522493
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 1710522493
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1710522493
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_66
timestamp 1710522493
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_78
timestamp 1710522493
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_91
timestamp 1710522493
transform 1 0 9476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_97
timestamp 1710522493
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1710522493
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_116
timestamp 1710522493
transform 1 0 11776 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_123
timestamp 1710522493
transform 1 0 12420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_135
timestamp 1710522493
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_139
timestamp 1710522493
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_152
timestamp 1710522493
transform 1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 1710522493
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_169
timestamp 1710522493
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_173
timestamp 1710522493
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_177
timestamp 1710522493
transform 1 0 17388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_189
timestamp 1710522493
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_197
timestamp 1710522493
transform 1 0 19228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_211
timestamp 1710522493
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_215
timestamp 1710522493
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1710522493
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_225
timestamp 1710522493
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_235
timestamp 1710522493
transform 1 0 22724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_247
timestamp 1710522493
transform 1 0 23828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_251
timestamp 1710522493
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_257
timestamp 1710522493
transform 1 0 24748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_272
timestamp 1710522493
transform 1 0 26128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1710522493
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1710522493
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1710522493
transform -1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1710522493
transform -1 0 24748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1710522493
transform -1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1710522493
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1710522493
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1710522493
transform -1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1710522493
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1710522493
transform -1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1710522493
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1710522493
transform -1 0 24104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1710522493
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1710522493
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1710522493
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1710522493
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1710522493
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1710522493
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1710522493
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1710522493
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1710522493
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1710522493
transform -1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1710522493
transform -1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1710522493
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1710522493
transform -1 0 3680 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1710522493
transform -1 0 5428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1710522493
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1710522493
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1710522493
transform 1 0 10120 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1710522493
transform 1 0 11868 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1710522493
transform -1 0 14628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1710522493
transform -1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1710522493
transform 1 0 27048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1710522493
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1710522493
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1710522493
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1710522493
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1710522493
transform -1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1710522493
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1710522493
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1710522493
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1710522493
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1710522493
transform -1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1710522493
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1710522493
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1710522493
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1710522493
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1710522493
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1710522493
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1710522493
transform 1 0 27232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1710522493
transform 1 0 27232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1710522493
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1710522493
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1710522493
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1710522493
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1710522493
transform 1 0 27232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1710522493
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1710522493
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1710522493
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1710522493
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1710522493
transform -1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1710522493
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1710522493
transform -1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1710522493
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1710522493
transform -1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1710522493
transform -1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1710522493
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1710522493
transform -1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1710522493
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1710522493
transform -1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1710522493
transform -1 0 26128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1710522493
transform -1 0 26864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1710522493
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1710522493
transform -1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1710522493
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1710522493
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1710522493
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1710522493
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1710522493
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1710522493
transform 1 0 27232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1710522493
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1710522493
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1710522493
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1710522493
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1710522493
transform -1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1710522493
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1710522493
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1710522493
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1710522493
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1710522493
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1710522493
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1710522493
transform -1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 1710522493
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1710522493
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 1710522493
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1710522493
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 1710522493
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1710522493
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 1710522493
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1710522493
transform -1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 1710522493
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1710522493
transform -1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 1710522493
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1710522493
transform -1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 1710522493
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1710522493
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 1710522493
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1710522493
transform -1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 1710522493
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1710522493
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 1710522493
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1710522493
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1710522493
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22
timestamp 1710522493
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1710522493
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp 1710522493
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 1710522493
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 1710522493
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp 1710522493
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp 1710522493
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 1710522493
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 1710522493
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_31
timestamp 1710522493
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_32
timestamp 1710522493
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_33
timestamp 1710522493
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_34
timestamp 1710522493
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_35
timestamp 1710522493
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1710522493
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1710522493
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1710522493
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1710522493
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1710522493
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_41
timestamp 1710522493
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 1710522493
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_43
timestamp 1710522493
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_44
timestamp 1710522493
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_45
timestamp 1710522493
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_46
timestamp 1710522493
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_47
timestamp 1710522493
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_48
timestamp 1710522493
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_49
timestamp 1710522493
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_50
timestamp 1710522493
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_51
timestamp 1710522493
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp 1710522493
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp 1710522493
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 1710522493
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 1710522493
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 1710522493
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1710522493
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_58
timestamp 1710522493
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_59
timestamp 1710522493
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_60
timestamp 1710522493
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_61
timestamp 1710522493
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1710522493
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1710522493
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_64
timestamp 1710522493
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 1710522493
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_66
timestamp 1710522493
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_67
timestamp 1710522493
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_68
timestamp 1710522493
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_69
timestamp 1710522493
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_70
timestamp 1710522493
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_71
timestamp 1710522493
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_72
timestamp 1710522493
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_73
timestamp 1710522493
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_74
timestamp 1710522493
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp 1710522493
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_76
timestamp 1710522493
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_77
timestamp 1710522493
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_78
timestamp 1710522493
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_79
timestamp 1710522493
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 4208 2128 4528 7664 0 FreeSans 1920 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4868 2128 5188 7664 0 FreeSans 1920 90 0 0 VSS
port 1 nsew ground bidirectional
rlabel metal1 14490 7072 14490 7072 0 VDD
rlabel metal1 14490 7616 14490 7616 0 VSS
rlabel metal1 22908 6766 22908 6766 0 _000_
rlabel metal2 11822 6052 11822 6052 0 _001_
rlabel metal1 4508 5338 4508 5338 0 _002_
rlabel metal1 3910 6392 3910 6392 0 _003_
rlabel metal1 11500 5338 11500 5338 0 _004_
rlabel metal1 4968 3570 4968 3570 0 _005_
rlabel metal1 7682 3094 7682 3094 0 _006_
rlabel metal1 6992 2618 6992 2618 0 _007_
rlabel metal1 9476 3570 9476 3570 0 _008_
rlabel metal1 8096 5882 8096 5882 0 _009_
rlabel metal1 10672 3162 10672 3162 0 _010_
rlabel metal1 11684 2890 11684 2890 0 _011_
rlabel metal1 14812 2618 14812 2618 0 _012_
rlabel metal1 16001 3706 16001 3706 0 _013_
rlabel metal1 17112 3094 17112 3094 0 _014_
rlabel metal1 19918 3128 19918 3128 0 _015_
rlabel metal1 22034 3570 22034 3570 0 _016_
rlabel metal1 6210 5338 6210 5338 0 _017_
rlabel metal1 8464 5270 8464 5270 0 _018_
rlabel metal1 3949 2822 3949 2822 0 _019_
rlabel metal1 15824 5882 15824 5882 0 _020_
rlabel metal1 19550 3400 19550 3400 0 _021_
rlabel metal1 14766 5338 14766 5338 0 _022_
rlabel metal2 14398 5916 14398 5916 0 _023_
rlabel metal1 13662 3162 13662 3162 0 _024_
rlabel via1 9886 6290 9886 6290 0 _025_
rlabel metal2 10534 6562 10534 6562 0 _026_
rlabel metal1 22448 4590 22448 4590 0 _027_
rlabel metal1 19422 5712 19422 5712 0 _028_
rlabel metal1 20286 5610 20286 5610 0 _029_
rlabel metal1 23230 3026 23230 3026 0 _030_
rlabel metal1 21022 6732 21022 6732 0 _031_
rlabel metal1 20010 6868 20010 6868 0 _032_
rlabel metal1 22448 4998 22448 4998 0 _033_
rlabel metal2 21482 5984 21482 5984 0 _034_
rlabel metal1 19412 4998 19412 4998 0 _035_
rlabel metal1 19044 5882 19044 5882 0 _036_
rlabel metal1 19780 5338 19780 5338 0 _037_
rlabel metal2 19458 6596 19458 6596 0 _038_
rlabel metal1 18906 4080 18906 4080 0 _039_
rlabel metal1 19964 4590 19964 4590 0 _040_
rlabel metal2 20470 5882 20470 5882 0 _041_
rlabel metal1 21022 5882 21022 5882 0 _042_
rlabel metal1 20930 5338 20930 5338 0 _043_
rlabel metal1 21114 5814 21114 5814 0 _044_
rlabel metal1 19550 6732 19550 6732 0 _045_
rlabel metal1 19274 5712 19274 5712 0 _046_
rlabel metal1 20010 5882 20010 5882 0 _047_
rlabel metal2 20470 7004 20470 7004 0 _048_
rlabel metal1 19504 6834 19504 6834 0 _049_
rlabel metal1 18032 4114 18032 4114 0 _050_
rlabel metal2 18262 4250 18262 4250 0 _051_
rlabel metal2 18354 4233 18354 4233 0 _052_
rlabel metal1 19458 3978 19458 3978 0 _053_
rlabel metal1 10810 5168 10810 5168 0 _054_
rlabel metal1 5106 6426 5106 6426 0 _055_
rlabel metal1 5750 4794 5750 4794 0 _056_
rlabel metal1 6532 6426 6532 6426 0 _057_
rlabel metal1 8740 5882 8740 5882 0 _058_
rlabel metal1 10120 5338 10120 5338 0 _059_
rlabel metal1 11408 6970 11408 6970 0 _060_
rlabel metal1 20930 2380 20930 2380 0 _061_
rlabel metal2 20102 3842 20102 3842 0 _062_
rlabel metal1 5060 4998 5060 4998 0 _063_
rlabel metal1 12558 5746 12558 5746 0 _064_
rlabel metal1 12190 5746 12190 5746 0 _065_
rlabel metal1 5566 5134 5566 5134 0 _066_
rlabel metal1 5014 5134 5014 5134 0 _067_
rlabel metal1 5750 4726 5750 4726 0 _068_
rlabel metal1 4738 6698 4738 6698 0 _069_
rlabel metal2 12098 4692 12098 4692 0 _070_
rlabel metal1 11684 5134 11684 5134 0 _071_
rlabel metal2 6854 5372 6854 5372 0 _072_
rlabel metal1 9568 6426 9568 6426 0 _073_
rlabel metal1 5152 4046 5152 4046 0 _074_
rlabel metal1 5566 3706 5566 3706 0 _075_
rlabel metal1 19642 5270 19642 5270 0 _076_
rlabel metal1 18722 3570 18722 3570 0 _077_
rlabel metal1 18768 3162 18768 3162 0 _078_
rlabel metal2 15410 5610 15410 5610 0 _079_
rlabel metal1 15042 5134 15042 5134 0 _080_
rlabel metal1 14996 5066 14996 5066 0 _081_
rlabel metal1 14260 6426 14260 6426 0 _082_
rlabel metal1 14168 2958 14168 2958 0 _083_
rlabel metal1 14030 3162 14030 3162 0 _084_
rlabel metal2 23322 6596 23322 6596 0 _085_
rlabel metal2 22218 4318 22218 4318 0 _086_
rlabel metal1 17204 7378 17204 7378 0 clk
rlabel metal2 3450 1384 3450 1384 0 comp_n
rlabel via1 7304 4590 7304 4590 0 counter\[0\]
rlabel metal1 21068 2550 21068 2550 0 counter\[10\]
rlabel metal1 21436 3502 21436 3502 0 counter\[11\]
rlabel metal2 17434 4437 17434 4437 0 counter\[1\]
rlabel metal2 7498 2587 7498 2587 0 counter\[2\]
rlabel metal1 7728 2414 7728 2414 0 counter\[3\]
rlabel metal1 9246 4080 9246 4080 0 counter\[4\]
rlabel metal1 11638 4794 11638 4794 0 counter\[5\]
rlabel metal1 13662 5236 13662 5236 0 counter\[6\]
rlabel metal1 17940 4250 17940 4250 0 counter\[7\]
rlabel metal1 17066 2482 17066 2482 0 counter\[8\]
rlabel metal1 19366 3060 19366 3060 0 counter\[9\]
rlabel metal1 23552 5882 23552 5882 0 counter_sample
rlabel metal1 22448 7446 22448 7446 0 debug_mux[0]
rlabel metal1 24334 7446 24334 7446 0 debug_mux[1]
rlabel metal1 26082 7412 26082 7412 0 debug_mux[2]
rlabel metal1 27186 7412 27186 7412 0 debug_mux[3]
rlabel metal1 20608 7378 20608 7378 0 en_offset_cal
rlabel metal1 14122 6766 14122 6766 0 net1
rlabel metal1 15686 7446 15686 7446 0 net10
rlabel metal2 19090 4148 19090 4148 0 net100
rlabel metal1 12926 6365 12926 6365 0 net101
rlabel metal1 13800 3706 13800 3706 0 net102
rlabel metal1 16330 6766 16330 6766 0 net103
rlabel metal1 15456 7174 15456 7174 0 net104
rlabel metal1 11546 6324 11546 6324 0 net105
rlabel metal1 21114 5678 21114 5678 0 net106
rlabel metal1 19274 3468 19274 3468 0 net107
rlabel metal1 13708 6698 13708 6698 0 net108
rlabel metal2 22770 7140 22770 7140 0 net11
rlabel metal1 5290 2618 5290 2618 0 net12
rlabel metal2 24058 2689 24058 2689 0 net13
rlabel metal1 6210 2856 6210 2856 0 net14
rlabel metal1 8970 2618 8970 2618 0 net15
rlabel metal1 10580 3910 10580 3910 0 net16
rlabel metal1 12742 4590 12742 4590 0 net17
rlabel metal1 13938 4794 13938 4794 0 net18
rlabel metal1 15318 3434 15318 3434 0 net19
rlabel metal2 20102 5678 20102 5678 0 net2
rlabel metal1 17710 2618 17710 2618 0 net20
rlabel metal1 19458 2618 19458 2618 0 net21
rlabel metal2 21942 2689 21942 2689 0 net22
rlabel metal1 15226 7412 15226 7412 0 net23
rlabel metal2 5842 7038 5842 7038 0 net24
rlabel metal1 1794 7412 1794 7412 0 net25
rlabel metal1 3726 6970 3726 6970 0 net26
rlabel metal1 5428 7378 5428 7378 0 net27
rlabel metal1 6716 6970 6716 6970 0 net28
rlabel metal1 8740 6970 8740 6970 0 net29
rlabel via2 18722 3451 18722 3451 0 net3
rlabel metal1 10212 6970 10212 6970 0 net30
rlabel metal1 11822 7378 11822 7378 0 net31
rlabel metal1 19274 6868 19274 6868 0 net32
rlabel metal2 2254 2465 2254 2465 0 net33
rlabel metal1 26910 2414 26910 2414 0 net34
rlabel metal2 25530 2414 25530 2414 0 net35
rlabel metal1 26542 2448 26542 2448 0 net36
rlabel via2 1794 2363 1794 2363 0 net37
rlabel metal2 24656 2788 24656 2788 0 net38
rlabel metal1 4646 2380 4646 2380 0 net39
rlabel metal1 18170 6120 18170 6120 0 net4
rlabel metal1 23506 2380 23506 2380 0 net40
rlabel metal2 6394 2618 6394 2618 0 net41
rlabel metal1 8142 2482 8142 2482 0 net42
rlabel metal2 9936 2414 9936 2414 0 net43
rlabel metal1 12236 2414 12236 2414 0 net44
rlabel metal1 13478 2414 13478 2414 0 net45
rlabel viali 15505 2414 15505 2414 0 net46
rlabel metal1 17342 2448 17342 2448 0 net47
rlabel metal2 19550 2618 19550 2618 0 net48
rlabel metal1 21022 2448 21022 2448 0 net49
rlabel metal2 18722 6052 18722 6052 0 net5
rlabel metal1 16054 1870 16054 1870 0 net50
rlabel metal2 2714 3536 2714 3536 0 net51
rlabel metal1 14214 2414 14214 2414 0 net52
rlabel metal2 2346 2720 2346 2720 0 net53
rlabel metal2 10350 6120 10350 6120 0 net54
rlabel metal2 2346 4063 2346 4063 0 net55
rlabel metal2 26542 6817 26542 6817 0 net56
rlabel metal1 15134 3706 15134 3706 0 net57
rlabel metal2 17066 2091 17066 2091 0 net58
rlabel via2 2622 5219 2622 5219 0 net59
rlabel metal2 19734 5678 19734 5678 0 net6
rlabel metal2 2346 4641 2346 4641 0 net60
rlabel metal2 2346 4947 2346 4947 0 net61
rlabel metal2 2254 7548 2254 7548 0 net62
rlabel metal1 1886 3468 1886 3468 0 net63
rlabel metal2 2070 5882 2070 5882 0 net64
rlabel metal2 1702 5729 1702 5729 0 net65
rlabel via2 2070 6307 2070 6307 0 net66
rlabel metal2 2438 5457 2438 5457 0 net67
rlabel metal1 1978 5304 1978 5304 0 net68
rlabel metal2 2668 5100 2668 5100 0 net69
rlabel metal1 20056 7310 20056 7310 0 net7
rlabel metal2 1702 7344 1702 7344 0 net70
rlabel metal2 2162 5491 2162 5491 0 net71
rlabel metal1 26082 2992 26082 2992 0 net72
rlabel metal1 26818 5236 26818 5236 0 net73
rlabel metal2 26174 2890 26174 2890 0 net74
rlabel metal1 26450 3094 26450 3094 0 net75
rlabel metal1 26634 3026 26634 3026 0 net76
rlabel metal1 27278 3060 27278 3060 0 net77
rlabel metal1 27002 3502 27002 3502 0 net78
rlabel metal1 26542 4080 26542 4080 0 net79
rlabel metal1 20884 5202 20884 5202 0 net8
rlabel metal1 27278 3468 27278 3468 0 net80
rlabel metal1 27278 4148 27278 4148 0 net81
rlabel metal1 26910 4556 26910 4556 0 net82
rlabel metal2 2944 2414 2944 2414 0 net83
rlabel metal1 1702 4624 1702 4624 0 net84
rlabel metal2 2622 2618 2622 2618 0 net85
rlabel metal1 2346 3026 2346 3026 0 net86
rlabel metal1 2116 3026 2116 3026 0 net87
rlabel metal1 1840 3026 1840 3026 0 net88
rlabel metal1 2162 3502 2162 3502 0 net89
rlabel metal2 25530 2822 25530 2822 0 net9
rlabel metal1 1702 3536 1702 3536 0 net90
rlabel metal1 2162 4114 2162 4114 0 net91
rlabel metal1 1702 4080 1702 4080 0 net92
rlabel metal1 2162 4590 2162 4590 0 net93
rlabel metal2 9154 6562 9154 6562 0 net94
rlabel metal1 9108 4182 9108 4182 0 net95
rlabel metal1 9614 6732 9614 6732 0 net96
rlabel metal1 15272 4998 15272 4998 0 net97
rlabel metal1 7314 2992 7314 2992 0 net98
rlabel metal1 14858 7412 14858 7412 0 net99
rlabel metal1 5382 6256 5382 6256 0 result\[0\]
rlabel metal2 19182 3111 19182 3111 0 result\[10\]
rlabel metal1 15364 6630 15364 6630 0 result\[11\]
rlabel metal1 5152 2822 5152 2822 0 result\[1\]
rlabel metal1 5888 5882 5888 5882 0 result\[2\]
rlabel metal1 8740 5746 8740 5746 0 result\[3\]
rlabel metal1 9752 4998 9752 4998 0 result\[4\]
rlabel metal2 10994 5474 10994 5474 0 result\[5\]
rlabel metal1 13248 6426 13248 6426 0 result\[6\]
rlabel metal1 12880 3910 12880 3910 0 result\[7\]
rlabel metal1 15548 5542 15548 5542 0 result\[8\]
rlabel metal1 14214 5202 14214 5202 0 result\[9\]
rlabel metal1 15640 7378 15640 7378 0 rst_z
rlabel metal1 18860 7378 18860 7378 0 start
rlabel metal1 21482 6154 21482 6154 0 state\[0\]
rlabel metal1 23414 4726 23414 4726 0 state\[1\]
rlabel metal2 22770 1452 22770 1452 0 vcm_o[10]
rlabel metal2 23690 1384 23690 1384 0 vcm_o_i[10]
rlabel metal2 8970 1384 8970 1384 0 vcm_o_i[2]
rlabel metal2 10810 1384 10810 1384 0 vcm_o_i[3]
rlabel metal2 12650 1384 12650 1384 0 vcm_o_i[4]
rlabel metal2 16330 1384 16330 1384 0 vcm_o_i[6]
rlabel metal2 18170 1384 18170 1384 0 vcm_o_i[7]
rlabel metal2 20010 1384 20010 1384 0 vcm_o_i[8]
rlabel metal2 21850 1384 21850 1384 0 vcm_o_i[9]
rlabel metal3 27608 7956 27608 7956 0 vin_n_sw_on
rlabel metal2 27462 4879 27462 4879 0 vref_z_n_o[0]
rlabel metal2 27462 7599 27462 7599 0 vref_z_n_o[10]
rlabel metal3 28114 5236 28114 5236 0 vref_z_n_o[1]
rlabel metal3 27930 5508 27930 5508 0 vref_z_n_o[2]
rlabel metal3 27746 5780 27746 5780 0 vref_z_n_o[3]
rlabel metal2 27462 5967 27462 5967 0 vref_z_n_o[4]
rlabel metal3 27746 6324 27746 6324 0 vref_z_n_o[5]
rlabel metal2 27462 6511 27462 6511 0 vref_z_n_o[6]
rlabel metal3 27930 6868 27930 6868 0 vref_z_n_o[7]
rlabel metal2 27462 7055 27462 7055 0 vref_z_n_o[8]
rlabel metal3 27746 7412 27746 7412 0 vref_z_n_o[9]
rlabel metal1 1564 7514 1564 7514 0 vref_z_p_o[10]
rlabel metal3 544 5236 544 5236 0 vref_z_p_o[1]
rlabel metal3 1096 5508 1096 5508 0 vref_z_p_o[2]
rlabel metal3 544 5780 544 5780 0 vref_z_p_o[3]
rlabel metal1 1702 6630 1702 6630 0 vref_z_p_o[5]
rlabel metal1 1150 6426 1150 6426 0 vref_z_p_o[6]
rlabel metal3 1372 6868 1372 6868 0 vref_z_p_o[7]
rlabel metal2 1518 7055 1518 7055 0 vref_z_p_o[8]
rlabel metal2 1886 7191 1886 7191 0 vref_z_p_o[9]
rlabel metal3 27700 4692 27700 4692 0 vss_n_o[10]
rlabel metal3 27562 2244 27562 2244 0 vss_n_o[1]
rlabel metal3 27424 2516 27424 2516 0 vss_n_o[2]
rlabel metal3 27746 2788 27746 2788 0 vss_n_o[3]
rlabel metal3 28114 3060 28114 3060 0 vss_n_o[4]
rlabel metal3 27930 3332 27930 3332 0 vss_n_o[5]
rlabel metal3 28229 3604 28229 3604 0 vss_n_o[6]
rlabel metal2 27462 3791 27462 3791 0 vss_n_o[7]
rlabel metal3 28114 4148 28114 4148 0 vss_n_o[8]
rlabel metal3 27930 4420 27930 4420 0 vss_n_o[9]
rlabel metal3 544 4692 544 4692 0 vss_p_o[10]
rlabel metal3 544 3060 544 3060 0 vss_p_o[4]
rlabel metal3 544 3604 544 3604 0 vss_p_o[6]
rlabel metal3 27372 1972 27372 1972 0 vss_n_o[0]
rlabel metal3 1071 1972 1071 1972 0 vss_p_o[0]
rlabel metal3 1025 2244 1025 2244 0 vss_p_o[1]
flabel metal3 s 28077 7896 28477 8016 0 FreeSans 480 0 0 0 vin_n_sw_on
port 49 nsew signal input
flabel metal3 s 28077 4904 28477 5024 0 FreeSans 480 0 0 0 vref_z_n_o[0]
port 51 nsew signal output
flabel metal3 s 28077 7624 28477 7744 0 FreeSans 480 0 0 0 vref_z_n_o[10]
port 52 nsew signal output
flabel metal3 s 28077 5176 28477 5296 0 FreeSans 480 0 0 0 vref_z_n_o[1]
port 53 nsew signal output
flabel metal3 s 28077 5448 28477 5568 0 FreeSans 480 0 0 0 vref_z_n_o[2]
port 54 nsew signal output
flabel metal3 s 28077 5720 28477 5840 0 FreeSans 480 0 0 0 vref_z_n_o[3]
port 55 nsew signal output
flabel metal3 s 28077 5992 28477 6112 0 FreeSans 480 0 0 0 vref_z_n_o[4]
port 56 nsew signal output
flabel metal3 s 28077 6264 28477 6384 0 FreeSans 480 0 0 0 vref_z_n_o[5]
port 57 nsew signal output
flabel metal3 s 28077 6536 28477 6656 0 FreeSans 480 0 0 0 vref_z_n_o[6]
port 58 nsew signal output
flabel metal3 s 28077 6808 28477 6928 0 FreeSans 480 0 0 0 vref_z_n_o[7]
port 59 nsew signal output
flabel metal3 s 28077 7080 28477 7200 0 FreeSans 480 0 0 0 vref_z_n_o[8]
port 60 nsew signal output
flabel metal3 s 28077 7352 28477 7472 0 FreeSans 480 0 0 0 vref_z_n_o[9]
port 61 nsew signal output
flabel metal3 s 28077 1912 28477 2032 0 FreeSans 480 0 0 0 vss_n_o[0]
port 73 nsew signal output
flabel metal3 s 28077 4632 28477 4752 0 FreeSans 480 0 0 0 vss_n_o[10]
port 74 nsew signal output
flabel metal3 s 28077 2184 28477 2304 0 FreeSans 480 0 0 0 vss_n_o[1]
port 75 nsew signal output
flabel metal3 s 28077 2456 28477 2576 0 FreeSans 480 0 0 0 vss_n_o[2]
port 76 nsew signal output
flabel metal3 s 28077 2728 28477 2848 0 FreeSans 480 0 0 0 vss_n_o[3]
port 77 nsew signal output
flabel metal3 s 28077 3000 28477 3120 0 FreeSans 480 0 0 0 vss_n_o[4]
port 78 nsew signal output
flabel metal3 s 28077 3272 28477 3392 0 FreeSans 480 0 0 0 vss_n_o[5]
port 79 nsew signal output
flabel metal3 s 28077 3544 28477 3664 0 FreeSans 480 0 0 0 vss_n_o[6]
port 80 nsew signal output
flabel metal3 s 28077 3816 28477 3936 0 FreeSans 480 0 0 0 vss_n_o[7]
port 81 nsew signal output
flabel metal3 s 28077 4088 28477 4208 0 FreeSans 480 0 0 0 vss_n_o[8]
port 82 nsew signal output
flabel metal3 s 28077 4360 28477 4480 0 FreeSans 480 0 0 0 vss_n_o[9]
port 83 nsew signal output
rlabel metal3 1012 4148 1012 4148 0 vss_p_o[8]
rlabel metal3 736 4964 736 4964 0 vref_z_p_o[0]
rlabel metal3 736 6052 736 6052 0 vref_z_p_o[4]
rlabel metal3 736 2788 736 2788 0 vss_p_o[3]
rlabel metal3 736 3332 736 3332 0 vss_p_o[5]
rlabel metal3 736 3876 736 3876 0 vss_p_o[7]
rlabel metal3 736 4420 736 4420 0 vss_p_o[9]
rlabel metal3 951 2516 951 2516 0 vss_p_o[2]
flabel metal3 s 480 4360 880 4480 0 FreeSans 480 0 0 0 vss_p_o[9]
port 94 nsew signal output
flabel metal3 s 480 4088 880 4208 0 FreeSans 480 0 0 0 vss_p_o[8]
port 93 nsew signal output
flabel metal3 s 480 3816 880 3936 0 FreeSans 480 0 0 0 vss_p_o[7]
port 92 nsew signal output
flabel metal3 s 480 3544 880 3664 0 FreeSans 480 0 0 0 vss_p_o[6]
port 91 nsew signal output
flabel metal3 s 480 3272 880 3392 0 FreeSans 480 0 0 0 vss_p_o[5]
port 90 nsew signal output
flabel metal3 s 480 3000 880 3120 0 FreeSans 480 0 0 0 vss_p_o[4]
port 89 nsew signal output
flabel metal3 s 480 2728 880 2848 0 FreeSans 480 0 0 0 vss_p_o[3]
port 88 nsew signal output
flabel metal3 s 480 2456 880 2576 0 FreeSans 480 0 0 0 vss_p_o[2]
port 87 nsew signal output
flabel metal3 s 480 2184 880 2304 0 FreeSans 480 0 0 0 vss_p_o[1]
port 86 nsew signal output
flabel metal3 s 480 4632 880 4752 0 FreeSans 480 0 0 0 vss_p_o[10]
port 85 nsew signal output
flabel metal3 s 480 1912 880 2032 0 FreeSans 480 0 0 0 vss_p_o[0]
port 84 nsew signal output
flabel metal3 s 480 7352 880 7472 0 FreeSans 480 0 0 0 vref_z_p_o[9]
port 72 nsew signal output
flabel metal3 s 480 7080 880 7200 0 FreeSans 480 0 0 0 vref_z_p_o[8]
port 71 nsew signal output
flabel metal3 s 480 6808 880 6928 0 FreeSans 480 0 0 0 vref_z_p_o[7]
port 70 nsew signal output
flabel metal3 s 480 6536 880 6656 0 FreeSans 480 0 0 0 vref_z_p_o[6]
port 69 nsew signal output
flabel metal3 s 480 6264 880 6384 0 FreeSans 480 0 0 0 vref_z_p_o[5]
port 68 nsew signal output
flabel metal3 s 480 5992 880 6112 0 FreeSans 480 0 0 0 vref_z_p_o[4]
port 67 nsew signal output
flabel metal3 s 480 5720 880 5840 0 FreeSans 480 0 0 0 vref_z_p_o[3]
port 66 nsew signal output
flabel metal3 s 480 5448 880 5568 0 FreeSans 480 0 0 0 vref_z_p_o[2]
port 65 nsew signal output
flabel metal3 s 480 5176 880 5296 0 FreeSans 480 0 0 0 vref_z_p_o[1]
port 64 nsew signal output
flabel metal3 s 480 7624 880 7744 0 FreeSans 480 0 0 0 vref_z_p_o[10]
port 63 nsew signal output
flabel metal3 s 480 4904 880 5024 0 FreeSans 480 0 0 0 vref_z_p_o[0]
port 62 nsew signal output
flabel metal3 s 480 7896 880 8016 0 FreeSans 480 0 0 0 vin_p_sw_on
port 50 nsew signal input
flabel metal2 s 3422 1360 3478 1760 0 FreeSans 224 90 0 0 comp_n
port 4 nsew signal input
flabel metal2 s 2502 1360 2558 1760 0 FreeSans 224 90 0 0 comp_p
port 5 nsew signal input
flabel metal2 s 1582 1360 1638 1760 0 FreeSans 224 90 0 0 en_comp
port 17 nsew signal output
flabel metal2 s 25502 1360 25558 1760 0 FreeSans 224 90 0 0 en_vcm_sw_o
port 20 nsew signal output
flabel metal2 s 26422 1360 26478 1760 0 FreeSans 224 90 0 0 en_vcm_sw_o_i
port 21 nsew signal input
flabel metal2 s 24582 1360 24638 1760 0 FreeSans 224 90 0 0 vcm_dummy_o
port 26 nsew signal output
flabel metal2 s 4342 1360 4398 1760 0 FreeSans 224 90 0 0 vcm_o[0]
port 27 nsew signal output
flabel metal2 s 22742 1360 22798 1760 0 FreeSans 224 90 0 0 vcm_o[10]
port 28 nsew signal output
flabel metal2 s 6182 1360 6238 1760 0 FreeSans 224 90 0 0 vcm_o[1]
port 29 nsew signal output
flabel metal2 s 8022 1360 8078 1760 0 FreeSans 224 90 0 0 vcm_o[2]
port 30 nsew signal output
flabel metal2 s 9862 1360 9918 1760 0 FreeSans 224 90 0 0 vcm_o[3]
port 31 nsew signal output
flabel metal2 s 11702 1360 11758 1760 0 FreeSans 224 90 0 0 vcm_o[4]
port 32 nsew signal output
flabel metal2 s 13542 1360 13598 1760 0 FreeSans 224 90 0 0 vcm_o[5]
port 33 nsew signal output
flabel metal2 s 15382 1360 15438 1760 0 FreeSans 224 90 0 0 vcm_o[6]
port 34 nsew signal output
flabel metal2 s 17222 1360 17278 1760 0 FreeSans 224 90 0 0 vcm_o[7]
port 35 nsew signal output
flabel metal2 s 19062 1360 19118 1760 0 FreeSans 224 90 0 0 vcm_o[8]
port 36 nsew signal output
flabel metal2 s 20902 1360 20958 1760 0 FreeSans 224 90 0 0 vcm_o[9]
port 37 nsew signal output
flabel metal2 s 5262 1360 5318 1760 0 FreeSans 224 90 0 0 vcm_o_i[0]
port 38 nsew signal input
flabel metal2 s 23662 1360 23718 1760 0 FreeSans 224 90 0 0 vcm_o_i[10]
port 39 nsew signal input
flabel metal2 s 7102 1360 7158 1760 0 FreeSans 224 90 0 0 vcm_o_i[1]
port 40 nsew signal input
flabel metal2 s 8942 1360 8998 1760 0 FreeSans 224 90 0 0 vcm_o_i[2]
port 41 nsew signal input
flabel metal2 s 10782 1360 10838 1760 0 FreeSans 224 90 0 0 vcm_o_i[3]
port 42 nsew signal input
flabel metal2 s 12622 1360 12678 1760 0 FreeSans 224 90 0 0 vcm_o_i[4]
port 43 nsew signal input
flabel metal2 s 14462 1360 14518 1760 0 FreeSans 224 90 0 0 vcm_o_i[5]
port 44 nsew signal input
flabel metal2 s 16302 1360 16358 1760 0 FreeSans 224 90 0 0 vcm_o_i[6]
port 45 nsew signal input
flabel metal2 s 18142 1360 18198 1760 0 FreeSans 224 90 0 0 vcm_o_i[7]
port 46 nsew signal input
flabel metal2 s 19982 1360 20038 1760 0 FreeSans 224 90 0 0 vcm_o_i[8]
port 47 nsew signal input
flabel metal2 s 21822 1360 21878 1760 0 FreeSans 224 90 0 0 vcm_o_i[9]
port 48 nsew signal input
flabel metal2 s 27066 1360 27122 1760 0 FreeSans 224 90 0 0 offset_cal_cycle
port 22 nsew signal output
rlabel metal2 27094 1775 27094 1775 0 offset_cal_cycle
flabel metal2 s 1040 1360 1096 1760 0 FreeSans 224 90 0 0 sample_o
port 24 nsew signal output
flabel metal2 s 27825 1360 27881 1760 0 FreeSans 224 90 0 0 en_offset_cal_o
port 19 nsew signal output
flabel metal2 s 17038 7580 17094 7980 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 1306 7580 1362 7980 0 FreeSans 224 90 0 0 clk_data
port 3 nsew signal output
flabel metal2 s 6550 7580 6606 7980 0 FreeSans 224 90 0 0 data[2]
port 8 nsew signal output
flabel metal2 s 8298 7580 8354 7980 0 FreeSans 224 90 0 0 data[3]
port 9 nsew signal output
flabel metal2 s 10046 7580 10102 7980 0 FreeSans 224 90 0 0 data[4]
port 10 nsew signal output
flabel metal2 s 11794 7580 11850 7980 0 FreeSans 224 90 0 0 data[5]
port 11 nsew signal output
flabel metal2 s 22282 7580 22338 7980 0 FreeSans 224 90 0 0 debug_mux[0]
port 12 nsew signal input
flabel metal2 s 24030 7580 24086 7980 0 FreeSans 224 90 0 0 debug_mux[1]
port 13 nsew signal input
flabel metal2 s 25778 7580 25834 7980 0 FreeSans 224 90 0 0 debug_mux[2]
port 14 nsew signal input
flabel metal2 s 27526 7580 27582 7980 0 FreeSans 224 90 0 0 debug_mux[3]
port 15 nsew signal input
flabel metal2 s 13542 7580 13598 7980 0 FreeSans 224 90 0 0 debug_out
port 16 nsew signal output
flabel metal2 s 20534 7580 20590 7980 0 FreeSans 224 90 0 0 en_offset_cal
port 18 nsew signal input
flabel metal2 s 15290 7580 15346 7980 0 FreeSans 224 90 0 0 rst_z
port 23 nsew signal input
flabel metal2 s 18786 7580 18842 7980 0 FreeSans 224 90 0 0 start
port 25 nsew signal input
flabel metal2 s 4709 7580 4765 7980 0 FreeSans 224 90 0 0 data[1]
port 7 nsew signal output
rlabel metal2 4740 7704 4740 7704 0 data[1]
flabel metal2 s 3146 7580 3202 7980 0 FreeSans 224 90 0 0 data[0]
port 6 nsew signal output
rlabel metal2 3170 7704 3170 7704 0 data[0]
rlabel metal2 1610 1616 1610 1616 0 en_comp
rlabel metal2 25530 1616 25530 1616 0 en_vcm_sw_o
rlabel metal2 24610 1616 24610 1616 0 vcm_dummy_o
rlabel metal2 6210 1616 6210 1616 0 vcm_o[1]
rlabel metal2 8050 1616 8050 1616 0 vcm_o[2]
rlabel metal2 9890 1616 9890 1616 0 vcm_o[3]
rlabel metal2 13570 1616 13570 1616 0 vcm_o[5]
rlabel metal2 15410 1616 15410 1616 0 vcm_o[6]
rlabel metal2 17250 1616 17250 1616 0 vcm_o[7]
rlabel metal2 19090 1616 19090 1616 0 vcm_o[8]
rlabel metal2 20930 1616 20930 1616 0 vcm_o[9]
rlabel metal2 7130 1616 7130 1616 0 vcm_o_i[1]
rlabel metal2 4370 1535 4370 1535 0 vcm_o[0]
rlabel metal2 11730 1535 11730 1535 0 vcm_o[4]
rlabel metal2 5290 1603 5290 1603 0 vcm_o_i[0]
rlabel metal2 14490 1603 14490 1603 0 vcm_o_i[5]
rlabel metal2 26450 1410 26450 1410 0 en_vcm_sw_o_i
rlabel metal2 27853 1410 27853 1410 0 en_offset_cal_o
rlabel metal2 2530 1390 2530 1390 0 comp_p
rlabel metal2 1068 1390 1068 1390 0 sample_o
rlabel metal3 728 7956 728 7956 0 vin_p_sw_on
rlabel metal2 13570 7838 13570 7838 0 debug_out
rlabel metal2 11822 7872 11822 7872 0 data[5]
rlabel metal2 10074 7872 10074 7872 0 data[4]
rlabel metal2 8326 7872 8326 7872 0 data[3]
rlabel metal2 6578 7872 6578 7872 0 data[2]
rlabel metal2 1334 7838 1334 7838 0 clk_data
<< properties >>
string FIXED_BBOX 0 0 29000 10000
<< end >>
