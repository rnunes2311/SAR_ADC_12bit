* NGSPICE file created from state_machine.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends


.subckt state_machine VDD VSS RST_Z START COMP_P COMP_N SAMPLE_O VCM_O[10] VCM_O[9] VCM_O[8] VCM_O[7] VCM_O[6] VCM_O[5] VCM_O[4] VCM_O[3] VCM_O[2]
+ VCM_O[1] VCM_O[0] EN_COMP VIN_P_SW_ON VIN_N_SW_ON VCM_DUMMY_O EN_VCM_SW_O EN_OFFSET_CAL OFFSET_CAL_CYCLE EN_OFFSET_CAL_O CLK_DATA DATA[5]
+ DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] DEBUG_MUX[3] DEBUG_MUX[2] DEBUG_MUX[1] DEBUG_MUX[0] DEBUG_OUT VSS_N_O[10] VSS_N_O[9] VSS_N_O[8]
+ VSS_N_O[7] VSS_N_O[6] VSS_N_O[5] VSS_N_O[4] VSS_N_O[3] VSS_N_O[2] VSS_N_O[1] VSS_N_O[0] VREF_Z_N_O[10] VREF_Z_N_O[9] VREF_Z_N_O[8]
+ VREF_Z_N_O[7] VREF_Z_N_O[6] VREF_Z_N_O[5] VREF_Z_N_O[4] VREF_Z_N_O[3] VREF_Z_N_O[2] VREF_Z_N_O[1] VREF_Z_N_O[0] VSS_P_O[10] VSS_P_O[9]
+ VSS_P_O[8] VSS_P_O[7] VSS_P_O[6] VSS_P_O[5] VSS_P_O[4] VSS_P_O[3] VSS_P_O[2] VSS_P_O[1] VSS_P_O[0] VREF_Z_P_O[10] VREF_Z_P_O[9]
+ VREF_Z_P_O[8] VREF_Z_P_O[7] VREF_Z_P_O[6] VREF_Z_P_O[5] VREF_Z_P_O[4] VREF_Z_P_O[3] VREF_Z_P_O[2] VREF_Z_P_O[1] VREF_Z_P_O[0] CLK EN_VCM_SW_O_I
+ VCM_O_I[10] VCM_O_I[9] VCM_O_I[8] VCM_O_I[7] VCM_O_I[6] VCM_O_I[5] VCM_O_I[4] VCM_O_I[3] VCM_O_I[2] VCM_O_I[1] VCM_O_I[0] SINGLE_ENDED
X_363_ net102 _139_ _140_ _135_ VSS VSS VDD VDD _141_ sky130_fd_sc_hd__a31o_1
X_432_ net116 _014_ net113 VSS VSS VDD VDD counter\[8\] sky130_fd_sc_hd__dfrtp_4
X_294_ _066_ _100_ VSS VSS VDD VDD net67 sky130_fd_sc_hd__or2_1
Xfanout105 net108 VSS VSS VDD VDD net105 sky130_fd_sc_hd__buf_2
XFILLER_0_1_152 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xfanout116 net117 VSS VSS VDD VDD net116 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_66 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ counter\[6\] net106 net101 net109 VSS VSS VDD VDD _170_ sky130_fd_sc_hd__and4bb_1
X_346_ counter\[7\] counter\[6\] counter\[5\] counter\[2\] VSS VSS VDD VDD _131_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_222 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_277_ result\[8\] _092_ VSS VSS VDD VDD _093_ sky130_fd_sc_hd__nor2_1
X_200_ result\[6\] result\[0\] net110 VSS VSS VDD VDD _051_ sky130_fd_sc_hd__mux2_1
X_329_ counter\[8\] net5 _047_ net6 VSS VSS VDD VDD _117_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_203 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_169 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
*XANTENNA_5 net75 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
Xoutput31 net31 VSS VSS VDD VDD data[4] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 VSS VSS VDD VDD vcm_o[1] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VSS VSS VDD VDD vss_p_o[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_35 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 VSS VSS VDD VDD vref_z_p_o[1] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VSS VSS VDD VDD vref_z_n_o[1] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VSS VSS VDD VDD vss_n_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_93 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_362_ counter\[10\] _074_ VSS VSS VDD VDD _140_ sky130_fd_sc_hd__or2_1
X_431_ net116 _013_ net113 VSS VSS VDD VDD counter\[7\] sky130_fd_sc_hd__dfrtp_1
X_293_ result\[5\] result\[4\] net104 VSS VSS VDD VDD _100_ sky130_fd_sc_hd__mux2_1
Xfanout106 net108 VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkbuf_2
Xfanout117 net1 VSS VSS VDD VDD net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_275 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_253 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_67 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ counter\[10\] net98 _071_ VSS VSS VDD VDD _092_ sky130_fd_sc_hd__a21oi_1
X_414_ _136_ result\[3\] _169_ VSS VSS VDD VDD _024_ sky130_fd_sc_hd__mux2_1
X_345_ counter\[1\] counter\[3\] counter\[11\] counter\[10\] VSS VSS VDD VDD _130_
+ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_4_Left_14 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_328_ counter\[9\] _046_ net4 _115_ VSS VSS VDD VDD _116_ sky130_fd_sc_hd__a31o_1
X_259_ net95 _084_ net55 VSS VSS VDD VDD net88 sky130_fd_sc_hd__o21ai_1
*XANTENNA_6 net76 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput32 net32 VSS VSS VDD VDD data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 VSS VSS VDD VDD vref_z_n_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_7_181 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput43 net43 VSS VSS VDD VDD vcm_o[2] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VSS VSS VDD VDD vss_p_o[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_36 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput76 net76 VSS VSS VDD VDD vss_n_o[2] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VSS VSS VDD VDD vref_z_p_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_5_129 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_361_ net106 _031_ VSS VSS VDD VDD _139_ sky130_fd_sc_hd__nand2_1
X_292_ _083_ _099_ VSS VSS VDD VDD net66 sky130_fd_sc_hd__or2_1
X_430_ net116 _012_ net113 VSS VSS VDD VDD counter\[6\] sky130_fd_sc_hd__dfrtp_4
Xfanout107 net108 VSS VSS VDD VDD net107 sky130_fd_sc_hd__clkbuf_2
X_344_ net12 _129_ _000_ VSS VSS VDD VDD _173_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_68 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_275_ result\[9\] _071_ VSS VSS VDD VDD net60 sky130_fd_sc_hd__nand2_1
X_413_ net100 _167_ _168_ _135_ VSS VSS VDD VDD _169_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_246 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_189_ result\[3\] VSS VSS VDD VDD _040_ sky130_fd_sc_hd__inv_2
X_258_ result\[3\] _083_ VSS VSS VDD VDD _084_ sky130_fd_sc_hd__nor2_1
X_327_ counter\[10\] _112_ VSS VSS VDD VDD _115_ sky130_fd_sc_hd__and2_1
Xoutput55 net55 VSS VSS VDD VDD vref_z_n_o[3] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VSS VSS VDD VDD debug_out sky130_fd_sc_hd__clkbuf_4
Xoutput66 net66 VSS VSS VDD VDD vref_z_p_o[3] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VSS VSS VDD VDD vcm_o[3] sky130_fd_sc_hd__buf_2
Xoutput88 net88 VSS VSS VDD VDD vss_p_o[3] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VSS VSS VDD VDD vss_n_o[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_37 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ result\[4\] result\[3\] net104 VSS VSS VDD VDD _099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_130 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_152 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_360_ result\[11\] _108_ _137_ _138_ net103 VSS VSS VDD VDD _001_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_266 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xfanout108 single_ended_reg VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_69 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _119_ _122_ _128_ _129_ _127_ VSS VSS VDD VDD net33 sky130_fd_sc_hd__o32a_1
X_274_ net95 _091_ net59 VSS VSS VDD VDD net92 sky130_fd_sc_hd__o21ai_1
X_412_ net105 counter\[3\] _034_ VSS VSS VDD VDD _168_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_85 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_326_ _109_ _110_ _113_ net6 VSS VSS VDD VDD _114_ sky130_fd_sc_hd__or4b_1
X_188_ result\[8\] VSS VSS VDD VDD _039_ sky130_fd_sc_hd__inv_2
X_257_ _059_ _082_ _065_ VSS VSS VDD VDD _083_ sky130_fd_sc_hd__o21a_1
X_309_ counter\[3\] _106_ VSS VSS VDD VDD net43 sky130_fd_sc_hd__nor2_1
XFILLER_0_1_42 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_8_106 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xoutput56 net56 VSS VSS VDD VDD vref_z_n_o[4] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VSS VSS VDD VDD vss_n_o[4] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VSS VSS VDD VDD vref_z_p_o[4] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VSS VSS VDD VDD vcm_o[4] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VSS VSS VDD VDD en_comp sky130_fd_sc_hd__buf_2
Xoutput89 net89 VSS VSS VDD VDD vss_p_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_38 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_186 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_290_ _080_ _098_ VSS VSS VDD VDD net65 sky130_fd_sc_hd__or2_1
XFILLER_0_1_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xfanout109 counter\[7\] VSS VSS VDD VDD net109 sky130_fd_sc_hd__buf_2
X_342_ state\[1\] state\[0\] VSS VSS VDD VDD _129_ sky130_fd_sc_hd__nor2_2
X_273_ result\[7\] _090_ VSS VSS VDD VDD _091_ sky130_fd_sc_hd__nor2_1
X_411_ net110 _082_ VSS VSS VDD VDD _167_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_53 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_5_281 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_187_ result\[2\] VSS VSS VDD VDD _038_ sky130_fd_sc_hd__inv_2
X_256_ net108 counter\[5\] VSS VSS VDD VDD _082_ sky130_fd_sc_hd__nand2_1
X_325_ _047_ _111_ _112_ counter\[6\] VSS VSS VDD VDD _113_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_8_Left_18 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_308_ counter\[2\] _106_ VSS VSS VDD VDD net42 sky130_fd_sc_hd__nor2_1
X_239_ _043_ _073_ net98 VSS VSS VDD VDD net83 sky130_fd_sc_hd__a21o_1
Xoutput57 net57 VSS VSS VDD VDD vref_z_n_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_162 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput46 net46 VSS VSS VDD VDD vcm_o[5] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VSS VSS VDD VDD en_offset_cal_o sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_2_39 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput79 net79 VSS VSS VDD VDD vss_n_o[5] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VSS VSS VDD VDD vref_z_p_o[5] sky130_fd_sc_hd__buf_2
X_341_ _048_ net6 _124_ _126_ VSS VSS VDD VDD _128_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_235 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_272_ counter\[9\] net98 _069_ VSS VSS VDD VDD _090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_190 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_410_ _166_ net3 _165_ VSS VSS VDD VDD _023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_76 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_324_ net5 net4 VSS VSS VDD VDD _112_ sky130_fd_sc_hd__nor2_1
X_255_ _042_ _065_ VSS VSS VDD VDD net55 sky130_fd_sc_hd__or2_1
X_186_ result\[7\] VSS VSS VDD VDD _037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_70 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_307_ counter\[1\] _106_ VSS VSS VDD VDD net40 sky130_fd_sc_hd__nor2_1
X_238_ net23 _072_ VSS VSS VDD VDD _073_ sky130_fd_sc_hd__nor2_1
Xoutput58 net58 VSS VSS VDD VDD vref_z_n_o[6] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VSS VSS VDD VDD vcm_o[6] sky130_fd_sc_hd__buf_2
Xoutput36 net36 VSS VSS VDD VDD en_vcm_sw_o sky130_fd_sc_hd__buf_2
Xoutput69 net69 VSS VSS VDD VDD vref_z_p_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_4_144 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_4_166 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_9_258 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_340_ _112_ _121_ VSS VSS VDD VDD _127_ sky130_fd_sc_hd__nand2_1
X_271_ result\[8\] _069_ VSS VSS VDD VDD net59 sky130_fd_sc_hd__nand2_1
X_254_ net95 _081_ net54 VSS VSS VDD VDD net87 sky130_fd_sc_hd__o21ai_1
X_185_ result\[1\] VSS VSS VDD VDD _036_ sky130_fd_sc_hd__inv_2
X_323_ counter\[2\] net5 VSS VSS VDD VDD _111_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_71 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ net103 net39 VSS VSS VDD VDD _106_ sky130_fd_sc_hd__nand2_4
X_237_ net107 counter\[10\] VSS VSS VDD VDD _072_ sky130_fd_sc_hd__nand2b_1
Xoutput26 net26 VSS VSS VDD VDD clk_data sky130_fd_sc_hd__clkbuf_4
Xoutput59 net59 VSS VSS VDD VDD vref_z_n_o[7] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VSS VSS VDD VDD vcm_o[7] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput37 net37 VSS VSS VDD VDD offset_cal_cycle sky130_fd_sc_hd__buf_2
XFILLER_0_7_11 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_178 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_40 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_248 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_270_ net95 _089_ net58 VSS VSS VDD VDD net91 sky130_fd_sc_hd__o21ai_1
X_399_ counter\[5\] _056_ _058_ _158_ VSS VSS VDD VDD _159_ sky130_fd_sc_hd__a211o_1
X_322_ counter\[0\] net5 net4 VSS VSS VDD VDD _110_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_72 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_253_ result\[2\] _080_ VSS VSS VDD VDD _081_ sky130_fd_sc_hd__nor2_1
X_184_ result\[6\] VSS VSS VDD VDD _035_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_287 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_236_ _041_ _071_ net98 VSS VSS VDD VDD net82 sky130_fd_sc_hd__a21o_1
X_305_ net103 _043_ net74 VSS VSS VDD VDD net63 sky130_fd_sc_hd__o21ai_1
X_219_ result\[1\] _062_ net95 VSS VSS VDD VDD net73 sky130_fd_sc_hd__o21ai_2
Xoutput27 net27 VSS VSS VDD VDD data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput38 net38 VSS VSS VDD VDD sample_o sky130_fd_sc_hd__clkbuf_4
Xoutput49 net49 VSS VSS VDD VDD vcm_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_7_45 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_4_135 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_41 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_398_ counter\[6\] net106 counter\[5\] VSS VSS VDD VDD _158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_24 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_73 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ net111 _046_ net4 VSS VSS VDD VDD _109_ sky130_fd_sc_hd__and3_1
X_252_ net110 net97 _064_ VSS VSS VDD VDD _080_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_20 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ net110 VSS VSS VDD VDD _034_ sky130_fd_sc_hd__inv_2
Xfanout95 _061_ VSS VSS VDD VDD net95 sky130_fd_sc_hd__buf_2
XFILLER_0_2_200 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_304_ _094_ _105_ VSS VSS VDD VDD net72 sky130_fd_sc_hd__or2_1
X_235_ net22 _070_ VSS VSS VDD VDD _071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_69 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_218_ net105 net13 counter\[1\] VSS VSS VDD VDD _062_ sky130_fd_sc_hd__or3b_1
Xoutput28 net28 VSS VSS VDD VDD data[1] sky130_fd_sc_hd__clkbuf_4
Xoutput39 net39 VSS VSS VDD VDD vcm_dummy_o sky130_fd_sc_hd__buf_2
XFILLER_0_7_57 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_9_217 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_42 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_250 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_150 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_397_ _136_ result\[7\] _157_ VSS VSS VDD VDD _019_ sky130_fd_sc_hd__mux2_1
X_320_ counter_sample _108_ VSS VSS VDD VDD _000_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_21 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ result\[3\] _064_ VSS VSS VDD VDD net54 sky130_fd_sc_hd__nand2_1
Xfanout96 _061_ VSS VSS VDD VDD net96 sky130_fd_sc_hd__dlymetal6s2s_1
X_182_ counter\[8\] VSS VSS VDD VDD _033_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_74 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_13 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_303_ result\[10\] result\[9\] net105 VSS VSS VDD VDD _105_ sky130_fd_sc_hd__mux2_1
X_234_ net107 counter\[9\] VSS VSS VDD VDD _070_ sky130_fd_sc_hd__nand2b_1
X_217_ net106 net39 VSS VSS VDD VDD _061_ sky130_fd_sc_hd__nand2_1
Xoutput29 net29 VSS VSS VDD VDD data[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_156 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_145 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_7_123 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_43 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_273 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_90 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_396_ _108_ _155_ _156_ _135_ VSS VSS VDD VDD _157_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_48 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_221 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_5_265 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_181_ counter\[9\] VSS VSS VDD VDD _032_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_22 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout97 _060_ VSS VSS VDD VDD net97 sky130_fd_sc_hd__buf_2
X_250_ net95 _079_ net53 VSS VSS VDD VDD net86 sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_75 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_379_ counter\[2\] net101 net99 counter\[1\] VSS VSS VDD VDD _007_ sky130_fd_sc_hd__a22o_1
X_233_ _039_ _069_ net97 VSS VSS VDD VDD net81 sky130_fd_sc_hd__a21o_1
X_302_ _092_ _104_ VSS VSS VDD VDD net71 sky130_fd_sc_hd__or2_1
X_216_ net106 net39 VSS VSS VDD VDD _060_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_26 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_44 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_395_ net109 net106 _033_ VSS VSS VDD VDD _156_ sky130_fd_sc_hd__or3_1
Xfanout98 _060_ VSS VSS VDD VDD net98 sky130_fd_sc_hd__buf_1
X_180_ counter\[11\] VSS VSS VDD VDD _031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_76 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_23 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_378_ counter\[1\] net101 net99 counter\[0\] VSS VSS VDD VDD _006_ sky130_fd_sc_hd__a22o_1
X_301_ result\[9\] result\[8\] net105 VSS VSS VDD VDD _104_ sky130_fd_sc_hd__mux2_1
X_232_ net107 _033_ net21 VSS VSS VDD VDD _069_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_6_55 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ _059_ VSS VSS VDD VDD net39 sky130_fd_sc_hd__inv_2
XFILLER_0_4_139 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_394_ _028_ _032_ counter\[8\] VSS VSS VDD VDD _155_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_201 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_245 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_77 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ state\[1\] state\[0\] VSS VSS VDD VDD _151_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_24 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 _151_ VSS VSS VDD VDD net99 sky130_fd_sc_hd__buf_2
X_446_ net1 _025_ net10 VSS VSS VDD VDD result\[6\] sky130_fd_sc_hd__dfrtp_2
X_300_ _090_ _103_ VSS VSS VDD VDD net70 sky130_fd_sc_hd__or2_1
X_231_ _037_ _068_ net97 VSS VSS VDD VDD net80 sky130_fd_sc_hd__a21o_1
X_429_ net117 _011_ net114 VSS VSS VDD VDD counter\[5\] sky130_fd_sc_hd__dfrtp_4
Xinput1 clk VSS VSS VDD VDD net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_214_ net24 net25 _058_ VSS VSS VDD VDD _059_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_6_56 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_110 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_393_ _154_ net3 _153_ VSS VSS VDD VDD _018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_29 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_78 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_25 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _136_ _150_ _149_ VSS VSS VDD VDD _005_ sky130_fd_sc_hd__mux2_1
X_445_ net115 _024_ net112 VSS VSS VDD VDD result\[3\] sky130_fd_sc_hd__dfrtp_4
X_230_ net20 net109 net103 VSS VSS VDD VDD _068_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_94 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_428_ net115 _010_ net112 VSS VSS VDD VDD counter\[4\] sky130_fd_sc_hd__dfrtp_1
X_359_ net100 _074_ _136_ VSS VSS VDD VDD _138_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_19 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xinput2 comp_n VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_1
X_213_ state\[0\] state\[1\] VSS VSS VDD VDD _058_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_6_57 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_149 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_2_73 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_3_130 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_166 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_392_ _038_ _107_ VSS VSS VDD VDD _154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_258 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_26 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_79 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ result\[0\] _108_ VSS VSS VDD VDD _150_ sky130_fd_sc_hd__and2_1
X_444_ net115 _023_ net112 VSS VSS VDD VDD result\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_73 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_427_ net115 _009_ net112 VSS VSS VDD VDD counter\[3\] sky130_fd_sc_hd__dfrtp_4
X_358_ net100 _074_ VSS VSS VDD VDD _137_ sky130_fd_sc_hd__nand2_1
X_289_ result\[3\] result\[2\] net104 VSS VSS VDD VDD _098_ sky130_fd_sc_hd__mux2_1
Xinput3 comp_p VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_58 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ state\[0\] state\[1\] VSS VSS VDD VDD _057_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_194 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_6_172 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_96 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_391_ net104 _030_ net110 net100 _152_ VSS VSS VDD VDD _153_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_0_27 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ net115 _022_ net112 VSS VSS VDD VDD result\[1\] sky130_fd_sc_hd__dfrtp_4
X_374_ net108 counter\[1\] _075_ _148_ _058_ VSS VSS VDD VDD _149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_30 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xinput4 debug_mux[0] VSS VSS VDD VDD net4 sky130_fd_sc_hd__clkbuf_2
X_357_ net3 _108_ VSS VSS VDD VDD _136_ sky130_fd_sc_hd__and2_1
X_426_ net117 _008_ net114 VSS VSS VDD VDD counter\[2\] sky130_fd_sc_hd__dfrtp_4
X_288_ _078_ _097_ VSS VSS VDD VDD net64 sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_59 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ result\[11\] _056_ net111 _044_ VSS VSS VDD VDD net32 sky130_fd_sc_hd__a2bb2o_1
X_409_ _044_ _107_ VSS VSS VDD VDD _166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_151 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_74 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_390_ net104 counter\[2\] counter\[3\] net100 VSS VSS VDD VDD _152_ sky130_fd_sc_hd__and4bb_1
X_442_ net117 _021_ net114 VSS VSS VDD VDD single_ended_reg sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_28 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_7 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_373_ counter\[0\] counter\[1\] VSS VSS VDD VDD _148_ sky130_fd_sc_hd__nand2b_1
Xinput5 debug_mux[1] VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkbuf_2
X_425_ net117 _007_ net114 VSS VSS VDD VDD counter\[1\] sky130_fd_sc_hd__dfrtp_4
X_356_ net102 _120_ _107_ VSS VSS VDD VDD net36 sky130_fd_sc_hd__a21o_1
X_287_ result\[2\] result\[1\] net104 VSS VSS VDD VDD _097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_108 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_210_ net105 net110 VSS VSS VDD VDD _056_ sky130_fd_sc_hd__or2_1
X_408_ counter\[6\] net103 _029_ net100 _164_ VSS VSS VDD VDD _165_ sky130_fd_sc_hd__a41o_1
X_339_ _046_ net101 _121_ _125_ VSS VSS VDD VDD _126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_122 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_199 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_372_ net3 _147_ _146_ VSS VSS VDD VDD _004_ sky130_fd_sc_hd__mux2_1
X_441_ net115 _020_ net112 VSS VSS VDD VDD result\[4\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_0_29 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ net100 _107_ VSS VSS VDD VDD _135_ sky130_fd_sc_hd__nor2_1
X_424_ net116 _006_ net113 VSS VSS VDD VDD counter\[0\] sky130_fd_sc_hd__dfrtp_1
X_286_ _076_ _096_ VSS VSS VDD VDD net62 sky130_fd_sc_hd__or2_1
Xinput6 debug_mux[2] VSS VSS VDD VDD net6 sky130_fd_sc_hd__buf_1
XFILLER_0_9_194 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_12 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_338_ net4 _108_ VSS VSS VDD VDD _125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_22 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_2_33 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_407_ net109 _027_ net106 net102 VSS VSS VDD VDD _164_ sky130_fd_sc_hd__and4_1
X_269_ result\[6\] _088_ VSS VSS VDD VDD _089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_60 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 vcm_o_i[6] VSS VSS VDD VDD net20 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_440_ net117 _019_ net10 VSS VSS VDD VDD result\[7\] sky130_fd_sc_hd__dfrtp_4
X_371_ _039_ _107_ VSS VSS VDD VDD _147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_251 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_55 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_423_ net115 _005_ net112 VSS VSS VDD VDD result\[0\] sky130_fd_sc_hd__dfrtp_1
X_285_ result\[1\] result\[0\] net104 VSS VSS VDD VDD _096_ sky130_fd_sc_hd__mux2_1
X_354_ net8 _120_ VSS VSS VDD VDD net37 sky130_fd_sc_hd__and2_1
Xinput7 debug_mux[3] VSS VSS VDD VDD net7 sky130_fd_sc_hd__buf_1
X_337_ net3 _046_ _047_ net2 _123_ VSS VSS VDD VDD _124_ sky130_fd_sc_hd__a221o_1
X_199_ net9 VSS VSS VDD VDD _050_ sky130_fd_sc_hd__inv_2
X_406_ _136_ result\[1\] _163_ VSS VSS VDD VDD _022_ sky130_fd_sc_hd__mux2_1
X_268_ counter\[8\] net98 _068_ VSS VSS VDD VDD _088_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_61 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 rst_z VSS VSS VDD VDD net10 sky130_fd_sc_hd__buf_1
Xinput21 vcm_o_i[7] VSS VSS VDD VDD net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_241 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_370_ counter\[8\] _058_ _070_ _145_ counter\[9\] VSS VSS VDD VDD _146_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_45 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_422_ net117 _004_ net114 VSS VSS VDD VDD result\[8\] sky130_fd_sc_hd__dfrtp_2
X_353_ net8 net113 VSS VSS VDD VDD net35 sky130_fd_sc_hd__and2_1
X_284_ _043_ net96 net52 VSS VSS VDD VDD net85 sky130_fd_sc_hd__o21ai_1
Xinput8 en_offset_cal VSS VSS VDD VDD net8 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_30 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ net8 VSS VSS VDD VDD _049_ sky130_fd_sc_hd__inv_2
X_405_ net100 _161_ _162_ _135_ VSS VSS VDD VDD _163_ sky130_fd_sc_hd__a31o_1
X_267_ result\[7\] _068_ VSS VSS VDD VDD net58 sky130_fd_sc_hd__nand2_1
X_336_ counter\[11\] net5 net4 VSS VSS VDD VDD _123_ sky130_fd_sc_hd__and3_1
Xinput11 single_ended VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_62 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 vcm_o_i[8] VSS VSS VDD VDD net22 sky130_fd_sc_hd__clkbuf_1
X_319_ state\[1\] state\[0\] VSS VSS VDD VDD _108_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_2_180 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_8_239 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_5_209 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_1_278 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_421_ net117 _003_ net114 VSS VSS VDD VDD result\[9\] sky130_fd_sc_hd__dfrtp_2
X_283_ net14 _074_ result\[11\] VSS VSS VDD VDD net52 sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_1_31 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ state\[1\] _050_ _129_ counter\[11\] VSS VSS VDD VDD net38 sky130_fd_sc_hd__a211oi_2
Xinput9 en_vcm_sw_o_i VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkbuf_1
X_197_ net7 VSS VSS VDD VDD _048_ sky130_fd_sc_hd__inv_2
X_335_ net5 net4 net34 _121_ VSS VSS VDD VDD _122_ sky130_fd_sc_hd__and4_1
X_266_ net95 _087_ net57 VSS VSS VDD VDD net90 sky130_fd_sc_hd__o21ai_1
X_404_ net105 counter\[1\] counter\[2\] VSS VSS VDD VDD _162_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_134 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_318_ state\[1\] state\[0\] VSS VSS VDD VDD _107_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_7_63 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 start VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 vcm_o_i[9] VSS VSS VDD VDD net23 sky130_fd_sc_hd__clkbuf_1
X_249_ result\[1\] _078_ VSS VSS VDD VDD _079_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_8_Right_8 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_80 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_420_ net115 _002_ net112 VSS VSS VDD VDD result\[10\] sky130_fd_sc_hd__dfrtp_1
X_351_ _029_ _058_ VSS VSS VDD VDD net26 sky130_fd_sc_hd__nor2_1
X_282_ net96 _095_ net61 VSS VSS VDD VDD net94 sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_32 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ net7 net6 VSS VSS VDD VDD _121_ sky130_fd_sc_hd__nor2_1
X_403_ net103 counter\[2\] _030_ VSS VSS VDD VDD _161_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_168 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_265_ result\[5\] _086_ VSS VSS VDD VDD _087_ sky130_fd_sc_hd__nor2_1
X_196_ net4 VSS VSS VDD VDD _047_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_179 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xinput24 vin_n_sw_on VSS VSS VDD VDD net24 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_64 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 vcm_o_i[0] VSS VSS VDD VDD net13 sky130_fd_sc_hd__clkbuf_1
X_179_ counter\[3\] VSS VSS VDD VDD _030_ sky130_fd_sc_hd__inv_2
X_317_ counter\[11\] _106_ VSS VSS VDD VDD net41 sky130_fd_sc_hd__nor2_1
X_248_ counter\[3\] net97 _063_ VSS VSS VDD VDD _078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_281_ result\[9\] _094_ VSS VSS VDD VDD _095_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_33 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _058_ _134_ _107_ counter_sample VSS VSS VDD VDD _174_ sky130_fd_sc_hd__a2bb2o_1
X_402_ net106 net11 _129_ VSS VSS VDD VDD _021_ sky130_fd_sc_hd__mux2_1
X_195_ net5 VSS VSS VDD VDD _046_ sky130_fd_sc_hd__inv_2
X_264_ net109 net97 _067_ VSS VSS VDD VDD _086_ sky130_fd_sc_hd__a21oi_1
X_333_ _049_ _120_ _058_ net116 VSS VSS VDD VDD net34 sky130_fd_sc_hd__a211oi_2
Xinput25 vin_p_sw_on VSS VSS VDD VDD net25 sky130_fd_sc_hd__clkbuf_1
X_316_ counter\[10\] _106_ VSS VSS VDD VDD net50 sky130_fd_sc_hd__nor2_1
Xinput14 vcm_o_i[10] VSS VSS VDD VDD net14 sky130_fd_sc_hd__buf_1
X_247_ result\[2\] _063_ VSS VSS VDD VDD net53 sky130_fd_sc_hd__nand2_1
X_178_ counter\[5\] VSS VSS VDD VDD _029_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_194 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7_275 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_4_212 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_49 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_280_ counter\[11\] net97 _073_ VSS VSS VDD VDD _094_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_34 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_401_ net3 _160_ _159_ VSS VSS VDD VDD _020_ sky130_fd_sc_hd__mux2_1
X_194_ net15 VSS VSS VDD VDD _045_ sky130_fd_sc_hd__inv_2
X_263_ result\[6\] _067_ VSS VSS VDD VDD net57 sky130_fd_sc_hd__nand2_1
X_332_ counter\[0\] counter\[1\] net107 VSS VSS VDD VDD _120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_115 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_177_ net108 VSS VSS VDD VDD _028_ sky130_fd_sc_hd__inv_2
Xinput15 vcm_o_i[1] VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkbuf_1
X_315_ counter\[9\] _106_ VSS VSS VDD VDD net49 sky130_fd_sc_hd__nor2_1
X_246_ net95 _077_ net51 VSS VSS VDD VDD net84 sky130_fd_sc_hd__o21ai_1
X_229_ _035_ _067_ net97 VSS VSS VDD VDD net79 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_45 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _116_ _118_ net7 _114_ VSS VSS VDD VDD _119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_71 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_400_ _042_ _107_ VSS VSS VDD VDD _160_ sky130_fd_sc_hd__nor2_1
X_262_ net56 _085_ VSS VSS VDD VDD net89 sky130_fd_sc_hd__nand2_1
X_193_ result\[5\] VSS VSS VDD VDD _044_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_193 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_314_ counter\[8\] _106_ VSS VSS VDD VDD net48 sky130_fd_sc_hd__nor2_1
Xinput16 vcm_o_i[2] VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkbuf_1
X_176_ counter\[6\] VSS VSS VDD VDD _027_ sky130_fd_sc_hd__inv_2
X_245_ result\[0\] _076_ VSS VSS VDD VDD _077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_141 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_228_ net19 counter\[6\] net103 VSS VSS VDD VDD _067_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_4_46 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_40 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_330_ net109 net5 net4 _117_ VSS VSS VDD VDD _118_ sky130_fd_sc_hd__a31o_1
X_192_ result\[10\] VSS VSS VDD VDD _043_ sky130_fd_sc_hd__inv_2
X_261_ result\[4\] _066_ net97 VSS VSS VDD VDD _085_ sky130_fd_sc_hd__o21ai_1
X_244_ _059_ _075_ _062_ VSS VSS VDD VDD _076_ sky130_fd_sc_hd__o21a_1
X_313_ net109 _106_ VSS VSS VDD VDD net47 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_1_Left_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xinput17 vcm_o_i[3] VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkbuf_1
X_175_ net109 VSS VSS VDD VDD _026_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_51 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_227_ result\[5\] _066_ net96 VSS VSS VDD VDD net78 sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_47 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_259 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_9_83 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_260_ net106 _029_ _044_ net18 VSS VSS VDD VDD net56 sky130_fd_sc_hd__or4_2
X_191_ result\[4\] VSS VSS VDD VDD _042_ sky130_fd_sc_hd__inv_2
X_389_ state\[1\] counter\[11\] net101 VSS VSS VDD VDD _017_ sky130_fd_sc_hd__a21o_1
Xinput18 vcm_o_i[4] VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkbuf_1
X_312_ counter\[6\] _106_ VSS VSS VDD VDD net46 sky130_fd_sc_hd__nor2_1
X_243_ net105 counter\[2\] VSS VSS VDD VDD _075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_132 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_226_ net106 _029_ net18 net95 _027_ VSS VSS VDD VDD _066_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_4_48 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _055_ VSS VSS VDD VDD net31 sky130_fd_sc_hd__inv_2
X_190_ result\[9\] VSS VSS VDD VDD _041_ sky130_fd_sc_hd__inv_2
X_388_ counter\[11\] net101 _151_ counter\[10\] VSS VSS VDD VDD _016_ sky130_fd_sc_hd__a22o_1
Xinput19 vcm_o_i[5] VSS VSS VDD VDD net19 sky130_fd_sc_hd__clkbuf_1
X_311_ counter\[5\] _106_ VSS VSS VDD VDD net45 sky130_fd_sc_hd__nor2_1
X_242_ _036_ _062_ VSS VSS VDD VDD net51 sky130_fd_sc_hd__or2_1
XFILLER_0_3_97 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_225_ result\[4\] _065_ net96 VSS VSS VDD VDD net77 sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_269 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_7_203 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_49 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ result\[10\] result\[4\] net110 VSS VSS VDD VDD _055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_85 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_387_ counter\[10\] net102 net99 counter\[9\] VSS VSS VDD VDD _015_ sky130_fd_sc_hd__a22o_1
X_310_ _056_ _059_ VSS VSS VDD VDD net44 sky130_fd_sc_hd__nor2_1
XFILLER_0_5_153 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_241_ result\[11\] net14 _074_ net96 VSS VSS VDD VDD net74 sky130_fd_sc_hd__o31ai_2
X_439_ net115 _018_ net112 VSS VSS VDD VDD result\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_43 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_224_ net105 _034_ net17 VSS VSS VDD VDD _065_ sky130_fd_sc_hd__or3_1
X_207_ _054_ VSS VSS VDD VDD net30 sky130_fd_sc_hd__inv_2
XFILLER_0_4_229 VDD VSS VDD VSS sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput90 net90 VSS VSS VDD VDD vss_p_o[5] sky130_fd_sc_hd__buf_2
X_386_ counter\[9\] net102 net99 counter\[8\] VSS VSS VDD VDD _014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_187 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_240_ net103 counter\[11\] VSS VSS VDD VDD _074_ sky130_fd_sc_hd__nand2_1
X_369_ net107 counter\[10\] net101 VSS VSS VDD VDD _145_ sky130_fd_sc_hd__nand3_1
X_438_ net117 _174_ net114 VSS VSS VDD VDD state\[1\] sky130_fd_sc_hd__dfrtp_4
Xfanout110 net111 VSS VSS VDD VDD net110 sky130_fd_sc_hd__clkbuf_4
X_223_ _040_ _064_ net97 VSS VSS VDD VDD net76 sky130_fd_sc_hd__a21o_1
XFILLER_0_6_271 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_206_ result\[9\] result\[3\] net110 VSS VSS VDD VDD _054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_45 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_50 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_119 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_6_33 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_385_ counter\[8\] net102 net99 net109 VSS VSS VDD VDD _013_ sky130_fd_sc_hd__a22o_1
Xoutput91 net91 VSS VSS VDD VDD vss_p_o[6] sky130_fd_sc_hd__buf_2
Xoutput80 net80 VSS VSS VDD VDD vss_n_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_5_111 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_144 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_177 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_299_ result\[8\] result\[7\] net104 VSS VSS VDD VDD _103_ sky130_fd_sc_hd__mux2_1
X_437_ net116 _173_ net113 VSS VSS VDD VDD state\[0\] sky130_fd_sc_hd__dfrtp_2
X_368_ net3 _144_ _143_ VSS VSS VDD VDD _003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_23 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_67 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_89 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
Xfanout111 counter\[4\] VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkbuf_2
Xfanout100 net102 VSS VSS VDD VDD net100 sky130_fd_sc_hd__buf_2
X_222_ net105 _030_ net16 VSS VSS VDD VDD _064_ sky130_fd_sc_hd__nor3_1
X_205_ _053_ VSS VSS VDD VDD net29 sky130_fd_sc_hd__inv_2
XFILLER_0_9_66 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_9_44 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_51 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_78 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_384_ net109 net101 net99 counter\[6\] VSS VSS VDD VDD _012_ sky130_fd_sc_hd__a22o_1
Xoutput70 net70 VSS VSS VDD VDD vref_z_p_o[7] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VSS VSS VDD VDD vss_p_o[7] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VSS VSS VDD VDD vss_n_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_5_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_436_ net116 _000_ net113 VSS VSS VDD VDD counter_sample sky130_fd_sc_hd__dfrtp_1
X_367_ _041_ _107_ VSS VSS VDD VDD _144_ sky130_fd_sc_hd__nor2_1
X_298_ _088_ _102_ VSS VSS VDD VDD net69 sky130_fd_sc_hd__or2_1
Xfanout112 net10 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_35 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
Xfanout101 net102 VSS VSS VDD VDD net101 sky130_fd_sc_hd__buf_2
X_221_ _038_ _063_ net97 VSS VSS VDD VDD net75 sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_9_Left_19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_419_ net115 _001_ net112 VSS VSS VDD VDD result\[11\] sky130_fd_sc_hd__dfrtp_1
X_204_ result\[8\] result\[2\] net110 VSS VSS VDD VDD _053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_69 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_0_257 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_52 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_1 net54 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
X_383_ counter\[6\] net100 net99 counter\[5\] VSS VSS VDD VDD _011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_7 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput60 net60 VSS VSS VDD VDD vref_z_n_o[8] sky130_fd_sc_hd__buf_2
Xoutput71 net71 VSS VSS VDD VDD vref_z_p_o[8] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VSS VSS VDD VDD vss_p_o[8] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VSS VSS VDD VDD vss_n_o[8] sky130_fd_sc_hd__buf_2
X_297_ result\[7\] result\[6\] net104 VSS VSS VDD VDD _102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_138 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_435_ net116 _017_ net113 VSS VSS VDD VDD counter\[11\] sky130_fd_sc_hd__dfrtp_4
X_366_ counter\[9\] _058_ _072_ _142_ counter\[10\] VSS VSS VDD VDD _143_ sky130_fd_sc_hd__o32a_1
Xfanout113 net114 VSS VSS VDD VDD net113 sky130_fd_sc_hd__clkbuf_4
Xfanout102 _057_ VSS VSS VDD VDD net102 sky130_fd_sc_hd__clkbuf_2
X_220_ net103 counter\[2\] _045_ VSS VSS VDD VDD _063_ sky130_fd_sc_hd__and3_1
X_418_ _172_ net3 _171_ VSS VSS VDD VDD _025_ sky130_fd_sc_hd__mux2_1
X_349_ _130_ _131_ _132_ _133_ VSS VSS VDD VDD _134_ sky130_fd_sc_hd__and4_1
X_203_ _052_ VSS VSS VDD VDD net28 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_53 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_2 net56 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_6_47 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput61 net61 VSS VSS VDD VDD vref_z_n_o[9] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VSS VSS VDD VDD vref_z_p_o[9] sky130_fd_sc_hd__buf_2
X_382_ net111 net99 net26 VSS VSS VDD VDD _010_ sky130_fd_sc_hd__a21o_1
Xoutput50 net50 VSS VSS VDD VDD vcm_o[9] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VSS VSS VDD VDD vss_p_o[9] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VSS VSS VDD VDD vss_n_o[9] sky130_fd_sc_hd__buf_2
X_434_ net116 _016_ net113 VSS VSS VDD VDD counter\[10\] sky130_fd_sc_hd__dfrtp_4
X_296_ _086_ _101_ VSS VSS VDD VDD net68 sky130_fd_sc_hd__or2_1
X_365_ net103 _031_ _058_ VSS VSS VDD VDD _142_ sky130_fd_sc_hd__or3_1
Xfanout114 net10 VSS VSS VDD VDD net114 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_0_Left_10 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xfanout103 _028_ VSS VSS VDD VDD net103 sky130_fd_sc_hd__buf_2
X_279_ result\[10\] _073_ VSS VSS VDD VDD net61 sky130_fd_sc_hd__nand2_1
X_417_ _035_ _107_ VSS VSS VDD VDD _172_ sky130_fd_sc_hd__nor2_1
X_348_ net107 counter\[0\] VSS VSS VDD VDD _133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_231 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_202_ result\[7\] result\[1\] net110 VSS VSS VDD VDD _052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_49 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_54 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
*XANTENNA_3 net57 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_8_156 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_381_ net111 net100 net99 counter\[3\] VSS VSS VDD VDD _009_ sky130_fd_sc_hd__a22o_1
Xoutput40 net40 VSS VSS VDD VDD vcm_o[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VSS VSS VDD VDD vss_p_o[0] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VSS VSS VDD VDD vss_n_o[0] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VSS VSS VDD VDD vref_z_p_o[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VSS VSS VDD VDD vref_z_n_o[0] sky130_fd_sc_hd__buf_2
X_433_ net116 _015_ net113 VSS VSS VDD VDD counter\[9\] sky130_fd_sc_hd__dfrtp_4
X_364_ _136_ result\[10\] _141_ VSS VSS VDD VDD _002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_107 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_295_ result\[6\] result\[5\] net104 VSS VSS VDD VDD _101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_240 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xfanout115 net1 VSS VSS VDD VDD net115 sky130_fd_sc_hd__buf_2
Xfanout104 net105 VSS VSS VDD VDD net104 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_65 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_278_ net95 _093_ net60 VSS VSS VDD VDD net93 sky130_fd_sc_hd__o21ai_1
X_347_ counter\[9\] counter\[8\] net111 VSS VSS VDD VDD _132_ sky130_fd_sc_hd__and3_1
X_416_ _026_ net107 counter\[8\] net101 _170_ VSS VSS VDD VDD _171_ sky130_fd_sc_hd__a41o_1
X_201_ _051_ VSS VSS VDD VDD net27 sky130_fd_sc_hd__inv_2
XFILLER_0_9_26 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
*XANTENNA_4 net73 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
Xoutput52 net52 VSS VSS VDD VDD vref_z_n_o[10] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VSS VSS VDD VDD data[3] sky130_fd_sc_hd__clkbuf_4
X_380_ counter\[3\] net101 net99 counter\[2\] VSS VSS VDD VDD _008_ sky130_fd_sc_hd__a22o_1
Xoutput41 net41 VSS VSS VDD VDD vcm_o[10] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VSS VSS VDD VDD vref_z_p_o[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VSS VSS VDD VDD vss_p_o[10] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VSS VSS VDD VDD vss_n_o[10] sky130_fd_sc_hd__buf_2
.ends

