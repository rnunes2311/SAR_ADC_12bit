magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -1951 845 -1889 851
rect -1823 845 -1761 851
rect -1695 845 -1633 851
rect -1567 845 -1505 851
rect -1439 845 -1377 851
rect -1311 845 -1249 851
rect -1183 845 -1121 851
rect -1055 845 -993 851
rect -927 845 -865 851
rect -799 845 -737 851
rect -671 845 -609 851
rect -543 845 -481 851
rect -415 845 -353 851
rect -287 845 -225 851
rect -159 845 -97 851
rect -31 845 31 851
rect 97 845 159 851
rect 225 845 287 851
rect 353 845 415 851
rect 481 845 543 851
rect 609 845 671 851
rect 737 845 799 851
rect 865 845 927 851
rect 993 845 1055 851
rect 1121 845 1183 851
rect 1249 845 1311 851
rect 1377 845 1439 851
rect 1505 845 1567 851
rect 1633 845 1695 851
rect 1761 845 1823 851
rect 1889 845 1951 851
rect -1951 811 -1939 845
rect -1823 811 -1811 845
rect -1695 811 -1683 845
rect -1567 811 -1555 845
rect -1439 811 -1427 845
rect -1311 811 -1299 845
rect -1183 811 -1171 845
rect -1055 811 -1043 845
rect -927 811 -915 845
rect -799 811 -787 845
rect -671 811 -659 845
rect -543 811 -531 845
rect -415 811 -403 845
rect -287 811 -275 845
rect -159 811 -147 845
rect -31 811 -19 845
rect 97 811 109 845
rect 225 811 237 845
rect 353 811 365 845
rect 481 811 493 845
rect 609 811 621 845
rect 737 811 749 845
rect 865 811 877 845
rect 993 811 1005 845
rect 1121 811 1133 845
rect 1249 811 1261 845
rect 1377 811 1389 845
rect 1505 811 1517 845
rect 1633 811 1645 845
rect 1761 811 1773 845
rect 1889 811 1901 845
rect -1951 805 -1889 811
rect -1823 805 -1761 811
rect -1695 805 -1633 811
rect -1567 805 -1505 811
rect -1439 805 -1377 811
rect -1311 805 -1249 811
rect -1183 805 -1121 811
rect -1055 805 -993 811
rect -927 805 -865 811
rect -799 805 -737 811
rect -671 805 -609 811
rect -543 805 -481 811
rect -415 805 -353 811
rect -287 805 -225 811
rect -159 805 -97 811
rect -31 805 31 811
rect 97 805 159 811
rect 225 805 287 811
rect 353 805 415 811
rect 481 805 543 811
rect 609 805 671 811
rect 737 805 799 811
rect 865 805 927 811
rect 993 805 1055 811
rect 1121 805 1183 811
rect 1249 805 1311 811
rect 1377 805 1439 811
rect 1505 805 1567 811
rect 1633 805 1695 811
rect 1761 805 1823 811
rect 1889 805 1951 811
<< nwell >>
rect -2151 -984 3611 984
<< pmoslvt >>
rect -1955 -836 -1885 764
rect -1827 -836 -1757 764
rect -1699 -836 -1629 764
rect -1571 -836 -1501 764
rect -1443 -836 -1373 764
rect -1315 -836 -1245 764
rect -1187 -836 -1117 764
rect -1059 -836 -989 764
rect -931 -836 -861 764
rect -803 -836 -733 764
rect -675 -836 -605 764
rect -547 -836 -477 764
rect -419 -836 -349 764
rect -291 -836 -221 764
rect -163 -836 -93 764
rect -35 -836 35 764
rect 93 -836 163 764
rect 221 -836 291 764
rect 349 -836 419 764
rect 477 -836 547 764
rect 605 -836 675 764
rect 733 -836 803 764
rect 861 -836 931 764
rect 989 -836 1059 764
rect 1117 -836 1187 764
rect 1245 -836 1315 764
rect 1373 -836 1443 764
rect 1501 -836 1571 764
rect 1629 -836 1699 764
rect 1757 -836 1827 764
rect 1885 -836 1955 764
<< pdiff >>
rect -2013 752 -1955 764
rect -2013 -824 -2001 752
rect -1967 -824 -1955 752
rect -2013 -836 -1955 -824
rect -1885 752 -1827 764
rect -1885 -824 -1873 752
rect -1839 -824 -1827 752
rect -1885 -836 -1827 -824
rect -1757 752 -1699 764
rect -1757 -824 -1745 752
rect -1711 -824 -1699 752
rect -1757 -836 -1699 -824
rect -1629 752 -1571 764
rect -1629 -824 -1617 752
rect -1583 -824 -1571 752
rect -1629 -836 -1571 -824
rect -1501 752 -1443 764
rect -1501 -824 -1489 752
rect -1455 -824 -1443 752
rect -1501 -836 -1443 -824
rect -1373 752 -1315 764
rect -1373 -824 -1361 752
rect -1327 -824 -1315 752
rect -1373 -836 -1315 -824
rect -1245 752 -1187 764
rect -1245 -824 -1233 752
rect -1199 -824 -1187 752
rect -1245 -836 -1187 -824
rect -1117 752 -1059 764
rect -1117 -824 -1105 752
rect -1071 -824 -1059 752
rect -1117 -836 -1059 -824
rect -989 752 -931 764
rect -989 -824 -977 752
rect -943 -824 -931 752
rect -989 -836 -931 -824
rect -861 752 -803 764
rect -861 -824 -849 752
rect -815 -824 -803 752
rect -861 -836 -803 -824
rect -733 752 -675 764
rect -733 -824 -721 752
rect -687 -824 -675 752
rect -733 -836 -675 -824
rect -605 752 -547 764
rect -605 -824 -593 752
rect -559 -824 -547 752
rect -605 -836 -547 -824
rect -477 752 -419 764
rect -477 -824 -465 752
rect -431 -824 -419 752
rect -477 -836 -419 -824
rect -349 752 -291 764
rect -349 -824 -337 752
rect -303 -824 -291 752
rect -349 -836 -291 -824
rect -221 752 -163 764
rect -221 -824 -209 752
rect -175 -824 -163 752
rect -221 -836 -163 -824
rect -93 752 -35 764
rect -93 -824 -81 752
rect -47 -824 -35 752
rect -93 -836 -35 -824
rect 35 752 93 764
rect 35 -824 47 752
rect 81 -824 93 752
rect 35 -836 93 -824
rect 163 752 221 764
rect 163 -824 175 752
rect 209 -824 221 752
rect 163 -836 221 -824
rect 291 752 349 764
rect 291 -824 303 752
rect 337 -824 349 752
rect 291 -836 349 -824
rect 419 752 477 764
rect 419 -824 431 752
rect 465 -824 477 752
rect 419 -836 477 -824
rect 547 752 605 764
rect 547 -824 559 752
rect 593 -824 605 752
rect 547 -836 605 -824
rect 675 752 733 764
rect 675 -824 687 752
rect 721 -824 733 752
rect 675 -836 733 -824
rect 803 752 861 764
rect 803 -824 815 752
rect 849 -824 861 752
rect 803 -836 861 -824
rect 931 752 989 764
rect 931 -824 943 752
rect 977 -824 989 752
rect 931 -836 989 -824
rect 1059 752 1117 764
rect 1059 -824 1071 752
rect 1105 -824 1117 752
rect 1059 -836 1117 -824
rect 1187 752 1245 764
rect 1187 -824 1199 752
rect 1233 -824 1245 752
rect 1187 -836 1245 -824
rect 1315 752 1373 764
rect 1315 -824 1327 752
rect 1361 -824 1373 752
rect 1315 -836 1373 -824
rect 1443 752 1501 764
rect 1443 -824 1455 752
rect 1489 -824 1501 752
rect 1443 -836 1501 -824
rect 1571 752 1629 764
rect 1571 -824 1583 752
rect 1617 -824 1629 752
rect 1571 -836 1629 -824
rect 1699 752 1757 764
rect 1699 -824 1711 752
rect 1745 -824 1757 752
rect 1699 -836 1757 -824
rect 1827 752 1885 764
rect 1827 -824 1839 752
rect 1873 -824 1885 752
rect 1827 -836 1885 -824
rect 1955 752 2013 764
rect 1955 -824 1967 752
rect 2001 -824 2013 752
rect 1955 -836 2013 -824
<< pdiffc >>
rect -2001 -824 -1967 752
rect -1873 -824 -1839 752
rect -1745 -824 -1711 752
rect -1617 -824 -1583 752
rect -1489 -824 -1455 752
rect -1361 -824 -1327 752
rect -1233 -824 -1199 752
rect -1105 -824 -1071 752
rect -977 -824 -943 752
rect -849 -824 -815 752
rect -721 -824 -687 752
rect -593 -824 -559 752
rect -465 -824 -431 752
rect -337 -824 -303 752
rect -209 -824 -175 752
rect -81 -824 -47 752
rect 47 -824 81 752
rect 175 -824 209 752
rect 303 -824 337 752
rect 431 -824 465 752
rect 559 -824 593 752
rect 687 -824 721 752
rect 815 -824 849 752
rect 943 -824 977 752
rect 1071 -824 1105 752
rect 1199 -824 1233 752
rect 1327 -824 1361 752
rect 1455 -824 1489 752
rect 1583 -824 1617 752
rect 1711 -824 1745 752
rect 1839 -824 1873 752
rect 1967 -824 2001 752
<< nsubdiff >>
rect -2115 914 -2019 948
rect 3509 914 3575 948
rect -2115 851 -2081 914
rect 3541 851 3575 914
rect -2115 -914 -2081 -851
rect 3541 -914 3575 -851
rect -2115 -948 -2019 -914
rect 3449 -948 3575 -914
<< nsubdiffcont >>
rect -2019 914 3509 948
rect -2115 -851 -2081 851
rect 3541 -851 3575 851
rect -2019 -948 3449 -914
<< poly >>
rect -1955 845 -1885 861
rect -1955 811 -1939 845
rect -1901 811 -1885 845
rect -1955 764 -1885 811
rect -1827 845 -1757 861
rect -1827 811 -1811 845
rect -1773 811 -1757 845
rect -1827 764 -1757 811
rect -1699 845 -1629 861
rect -1699 811 -1683 845
rect -1645 811 -1629 845
rect -1699 764 -1629 811
rect -1571 845 -1501 861
rect -1571 811 -1555 845
rect -1517 811 -1501 845
rect -1571 764 -1501 811
rect -1443 845 -1373 861
rect -1443 811 -1427 845
rect -1389 811 -1373 845
rect -1443 764 -1373 811
rect -1315 845 -1245 861
rect -1315 811 -1299 845
rect -1261 811 -1245 845
rect -1315 764 -1245 811
rect -1187 845 -1117 861
rect -1187 811 -1171 845
rect -1133 811 -1117 845
rect -1187 764 -1117 811
rect -1059 845 -989 861
rect -1059 811 -1043 845
rect -1005 811 -989 845
rect -1059 764 -989 811
rect -931 845 -861 861
rect -931 811 -915 845
rect -877 811 -861 845
rect -931 764 -861 811
rect -803 845 -733 861
rect -803 811 -787 845
rect -749 811 -733 845
rect -803 764 -733 811
rect -675 845 -605 861
rect -675 811 -659 845
rect -621 811 -605 845
rect -675 764 -605 811
rect -547 845 -477 861
rect -547 811 -531 845
rect -493 811 -477 845
rect -547 764 -477 811
rect -419 845 -349 861
rect -419 811 -403 845
rect -365 811 -349 845
rect -419 764 -349 811
rect -291 845 -221 861
rect -291 811 -275 845
rect -237 811 -221 845
rect -291 764 -221 811
rect -163 845 -93 861
rect -163 811 -147 845
rect -109 811 -93 845
rect -163 764 -93 811
rect -35 845 35 861
rect -35 811 -19 845
rect 19 811 35 845
rect -35 764 35 811
rect 93 845 163 861
rect 93 811 109 845
rect 147 811 163 845
rect 93 764 163 811
rect 221 845 291 861
rect 221 811 237 845
rect 275 811 291 845
rect 221 764 291 811
rect 349 845 419 861
rect 349 811 365 845
rect 403 811 419 845
rect 349 764 419 811
rect 477 845 547 861
rect 477 811 493 845
rect 531 811 547 845
rect 477 764 547 811
rect 605 845 675 861
rect 605 811 621 845
rect 659 811 675 845
rect 605 764 675 811
rect 733 845 803 861
rect 733 811 749 845
rect 787 811 803 845
rect 733 764 803 811
rect 861 845 931 861
rect 861 811 877 845
rect 915 811 931 845
rect 861 764 931 811
rect 989 845 1059 861
rect 989 811 1005 845
rect 1043 811 1059 845
rect 989 764 1059 811
rect 1117 845 1187 861
rect 1117 811 1133 845
rect 1171 811 1187 845
rect 1117 764 1187 811
rect 1245 845 1315 861
rect 1245 811 1261 845
rect 1299 811 1315 845
rect 1245 764 1315 811
rect 1373 845 1443 861
rect 1373 811 1389 845
rect 1427 811 1443 845
rect 1373 764 1443 811
rect 1501 845 1571 861
rect 1501 811 1517 845
rect 1555 811 1571 845
rect 1501 764 1571 811
rect 1629 845 1699 861
rect 1629 811 1645 845
rect 1683 811 1699 845
rect 1629 764 1699 811
rect 1757 845 1827 861
rect 1757 811 1773 845
rect 1811 811 1827 845
rect 1757 764 1827 811
rect 1885 845 1955 861
rect 1885 811 1901 845
rect 1939 811 1955 845
rect 1885 764 1955 811
rect -1955 -862 -1885 -836
rect -1827 -862 -1757 -836
rect -1699 -862 -1629 -836
rect -1571 -862 -1501 -836
rect -1443 -862 -1373 -836
rect -1315 -862 -1245 -836
rect -1187 -862 -1117 -836
rect -1059 -862 -989 -836
rect -931 -862 -861 -836
rect -803 -862 -733 -836
rect -675 -862 -605 -836
rect -547 -862 -477 -836
rect -419 -862 -349 -836
rect -291 -862 -221 -836
rect -163 -862 -93 -836
rect -35 -862 35 -836
rect 93 -862 163 -836
rect 221 -862 291 -836
rect 349 -862 419 -836
rect 477 -862 547 -836
rect 605 -862 675 -836
rect 733 -862 803 -836
rect 861 -862 931 -836
rect 989 -862 1059 -836
rect 1117 -862 1187 -836
rect 1245 -862 1315 -836
rect 1373 -862 1443 -836
rect 1501 -862 1571 -836
rect 1629 -862 1699 -836
rect 1757 -862 1827 -836
rect 1885 -862 1955 -836
<< polycont >>
rect -1939 811 -1901 845
rect -1811 811 -1773 845
rect -1683 811 -1645 845
rect -1555 811 -1517 845
rect -1427 811 -1389 845
rect -1299 811 -1261 845
rect -1171 811 -1133 845
rect -1043 811 -1005 845
rect -915 811 -877 845
rect -787 811 -749 845
rect -659 811 -621 845
rect -531 811 -493 845
rect -403 811 -365 845
rect -275 811 -237 845
rect -147 811 -109 845
rect -19 811 19 845
rect 109 811 147 845
rect 237 811 275 845
rect 365 811 403 845
rect 493 811 531 845
rect 621 811 659 845
rect 749 811 787 845
rect 877 811 915 845
rect 1005 811 1043 845
rect 1133 811 1171 845
rect 1261 811 1299 845
rect 1389 811 1427 845
rect 1517 811 1555 845
rect 1645 811 1683 845
rect 1773 811 1811 845
rect 1901 811 1939 845
<< locali >>
rect -2115 914 -2019 948
rect 3509 914 3575 948
rect -2115 851 -2081 914
rect 3541 851 3575 914
rect -1955 811 -1939 845
rect -1901 811 -1885 845
rect -1827 811 -1811 845
rect -1773 811 -1757 845
rect -1699 811 -1683 845
rect -1645 811 -1629 845
rect -1571 811 -1555 845
rect -1517 811 -1501 845
rect -1443 811 -1427 845
rect -1389 811 -1373 845
rect -1315 811 -1299 845
rect -1261 811 -1245 845
rect -1187 811 -1171 845
rect -1133 811 -1117 845
rect -1059 811 -1043 845
rect -1005 811 -989 845
rect -931 811 -915 845
rect -877 811 -861 845
rect -803 811 -787 845
rect -749 811 -733 845
rect -675 811 -659 845
rect -621 811 -605 845
rect -547 811 -531 845
rect -493 811 -477 845
rect -419 811 -403 845
rect -365 811 -349 845
rect -291 811 -275 845
rect -237 811 -221 845
rect -163 811 -147 845
rect -109 811 -93 845
rect -35 811 -19 845
rect 19 811 35 845
rect 93 811 109 845
rect 147 811 163 845
rect 221 811 237 845
rect 275 811 291 845
rect 349 811 365 845
rect 403 811 419 845
rect 477 811 493 845
rect 531 811 547 845
rect 605 811 621 845
rect 659 811 675 845
rect 733 811 749 845
rect 787 811 803 845
rect 861 811 877 845
rect 915 811 931 845
rect 989 811 1005 845
rect 1043 811 1059 845
rect 1117 811 1133 845
rect 1171 811 1187 845
rect 1245 811 1261 845
rect 1299 811 1315 845
rect 1373 811 1389 845
rect 1427 811 1443 845
rect 1501 811 1517 845
rect 1555 811 1571 845
rect 1629 811 1645 845
rect 1683 811 1699 845
rect 1757 811 1773 845
rect 1811 811 1827 845
rect 1885 811 1901 845
rect 1939 811 1955 845
rect -2001 752 -1967 768
rect -2001 -840 -1967 -824
rect -1873 752 -1839 768
rect -1873 -840 -1839 -824
rect -1745 752 -1711 768
rect -1745 -840 -1711 -824
rect -1617 752 -1583 768
rect -1617 -840 -1583 -824
rect -1489 752 -1455 768
rect -1489 -840 -1455 -824
rect -1361 752 -1327 768
rect -1361 -840 -1327 -824
rect -1233 752 -1199 768
rect -1233 -840 -1199 -824
rect -1105 752 -1071 768
rect -1105 -840 -1071 -824
rect -977 752 -943 768
rect -977 -840 -943 -824
rect -849 752 -815 768
rect -849 -840 -815 -824
rect -721 752 -687 768
rect -721 -840 -687 -824
rect -593 752 -559 768
rect -593 -840 -559 -824
rect -465 752 -431 768
rect -465 -840 -431 -824
rect -337 752 -303 768
rect -337 -840 -303 -824
rect -209 752 -175 768
rect -209 -840 -175 -824
rect -81 752 -47 768
rect -81 -840 -47 -824
rect 47 752 81 768
rect 47 -840 81 -824
rect 175 752 209 768
rect 175 -840 209 -824
rect 303 752 337 768
rect 303 -840 337 -824
rect 431 752 465 768
rect 431 -840 465 -824
rect 559 752 593 768
rect 559 -840 593 -824
rect 687 752 721 768
rect 687 -840 721 -824
rect 815 752 849 768
rect 815 -840 849 -824
rect 943 752 977 768
rect 943 -840 977 -824
rect 1071 752 1105 768
rect 1071 -840 1105 -824
rect 1199 752 1233 768
rect 1199 -840 1233 -824
rect 1327 752 1361 768
rect 1327 -840 1361 -824
rect 1455 752 1489 768
rect 1455 -840 1489 -824
rect 1583 752 1617 768
rect 1583 -840 1617 -824
rect 1711 752 1745 768
rect 1711 -840 1745 -824
rect 1839 752 1873 768
rect 1839 -840 1873 -824
rect 1967 752 2001 768
rect 1967 -840 2001 -824
rect -2115 -914 -2081 -851
rect 3541 -914 3575 -851
rect -2115 -948 -2019 -914
rect 3449 -948 3575 -914
<< viali >>
rect -1939 811 -1901 845
rect -1811 811 -1773 845
rect -1683 811 -1645 845
rect -1555 811 -1517 845
rect -1427 811 -1389 845
rect -1299 811 -1261 845
rect -1171 811 -1133 845
rect -1043 811 -1005 845
rect -915 811 -877 845
rect -787 811 -749 845
rect -659 811 -621 845
rect -531 811 -493 845
rect -403 811 -365 845
rect -275 811 -237 845
rect -147 811 -109 845
rect -19 811 19 845
rect 109 811 147 845
rect 237 811 275 845
rect 365 811 403 845
rect 493 811 531 845
rect 621 811 659 845
rect 749 811 787 845
rect 877 811 915 845
rect 1005 811 1043 845
rect 1133 811 1171 845
rect 1261 811 1299 845
rect 1389 811 1427 845
rect 1517 811 1555 845
rect 1645 811 1683 845
rect 1773 811 1811 845
rect 1901 811 1939 845
rect -2001 -824 -1967 752
rect -1873 -824 -1839 752
rect -1745 -824 -1711 752
rect -1617 -824 -1583 752
rect -1489 -824 -1455 752
rect -1361 -824 -1327 752
rect -1233 -824 -1199 752
rect -1105 -824 -1071 752
rect -977 -824 -943 752
rect -849 -824 -815 752
rect -721 -824 -687 752
rect -593 -824 -559 752
rect -465 -824 -431 752
rect -337 -824 -303 752
rect -209 -824 -175 752
rect -81 -824 -47 752
rect 47 -824 81 752
rect 175 -824 209 752
rect 303 -824 337 752
rect 431 -824 465 752
rect 559 -824 593 752
rect 687 -824 721 752
rect 815 -824 849 752
rect 943 -824 977 752
rect 1071 -824 1105 752
rect 1199 -824 1233 752
rect 1327 -824 1361 752
rect 1455 -824 1489 752
rect 1583 -824 1617 752
rect 1711 -824 1745 752
rect 1839 -824 1873 752
rect 1967 -824 2001 752
<< metal1 >>
rect -1951 845 -1889 851
rect -1951 811 -1939 845
rect -1901 811 -1889 845
rect -1951 805 -1889 811
rect -1823 845 -1761 851
rect -1823 811 -1811 845
rect -1773 811 -1761 845
rect -1823 805 -1761 811
rect -1695 845 -1633 851
rect -1695 811 -1683 845
rect -1645 811 -1633 845
rect -1695 805 -1633 811
rect -1567 845 -1505 851
rect -1567 811 -1555 845
rect -1517 811 -1505 845
rect -1567 805 -1505 811
rect -1439 845 -1377 851
rect -1439 811 -1427 845
rect -1389 811 -1377 845
rect -1439 805 -1377 811
rect -1311 845 -1249 851
rect -1311 811 -1299 845
rect -1261 811 -1249 845
rect -1311 805 -1249 811
rect -1183 845 -1121 851
rect -1183 811 -1171 845
rect -1133 811 -1121 845
rect -1183 805 -1121 811
rect -1055 845 -993 851
rect -1055 811 -1043 845
rect -1005 811 -993 845
rect -1055 805 -993 811
rect -927 845 -865 851
rect -927 811 -915 845
rect -877 811 -865 845
rect -927 805 -865 811
rect -799 845 -737 851
rect -799 811 -787 845
rect -749 811 -737 845
rect -799 805 -737 811
rect -671 845 -609 851
rect -671 811 -659 845
rect -621 811 -609 845
rect -671 805 -609 811
rect -543 845 -481 851
rect -543 811 -531 845
rect -493 811 -481 845
rect -543 805 -481 811
rect -415 845 -353 851
rect -415 811 -403 845
rect -365 811 -353 845
rect -415 805 -353 811
rect -287 845 -225 851
rect -287 811 -275 845
rect -237 811 -225 845
rect -287 805 -225 811
rect -159 845 -97 851
rect -159 811 -147 845
rect -109 811 -97 845
rect -159 805 -97 811
rect -31 845 31 851
rect -31 811 -19 845
rect 19 811 31 845
rect -31 805 31 811
rect 97 845 159 851
rect 97 811 109 845
rect 147 811 159 845
rect 97 805 159 811
rect 225 845 287 851
rect 225 811 237 845
rect 275 811 287 845
rect 225 805 287 811
rect 353 845 415 851
rect 353 811 365 845
rect 403 811 415 845
rect 353 805 415 811
rect 481 845 543 851
rect 481 811 493 845
rect 531 811 543 845
rect 481 805 543 811
rect 609 845 671 851
rect 609 811 621 845
rect 659 811 671 845
rect 609 805 671 811
rect 737 845 799 851
rect 737 811 749 845
rect 787 811 799 845
rect 737 805 799 811
rect 865 845 927 851
rect 865 811 877 845
rect 915 811 927 845
rect 865 805 927 811
rect 993 845 1055 851
rect 993 811 1005 845
rect 1043 811 1055 845
rect 993 805 1055 811
rect 1121 845 1183 851
rect 1121 811 1133 845
rect 1171 811 1183 845
rect 1121 805 1183 811
rect 1249 845 1311 851
rect 1249 811 1261 845
rect 1299 811 1311 845
rect 1249 805 1311 811
rect 1377 845 1439 851
rect 1377 811 1389 845
rect 1427 811 1439 845
rect 1377 805 1439 811
rect 1505 845 1567 851
rect 1505 811 1517 845
rect 1555 811 1567 845
rect 1505 805 1567 811
rect 1633 845 1695 851
rect 1633 811 1645 845
rect 1683 811 1695 845
rect 1633 805 1695 811
rect 1761 845 1823 851
rect 1761 811 1773 845
rect 1811 811 1823 845
rect 1761 805 1823 811
rect 1889 845 1951 851
rect 1889 811 1901 845
rect 1939 811 1951 845
rect 1889 805 1951 811
rect -2007 752 -1961 764
rect -2007 -824 -2001 752
rect -1967 -824 -1961 752
rect -2007 -836 -1961 -824
rect -1879 752 -1833 764
rect -1879 -824 -1873 752
rect -1839 -824 -1833 752
rect -1879 -836 -1833 -824
rect -1751 752 -1705 764
rect -1751 -824 -1745 752
rect -1711 -824 -1705 752
rect -1751 -836 -1705 -824
rect -1623 752 -1577 764
rect -1623 -824 -1617 752
rect -1583 -824 -1577 752
rect -1623 -836 -1577 -824
rect -1495 752 -1449 764
rect -1495 -824 -1489 752
rect -1455 -824 -1449 752
rect -1495 -836 -1449 -824
rect -1367 752 -1321 764
rect -1367 -824 -1361 752
rect -1327 -824 -1321 752
rect -1367 -836 -1321 -824
rect -1239 752 -1193 764
rect -1239 -824 -1233 752
rect -1199 -824 -1193 752
rect -1239 -836 -1193 -824
rect -1111 752 -1065 764
rect -1111 -824 -1105 752
rect -1071 -824 -1065 752
rect -1111 -836 -1065 -824
rect -983 752 -937 764
rect -983 -824 -977 752
rect -943 -824 -937 752
rect -983 -836 -937 -824
rect -855 752 -809 764
rect -855 -824 -849 752
rect -815 -824 -809 752
rect -855 -836 -809 -824
rect -727 752 -681 764
rect -727 -824 -721 752
rect -687 -824 -681 752
rect -727 -836 -681 -824
rect -599 752 -553 764
rect -599 -824 -593 752
rect -559 -824 -553 752
rect -599 -836 -553 -824
rect -471 752 -425 764
rect -471 -824 -465 752
rect -431 -824 -425 752
rect -471 -836 -425 -824
rect -343 752 -297 764
rect -343 -824 -337 752
rect -303 -824 -297 752
rect -343 -836 -297 -824
rect -215 752 -169 764
rect -215 -824 -209 752
rect -175 -824 -169 752
rect -215 -836 -169 -824
rect -87 752 -41 764
rect -87 -824 -81 752
rect -47 -824 -41 752
rect -87 -836 -41 -824
rect 41 752 87 764
rect 41 -824 47 752
rect 81 -824 87 752
rect 41 -836 87 -824
rect 169 752 215 764
rect 169 -824 175 752
rect 209 -824 215 752
rect 169 -836 215 -824
rect 297 752 343 764
rect 297 -824 303 752
rect 337 -824 343 752
rect 297 -836 343 -824
rect 425 752 471 764
rect 425 -824 431 752
rect 465 -824 471 752
rect 425 -836 471 -824
rect 553 752 599 764
rect 553 -824 559 752
rect 593 -824 599 752
rect 553 -836 599 -824
rect 681 752 727 764
rect 681 -824 687 752
rect 721 -824 727 752
rect 681 -836 727 -824
rect 809 752 855 764
rect 809 -824 815 752
rect 849 -824 855 752
rect 809 -836 855 -824
rect 937 752 983 764
rect 937 -824 943 752
rect 977 -824 983 752
rect 937 -836 983 -824
rect 1065 752 1111 764
rect 1065 -824 1071 752
rect 1105 -824 1111 752
rect 1065 -836 1111 -824
rect 1193 752 1239 764
rect 1193 -824 1199 752
rect 1233 -824 1239 752
rect 1193 -836 1239 -824
rect 1321 752 1367 764
rect 1321 -824 1327 752
rect 1361 -824 1367 752
rect 1321 -836 1367 -824
rect 1449 752 1495 764
rect 1449 -824 1455 752
rect 1489 -824 1495 752
rect 1449 -836 1495 -824
rect 1577 752 1623 764
rect 1577 -824 1583 752
rect 1617 -824 1623 752
rect 1577 -836 1623 -824
rect 1705 752 1751 764
rect 1705 -824 1711 752
rect 1745 -824 1751 752
rect 1705 -836 1751 -824
rect 1833 752 1879 764
rect 1833 -824 1839 752
rect 1873 -824 1879 752
rect 1833 -836 1879 -824
rect 1961 752 2007 764
rect 1961 -824 1967 752
rect 2001 -824 2007 752
rect 1961 -836 2007 -824
rect 3530 -916 3580 984
rect 3510 -986 3580 -916
<< properties >>
string FIXED_BBOX -2098 -931 2098 931
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8 l 0.35 m 1 nf 31 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
