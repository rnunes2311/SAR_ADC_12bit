* SPICE3 file created from SAR_ADC_12bit_flat.ext - technology: sky130A
* Changed subckt name from SAR_ADC_12bit_flat to SAR_ADC_12bit

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START
+ EN_OFFSET_CAL CLK VREF_GND SINGLE_ENDED
X0 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1 a_13076_44458# a_13259_45724# a_13296_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4 VSS a_12427_45724# a_10490_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X9 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=361.2627 ps=3.22652k w=10 l=10
X10 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X11 VDD a_2903_42308# a_3080_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X13 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X14 VDD a_12861_44030# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VSS a_1209_43370# a_n1557_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X17 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X18 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X19 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X20 a_16237_45028# a_16147_45260# a_16019_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VDD a_n755_45592# a_1176_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X23 a_6756_44260# a_5937_45572# a_6453_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X24 a_n1533_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X25 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X26 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X27 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X28 a_15868_43402# a_15681_43442# a_15781_43660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X29 a_8103_44636# a_8375_44464# a_8333_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X31 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X32 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X33 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X34 VSS a_16327_47482# a_16377_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 a_2437_43646# a_n443_46116# a_2437_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X37 a_n2810_45028# a_n2840_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X38 a_2113_38308# VDAC_Ni a_2112_39137# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X39 VDD a_3626_43646# a_19647_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X40 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X41 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X42 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X43 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X44 VSS a_10334_44484# a_10440_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X45 a_1576_42282# a_1755_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X46 a_10933_46660# a_10554_47026# a_10861_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X47 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X48 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X49 a_16867_43762# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X50 a_14021_43940# a_13483_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X51 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X52 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X53 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X54 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X56 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X57 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X58 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X59 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X61 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X62 a_n2840_43370# a_n2661_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X63 a_3457_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X64 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 VSS a_9672_43914# a_2107_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X66 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X67 a_14180_46482# a_14035_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X68 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X69 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X70 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X71 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 VSS a_18989_43940# a_19006_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X73 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X74 a_20749_43396# a_12549_44172# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X75 a_n2104_42282# a_n1925_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X76 VSS a_10695_43548# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X77 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X78 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X79 VDD a_3877_44458# a_2382_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X80 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X81 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X82 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X83 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X84 a_n1699_44726# a_n1917_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X85 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X86 VDD a_12883_44458# a_n2293_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X87 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X88 a_9241_45822# a_5066_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X89 a_11909_44484# a_3232_43370# a_11827_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X90 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X91 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X92 a_835_46155# a_584_46384# a_376_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X93 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X94 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X95 a_5210_46155# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X96 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X97 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X98 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X99 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X100 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X101 VDD a_167_45260# a_1609_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X102 VSS a_526_44458# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X103 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X104 a_19268_43646# a_19319_43548# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X105 VSS a_22959_44484# a_19237_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X107 a_n2216_39072# a_n2312_39304# a_n2302_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X108 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X109 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X110 a_19987_42826# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X111 a_6151_47436# a_14311_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X112 a_8145_46902# a_7927_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X113 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X114 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X115 a_14275_46494# a_13925_46122# a_14180_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X116 a_20512_43084# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X117 a_14539_43914# a_17701_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X118 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X119 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X121 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X122 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X123 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X124 a_644_44056# a_626_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X125 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X126 a_10949_43914# a_12429_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X127 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X128 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X130 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X131 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X132 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X133 VDD a_3699_46634# a_3686_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X134 VSS a_21811_47423# a_20916_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X135 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X136 a_5691_45260# a_5111_44636# a_5837_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X137 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X138 a_18249_42858# a_18083_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X139 a_8035_47026# a_7411_46660# a_7927_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X140 VDD a_1307_43914# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X141 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X142 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X143 VDD a_104_43370# a_n971_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X144 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X145 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X146 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X147 VSS a_n3565_39590# a_n3607_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X148 a_n1331_43914# a_n1549_44318# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X149 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X150 a_3363_44484# a_1823_45246# a_3232_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X152 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X153 VSS a_12281_43396# a_12563_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X154 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X155 VSS a_22400_42852# a_22780_40081# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X156 VSS a_18780_47178# a_13661_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X158 a_n4318_39768# a_n2840_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X160 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X161 a_15004_44636# a_11691_44458# a_15146_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X162 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X163 VDD a_8049_45260# a_22959_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X164 a_7230_45938# a_6472_45840# a_6667_45809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X165 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X166 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X167 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X168 a_8746_45002# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X169 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X171 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X172 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X173 a_17124_42282# a_17303_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X174 a_16223_45938# a_15599_45572# a_16115_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X175 a_n809_44244# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X176 VSS a_3065_45002# a_2680_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X178 a_5193_42852# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X179 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X180 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X181 VDD a_6969_46634# a_6999_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X182 VDD a_10623_46897# a_10554_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X183 a_16137_43396# a_15781_43660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X184 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X185 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X187 VDD a_n2472_46634# a_n2442_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X188 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X190 VDD a_4185_45028# a_22959_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X191 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X192 a_15225_45822# a_15037_45618# a_15143_45578# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X193 VSS a_3537_45260# a_4640_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X194 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X195 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X196 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X197 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X199 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X200 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X201 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X202 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X203 a_n2012_43396# a_n2129_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X204 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X205 VDD a_n13_43084# a_n1853_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X206 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X207 a_5068_46348# a_n1151_42308# a_5210_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X208 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X209 a_873_42968# a_685_42968# a_791_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X211 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X212 VDD a_22485_44484# a_20974_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 a_17730_32519# a_22591_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X214 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X215 a_n1021_46688# a_n1151_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X217 VSS a_11599_46634# a_11735_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X218 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X219 a_13163_45724# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X220 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X221 a_n2012_44484# a_n2129_44697# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X222 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X223 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X225 a_8487_44056# a_4223_44672# a_8415_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X226 a_13940_44484# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X227 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X228 VSS a_1414_42308# a_1525_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X230 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X231 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X233 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X234 a_16434_46660# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X235 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X236 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X237 a_3315_47570# a_n1151_42308# a_2952_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X238 a_2680_45002# a_1823_45246# a_2903_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X239 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X240 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X241 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X242 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X243 a_22731_47423# SMPL_ON_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X244 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X245 VDD a_1307_43914# a_3681_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X246 a_n863_45724# a_1667_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X247 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X248 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X249 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X250 a_22521_40599# COMP_P VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X252 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X253 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X254 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X255 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X256 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X257 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X258 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X259 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=218.18214 ps=2.11206k w=0.55 l=0.59
X260 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X261 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X262 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X265 a_10467_46802# a_11599_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X266 VDD a_13747_46662# a_19862_44208# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X267 a_n2946_39866# a_n2956_39768# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X269 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X270 VSS a_15279_43071# a_14579_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X271 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X272 a_7584_44260# a_7542_44172# a_7281_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X273 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X274 VSS a_8049_45260# a_22959_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X276 a_n97_42460# a_19700_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X277 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X278 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X280 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X281 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X282 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X283 VDD a_19647_42308# a_13258_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X284 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X285 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X286 a_3754_39466# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X287 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X288 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X289 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X290 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X291 VDD a_16751_45260# a_6171_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X292 VSS a_2952_47436# a_2747_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X293 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X294 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X295 a_18326_43940# a_18079_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X296 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X297 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X298 VDAC_N C0_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X299 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X300 a_9248_44260# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X301 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X302 a_3503_45724# a_3775_45552# a_3733_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X303 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X304 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X305 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X307 a_n2017_45002# a_19987_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X309 a_288_46660# a_171_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X310 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X311 VDD a_196_42282# a_n3674_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X312 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X313 a_10037_46155# a_9804_47204# a_9823_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X314 a_20075_46420# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X315 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X316 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X317 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X318 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X319 a_1149_42558# a_961_42354# a_1067_42314# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X321 VSS a_14513_46634# a_14447_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X322 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X323 a_13569_47204# a_13381_47204# a_13487_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X324 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X325 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X326 VDD a_14840_46494# a_15015_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X328 C6_P_btm a_n3565_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X329 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X330 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X331 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X332 a_14537_43396# a_14358_43442# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X333 VDD a_14955_47212# a_10227_46804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X334 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X335 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X336 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X337 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X338 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X339 a_n901_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X340 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X341 a_17668_45572# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X342 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X343 a_7309_43172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X344 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X345 a_15493_43396# a_14955_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X346 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X347 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X348 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X349 VDD a_1138_42852# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X350 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X351 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X352 a_1427_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X353 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X354 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X355 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X356 a_18184_42460# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X357 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X358 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X359 VDD a_13351_46090# a_10903_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X360 VDD a_9290_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X361 a_8379_46155# a_8128_46384# a_7920_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X362 VSS a_3483_46348# a_17325_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X363 a_18310_42308# a_10193_42453# a_18220_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X364 VSS a_11823_42460# a_14358_43442# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X365 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X367 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X368 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X369 VDD a_n2288_47178# a_n2312_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X372 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X373 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X374 a_17719_45144# a_16375_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X376 VDD a_5891_43370# a_5147_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X377 a_22609_38406# a_22469_39537# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X378 a_7287_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X379 a_11173_44260# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X381 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X382 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X383 a_11897_42308# a_11823_42460# a_11551_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X384 a_19466_46812# a_19778_44110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X385 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X386 a_9049_44484# a_8701_44490# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X387 VDD a_12861_44030# a_13759_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X388 VDD a_16588_47582# a_16763_47508# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X389 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X390 a_9396_43370# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X391 C0_P_btm a_n784_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X392 a_n1736_42282# a_n1557_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X393 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X394 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X397 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X398 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X399 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X400 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X401 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X402 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X403 VDD a_14113_42308# a_16522_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X404 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X405 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X406 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X407 a_10651_43940# a_3090_45724# a_10555_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X408 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X409 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X410 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X411 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X412 VDD a_8667_46634# a_n237_47217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X413 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X415 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X416 a_6123_31319# a_7227_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X417 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X418 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X419 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X420 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X421 VSS a_n755_45592# a_1145_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X422 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X423 C7_P_btm a_5534_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X424 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X425 VSS a_n4064_37984# a_n2302_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X426 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X427 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X428 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 a_n3674_38680# a_n2840_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X431 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X432 a_3581_42558# a_3539_42460# a_3497_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X434 VSS a_5907_45546# a_5937_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 a_18783_43370# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X436 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X437 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X438 VSS a_1799_45572# a_1983_46706# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X439 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X440 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X441 VDD a_22959_46660# a_21076_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X442 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X443 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X444 VDD a_1736_39043# a_1239_39043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X445 a_13467_32519# a_21487_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X446 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X447 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X448 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X449 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X450 a_2864_46660# a_2747_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X451 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X452 a_8199_44636# a_10355_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X453 a_14403_45348# a_13259_45724# a_14309_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X454 a_556_44484# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X455 VSS a_15433_44458# a_15367_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X456 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X457 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X458 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X459 a_n1630_35242# a_564_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X460 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X461 a_n2840_43370# a_n2661_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X462 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X463 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X464 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X465 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X466 VSS a_13747_46662# a_13693_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X467 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X468 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X469 a_18245_44484# a_17767_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X470 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X471 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X472 a_13113_42826# a_12895_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X473 a_16855_43396# a_16409_43396# a_16759_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X474 a_19741_43940# a_19862_44208# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_n1079_45724# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X476 VSS a_22365_46825# a_20202_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X477 a_19386_47436# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X478 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X479 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X480 a_1176_45822# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X481 a_13887_32519# a_22223_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X482 a_n89_47570# a_n237_47217# a_n452_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X483 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X484 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=10.615 ps=76.96 w=3.75 l=15
X485 a_10341_43396# a_9803_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X486 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X487 a_5111_42852# a_4905_42826# a_5193_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X488 VDD a_n4209_38502# a_n4334_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X489 a_5437_45600# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X490 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X491 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X492 a_18953_45572# a_18909_45814# a_18787_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X493 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X494 a_n3607_39616# a_n3674_39768# a_n3690_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X495 VDD a_3429_45260# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X496 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X497 VDD a_4791_45118# a_6165_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X498 a_4842_47570# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X499 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X500 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X501 a_1337_46116# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X502 a_n2661_42834# a_10809_44734# a_12189_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X503 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X504 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X505 a_11136_45572# a_11322_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X506 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X507 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X508 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X510 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X511 VREF_GND a_n3420_39072# C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X512 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X513 VSS a_10249_46116# a_11186_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X514 a_16655_46660# a_n743_46660# a_16292_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X515 a_n1991_46122# a_n2157_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X516 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X517 VDD a_1576_42282# a_1606_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X518 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X519 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X520 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X521 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X522 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X523 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X524 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X525 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X526 a_5159_47243# a_n443_46116# a_4700_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X527 VSS a_5891_43370# a_8375_44464# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X528 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X529 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X530 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X531 VSS a_14539_43914# a_14485_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X533 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X534 VDD a_13076_44458# a_12883_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X535 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X536 VDD en_comp a_1177_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X538 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X539 C0_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X540 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X541 a_15297_45822# a_11823_42460# a_15225_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X542 a_8103_44636# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X543 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X544 a_1423_45028# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X545 a_n1899_43946# a_n2065_43946# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X546 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X547 a_18479_47436# a_20075_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X548 a_2382_45260# a_3877_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X549 a_6765_43638# a_6547_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X550 a_n2293_43922# a_12741_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X551 a_945_42968# a_n1059_45260# a_873_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X552 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X553 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X554 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X555 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X556 VDD a_3785_47178# a_3815_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 VDD a_14084_46812# a_14035_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X558 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X559 a_765_45546# a_12549_44172# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X560 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X561 VDD a_20974_43370# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X562 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X563 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X564 a_14275_46494# a_13759_46122# a_14180_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X565 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X566 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X567 a_17517_44484# a_16979_44734# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X568 a_1609_45822# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X569 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X570 VDD a_4915_47217# a_12891_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X572 a_20679_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X574 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X576 a_13921_42308# a_13259_45724# a_13575_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X577 VSS a_1423_45028# a_9838_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X578 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X579 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X580 VCM a_n784_42308# C0_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X581 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X582 VSS a_11599_46634# a_13759_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X583 a_14127_45572# a_11823_42460# a_14033_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X584 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X585 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X586 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X587 a_13569_43230# a_12379_42858# a_13460_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X588 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X589 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X590 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X591 a_5072_46660# a_4955_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X593 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X594 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X595 a_8037_42858# a_7871_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X596 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X597 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X598 VSS a_22591_46660# a_20820_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X599 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X600 a_3686_47026# a_2609_46660# a_3524_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X601 a_9672_43914# a_10057_43914# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X602 VDD a_18429_43548# a_16823_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X603 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X604 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X605 a_17339_46660# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X606 VSS a_1606_42308# a_2351_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X607 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X608 a_16409_43396# a_16243_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X609 VDD a_n4209_37414# a_n4334_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X610 VSS a_9625_46129# a_10044_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X611 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X612 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X613 a_13468_44734# a_768_44030# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X615 a_2124_47436# a_584_46384# a_2266_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X616 VDD a_n971_45724# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X617 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X618 a_10809_44734# a_2063_45854# a_10809_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X619 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X620 a_7577_46660# a_7411_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X621 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X622 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X623 a_4921_42308# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X625 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X627 a_16023_47582# a_15507_47210# a_15928_47570# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X628 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X629 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X630 a_10193_42453# a_20712_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X631 a_12791_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X632 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X633 a_6481_42558# a_n913_45002# a_1755_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X634 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X635 VSS a_n881_46662# a_n659_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X636 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X637 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X638 a_14955_43940# a_14537_43396# a_15037_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X639 VSS C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X640 a_n2956_38680# a_n2472_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X641 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X642 VREF_GND a_14097_32519# C4_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X643 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X644 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X645 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X646 VDD a_21188_45572# a_21363_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X647 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X648 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X649 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X651 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X652 a_18907_42674# a_18727_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X653 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X654 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X655 a_12545_42858# a_12379_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X656 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X657 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X658 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X659 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X660 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X662 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X663 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X664 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X666 a_15125_43396# a_15095_43370# a_15037_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X667 VREF a_20692_30879# C6_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X668 a_13720_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X669 a_20974_43370# a_22485_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X670 a_18548_42308# a_18494_42460# a_18057_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X671 a_2998_44172# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X673 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X674 a_n875_44318# a_n2065_43946# a_n984_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X675 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X676 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X677 a_n2293_42834# a_8049_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X678 VSS a_4743_44484# a_4791_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X680 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X681 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X682 a_3626_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X684 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X686 VSS a_n2438_43548# a_n2433_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X687 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X688 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X689 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X690 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X691 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X692 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X693 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X694 VDD a_17973_43940# a_18079_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X695 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X696 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X697 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X698 VREF_GND a_17538_32519# C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X699 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X700 VDD a_22223_46124# a_20205_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X701 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X702 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X703 a_4704_46090# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X704 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X705 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X706 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X707 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X708 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X709 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X710 a_17478_45572# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X711 a_5815_47464# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X712 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X713 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X714 a_22609_38406# a_22521_39511# CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X715 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X716 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X717 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X718 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X719 VSS a_19864_35138# a_21589_35634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 VSS a_n3420_39616# a_n2946_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VDAC_P C0_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X722 a_17034_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X723 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X724 a_133_42852# a_n97_42460# a_n13_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X725 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X726 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X727 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X728 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X729 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X731 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X732 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X733 a_n1925_46634# a_8162_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X734 a_21350_47026# a_20273_46660# a_21188_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X735 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X736 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X737 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X738 VDD a_2713_42308# a_2903_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X740 a_n3674_39304# a_n2840_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X741 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X742 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X744 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_13565_43940# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X746 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X747 VDD a_1823_45246# a_2202_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X748 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X749 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X750 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X751 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X752 a_2211_45572# a_2063_45854# a_1848_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X753 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X754 VSS a_16112_44458# a_14673_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X755 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X756 VSS a_3316_45546# a_3260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X757 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X758 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X759 VDD a_n443_46116# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X761 a_21177_47436# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X762 VSS a_9290_44172# a_13943_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X763 a_n3674_37592# a_196_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X764 a_n310_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X766 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X767 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X768 a_421_43172# a_n97_42460# a_n13_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X769 a_18780_47178# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X770 VSS a_8791_42308# a_5934_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X771 VDD a_17339_46660# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X772 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 VSS a_n2840_46090# a_n2956_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X774 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X775 a_n2661_43370# a_10907_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X776 a_9396_43370# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X777 VDD a_19333_46634# a_19123_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X778 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X779 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X780 a_5755_42852# a_n97_42460# a_5837_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X781 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X782 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X783 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X784 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X785 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X786 a_n4251_39392# a_n4318_39304# a_n4334_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X787 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X788 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X789 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X790 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X791 a_805_46414# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X792 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X793 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X794 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X795 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X796 VDD a_n1076_43230# a_n901_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X798 VDD a_4520_42826# a_4093_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X799 a_21845_43940# a_12549_44172# a_19692_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X800 a_15415_45028# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X801 a_12469_46902# a_12251_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X802 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X803 a_19479_31679# a_22223_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X804 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X805 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X806 VSS a_22165_42308# a_22223_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X807 a_7542_44172# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X809 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X810 a_3080_42308# a_2903_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X811 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X812 VDD a_10249_46116# a_11186_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X813 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X814 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X815 a_3905_42558# a_2382_45260# a_3823_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X816 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X817 a_12347_46660# a_11901_46660# a_12251_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X818 VSS a_16137_43396# a_16414_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X819 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X820 a_5066_45546# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X821 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X822 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X823 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X824 VSS C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X825 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X826 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X827 a_14581_44484# a_13249_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X828 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X829 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X831 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X832 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X833 a_2113_38308# a_1343_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X834 a_n473_42460# a_n755_45592# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X835 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X836 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X837 VDD a_n1699_43638# a_n1809_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X839 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X840 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X841 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X842 a_13759_47204# a_13717_47436# a_13675_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X844 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X845 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X846 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X847 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X848 C4_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X849 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X850 a_2779_44458# a_1423_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X851 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X852 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X853 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X854 VDD a_19319_43548# a_19268_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X855 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X856 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X857 a_1123_46634# a_948_46660# a_1302_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X858 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X859 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X860 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X861 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X862 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X864 a_5807_45002# a_16763_47508# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X865 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X866 a_6293_42852# a_5755_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X867 a_2952_47436# a_3160_47472# a_3094_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X868 a_8120_45572# a_8034_45724# a_n1925_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X869 a_11541_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X870 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X871 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X873 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X874 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X875 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X876 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X877 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X878 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X879 a_4880_45572# a_5066_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X880 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X881 VIN_P EN_VIN_BSTR_P C0_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X882 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X883 a_5257_43370# a_5907_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X884 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X885 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X886 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X887 a_3497_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X888 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X889 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X890 a_16223_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X891 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X892 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X893 a_2711_45572# a_768_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X894 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X895 a_4883_46098# a_21363_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X896 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X897 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X898 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X899 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X900 VSS a_2553_47502# a_2487_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X901 VDD a_12469_46902# a_12359_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X902 a_6453_43914# a_6109_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X903 a_7765_42852# a_7227_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X904 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X905 a_18450_45144# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X907 a_17786_45822# a_15861_45028# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X908 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X909 a_6765_43638# a_6547_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X910 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X911 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X912 a_12089_42308# a_11551_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X913 a_16547_43609# a_16414_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X914 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X916 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X917 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X918 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X919 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X920 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X921 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X922 a_3221_46660# a_3177_46902# a_3055_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X923 a_6667_45809# a_6472_45840# a_6977_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X924 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X926 a_6643_43396# a_6197_43396# a_6547_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X927 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X928 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X929 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X930 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X932 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X933 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X934 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X935 a_5837_45348# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X936 a_5565_43396# a_4905_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X937 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X938 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X939 a_7418_45067# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X940 a_1793_42852# a_742_44458# a_1709_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X942 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X943 VDD a_10227_46804# a_10083_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X944 a_11301_43218# a_10922_42852# a_11229_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X945 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X946 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X947 VSS C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X948 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X949 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X950 VSS a_13291_42460# a_13249_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X951 a_18341_45572# a_18175_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X952 a_19113_45348# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X953 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X954 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X955 a_8696_44636# a_16855_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X956 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X957 a_12189_44484# a_8975_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X958 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X959 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X961 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X962 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X963 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X964 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X965 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X966 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X967 a_n1736_46482# a_n1853_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X968 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X969 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X970 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X971 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X972 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X973 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X974 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X975 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X976 a_1239_47204# a_1209_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X977 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X978 a_1606_42308# a_1576_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X979 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X980 VDD VDAC_Ni a_6886_37412# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X981 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X982 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X983 VDD a_n443_42852# a_6481_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X985 a_16795_42852# a_n97_42460# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X986 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X987 a_18315_45260# a_18587_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X988 VSS a_768_44030# a_3600_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X989 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X990 VDD a_12005_46116# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X991 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X993 VDD a_4958_30871# a_17531_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X995 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X996 a_17973_43940# a_17737_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X997 a_18900_46660# a_18834_46812# a_18285_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X998 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X999 VSS a_22821_38993# a_22876_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1000 a_6419_46155# a_5257_43370# a_6347_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1001 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1002 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1003 a_18597_46090# a_19431_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1004 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1005 a_3737_43940# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1006 VDD a_1823_45246# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1007 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1009 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1010 EN_VIN_BSTR_P VDD a_n1386_35608# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X1011 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1012 VSS a_21496_47436# a_13507_46334# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1013 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1014 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1015 VSS a_10723_42308# a_5742_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1017 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1018 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1019 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1020 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1021 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1022 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1023 VSS a_n4209_38216# a_n4251_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1024 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1025 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1026 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1027 a_12891_46348# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1028 VSS a_20679_44626# a_20640_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1029 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1030 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1031 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1032 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1033 a_21115_43940# a_20935_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1034 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1035 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1036 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1037 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1038 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1040 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1041 VDD a_10951_45334# a_10775_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1042 a_20850_46155# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1043 VDD a_13661_43548# a_18587_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1044 a_11649_44734# a_3232_43370# a_n2661_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X1045 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1046 a_17364_32525# a_22959_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1047 a_20820_30879# a_22591_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1048 VSS a_21359_45002# a_21101_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1049 EN_VIN_BSTR_P VDD a_n83_35174# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1050 a_18989_43940# a_18451_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1051 a_6197_43396# a_6031_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1052 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1053 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1054 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1055 VDD a_12891_46348# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1056 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1057 VREF_GND a_13467_32519# C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1058 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1059 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1060 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1061 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1062 a_8873_43396# a_5891_43370# a_8791_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 VDD a_584_46384# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X1064 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1065 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1066 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1067 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1068 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1069 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1070 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1071 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1072 C6_N_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1073 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1074 a_10809_44484# a_10057_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1075 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1076 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1077 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1078 a_n4318_38216# a_n2472_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1079 VSS C0_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1080 a_6545_47178# a_6419_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X1081 a_6109_44484# a_5518_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1082 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1083 a_13258_32519# a_19647_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1084 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1085 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1086 VDD a_11599_46634# a_18819_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1087 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1088 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1089 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1090 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1091 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1092 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1094 a_n1435_47204# a_n1605_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1095 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1096 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1097 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1098 a_14113_42308# a_13575_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1099 VSS a_4646_46812# a_4651_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1100 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1101 VSS a_n2472_46090# a_n2956_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1103 a_4958_30871# a_17124_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1104 VSS a_22223_42860# a_22400_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 a_13381_47204# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1106 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1107 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1108 C0_P_btm a_n3565_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1109 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1110 VDD a_1208_46090# a_472_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1111 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 VSS a_18479_47436# a_19452_47524# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1114 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1115 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1116 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1117 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1118 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1119 a_22545_38993# a_22459_39145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X1121 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1122 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1123 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1124 a_20623_45572# a_20107_45572# a_20528_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1125 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1126 VSS a_n3565_39304# a_n3607_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1127 a_12281_43396# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1128 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1129 a_15486_42560# a_15764_42576# a_15720_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1130 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1131 C1_P_btm a_n4209_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1132 VSS a_n1613_43370# a_8649_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1133 a_15765_45572# a_15599_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1134 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1135 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1136 VCM a_5932_42308# C3_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1137 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1138 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1139 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1140 VSS a_14495_45572# a_n881_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1141 a_10617_44484# a_10440_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1142 VDD a_5111_44636# a_8487_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1143 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1144 VSS a_1847_42826# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1145 a_n2267_44484# a_n2433_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1146 a_20708_46348# a_15227_44166# a_20850_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1147 a_1115_44172# a_453_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1148 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1149 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1150 VSS COMP_P a_n1329_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1151 VSS a_15861_45028# a_17023_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1152 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1153 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1155 a_16292_46812# a_5807_45002# a_16434_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1156 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X1157 a_17325_44484# a_15227_44166# a_16979_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 a_5534_30871# a_12563_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1159 a_15803_42450# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1160 VSS a_3381_47502# a_3315_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1162 VDD a_9863_46634# a_2063_45854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1163 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1164 VIN_N EN_VIN_BSTR_N C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1165 VSS a_584_46384# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1166 a_3863_42891# a_3681_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1167 VDD a_n2840_43370# a_n4318_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1168 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1169 VDD a_9049_44484# a_9313_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X1170 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1171 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1172 a_11541_44484# a_11453_44696# a_n2661_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1173 VDD a_376_46348# a_171_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1174 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1175 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1176 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1177 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1178 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1179 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1181 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1182 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1184 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1185 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1186 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1188 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1189 a_21589_35634# a_19864_35138# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1191 a_19553_46090# a_19335_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1192 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1193 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1194 a_18727_42674# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1195 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1196 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1197 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1198 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1199 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1200 a_n1925_42282# a_4185_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1201 VDD a_19164_43230# a_19339_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1202 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1204 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1205 VSS a_4361_42308# a_21855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1206 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1207 a_2479_44172# a_2905_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X1208 VDD a_8103_44636# a_7640_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1209 a_n1741_47186# a_12891_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1211 a_8192_45572# a_8162_45546# a_8120_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1212 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1213 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1214 a_5009_45028# a_3090_45724# a_4927_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1215 a_12549_44172# a_20567_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1216 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1217 VSS a_n2840_42282# a_n3674_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1218 a_5129_47502# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1219 a_14840_46494# a_13759_46122# a_14493_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1220 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1221 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1222 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1223 VSS a_n913_45002# a_2713_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1225 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1226 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1227 VDD a_n863_45724# a_1221_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1228 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1229 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1230 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1231 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1232 a_2307_45899# a_n237_47217# a_1848_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1233 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1234 VDD a_n4209_39304# a_n4334_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1235 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1236 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1237 a_8601_46660# a_7411_46660# a_8492_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1238 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1239 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1240 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1243 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1244 a_n2946_39072# a_n2956_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1246 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1247 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1248 a_15861_45028# a_15595_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1249 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1250 VSS a_n1613_43370# a_3221_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1251 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1252 a_1756_43548# a_768_44030# a_1987_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1253 a_3754_39134# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1254 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1255 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1256 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1257 a_n4318_40392# a_n2840_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1258 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1259 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1260 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1261 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1263 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1266 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1267 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1269 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1270 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1271 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1272 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1273 a_19332_42282# a_19511_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1274 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1275 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1276 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1277 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1278 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1279 VSS a_17583_46090# a_13259_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1280 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1281 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1282 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1283 a_20623_43914# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1284 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1285 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1286 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 a_n2661_46634# a_13017_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1288 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1289 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1290 a_4185_45348# a_3065_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1291 VDD a_19321_45002# a_20567_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1292 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1293 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1294 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1295 VDD a_6545_47178# a_6575_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1296 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1297 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1298 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1299 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1300 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1301 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1302 VDD a_18285_46348# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X1303 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1304 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1307 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1308 a_2864_46660# a_2747_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1309 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1310 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1311 VDD a_1307_43914# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1312 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1313 a_18374_44850# a_18248_44752# a_17970_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1314 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1315 a_13351_46090# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X1316 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1317 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1318 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1319 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1320 a_13657_42308# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1321 a_3090_45724# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1322 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1323 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1324 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1325 a_375_42282# a_413_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1326 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1327 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1328 VSS a_10903_43370# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1329 a_10334_44484# a_10157_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1330 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X1331 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1332 VSS a_22959_46124# a_20692_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1333 a_n3674_39768# a_n2472_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1334 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1335 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1336 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1337 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1338 VREF a_n4209_39304# C7_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1339 VSS a_20107_42308# a_7174_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1340 VSS a_n2438_43548# a_n133_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1342 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1344 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1345 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1346 VDAC_N C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1347 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1348 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1349 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1350 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1351 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1352 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1353 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1354 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1355 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1356 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1357 a_20301_43646# a_19692_46634# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1358 VDD a_n901_46420# a_n914_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1359 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1360 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1361 a_n971_45724# a_104_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1362 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1363 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1364 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1365 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1366 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1367 a_20447_31679# a_22959_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1368 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1369 a_n4334_38304# a_n4318_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1370 VSS a_13348_45260# a_13159_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1371 a_8685_42308# a_8515_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1372 VSS a_n881_46662# a_6517_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1373 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X1374 VDD a_14493_46090# a_14383_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1375 VSS a_6491_46660# a_6851_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1376 a_n327_42308# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X1377 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1378 a_22485_44484# a_22315_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1379 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1380 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1381 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1382 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1383 a_8605_42826# a_8387_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1384 a_15673_47210# a_15507_47210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1385 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1386 a_1709_42852# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1387 VDD a_n1736_42282# a_n4318_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1388 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1389 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1390 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1391 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1393 VREF a_19721_31679# C2_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1394 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1397 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1398 VSS a_895_43940# a_2537_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1399 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1400 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1401 a_13249_42308# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1402 a_8945_43396# a_3537_45260# a_8873_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1403 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1404 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1405 a_17609_46634# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1406 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1407 VDD a_11599_46634# a_18175_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1408 a_601_46902# a_383_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1409 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1410 a_4640_45348# a_4574_45260# a_4558_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1411 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1412 a_n467_45028# a_n745_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1413 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1415 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1417 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1418 a_1208_46090# a_765_45546# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1419 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1420 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1421 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1423 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1424 VSS a_n863_45724# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1425 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1426 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1427 a_3820_44260# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X1428 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1429 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1431 C5_P_btm a_n4064_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1432 VSS a_16721_46634# a_16655_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1433 a_21588_30879# a_22223_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1434 a_16877_42852# a_16823_43084# a_16795_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1435 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1436 VSS a_17715_44484# a_17737_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1437 a_16241_47178# a_16023_47582# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1438 a_17665_42852# a_17595_43084# a_14539_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1439 VSS a_n2438_43548# a_n2157_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1440 a_16759_43396# a_16409_43396# a_16664_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1441 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1442 a_22876_39857# a_22545_38993# a_22780_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1443 a_12359_47026# a_11735_46660# a_12251_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1444 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1445 a_5883_43914# a_8333_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1446 VDD a_n3565_39590# a_n3690_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1447 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1448 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1449 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1450 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1451 a_1990_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1452 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1453 a_5072_46660# a_4955_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1454 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1455 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1456 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1457 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1458 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1459 VDD a_3357_43084# a_22591_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1460 VSS a_3815_47204# a_4007_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1462 a_1736_39587# a_1736_39043# a_2112_39137# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1463 a_15803_42450# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1464 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1465 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1466 a_20528_46660# a_20411_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1467 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1468 a_n3607_39392# a_n3674_39304# a_n3690_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X1469 a_21421_42336# a_16327_47482# a_21335_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1470 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1471 VDD a_n4064_39616# a_n2216_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1472 a_n1838_35608# a_n1386_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1473 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1474 a_6655_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1475 a_14371_46494# a_13925_46122# a_14275_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1476 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1477 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1478 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1479 VDD a_3503_45724# a_3218_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1480 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1481 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1482 VDD a_n2840_43914# a_n4318_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1483 a_15037_43940# a_13556_45296# a_14955_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1484 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1485 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1486 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1487 VDD a_10467_46802# a_10428_46928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1488 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1489 a_15060_45348# a_13661_43548# a_14976_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X1490 a_9895_44260# a_9290_44172# a_9801_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1491 VDD a_6171_42473# a_5379_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1492 a_5009_45028# a_5147_45002# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1493 a_13904_45546# a_10903_43370# a_14127_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1494 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1496 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1497 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1499 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1500 VDD a_8696_44636# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1501 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1502 a_19900_46494# a_18985_46122# a_19553_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1503 a_3935_42891# a_3905_42865# a_3863_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1504 VSS a_n881_46662# a_11117_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1505 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1506 C3_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1507 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1508 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1509 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1510 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1511 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1512 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1513 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1514 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1515 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1516 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1517 a_1057_46660# a_n133_46660# a_948_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1518 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1519 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1520 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1521 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1522 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1523 VSS a_2982_43646# a_21487_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1524 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1525 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1526 a_21363_45546# a_21188_45572# a_21542_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1527 a_18204_44850# a_17767_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1528 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1529 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1530 VSS a_11823_42460# a_11322_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 a_n447_43370# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1532 VSS a_n4064_38528# a_n2302_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 a_17324_43396# a_16409_43396# a_16977_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1534 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1535 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1536 a_15095_43370# a_15567_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1537 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1539 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1540 a_10150_46912# a_10428_46928# a_10384_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1541 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1542 VSS a_n2472_42282# a_n4318_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1543 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1544 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1545 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1546 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1547 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1548 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1549 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1550 a_8492_46660# a_7577_46660# a_8145_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1551 a_5649_42852# a_5111_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1552 VDD a_18287_44626# a_18248_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1553 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1554 a_20894_47436# a_20990_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1555 a_19636_46660# a_19594_46812# a_19333_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1556 a_10249_46116# a_9823_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1557 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1558 a_739_46482# a_n743_46660# a_376_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1559 VSS a_10775_45002# a_10180_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 a_2896_43646# a_2479_44172# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X1561 a_10227_46804# a_14955_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1562 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1563 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1564 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1565 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1566 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1567 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1568 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1569 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1570 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1571 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1572 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1575 a_12791_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1576 VSS a_5807_45002# a_11691_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1577 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1578 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1579 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1580 VSS a_2382_45260# a_2304_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1581 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1582 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1583 VSS a_3357_43084# a_22591_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1584 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1585 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1586 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1587 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1588 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1589 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1590 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1592 VDD a_2277_45546# a_2307_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1593 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1594 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1595 a_10053_45546# a_8746_45002# a_10306_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1596 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1597 a_n2956_39768# a_n2840_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1598 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1599 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1600 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1601 VDD a_4361_42308# a_21855_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1602 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1603 VSS a_6945_45028# a_22223_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1604 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1605 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1606 VDD a_5257_43370# a_5263_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1607 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1608 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1609 a_18494_42460# a_18907_42674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1610 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1611 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1612 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1613 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1615 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1616 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1617 a_n1151_42308# a_n1329_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1618 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1619 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1620 a_16763_47508# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1621 a_21259_43561# a_4190_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1622 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1623 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1625 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1626 a_8349_46414# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1627 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1628 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1629 a_17970_44736# a_18287_44626# a_18245_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1630 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1631 a_1123_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1632 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1633 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1634 a_n237_47217# a_8667_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1635 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1636 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1638 a_5837_42852# a_3537_45260# a_5755_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1639 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1640 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1641 VSS a_19692_46634# a_19636_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1642 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1643 a_8697_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1644 a_1145_45348# a_n863_45724# a_626_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1645 VSS a_5934_30871# a_8515_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1646 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1647 VSS a_1239_47204# a_1431_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1648 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1649 a_22705_38406# a_22521_40055# a_22609_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1650 a_11173_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X1651 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1652 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1653 a_22165_42308# a_21887_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1654 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1655 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1656 VDD a_8952_43230# a_9127_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1657 VSS a_n4064_37440# a_n2302_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1658 a_5244_44056# a_5147_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1659 VSS a_2127_44172# a_n2661_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1661 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1662 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1663 a_n2956_37592# a_n2472_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1664 VSS a_15493_43940# a_22959_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1665 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1666 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1667 a_19339_43156# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1668 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1669 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1670 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1671 VDD a_n1177_44458# a_n1190_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1672 VDD a_n1920_47178# a_n2312_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1673 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1675 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1676 VDD a_16292_46812# a_15811_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1677 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1679 a_5164_46348# a_4927_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1680 a_9482_43914# a_9838_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1681 a_20835_44721# a_20679_44626# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1682 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1683 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1684 a_5837_42852# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1685 VSS a_5937_45572# a_8781_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1686 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1687 a_7221_43396# a_6031_43396# a_7112_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1688 a_10037_47542# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1689 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1690 C7_N_btm a_20820_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1691 VSS a_5937_45572# a_8560_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1692 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1693 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1694 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1695 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1696 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1697 VSS a_15559_46634# a_13059_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1699 a_5385_46902# a_5167_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1700 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1701 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1702 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1703 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1704 VDD a_10334_44484# a_10440_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1705 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1706 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1707 a_19597_46482# a_19553_46090# a_19431_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1708 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1709 a_18051_46116# a_18189_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1710 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1711 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1712 a_16414_43172# a_n1059_45260# a_16328_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1713 a_15493_43940# a_14955_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1714 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1715 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1716 a_21297_46660# a_20107_46660# a_21188_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1717 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1718 a_11813_46116# a_11387_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X1719 VSS SMPL_ON_P a_n1605_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1720 VDD a_4699_43561# a_3539_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1721 VSS a_n3420_39072# a_n2946_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1722 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1723 a_5894_47026# a_4817_46660# a_5732_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1724 VDD a_n97_42460# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1725 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1726 VDD a_13163_45724# a_11962_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1727 a_15433_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1728 VDD a_16327_47482# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1729 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1730 a_18114_32519# a_22223_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1731 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1732 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1733 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1734 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1735 a_n452_44636# a_n1151_42308# a_n310_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1737 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1738 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1739 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1740 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1741 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1742 VDD a_22959_43396# a_17364_32525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1743 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1744 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1745 VSS a_n357_42282# a_7573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1746 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1747 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1748 VDD a_1307_43914# a_4149_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X1749 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1750 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1751 VDD a_9863_47436# a_9804_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1752 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1753 a_22821_38993# a_22400_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1754 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1755 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1756 a_3754_39134# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1757 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1758 a_4649_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1759 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1761 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1762 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1763 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1764 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1766 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1767 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1768 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1769 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1770 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1771 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1772 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1773 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1774 VSS a_1848_45724# a_1799_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1775 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1776 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1777 a_20885_45572# a_20841_45814# a_20719_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1778 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1779 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1780 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1781 a_10554_47026# a_10428_46928# a_10150_46912# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1782 a_n746_45260# a_n1177_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1783 a_7_44811# a_n1151_42308# a_n452_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1784 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1785 VDD a_10355_46116# a_8199_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1786 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1787 a_4181_43396# a_4093_43548# a_n2661_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 a_21005_45260# a_21101_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1789 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1790 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1791 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1792 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1793 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1794 VDD a_2437_43646# a_22223_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1795 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1796 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1797 a_3754_38802# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1798 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1799 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1800 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1801 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1802 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1803 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1804 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1805 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1806 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1807 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1809 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1810 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1811 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1812 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1813 VDD a_n2840_45002# a_n2810_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1814 VSS a_12861_44030# a_17339_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1815 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1816 a_10057_43914# a_10807_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1817 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1818 a_5343_44458# a_7963_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1819 a_n1423_42826# a_n1641_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1820 VDD a_11827_44484# a_22223_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1821 VDD a_n2472_43914# a_n3674_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1822 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1823 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1824 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1826 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1827 a_6945_45028# a_5937_45572# a_6945_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1828 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1829 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1830 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1831 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1832 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1833 a_20301_43646# a_13661_43548# a_743_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1835 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1836 a_n2216_39866# a_n2442_46660# a_n2302_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1837 VDD a_22000_46634# a_15227_44166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1838 a_n3674_38216# a_n2104_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1839 VSS a_2889_44172# a_413_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1840 VSS a_n97_42460# a_n144_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1841 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1842 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1843 a_133_42852# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1844 a_16321_45348# a_1307_43914# a_16019_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X1845 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1846 VDD a_9290_44172# a_13070_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1847 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1848 VDD a_22465_38105# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1849 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X1850 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1851 a_n2860_38778# a_n2956_38680# a_n2946_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1852 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1853 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1854 a_10555_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1855 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1856 a_6517_45366# a_5937_45572# a_6431_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1857 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1858 a_14401_32519# a_22223_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1859 VDD a_5111_44636# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1860 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1861 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1862 VSS a_9290_44172# a_13070_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1864 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1865 VDD a_9290_44172# a_10586_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1866 a_16751_45260# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1867 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1868 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1869 VSS a_5068_46348# a_4955_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1870 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1871 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1872 a_1736_39587# a_1736_39043# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X1873 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1874 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1875 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1876 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1877 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1878 VSS a_11599_46634# a_15507_47210# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1879 VSS a_768_44030# a_644_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1880 VDD a_n357_42282# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1881 a_5193_43172# a_3905_42865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1882 VSS a_18783_43370# a_18525_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1883 a_12465_44636# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1884 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1885 a_3540_43646# a_1414_42308# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X1886 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1887 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1888 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1890 a_5421_42558# a_5379_42460# a_5337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1891 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1892 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1893 a_21363_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1894 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1895 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1896 VDD a_12861_44030# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1897 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1898 a_n2956_38216# a_n2472_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1899 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1900 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1901 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1902 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1903 a_13885_46660# a_13607_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1904 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1905 a_2232_45348# a_1609_45822# a_n2293_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X1906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1907 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1908 a_5691_45260# a_6171_45002# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1909 a_9801_44260# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1910 VCM a_3080_42308# C2_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1911 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1912 a_15743_43084# a_19339_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1913 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1914 VSS a_22591_43396# a_14209_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1915 a_327_44734# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1916 VSS a_7499_43078# a_8746_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1917 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1918 VSS a_2437_43646# a_22223_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1919 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1920 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1921 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1922 a_6547_43396# a_6197_43396# a_6452_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1923 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1924 a_20556_43646# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1925 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1926 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1927 a_1987_43646# a_742_44458# a_1891_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1929 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1930 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1931 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1932 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1933 a_648_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X1934 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1935 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1936 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1937 VDD a_n23_47502# a_7_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1938 a_17609_46634# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1939 a_3602_45348# a_3537_45260# a_3495_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X1940 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1941 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1942 VDD a_2982_43646# a_21487_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1943 a_13661_43548# a_18780_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1944 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1945 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1946 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1947 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1948 a_11323_42473# a_5742_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1949 a_9313_44734# a_3232_43370# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1950 C6_P_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1951 a_14383_46116# a_13759_46122# a_14275_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1952 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1953 a_2813_43396# a_2479_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1955 a_16721_46634# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1957 VREF a_20820_30879# C7_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1958 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1959 VDD a_526_44458# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1960 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1961 VDD a_15681_43442# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1962 a_6125_45348# a_3232_43370# a_5691_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1963 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1964 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1965 a_10907_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1966 a_14955_43396# a_9145_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1967 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1968 a_3429_45260# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1969 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1970 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1971 a_8128_46384# a_7903_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1972 VDD a_15227_44166# a_17969_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X1973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1974 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1975 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1976 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1977 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1978 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1979 VSS C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1980 a_n2860_37690# a_n2956_37592# a_n2946_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1981 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1982 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1983 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1984 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1985 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1986 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1987 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1989 C4_P_btm a_n3420_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1990 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1991 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1993 a_18599_43230# a_18083_42858# a_18504_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1994 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1995 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1996 a_18057_42282# a_18494_42460# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1997 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1998 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1999 a_11117_47542# a_4915_47217# a_11031_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2000 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2001 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2002 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2003 VDD a_22400_42852# a_22521_40599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2004 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2005 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2006 a_7112_43396# a_6197_43396# a_6765_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2007 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2008 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2009 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2010 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2011 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2012 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2013 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2014 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2015 a_19240_46482# a_19123_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2016 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2017 VCM a_5742_30871# C6_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2018 VSS a_10193_42453# a_10149_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2019 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2020 VDD a_10193_42453# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2021 a_564_42282# a_743_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2022 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2023 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2024 VSS a_n967_45348# a_n961_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2025 a_21195_42852# a_20922_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2026 VDD a_6575_47204# a_9067_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2027 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2028 a_22612_30879# a_22959_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2029 a_21188_46660# a_20273_46660# a_20841_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2030 a_13749_43396# a_13661_43548# a_13667_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2031 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2032 VSS a_n2840_45546# a_n2810_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2033 a_13490_45394# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2034 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2035 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2036 a_n2840_43914# a_n2661_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2037 a_n822_43940# a_n1899_43946# a_n984_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2038 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2040 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2041 a_21613_42308# a_21335_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2042 a_14537_43396# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2043 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2044 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2045 a_7112_43396# a_6031_43396# a_6765_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2046 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2047 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2048 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2049 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2051 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2052 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2053 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2054 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2055 a_n23_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2056 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2057 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2058 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2059 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2060 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2061 a_14543_43071# a_5534_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2062 VDD a_7227_45028# a_7230_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2063 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2064 VDD a_19900_46494# a_20075_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2065 VSS a_16327_47482# a_19597_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2066 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2067 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2068 a_9823_46155# a_n743_46660# a_9751_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2069 a_18214_42558# a_16137_43396# a_18057_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2070 VDD a_22959_43948# a_17538_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2071 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2072 a_n3690_38304# a_n3674_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2073 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2074 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2075 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2076 a_15009_46634# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2077 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2078 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2079 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2080 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2081 VSS a_10227_46804# a_15521_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2082 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2083 a_17591_47464# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2084 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2085 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2086 a_22485_44484# a_22315_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2087 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2088 a_n1644_44306# a_n1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2090 VDD a_n1329_42308# a_n1151_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2091 VDD RST_Z a_8530_39574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2092 VSS a_13507_46334# a_18184_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2093 a_n630_44306# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2095 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2096 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2097 a_18783_43370# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2098 VSS C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2099 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2100 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2101 a_8325_42308# a_n913_45002# a_8337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2102 VSS a_22521_40599# a_22469_40625# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2103 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2104 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2105 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2106 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2107 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2108 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2109 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2110 a_21973_42336# a_20202_43084# a_21887_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2111 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2112 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2113 VSS a_n1613_43370# a_645_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2114 a_10341_42308# a_9803_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2115 VSS a_10807_43548# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2116 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2117 VSS a_16327_47482# a_20885_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2118 a_n1920_47178# a_n1741_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2119 a_9127_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2120 VSS a_5257_43370# a_3905_42865# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2122 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2123 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2124 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2125 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2126 VDD a_n2472_45002# a_n2956_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2127 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2128 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2129 a_13259_45724# a_17583_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2130 VSS a_10586_45546# a_10544_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2131 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2132 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2133 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2134 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2135 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2136 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2137 a_16751_45260# a_17023_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2139 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2140 VSS a_n4209_38502# a_n4251_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2141 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2142 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2143 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2144 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2145 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2146 a_n2840_42826# a_n2661_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2147 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2148 VSS a_7227_42308# a_6123_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2149 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2150 a_1302_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2151 a_5907_45546# a_6194_45824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2152 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2153 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2154 a_n2302_37984# a_n2810_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_13059_46348# a_15559_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2156 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2157 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2158 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2159 VREF_GND a_14209_32519# C5_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2161 a_3065_45002# a_3318_42354# a_3581_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2162 a_16023_47582# a_15673_47210# a_15928_47570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2163 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2164 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2165 VSS a_n881_46662# a_n935_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 VDD a_21487_43396# a_13467_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2167 C6_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2168 VDD a_n443_42852# a_997_45618# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2169 a_2553_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2170 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2171 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2172 a_13635_43156# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2173 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2174 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2175 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2176 a_8568_45546# a_8199_44636# a_8791_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2177 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2178 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2179 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2180 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2181 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2182 VDD a_564_42282# a_n1630_35242# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2183 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2184 a_n473_42460# a_n971_45724# a_n327_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X2185 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2186 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2187 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2188 a_16335_44484# a_13661_43548# a_16241_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2190 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2191 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2192 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2193 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2194 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2195 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2196 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2197 VDD a_15861_45028# a_17023_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2198 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2199 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2200 a_5205_44734# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2201 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X2202 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2203 VSS a_1123_46634# a_1057_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2204 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2205 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2206 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2207 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2208 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2209 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2210 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2211 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2212 VSS a_13259_45724# a_18315_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2213 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2214 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2215 VSS a_22223_43396# a_13887_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2217 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2218 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2219 a_11682_45822# a_11322_45546# a_11525_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2220 VDD a_22591_45572# a_19963_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2221 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2222 a_18429_43548# a_18525_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2223 a_5934_30871# a_8791_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2224 a_509_45822# a_n1099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2225 a_4190_30871# a_19332_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2226 a_20980_44850# a_20766_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2227 a_3381_47502# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2228 VDD a_3537_45260# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2229 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2230 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2231 VDD a_1423_45028# a_9838_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2233 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2234 a_6682_46660# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2235 a_20273_45572# a_20107_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2236 VDD a_11963_45334# a_11787_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2237 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2238 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2239 a_19256_45572# a_18175_45572# a_18909_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2240 VSS a_5937_45572# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2241 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2242 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2243 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2244 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2245 VSS a_3699_46634# a_3633_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2246 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2247 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2248 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2249 VSS a_n2438_43548# a_n2157_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2250 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2251 a_14226_46987# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2253 a_n722_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2254 a_n2840_45002# a_n2661_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2255 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2256 VSS a_8953_45546# a_9241_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 a_12005_46436# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2258 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2259 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2260 a_9885_43396# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2261 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2262 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2263 VSS a_n4209_37414# a_n4251_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2265 a_18817_42826# a_18599_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2266 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2267 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2268 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2269 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2270 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2271 VDD a_167_45260# a_1423_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2272 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2273 VSS a_4704_46090# a_1823_45246# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2274 a_16886_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X2275 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2276 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2277 VSS C0_dummy_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2278 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2279 a_11688_45572# a_11652_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2280 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2281 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2282 a_4520_42826# a_1823_45246# a_4743_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2283 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2284 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2285 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2286 VDD a_n2104_42282# a_n3674_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2287 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2288 VDD RST_Z a_14311_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2289 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2290 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2291 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2292 a_19339_43156# a_19164_43230# a_19518_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2293 a_19721_31679# a_22959_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2294 a_458_43396# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X2295 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2296 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2298 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2299 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2300 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2301 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2302 a_11453_44696# a_17719_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2303 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2304 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2306 a_22717_36887# a_22459_39145# a_22609_37990# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2307 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2308 VDD a_n3420_37984# a_n2860_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2309 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2310 a_13711_45394# a_12891_46348# a_13348_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2312 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2313 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2314 a_1138_42852# a_791_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2315 a_16664_43396# a_16547_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2316 a_21259_43561# a_4190_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2317 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2318 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2319 a_10586_45546# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2320 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2321 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2322 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2323 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2324 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2325 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2326 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2327 VSS a_11599_46634# a_15599_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2328 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2329 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2330 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X2331 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2332 a_196_42282# a_375_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2333 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2334 VSS a_n881_46662# a_7989_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2335 a_7832_46660# a_7715_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2336 VDD a_n2109_45247# en_comp VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2337 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2338 a_3633_46660# a_2443_46660# a_3524_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2339 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2340 a_15928_47570# a_15811_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2341 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2342 a_2127_44172# a_2675_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2343 a_9885_43646# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2344 VSS a_n2472_45546# a_n2956_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 a_n2472_43914# a_n2293_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2346 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2347 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2348 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2349 VDD a_12991_46634# a_12978_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2350 VDD a_1667_45002# a_n863_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2351 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2352 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2353 a_5837_45028# a_3232_43370# a_5691_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X2354 VDD a_21195_42852# a_21671_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2355 a_14084_46812# a_n1151_42308# a_14226_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2356 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2357 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2358 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2359 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2360 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2361 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2362 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2363 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2364 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2365 VSS a_n913_45002# a_4921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2367 a_14209_32519# a_22591_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2368 a_12427_45724# a_12791_45546# a_12749_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2369 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2370 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2372 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2373 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2374 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2375 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2376 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2377 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2378 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2379 a_12553_44484# a_12465_44636# a_n2661_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2381 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2382 a_5829_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2383 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2384 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2385 a_16237_45028# a_n743_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2386 VDD a_22959_45036# a_19721_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2388 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2389 a_14761_44260# a_14673_44172# a_n2293_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2390 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2391 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2393 VSS a_n1613_43370# a_5429_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2394 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2395 VDD a_n452_45724# a_n1853_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2396 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2397 VSS a_21363_46634# a_21297_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2398 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2399 VDD a_584_46384# a_2998_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2400 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2401 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2402 VDD a_15959_42545# a_15890_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2403 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2405 VSS a_4699_43561# a_3539_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2406 VSS a_10227_46804# a_13157_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2407 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2408 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2409 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2410 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2411 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2412 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2413 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2414 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2415 a_n144_43396# a_n971_45724# a_n447_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2416 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2417 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2418 a_17538_32519# a_22959_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2419 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2421 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2422 a_16680_45572# a_15599_45572# a_16333_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2423 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2424 VSS a_5937_45572# a_6101_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2425 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2426 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2427 a_8387_43230# a_7871_42858# a_8292_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2428 a_15231_43396# a_9145_43396# a_15125_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2429 a_9672_43914# a_8199_44636# a_9895_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2431 VDD a_22731_47423# a_13717_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2432 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2433 VDD a_9290_44172# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2434 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2435 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2436 VDD a_17767_44458# a_17715_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X2437 VDD a_7845_44172# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2438 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2439 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2440 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2441 VDD a_10903_43370# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X2442 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2443 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2444 a_n2840_44458# a_n2661_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2445 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2446 VDD a_n863_45724# a_945_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2447 a_22400_42852# a_22223_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2448 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2449 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2450 VDD a_12549_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X2451 a_4933_42558# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2452 VSS a_9482_43914# a_10157_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2453 a_19333_46634# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2454 a_13565_44260# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2455 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2456 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2457 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2458 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2459 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2460 a_n2293_46098# a_5663_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X2461 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2462 VSS a_11453_44696# a_22959_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2463 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2464 VSS a_12563_42308# a_5534_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2465 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2466 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2467 a_n2472_42826# a_n2293_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2468 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2469 a_n13_43084# a_n443_42852# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2470 a_7920_46348# a_8128_46384# a_8062_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2471 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2472 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2473 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2474 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2475 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2476 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2477 a_2698_46116# a_2521_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2478 a_15785_43172# a_15743_43084# a_15095_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2479 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2480 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2481 a_8654_47026# a_7577_46660# a_8492_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2482 VDD a_21363_46634# a_21350_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2483 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2484 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2485 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2486 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2487 VDD a_n809_44244# a_n822_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2488 a_766_43646# a_626_44172# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X2489 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2490 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2491 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2492 a_n784_42308# a_n961_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2493 a_12895_43230# a_12379_42858# a_12800_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2494 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2495 VSS a_8191_45002# a_8137_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2496 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2497 a_15959_42545# a_15803_42450# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2499 VSS a_805_46414# a_739_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2500 a_11341_43940# a_3232_43370# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X2501 a_5210_46482# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2502 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2503 VDD a_7705_45326# a_7735_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2504 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2505 a_13720_44458# a_13661_43548# a_13940_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2506 a_2162_46660# a_2107_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2507 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2508 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2509 a_n1423_42826# a_n1641_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2510 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2511 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2512 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2513 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2514 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2515 a_n2956_39304# a_n2840_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2516 VDD a_11415_45002# a_n2661_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2517 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2518 a_15037_43940# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2519 VDD a_1606_42308# a_2351_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2520 a_2277_45546# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2521 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2522 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2523 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2524 VDD a_14180_45002# a_13017_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2525 a_3232_43370# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2526 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2527 a_6903_46660# a_6755_46942# a_6540_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2528 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2529 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2530 a_22521_40055# en_comp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2532 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2533 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2534 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2535 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2536 a_1576_42282# a_1755_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2537 VDD a_8199_44636# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2538 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2539 VSS a_21855_43396# a_13678_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2540 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2541 a_7573_43172# a_7499_43078# a_7227_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2542 VDD a_18989_43940# a_19006_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2543 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2544 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2545 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2546 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2547 VSS a_6540_46812# a_6491_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2548 VDD a_22223_45572# a_19479_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2549 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2550 VIN_N EN_VIN_BSTR_N C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2551 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2552 VSS a_2903_42308# a_3080_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2553 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2554 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2555 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2556 VSS a_n863_45724# a_n906_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2557 a_3823_42558# a_3065_45002# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2558 a_n2840_44458# a_n2661_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2559 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2560 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2561 VSS a_5263_45724# a_5204_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2562 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2563 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2564 VDD a_2124_47436# a_1209_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2565 VSS a_2957_45546# a_2905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2566 a_12925_46660# a_11735_46660# a_12816_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2567 a_376_46348# a_n743_46660# a_518_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2568 a_11415_45002# a_4915_47217# a_14581_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2569 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2570 a_n2104_42282# a_n1925_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2571 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2573 a_n2472_45002# a_n2293_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2574 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2575 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2576 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2577 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2578 a_21398_44850# a_20679_44626# a_20835_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2580 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2581 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2582 VDD a_22521_40599# a_22705_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2583 VSS a_8685_43396# a_15231_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2584 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2585 VDD a_16333_45814# a_16223_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2586 a_16241_44484# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X2587 a_3905_42865# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2588 a_13485_45572# a_12549_44172# a_13385_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X2589 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2590 C3_P_btm a_n4209_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2591 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2592 VSS a_10623_46897# a_10554_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2593 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2594 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2595 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2596 VSS a_22959_45572# a_20447_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2597 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2598 a_19120_35138# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2599 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2600 VDD a_19987_42826# a_n2017_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X2601 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2602 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2603 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2604 a_9028_43914# a_9482_43914# a_9420_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2605 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2606 a_n2860_39072# a_n2956_39304# a_n2946_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2607 VSS a_17973_43940# a_18079_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2608 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2609 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2610 a_3059_42968# a_742_44458# a_2987_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2611 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2612 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2613 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2616 a_n452_44636# a_n467_45028# a_n310_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2617 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2619 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2620 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2622 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2623 VDD a_768_44030# a_2711_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2624 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2625 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2627 VDAC_N C0_dummy_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2628 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2629 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2630 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2631 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2632 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2633 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2634 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2635 VDD a_12281_43396# a_12563_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2636 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2637 VDD a_12741_44636# a_22959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2638 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2639 a_8333_44734# a_3537_45260# a_8238_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2640 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2641 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2642 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2643 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2644 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2645 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2646 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2647 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2648 a_17124_42282# a_17303_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2649 a_12156_46660# a_11813_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2650 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2651 VDD a_n447_43370# a_n2129_43609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2652 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2653 VDD a_10809_44734# a_22959_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2654 VSS a_1115_44172# a_n2293_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X2655 a_5013_44260# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2656 a_3357_43084# a_5257_43370# a_5565_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2658 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2659 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2660 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2661 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2662 a_1568_43370# a_1847_42826# a_1793_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2663 a_11682_45822# a_10586_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2664 a_n2012_44484# a_n2129_44697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2665 a_18315_45260# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X2666 a_14543_43071# a_5534_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2667 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2668 a_16147_45260# a_17478_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2670 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2671 a_19963_31679# a_22591_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2672 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2673 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2674 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2675 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2676 a_n967_45348# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2677 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2678 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2679 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2680 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2681 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2682 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2684 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2685 VSS a_7276_45260# a_7227_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2686 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2687 a_1241_44260# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X2688 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2689 VDD a_11599_46634# a_20107_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2690 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2691 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2692 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2693 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2694 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2695 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2696 a_n4334_40480# a_n4318_40392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2697 VSS a_n815_47178# a_n785_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2698 a_3175_45822# a_3090_45724# a_2957_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2699 a_14621_43646# a_14579_43548# a_14537_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2700 VDD a_n1386_35608# a_n1838_35608# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2701 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2702 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2703 VREF a_20205_31679# C4_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2704 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2705 VSS a_15227_44166# a_18900_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2706 a_n310_44811# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2707 VDD a_16977_43638# a_16867_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2708 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2709 VDD a_15227_44166# a_17749_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2710 a_3147_46376# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2711 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2712 a_12638_46436# a_12594_46348# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2713 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2714 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2715 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2716 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2717 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2718 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2719 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2720 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2721 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2722 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2723 a_21071_46482# a_15227_44166# a_20708_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2724 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2725 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2726 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2727 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2728 a_9127_43156# a_8952_43230# a_9306_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2729 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2730 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2731 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2732 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2733 VDD a_1343_38525# a_2684_37794# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2734 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2735 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2736 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2737 a_961_42354# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2738 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2739 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2740 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2741 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2742 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2743 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2744 VSS a_8349_46414# a_8283_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2745 VSS a_11787_45002# a_11652_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X2746 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2747 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2748 VSS a_12741_44636# a_22959_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2750 a_4223_44672# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2751 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2752 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2753 a_509_45822# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2754 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2755 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2756 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2757 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2758 a_16119_47582# a_15673_47210# a_16023_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2759 a_6452_43396# a_6293_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2761 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2762 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2763 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2764 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2766 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2767 a_6194_45824# a_6472_45840# a_6428_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2768 a_3754_38802# a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X2769 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2770 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2771 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2772 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2773 VDD a_n881_46662# a_11031_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2774 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2775 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2776 VSS a_1209_47178# a_1239_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2777 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2778 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2779 a_12429_44172# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2780 a_15559_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X2781 a_11229_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2782 a_16020_45572# a_15903_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2783 a_10149_42308# a_9290_44172# a_9803_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2784 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2785 C3_P_btm a_5932_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2786 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2787 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2788 a_10793_43218# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2789 VSS a_20708_46348# a_20411_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2790 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2791 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2792 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2793 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2794 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2795 a_13635_43156# a_13460_43230# a_13814_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2796 a_n863_45724# a_1667_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2797 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2798 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2799 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2800 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2801 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2802 a_12379_46436# a_12594_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2803 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2804 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2805 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2806 a_1209_43370# a_1049_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2807 a_2982_43646# a_3232_43370# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2809 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2810 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2811 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2812 a_21542_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2813 VSS a_19647_42308# a_13258_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2814 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2815 a_18985_46122# a_18819_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2816 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2817 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2818 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2819 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2821 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2822 a_12839_46116# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2823 VDD a_n2438_43548# a_2443_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2824 VDD a_9028_43914# a_8975_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2825 VDD a_17124_42282# a_4958_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2826 VSS a_10053_45546# a_9625_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X2827 VSS a_380_45546# a_n356_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2828 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2829 VSS a_20193_45348# a_21973_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2830 VSS a_196_42282# a_n3674_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2831 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2832 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2833 a_17639_46660# a_17609_46634# a_765_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2834 VDD a_5257_43370# a_5826_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2835 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2836 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2837 a_9803_42558# a_n97_42460# a_9885_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2839 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2840 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2841 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2843 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2844 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2845 VSS a_10227_46804# a_10553_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2846 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2847 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2848 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2849 VSS a_n913_45002# a_12281_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2850 VSS a_18597_46090# a_16375_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2852 a_12816_46660# a_11901_46660# a_12469_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2853 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2854 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2855 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2856 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2857 a_20205_45028# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2858 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2859 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2860 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2861 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2862 VDD a_13259_45724# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X2863 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2864 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2866 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2867 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2868 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2869 a_n1736_42282# a_n1557_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2870 a_13747_46662# a_19386_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2871 VSS a_4791_45118# a_6165_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2872 a_261_44278# a_n863_45724# a_175_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2873 a_8325_42308# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2874 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2875 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2876 a_10623_46897# a_10467_46802# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2877 a_2675_43914# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2878 a_18695_43230# a_18249_42858# a_18599_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2879 a_17957_46116# a_765_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X2880 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2881 a_17613_45144# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2882 a_n4318_39304# a_n2840_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2883 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2884 a_18799_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2885 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2886 VSS a_19862_44208# a_20922_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X2887 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2888 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2889 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2890 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2891 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2892 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2893 a_6151_47436# a_14311_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2894 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2895 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2896 VSS a_5129_47502# a_5063_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2897 VSS a_167_45260# a_2521_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2898 a_16333_45814# a_16115_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2899 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2900 a_3733_45822# a_n755_45592# a_3638_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2901 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2902 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2903 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2904 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2905 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2907 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2908 a_13163_45724# a_13527_45546# a_13485_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2909 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2910 a_8605_42826# a_8387_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2911 a_1337_46116# a_1176_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2912 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2913 a_n83_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2914 VDD a_4419_46090# a_n1925_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2915 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2916 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2917 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2918 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2919 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2920 a_20712_42282# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2921 a_1241_43940# a_1467_44172# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2922 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2923 VDD a_n961_42308# a_n784_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2924 a_7227_42852# a_n97_42460# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2925 a_9145_43396# a_8791_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2926 a_14976_45348# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2927 a_9863_47436# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2928 a_743_42282# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2929 VSS a_12891_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2930 a_4915_47217# a_12991_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2933 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2934 a_n3674_38680# a_n2840_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2935 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2936 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2937 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2938 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2939 VSS a_3539_42460# a_3065_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2940 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2941 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2942 a_17801_45144# a_17613_45144# a_17719_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X2943 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2944 VDD a_n4209_39590# a_n4334_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2945 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2946 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2947 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2948 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2949 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2950 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2951 a_18787_45572# a_18341_45572# a_18691_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2952 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2953 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2955 a_10922_42852# a_10796_42968# a_10518_42984# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2957 a_3754_39964# a_7754_40130# VSS sky130_fd_pr__res_high_po_0p35 l=18
X2958 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2959 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2961 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2962 VDD a_526_44458# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2963 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2964 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2965 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2966 a_n1630_35242# a_564_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2967 a_167_45260# a_2202_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2968 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2969 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2970 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2971 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2972 VDD a_11967_42832# a_20512_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2974 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2975 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2976 VDD a_16019_45002# a_15903_45785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2977 a_2896_43646# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2978 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2979 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2980 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2981 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2982 a_12005_46116# a_10903_43370# a_12005_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2983 a_n2312_38680# a_n2104_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2984 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2985 a_14097_32519# a_22959_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2986 a_n2288_47178# a_n2109_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2987 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2988 a_6999_46987# a_3877_44458# a_6540_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2989 a_8199_44636# a_10355_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2990 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2991 a_3429_45260# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2992 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2993 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2995 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2996 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2997 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2998 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2999 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3000 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3001 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3002 C8_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3003 a_9293_42558# a_9223_42460# a_8953_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X3004 a_4338_37500# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X3005 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3006 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3007 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3009 VDD a_n452_47436# a_n815_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3010 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3011 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3012 a_13807_45067# a_13556_45296# a_13348_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3013 a_14309_45348# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3014 a_1176_45822# a_997_45618# a_1260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X3015 VDD a_13159_45002# a_n2661_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3016 VSS a_20269_44172# a_19319_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3017 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3018 a_16104_42674# a_15890_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3019 a_2981_46116# a_2804_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3020 a_4185_45028# a_3877_44458# a_4185_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3021 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3023 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3024 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3025 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3026 a_22731_47423# SMPL_ON_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3027 a_n722_46482# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3028 VSS a_n443_42852# a_997_45618# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X3029 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3030 a_6945_45348# a_5205_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3031 a_4791_45118# a_4743_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3032 a_21513_45002# a_21363_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3034 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3035 VSS a_1576_42282# a_1606_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3036 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3037 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3038 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3039 a_15227_44166# a_22000_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3040 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3041 VDAC_P C0_dummy_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3042 VSS en_comp a_1177_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3043 a_n743_46660# a_n1021_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3044 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3045 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3046 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3047 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3048 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3049 VSS a_5205_44484# a_6756_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3051 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3052 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3053 VDD a_19321_45002# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X3054 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3055 VSS a_3483_46348# a_13829_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3056 VDD a_327_44734# a_375_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3057 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3058 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3059 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3060 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3061 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3062 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3063 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3064 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3065 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3066 VDD a_5937_45572# a_6671_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3067 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3068 VDD a_n863_45724# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X3069 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3070 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3071 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3072 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3073 VDD a_1756_43548# a_1467_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X3074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3075 a_20269_44172# a_20365_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X3076 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3077 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3078 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3079 VDD a_4791_45118# a_5066_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3080 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3081 VDD a_14976_45028# a_15227_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3082 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3083 VSS a_13904_45546# a_12594_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3084 VSS a_8953_45546# a_8568_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3085 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3087 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3088 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3089 a_16112_44458# a_15227_44166# a_16335_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3090 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3091 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3092 VSS a_20974_43370# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3093 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3095 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3096 VSS a_16327_47482# a_17021_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3097 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3098 a_16388_46812# a_17957_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X3099 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3100 a_n4318_37592# a_n1736_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3101 VSS a_20159_44458# a_19321_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3103 VDD a_9672_43914# a_2107_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3104 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3105 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3107 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3108 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3109 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3110 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3111 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3112 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3113 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3114 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3115 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3116 VSS a_6151_47436# a_8189_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3117 VDD a_12549_44172# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3118 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3119 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3121 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3122 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3123 a_6229_45572# a_6194_45824# a_5907_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3124 VDD a_19700_43370# a_n97_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3125 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3126 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3127 a_6851_47204# a_6491_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3128 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3129 a_8423_43396# a_n443_42852# a_8317_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3130 VDD a_19615_44636# a_18579_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3131 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3132 a_1755_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3133 a_18799_45938# a_18175_45572# a_18691_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3134 VDD a_7499_43078# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3135 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3136 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3137 VDD a_6765_43638# a_6655_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3138 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3139 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3140 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3141 a_n1741_47186# a_12005_46116# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3142 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3143 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3144 VDD a_22223_47212# a_21588_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3145 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3146 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3147 a_685_42968# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3148 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3149 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3150 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3151 a_10467_46802# a_11599_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3152 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3153 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3154 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3155 a_17749_42852# a_17701_42308# a_17665_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3156 VDD a_n443_42852# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X3157 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3158 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3159 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3161 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3162 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3163 a_18599_43230# a_18249_42858# a_18504_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3164 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3165 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3166 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3167 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3168 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3169 VDD a_7920_46348# a_7715_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3170 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3171 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3172 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3173 a_2809_45028# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3174 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3175 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3176 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3177 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3178 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3179 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3180 a_7832_46660# a_7715_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3181 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3182 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3183 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3184 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3185 VSS a_4905_42826# a_4520_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3186 a_3873_46454# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X3187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3188 VSS a_20202_43084# a_21421_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3189 a_6709_45028# a_6431_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3190 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3191 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3192 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3193 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3194 a_20623_43914# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3195 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3196 a_20193_45348# a_18494_42460# a_20205_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3197 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3198 VSS a_9313_45822# a_11459_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3199 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3200 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3201 a_n4318_39768# a_n2840_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3202 VSS a_22469_40625# a_22717_36887# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3203 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3204 a_6428_45938# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3205 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3206 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3207 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3208 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3209 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3210 a_n2104_46634# a_n1925_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3211 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3212 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3213 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 EN_VIN_BSTR_N VDD a_19120_35138# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X3215 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3216 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3217 a_2987_42968# a_1847_42826# a_2905_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3218 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3219 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3220 a_11031_47542# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3221 VSS a_12991_46634# a_12925_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3222 VDAC_Ni a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3223 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3225 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3226 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3227 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3228 VSS a_20894_47436# a_20843_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3230 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3231 a_10752_42852# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3232 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3233 a_13076_44458# a_9482_43914# a_13468_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3234 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3235 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3236 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3237 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3238 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3239 a_17970_44736# a_18248_44752# a_18204_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3240 a_5663_43940# a_5883_43914# a_5841_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3242 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3243 a_n2302_38778# a_n2312_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3244 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3246 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3248 a_16588_47582# a_15507_47210# a_16241_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3249 VSS a_4099_45572# a_3483_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3250 VSS a_14539_43914# a_16112_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3251 a_16867_43762# a_16243_43396# a_16759_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3252 a_n745_45366# a_n746_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3253 a_10518_42984# a_10835_43094# a_10793_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3254 C2_P_btm a_n3420_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3255 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3256 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3257 VIN_P EN_VIN_BSTR_P C5_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3258 a_n37_45144# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3259 VSS a_11341_43940# a_22223_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3260 VSS a_8530_39574# a_3754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3261 a_18287_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3264 a_20159_44458# a_20362_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3265 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3266 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3267 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3269 a_6969_46634# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3270 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3271 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3272 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3273 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3274 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3275 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3276 a_18861_43218# a_18817_42826# a_18695_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3277 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3278 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3280 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3281 a_11322_45546# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3282 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3283 a_n3674_37592# a_196_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3284 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3285 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3286 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3287 a_n1809_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3288 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3289 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3290 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3291 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3292 a_4419_46090# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3293 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3294 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3295 VDD a_11189_46129# a_11133_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X3296 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3297 a_15959_42545# a_15764_42576# a_16269_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3298 VIN_P EN_VIN_BSTR_P a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3299 VSS a_7640_43914# a_7584_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3300 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3301 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3302 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3303 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3304 a_16375_45002# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3305 a_4235_43370# a_3935_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3306 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3307 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3308 VDD a_n1699_44726# a_n1809_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3309 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3310 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3311 a_21177_47436# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X3312 a_7418_45394# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3313 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3314 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3315 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3316 a_22000_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3317 VDD a_7542_44172# a_7499_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3318 a_11309_47204# a_11031_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3319 VDD a_1307_43914# a_3353_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3321 a_3905_42308# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3322 a_8483_43230# a_8037_42858# a_8387_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3323 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3324 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3325 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3326 a_n2104_46634# a_n1925_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3327 a_7281_43914# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3328 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3329 a_9028_43914# a_9290_44172# a_9248_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3330 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3331 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3332 a_453_43940# a_175_44278# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3333 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3334 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3335 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3336 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3337 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3338 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3339 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3340 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3341 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3342 a_15521_42308# a_15486_42560# a_15051_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3344 VDD a_4700_47436# a_3785_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3345 a_18909_45814# a_18691_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3346 a_11551_42558# a_n97_42460# a_11633_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3347 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3348 VDD a_15227_44166# a_15415_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3349 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3350 VSS a_16327_47482# a_20397_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3351 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3352 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3353 VDD a_8270_45546# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3354 a_n809_44244# a_n984_44318# a_n630_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3355 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3356 VDD a_948_46660# a_1123_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3357 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3358 a_20766_44850# a_20679_44626# a_20362_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3359 VDD a_15009_46634# a_14180_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3360 a_13385_45572# a_10903_43370# a_13297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3361 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3362 VDD a_13777_45326# a_13807_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3363 VSS a_n755_45592# a_n39_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3364 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3365 a_14976_45028# a_14797_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3367 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3368 a_6886_37412# VDAC_Pi VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X3369 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3371 a_6419_46482# a_6165_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3372 a_n2302_37690# a_n2810_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3373 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3374 VSS a_768_44030# a_5244_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3375 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3376 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3377 a_20623_45572# a_20273_45572# a_20528_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3378 VDD a_8199_44636# a_8336_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3379 VSS a_9396_43370# a_5111_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3380 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3381 a_743_42282# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3382 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3383 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3384 a_20009_46494# a_18819_46122# a_19900_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3385 a_7309_42852# a_5891_43370# a_7227_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3386 a_n2312_39304# a_n1920_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3388 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3389 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3390 VSS a_n4064_40160# a_n2302_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3391 a_12991_43230# a_12545_42858# a_12895_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3393 a_22397_42558# a_n913_45002# a_17303_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3394 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3395 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3396 VSS a_3905_42865# a_5013_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3397 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3398 VSS C0_dummy_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3400 a_22765_42852# a_15743_43084# a_18184_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3401 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3402 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3403 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3405 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3406 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3407 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3408 a_7705_45326# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3409 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3410 a_3065_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3411 VSS a_10405_44172# a_8016_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3412 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3413 a_742_44458# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3414 VDD a_526_44458# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3415 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3417 a_310_45028# a_n37_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X3418 VDD a_3232_43370# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3419 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3420 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3421 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3422 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3423 VSS a_18184_42460# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X3424 a_19466_46812# a_13747_46662# a_19929_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3425 VDD a_16241_47178# a_16131_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3426 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3427 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3428 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3429 VSS a_768_44030# a_9028_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X3430 a_20850_46482# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3431 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3432 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3434 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3435 a_12089_42308# a_11551_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3436 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3437 a_11173_43940# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3438 a_3457_43396# a_1414_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3440 a_8034_45724# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3441 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3442 VDD a_5907_46634# a_5894_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3443 a_22000_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3444 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3445 a_5841_46660# a_4651_46660# a_5732_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3446 VSS a_3699_46348# a_3160_47472# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3447 VSS a_22223_45036# a_18114_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3448 a_2437_43396# a_1568_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3450 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3451 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3452 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3453 a_2448_45028# a_2382_45260# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3454 VDD a_n2104_46634# a_n2312_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3455 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3456 a_21167_46155# a_20916_46384# a_20708_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3457 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3459 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3461 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3462 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3463 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3464 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3465 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3466 a_5205_44484# a_5343_44458# a_5289_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3467 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3468 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3469 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3470 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3471 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3472 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3473 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3474 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3475 a_948_46660# a_33_46660# a_601_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3476 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3477 VSS a_21005_45260# a_19778_44110# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3478 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3479 a_9241_46436# a_n237_47217# a_8049_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3480 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3481 a_15015_46420# a_14840_46494# a_15194_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3482 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3483 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3484 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3485 VDD a_20567_45036# a_12549_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3486 a_22717_37285# a_22459_39145# a_22609_38406# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3487 a_21398_44850# a_20640_44752# a_20835_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3488 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3489 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3490 a_5527_46155# a_5204_45822# a_5068_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3491 a_1823_45246# a_4704_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3492 a_1606_42308# a_1576_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3493 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3494 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3496 VSS a_4235_43370# a_4181_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3497 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3498 VSS a_18194_35068# a_19120_35138# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3499 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3500 VDD a_18783_43370# a_18525_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3501 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3502 VCM a_5534_30871# C7_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3503 a_n881_46662# a_14495_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3504 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3505 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3506 a_21188_45572# a_20107_45572# a_20841_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3507 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3508 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3509 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3510 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3511 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3512 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3513 VSS a_8270_45546# a_8192_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3514 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3515 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3516 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3517 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3518 VDD a_n863_45724# a_3059_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3519 VDD a_17609_46634# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3520 VSS a_n755_45592# a_3503_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3521 a_19237_31679# a_22959_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3522 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3523 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3524 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3525 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3526 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3527 a_n4334_38528# a_n4318_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3528 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3529 a_12156_46660# a_11813_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3530 a_n901_43156# a_n1076_43230# a_n722_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3531 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3532 a_n2810_45028# a_n2840_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3533 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3534 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3535 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3536 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3539 a_16333_45814# a_16115_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3540 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3541 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3542 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3543 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3544 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3545 a_16795_42852# a_n97_42460# a_16877_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3546 a_6905_45572# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3547 VDD a_21188_46660# a_21363_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3549 VDD a_5934_30871# a_8515_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3550 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3551 a_14180_45002# a_13059_46348# a_14403_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3552 a_16405_45348# a_16375_45002# a_16321_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3553 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3554 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=10.615 ps=76.96 w=3.75 l=15
X3555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3556 VREF a_19963_31679# C3_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3557 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3558 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3559 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3560 VDD a_3422_30871# a_22315_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3561 a_2123_42473# a_n784_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3562 VSS a_n1613_43370# a_n1287_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3563 VSS a_22223_43948# a_14401_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3564 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3565 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3566 a_19518_43218# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3568 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3569 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3570 VSS a_20075_46420# a_20009_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3571 VSS a_16922_45042# a_16751_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3573 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3574 a_1049_43396# a_458_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3575 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3576 VDD a_3232_43370# a_11341_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X3577 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3578 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3579 VDD a_n237_47217# a_8270_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3580 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3581 a_1848_45724# a_n237_47217# a_1990_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3582 VDD a_14539_43914# a_12465_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3583 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3584 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3585 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3586 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3587 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3588 VDD a_n881_46662# a_7903_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3590 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3591 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3592 VDD a_n1423_46090# a_n1533_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3593 VDD a_5111_44636# a_5421_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3594 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3595 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3596 a_11778_45572# a_10193_42453# a_11688_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3597 a_20623_46660# a_20107_46660# a_20528_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3598 a_6347_46155# a_6165_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3599 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3600 VDD a_21359_45002# a_21101_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3601 a_4700_47436# a_n443_46116# a_4842_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3602 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3603 C4_P_btm a_n3565_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3605 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3606 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3607 VDD a_5755_42308# a_5932_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3608 a_14113_42308# a_13575_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3609 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3610 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3611 a_17333_42852# a_16795_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3613 a_10695_43548# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3615 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3616 a_4958_30871# a_17124_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3617 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3619 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3620 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3621 VSS a_19339_43156# a_19273_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3622 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3623 a_8387_43230# a_8037_42858# a_8292_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3624 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3625 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3626 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3627 VSS a_16327_47482# a_18861_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3628 VDD a_n2840_44458# a_n4318_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3629 VDD a_15004_44636# a_14815_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3630 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3631 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3632 VSS a_1823_45246# a_3602_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3633 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3635 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3636 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3638 a_n4334_37440# a_n4318_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3639 VDD a_18780_47178# a_13661_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3640 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3641 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3642 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3643 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3644 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3645 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3646 a_2455_43940# a_895_43940# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3647 a_13667_43396# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3648 CAL_P a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3649 a_2680_45002# a_3065_45002# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3650 a_21381_43940# a_21115_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3651 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3652 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3653 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3654 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3655 VSS a_22521_39511# a_22469_39537# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3656 a_15781_43660# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3657 a_380_45546# a_765_45546# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3659 a_16019_45002# a_16147_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X3660 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3662 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3663 a_5534_30871# a_12563_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3664 a_12741_44636# a_6755_46942# a_16789_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3665 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3667 VDD a_3537_45260# a_4558_45348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3668 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3669 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3670 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3671 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3672 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3673 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3675 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3676 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3677 VDD a_n473_42460# a_n1761_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3679 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3680 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3681 a_12895_43230# a_12545_42858# a_12800_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3682 a_20836_43172# a_20193_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3683 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3684 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3685 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3686 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3687 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3688 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3689 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3690 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3691 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3692 a_726_44056# a_626_44172# a_644_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3693 a_6655_43762# a_6031_43396# a_6547_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3695 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3696 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3697 VDD a_3232_43370# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3698 a_5343_44458# a_7963_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3699 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3700 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3701 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3702 a_2889_44172# a_1414_42308# a_3052_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3703 a_9313_44734# a_5883_43914# a_9241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3705 a_3483_46348# a_4099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3706 a_2809_45028# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3707 VDD a_6171_45002# a_11827_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3708 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3709 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3710 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3711 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3712 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3713 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3714 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3715 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3716 VDD a_9625_46129# a_9569_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X3717 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3718 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3719 a_15567_42826# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3720 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3721 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3722 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3723 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3724 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3725 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X3726 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3727 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3728 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3729 a_n2810_45572# a_n2840_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3732 a_7_45899# a_n443_46116# a_n452_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3733 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3734 VDD a_13259_45724# a_22397_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3735 a_5708_44484# a_3483_46348# a_5608_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3736 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3737 a_5732_46660# a_4817_46660# a_5385_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3738 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3740 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3741 VDD a_13507_46334# a_22765_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3742 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X3743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3744 VSS a_22521_40055# a_22459_39145# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3745 a_13678_32519# a_21855_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3746 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3747 a_5365_45348# a_5111_44636# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3748 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3749 a_17021_43396# a_16977_43638# a_16855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3750 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3751 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3752 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3753 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3754 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3755 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3756 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3757 a_7989_47542# a_n237_47217# a_7903_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3758 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3759 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3760 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3761 a_19332_42282# a_19511_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3762 VSS a_6851_47204# a_7227_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3763 a_13607_46688# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3764 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3765 a_4880_45572# a_526_44458# a_4808_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3766 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3767 a_20922_43172# a_10193_42453# a_20836_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3768 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3769 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3770 a_12978_47026# a_11901_46660# a_12816_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3771 VDD a_13720_44458# a_12607_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3772 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3773 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3774 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3775 VDD a_2952_47436# a_2747_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3776 a_5147_45002# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3777 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3778 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3779 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3780 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3781 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3782 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3783 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3784 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3785 VDD a_14513_46634# a_14543_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3786 VDD a_21259_43561# a_16922_45042# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3787 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3788 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3789 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3790 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3791 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3792 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3793 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3794 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3795 VDD a_21137_46414# a_21167_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3796 a_3905_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3797 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3798 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3799 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3800 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3801 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3802 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3803 VSS a_22959_47212# a_22612_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3804 VSS a_6755_46942# a_13556_45296# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3805 a_383_46660# a_33_46660# a_288_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3806 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3807 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3808 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3809 a_17061_44734# a_11691_44458# a_16979_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3810 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3811 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3812 a_4149_42891# a_2382_45260# a_3935_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X3813 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3814 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3815 VDD a_n755_45592# a_3318_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3816 VDD a_n443_46116# a_1427_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3817 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3818 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3819 VDD a_5497_46414# a_5527_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3821 a_5937_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3822 a_11323_42473# a_5742_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3823 VSS a_4921_42308# a_5755_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3824 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3826 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3827 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3828 a_21076_30879# a_22959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3829 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3830 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3831 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3832 VSS a_n755_45592# a_3318_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X3833 VDD a_17583_46090# a_13259_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3835 a_3699_46634# a_3524_46660# a_3878_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3836 VSS a_3600_43914# a_3499_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X3837 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3838 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3839 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3840 a_17595_43084# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3841 a_5111_44636# a_9396_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3842 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3843 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3844 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3845 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3846 a_13829_44260# a_13059_46348# a_13483_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3847 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3848 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3849 a_18341_45572# a_18175_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3850 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3851 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3852 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3854 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3855 a_12991_46634# a_12816_46660# a_13170_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3856 VSS a_2277_45546# a_2211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3857 a_18429_43548# a_18525_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X3858 VSS a_6453_43914# a_n2661_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3859 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3860 a_6773_42558# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3861 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3862 a_2253_44260# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X3863 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3864 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3865 a_9885_42558# a_7499_43078# a_9803_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3866 a_16414_43172# a_16137_43396# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X3867 a_3726_37500# a_6886_37412# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3868 a_2304_45348# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3869 a_21811_47423# SINGLE_ENDED VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3871 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3872 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3873 a_13351_46090# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3874 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3875 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3876 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3877 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3878 a_n1435_47204# a_n1605_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3879 a_n935_46688# a_n1151_42308# a_n1021_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3880 VSS a_12549_44172# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X3881 a_6977_45572# a_6598_45938# a_6905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X3882 a_11530_34132# EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3883 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3884 VSS a_n1177_43370# a_n1243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3885 VSS a_n23_44458# a_n89_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3886 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3887 VDD a_13460_43230# a_13635_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3888 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3889 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3890 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3891 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3892 VSS a_n913_45002# a_n967_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3893 VDD a_11525_45546# a_11189_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3894 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3895 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3896 VDD a_n755_45592# a_626_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3897 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3898 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3899 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3900 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3901 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3902 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3903 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3904 VDD a_10227_46804# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3905 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3907 a_895_43940# a_644_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3908 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3909 a_11136_42852# a_10922_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3910 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3911 a_n699_43396# a_n1177_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3913 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3914 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3915 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3916 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3917 VDD a_8568_45546# a_8162_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3918 a_11551_42558# a_n97_42460# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3919 a_6293_42852# a_5755_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3920 a_n2840_42826# a_n2661_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3921 a_14033_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3923 VSS a_n1736_42282# a_n4318_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3924 a_16131_47204# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3925 a_5289_44734# a_4223_44672# a_5205_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3926 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3927 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3928 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3929 VSS a_5147_45002# a_5708_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3930 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3931 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3932 VDD a_11415_45002# a_22591_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3933 VIN_N EN_VIN_BSTR_N C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3934 VSS a_6886_37412# a_4338_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3935 VDD a_13259_45724# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3936 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3937 a_10053_45546# a_10490_45724# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3938 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3939 VDD a_19332_42282# a_4190_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3940 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3941 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3942 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3943 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3944 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3945 a_n998_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3946 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3947 a_6671_43940# a_6109_44484# a_6453_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3948 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3949 a_3090_45724# a_18911_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X3950 VSS a_18287_44626# a_18248_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3951 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3952 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3953 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3954 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3955 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3956 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3957 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3958 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3959 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3960 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3961 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3962 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3963 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3964 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3965 a_16131_47204# a_15507_47210# a_16023_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3966 a_11750_44172# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3967 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3968 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3969 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3970 a_n23_44458# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3971 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3972 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3973 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3974 VIN_N EN_VIN_BSTR_N C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3975 a_7845_44172# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3976 VSS a_6123_31319# a_7963_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3977 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3978 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3979 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3980 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3981 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3982 a_8560_45348# a_8746_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3983 a_5907_46634# a_5732_46660# a_6086_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3984 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3985 a_19095_43396# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X3986 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3987 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3988 a_21363_46634# a_21188_46660# a_21542_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3989 VSS a_n4315_30879# a_n4251_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3990 VSS a_n4064_39616# a_n2302_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3991 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3992 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3993 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3994 a_14180_46482# a_14035_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3995 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3996 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3997 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3998 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3999 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4000 a_18315_45260# a_18587_45118# a_18545_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4001 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4002 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4003 a_8349_46414# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4004 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4005 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4006 VSS a_3499_42826# a_3445_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4007 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4008 a_2537_44260# a_2479_44172# a_2127_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4009 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4010 VDD a_3815_47204# a_4007_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4011 a_9306_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4012 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4013 VDD a_6667_45809# a_6598_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4014 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4015 a_7230_45938# a_6511_45714# a_6667_45809# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X4016 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4017 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4018 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4019 a_8685_43396# a_8147_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X4020 VDD a_1343_38525# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4021 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4022 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4023 VSS VSS a_3726_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X4024 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4025 a_8270_45546# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4026 a_3992_43940# a_768_44030# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4027 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4028 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4029 a_15765_45572# a_15599_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4031 a_3815_47204# a_3785_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4032 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4033 a_2063_45854# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4034 VDD a_19431_45546# a_19418_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4035 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4036 VSS a_14021_43940# a_22959_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4037 VSS a_11415_45002# a_22591_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4038 a_6755_46942# a_15015_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4039 a_19328_44172# a_19478_44306# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X4040 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4041 VDD a_768_44030# a_726_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4042 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4043 VSS a_10227_46804# a_14537_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4044 a_21073_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4045 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4046 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4047 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4048 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4049 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4051 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4052 VDD a_13059_46348# a_15297_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X4053 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4054 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4056 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4057 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4058 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4059 VSS a_12465_44636# a_22223_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4060 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4061 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4062 a_19164_43230# a_18083_42858# a_18817_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4063 VDD a_n1352_43396# a_n1177_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4064 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4065 VSS a_n863_45724# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4066 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4067 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4068 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4069 a_383_46660# a_n133_46660# a_288_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4070 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4071 a_13814_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4072 VSS a_9127_43156# a_9061_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4073 a_3524_46660# a_2443_46660# a_3177_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4075 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4076 VDD a_9482_43914# a_10157_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4077 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4078 VSS a_12607_44458# a_12553_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4079 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4080 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4081 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4082 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4083 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4084 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4085 VSS a_17499_43370# a_17433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4086 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4087 VSS a_10903_43370# a_11963_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4088 C1_P_btm a_1606_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4089 VSS a_14815_43914# a_14761_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4090 a_13213_44734# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4091 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4092 VDD a_12427_45724# a_10490_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4094 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4095 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4096 VSS a_11323_42473# a_10807_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4097 a_12513_46660# a_12469_46902# a_12347_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4098 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4099 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4100 VDD a_1209_43370# a_n1557_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4101 a_18989_43940# a_18451_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4102 VSS a_8667_46634# a_8601_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4104 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4105 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4107 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4108 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4109 a_2889_44172# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X4110 VSS a_7281_43914# a_7229_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4111 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4112 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4113 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4114 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4115 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4116 VSS a_21195_42852# a_21671_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4118 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4119 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4120 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4121 VSS a_n699_43396# a_4743_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X4122 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4123 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4124 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4125 VDD a_n443_46116# a_2437_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4126 a_n2956_38680# a_n2472_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4127 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4128 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4129 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4130 a_10553_43218# a_10518_42984# a_10083_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4131 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4132 VSS a_13635_43156# a_13569_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4133 a_16789_44484# a_14537_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4134 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4135 a_18834_46812# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4136 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4137 a_n1151_42308# a_n1329_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4138 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4139 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4140 a_10405_44172# a_7499_43078# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X4141 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4142 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4143 VSS a_18315_45260# a_18189_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X4144 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4145 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4146 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4147 VDD a_17499_43370# a_17486_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4148 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4149 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4150 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4151 VDD a_22223_42860# a_22400_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4153 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4154 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4155 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4156 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4157 VDD a_3524_46660# a_3699_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4158 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4160 a_10765_43646# a_10695_43548# a_10057_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X4161 a_15890_42674# a_15803_42450# a_15486_42560# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD a_12549_44172# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4163 VSS a_12861_44030# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4164 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4165 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4166 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4167 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4168 a_17433_43396# a_16243_43396# a_17324_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4169 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4170 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4171 a_11827_44484# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4172 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4173 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4174 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4175 a_1847_42826# a_2351_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4176 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4177 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4178 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4179 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4180 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4181 VSS a_6151_47436# a_14955_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4182 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4183 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4184 a_20205_31679# a_22223_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4185 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4187 VSS a_15227_44166# a_15785_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4188 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4190 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4191 VDD a_8667_46634# a_8654_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4192 a_n452_45724# a_n443_46116# a_n310_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4193 VDD a_1239_47204# a_1431_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4194 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4195 a_700_44734# a_n746_45260# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X4196 a_19862_44208# a_13747_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4197 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4199 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4200 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4201 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4202 a_10775_45002# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X4203 a_1115_44172# a_453_43940# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4205 a_3232_43370# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4206 VDD a_22959_44484# a_19237_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4207 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4208 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4209 a_n3690_38528# a_n3674_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4210 a_484_44484# a_n863_45724# a_327_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X4211 VDD a_14543_43071# a_13291_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4212 VSS a_12549_44172# a_21205_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4213 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4214 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4215 a_20512_43084# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4216 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4217 a_20256_43172# a_20202_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X4218 a_6761_42308# a_n913_45002# a_6773_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4219 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4220 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4221 a_n2840_42282# a_n2661_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4222 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4223 VDD a_19864_35138# a_21589_35634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4224 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4225 a_n2661_46098# a_1983_46706# a_2162_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4226 VDD a_8685_43396# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X4227 VSS a_15368_46634# a_15312_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4228 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4229 a_5429_46660# a_5385_46902# a_5263_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4230 VDD a_16855_45546# a_16842_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4231 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4232 a_1221_42558# a_1184_42692# a_1149_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X4233 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4234 a_11315_46155# a_11133_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4235 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4236 a_16522_42674# a_15803_42450# a_15959_42545# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X4237 a_n923_35174# EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4238 a_20885_46660# a_20841_46902# a_20719_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4239 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4240 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4242 a_14456_42282# a_14635_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4243 a_20719_45572# a_20273_45572# a_20623_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4244 a_1756_43548# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X4245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4246 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4248 a_n2472_42826# a_n2293_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4249 a_7276_45260# a_6709_45028# a_7418_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4250 VDD a_1823_45246# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4251 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4253 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4254 VDD a_22400_42852# a_22521_40055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4255 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4256 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4257 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4258 VSS a_3422_30871# a_22315_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4259 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4260 VDD a_10341_42308# a_11554_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X4261 a_n2497_47436# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4262 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4264 a_3260_45572# a_3218_45724# a_2957_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4265 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4266 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4267 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4269 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4270 a_11280_45822# a_2063_45854# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X4271 a_603_45572# a_310_45028# a_509_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4272 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4273 a_8746_45002# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4274 a_15002_46116# a_13925_46122# a_14840_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4275 a_2479_44172# a_2905_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4276 a_11064_45572# a_10903_43370# a_10907_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X4277 a_n906_45572# a_n971_45724# a_n1013_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X4278 a_21205_44306# a_20935_43940# a_21115_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4279 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4280 VDD a_n2840_46090# a_n2956_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4281 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4282 VDD a_6945_45028# a_22223_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4283 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4284 a_13556_45296# a_6755_46942# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4285 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4286 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4287 VCM a_7174_31319# C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4288 VDD a_8199_44636# a_9377_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4289 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4290 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4291 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4292 a_n4334_39392# a_n4318_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4293 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X4294 a_12710_44260# a_10903_43370# a_12603_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X4295 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4296 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4297 a_13777_45326# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4299 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4300 a_16522_42674# a_15764_42576# a_15959_42545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4301 a_14205_43396# a_13667_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X4302 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4303 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4304 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4307 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4309 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4310 a_6419_46155# a_5807_45002# a_6419_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4312 VDD a_5732_46660# a_5907_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4313 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4314 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4315 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4316 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4317 a_n2860_39866# a_n2956_39768# a_n2946_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4318 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4319 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X4320 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4321 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4322 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4323 a_18533_44260# a_18326_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4324 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4325 VDD a_13556_45296# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4326 a_5066_45546# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4327 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4328 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X4329 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4330 a_n901_46420# a_n1076_46494# a_n722_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4331 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4332 VSS a_11599_46634# a_18175_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4333 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4334 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4335 VSS a_11599_46634# a_18819_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4336 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4337 a_n3690_37440# a_n3674_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4338 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4339 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4340 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4341 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4342 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4344 a_n2442_46660# a_n2472_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4345 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4346 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4347 VSS a_n1435_47204# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X4348 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4349 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4350 a_8317_43396# a_n755_45592# a_8229_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4351 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4352 a_n3674_38216# a_n2104_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4353 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4354 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4355 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4356 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4357 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4358 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4359 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4360 a_n2312_40392# a_n2288_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4361 VSS a_22591_44484# a_17730_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4362 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4363 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4364 VDD a_n1079_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X4365 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4367 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4368 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4369 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4370 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4371 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4372 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4373 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4374 a_n97_42460# a_19700_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4376 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4377 a_3877_44458# a_3699_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4378 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4379 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4380 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4381 a_15368_46634# a_15143_45578# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4382 a_11206_38545# CAL_N a_4338_37500# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4383 a_4905_42826# a_5379_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4384 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4385 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4386 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4387 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4388 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4389 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4390 VSS a_10467_46802# a_10428_46928# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4391 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4392 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4393 a_9313_45822# a_9049_44484# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4394 a_21145_44484# a_20766_44850# a_21073_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4395 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4396 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4397 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4398 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4400 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4401 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4402 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4403 VSS a_22521_40599# a_22717_37285# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4404 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4405 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4406 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4407 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4408 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4409 VSS a_2680_45002# a_2274_45254# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4410 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4411 a_10768_47026# a_10554_47026# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X4412 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4413 VSS a_21671_42860# a_3422_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4415 a_5837_45028# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4416 C0_dummy_P_btm a_7174_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4417 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4418 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4419 a_n785_47204# a_n815_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4420 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4421 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4423 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4424 a_14537_43396# a_14358_43442# a_14621_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X4425 a_n1736_43218# a_n1853_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X4426 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4427 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4428 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4429 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4430 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4431 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4432 a_16877_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4433 a_6640_46482# a_5257_43370# a_6419_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4434 VDD a_3090_45724# a_17786_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X4435 a_15493_43396# a_14955_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4436 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4437 a_9823_46482# a_9569_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4438 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4439 VDD a_14021_43940# a_22959_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4440 VDD a_n3420_38528# a_n2860_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4441 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4442 VSS a_10227_46804# a_12513_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4443 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4444 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4445 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4446 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4447 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4448 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4449 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4450 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4451 VDD a_3483_46348# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4452 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4453 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4454 VSS a_17339_46660# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4455 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4456 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4457 VSS a_n1532_35090# a_n83_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4459 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4461 a_3699_46348# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X4462 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4463 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4464 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4465 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4466 VSS a_10533_42308# a_10723_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4467 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4468 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4469 a_18214_42558# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4470 VSS a_3537_45260# a_4223_44672# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4471 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4472 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4473 VSS a_14537_43396# a_14180_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4474 a_16501_45348# a_10193_42453# a_16405_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4475 VSS a_21259_43561# a_16922_45042# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4476 VSS a_15743_43084# a_15567_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4477 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4478 VDD a_22821_38993# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4479 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4480 VSS a_n2840_46634# a_n2956_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4481 a_9049_44484# a_8701_44490# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4482 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4483 VDD a_2382_45260# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4484 VDD a_n967_45348# a_n961_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4485 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4486 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4487 a_19615_44636# a_12861_44030# a_19789_44512# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4488 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4489 a_9863_46634# a_10150_46912# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X4490 VDD a_n881_46662# a_n745_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4491 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4492 a_n2109_45247# a_n2017_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4493 VDD a_21496_47436# a_13507_46334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4494 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4495 VSS a_n143_45144# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4496 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4497 a_19418_45938# a_18341_45572# a_19256_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4498 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4499 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4500 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4501 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4502 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4503 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4504 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4505 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4507 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4508 VDD a_n2438_43548# a_n2433_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4510 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4511 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4512 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4513 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4514 VDD a_5907_45546# a_5937_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X4515 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4516 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4517 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4518 C5_P_btm a_n4209_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4519 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4520 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4521 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4522 VSS a_n452_44636# a_n2129_44697# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4523 a_n4318_38680# a_n2472_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4524 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4525 a_n2472_42282# a_n2293_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4526 a_5608_44484# a_5111_44636# a_5518_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X4527 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4528 VDD a_742_44458# a_700_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4529 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4530 VSS a_7287_43370# a_7221_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4532 VSS a_768_44030# a_13720_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4533 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4534 a_n89_44484# a_n467_45028# a_n452_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4535 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4536 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4537 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4538 a_2609_46660# a_2443_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4539 VDD a_9290_44172# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4540 VSS a_n1613_43370# a_6809_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4541 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4542 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4543 a_556_44484# a_526_44458# a_484_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4544 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4545 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4546 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4547 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4549 a_2112_39137# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4550 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4551 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4552 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4553 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4554 VSS a_19328_44172# a_19279_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X4555 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4556 VDD a_n3420_37440# a_n2860_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4557 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4558 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4559 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X4560 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4561 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4562 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4563 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4564 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4565 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4568 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4569 a_13887_32519# a_22223_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4570 a_11387_46155# a_n1151_42308# a_11315_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4571 a_10341_43396# a_9803_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4573 a_10554_47026# a_10467_46802# a_10150_46912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X4574 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4576 VSS a_16137_43396# a_18548_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X4577 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4578 C0_P_btm a_n3420_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4579 VSS a_10227_46804# a_20885_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4580 VIN_P EN_VIN_BSTR_P C2_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4581 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4582 a_n452_45724# a_n743_46660# a_n310_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4583 a_11682_45822# a_11652_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X4584 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4585 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4586 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4587 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4588 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4589 VDD a_n2472_46090# a_n2956_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4590 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X4591 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4592 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4593 VSS a_13747_46662# a_14495_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X4594 VDD a_10809_44734# a_n2661_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4595 C0_dummy_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4596 VDD a_11322_45546# a_11280_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4597 VSS a_n1329_42308# a_n1151_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4598 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4599 VSS a_n4209_39590# a_n4251_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X4600 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4601 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4602 a_5649_42852# a_5111_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4603 VDD a_18479_47436# a_13747_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4605 a_3381_47502# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4606 VSS a_n746_45260# a_261_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4607 VDAC_P C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4608 VSS a_n913_45002# a_8325_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4609 a_17486_43762# a_16409_43396# a_17324_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4610 a_11136_45572# a_3483_46348# a_11064_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4611 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4612 VSS a_13249_42308# a_13904_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4613 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4614 VSS a_1307_43914# a_2675_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4615 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4617 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4618 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4619 VSS a_n1532_35090# a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4620 VSS a_13259_45724# a_14797_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X4621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4622 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4623 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4625 a_3699_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4626 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4627 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4628 VIN_N EN_VIN_BSTR_N C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X4629 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4630 a_20841_45814# a_20623_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4631 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4632 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4633 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4635 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4636 a_10341_42308# a_9803_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4637 a_17639_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4638 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4639 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4640 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4641 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4642 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4643 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4644 a_20397_44484# a_20362_44736# a_20159_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4646 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4647 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4648 a_1260_45572# a_n755_45592# a_1176_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X4649 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4650 a_12991_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4651 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4652 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4653 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4654 a_518_46155# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4655 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4656 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4657 VDD a_20841_45814# a_20731_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4658 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4659 a_9751_46155# a_9569_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4660 a_1443_43940# a_1414_42308# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4661 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X4662 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4663 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4664 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4665 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4666 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4667 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4668 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4669 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4670 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4671 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4672 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4673 VDD a_11823_42460# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4675 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4676 VSS a_n2840_42826# a_n3674_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4677 VSS a_3537_45260# a_5365_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X4678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4679 a_21589_35634# a_19864_35138# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4680 a_3065_45002# a_3318_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4681 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4682 C8_P_btm a_n3420_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4683 a_n310_45899# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4684 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4685 VDD a_22591_46660# a_20820_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4686 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4687 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4688 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4689 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4690 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4691 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4692 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4693 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4695 a_8337_42558# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4696 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4697 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4698 VDD a_n1331_43914# a_n1441_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4699 VDD a_4646_46812# a_7411_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4700 VSS a_3877_44458# a_2382_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4701 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4702 a_11186_47026# a_10428_46928# a_10623_46897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4703 a_20273_46660# a_20107_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4704 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4705 VDD a_10835_43094# a_10796_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4706 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4707 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4708 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4709 VSS a_12883_44458# a_12829_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4710 a_11341_43940# a_10729_43914# a_11257_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X4711 VSS a_564_42282# a_n1630_35242# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4712 VSS a_5066_45546# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4713 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4714 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4715 a_12549_44172# a_20567_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4716 VDD a_14456_42282# a_5342_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4717 VDD a_2063_45854# a_10809_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4718 VDD a_10227_46804# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X4719 a_645_46660# a_601_46902# a_479_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4720 VDD a_2127_44172# a_n2661_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X4721 a_n2840_46090# a_n2661_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4722 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X4723 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X4724 a_14513_46634# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4725 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4726 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4727 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4728 a_14635_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4729 a_21137_46414# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4730 a_1609_45822# a_167_45260# a_1609_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4731 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4732 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4733 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4734 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4735 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4736 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4737 a_10544_45572# a_10490_45724# a_10053_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4738 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4739 a_10555_44260# a_10949_43914# a_10405_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4740 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4741 C2_P_btm a_n3565_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4742 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4743 a_8952_43230# a_7871_42858# a_8605_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4744 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4745 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4746 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4747 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4748 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4749 VDD a_1736_39587# a_1239_39587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4750 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4751 a_9377_42558# a_8685_42308# a_9293_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4752 a_3067_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4753 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4754 a_4190_30871# a_19332_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4755 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4756 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4757 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4758 a_15861_45028# a_15595_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4759 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4760 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4761 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4762 a_13720_44458# a_9482_43914# a_14112_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X4763 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4764 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4765 a_16245_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X4766 a_6469_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X4767 VSS a_n357_42282# a_6101_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4768 a_15194_46482# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4769 a_15493_43940# a_14955_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4770 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4771 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4772 a_20692_30879# a_22959_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4774 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4775 a_5497_46414# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4776 VSS a_104_43370# a_n971_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4777 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4778 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4779 a_5907_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4780 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4781 a_3177_46902# a_2959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4782 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4783 VREF_GND a_13258_32519# C0_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4784 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4785 VDD a_4743_44484# a_4791_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4786 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4787 a_19700_43370# a_18579_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4788 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X4789 a_21363_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4790 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4791 VSS a_n443_42852# a_15940_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X4792 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4793 a_12427_45724# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X4794 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4795 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4796 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4798 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4799 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4800 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4801 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4802 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4803 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4804 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4805 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4806 a_n1920_47178# a_n1741_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4807 a_10903_43370# a_13351_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4808 a_n955_45028# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4809 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4810 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4811 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4812 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4813 VDD a_n357_42282# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4814 a_4185_45028# a_3065_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4815 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4816 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4817 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4818 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4819 a_18596_45572# a_18479_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4820 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4821 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4822 a_16137_43396# a_15781_43660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X4823 a_6575_47204# a_6545_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4824 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4826 a_4649_42852# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4827 VSS a_n2472_46634# a_n2442_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4828 VSS a_2711_45572# a_20107_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4829 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4831 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4832 VSS a_n2104_42282# a_n3674_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4833 VIN_N EN_VIN_BSTR_N a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4834 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4835 VSS a_15015_46420# a_14949_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4836 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4837 VSS a_5691_45260# a_n2109_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4838 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4839 a_17730_32519# a_22591_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4840 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4841 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4842 a_3600_43914# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4843 a_17583_46090# a_17715_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X4844 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4845 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4846 a_13925_46122# a_13759_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4847 VDD a_n901_43156# a_n914_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4848 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4849 a_8191_45002# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4850 a_n310_44484# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4851 a_21125_42558# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4852 VDD a_22959_46124# a_20692_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4854 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4855 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4856 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4857 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4858 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4859 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4860 VSS a_14543_43071# a_13291_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4861 a_5932_42308# a_5755_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4862 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4863 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4864 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4865 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4866 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4867 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4868 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4869 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4870 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4871 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4872 VDD a_16112_44458# a_14673_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X4873 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4875 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4876 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4877 a_3175_45822# a_3316_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4878 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4879 VSS a_16763_47508# a_5807_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4880 VREF a_20447_31679# C5_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4881 a_14226_46660# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4882 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4883 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4884 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4885 VDD a_13348_45260# a_13159_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4886 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4887 VDD a_6491_46660# a_6851_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4888 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4890 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4891 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4892 a_6511_45714# a_4646_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4893 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4894 a_3422_30871# a_21671_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4895 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4896 VDD a_2889_44172# a_413_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X4897 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4898 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4899 VSS a_16763_47508# a_16697_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4900 VSS a_n443_42852# a_1755_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4901 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4902 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4903 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4904 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4905 a_10405_44172# a_10729_43914# a_10651_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4907 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4908 a_n2840_45546# a_n2661_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4909 a_14401_32519# a_22223_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4910 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4911 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4913 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4914 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4916 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4917 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4918 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4919 a_4558_45348# a_4574_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4920 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4921 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4923 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4924 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4926 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4927 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4928 a_5193_42852# a_3905_42865# a_5111_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4929 a_18143_47464# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4930 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4931 a_10533_42308# a_n913_45002# a_10545_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4932 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4933 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4934 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4935 VDD a_16721_46634# a_16751_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4936 a_18909_45814# a_18691_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4937 a_n2840_45002# a_n2661_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4938 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4939 a_948_46660# a_n133_46660# a_601_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4940 a_117_45144# a_n443_42852# a_45_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X4941 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4942 a_11415_45002# a_13249_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4943 a_3699_46348# a_3877_44458# a_3873_46454# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4944 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4945 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4946 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4947 a_15681_43442# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4948 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4949 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4950 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X4951 VDD a_n1059_45260# a_18727_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4952 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4953 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4955 a_n4251_38304# a_n4318_38216# a_n4334_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4956 VSS a_5013_44260# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4957 a_9801_43940# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4958 a_22521_39511# a_22545_38993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X4959 VSS a_10193_42453# a_18797_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4960 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4961 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4962 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4963 a_19789_44512# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X4964 VDD a_18057_42282# a_n356_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4965 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4966 a_2779_44458# a_1423_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4967 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4968 a_13113_42826# a_12895_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4969 a_16197_42308# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4970 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4971 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4972 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4974 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4975 VDD a_8034_45724# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4976 VDD a_11691_44458# a_11649_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4977 a_15761_42308# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X4978 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4979 a_n3690_39392# a_n3674_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4980 VSS a_1568_43370# a_1512_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4981 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4982 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4983 a_16680_45572# a_15765_45572# a_16333_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4985 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4986 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4987 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4989 VDD a_5066_45546# a_5024_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4990 VSS a_n809_44244# a_n875_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4991 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4993 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4994 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4995 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4996 a_10518_42984# a_10796_42968# a_10752_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X4997 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4998 a_n2267_43396# a_n2433_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4999 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5000 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5001 a_8189_46660# a_8145_46902# a_8023_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5002 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5003 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5004 VSS a_n4064_39072# a_n2302_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X5005 VDD a_13661_43548# a_14976_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X5006 a_11691_44458# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5007 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5008 VSS a_5891_43370# a_5837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5009 a_20062_46116# a_18985_46122# a_19900_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5010 a_20269_44172# a_20365_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X5011 VSS a_n2472_42826# a_n4318_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5012 a_18707_42852# a_18083_42858# a_18599_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5013 VSS a_7754_38470# a_7754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5014 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5015 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5016 a_n784_42308# a_n961_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5017 a_12638_46436# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5018 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5019 a_13157_43218# a_13113_42826# a_12991_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5020 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5021 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5023 VDD a_15015_46420# a_15002_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5024 VDD a_16327_47482# a_20159_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5025 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5026 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5027 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5028 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5029 VSS a_n785_47204# a_327_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X5030 a_18834_46812# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5031 a_n2840_45546# a_n2661_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5032 VSS a_21177_47436# a_20990_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5034 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5035 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5036 VSS a_7499_43078# a_11816_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5037 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5038 a_6761_42308# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5040 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5041 a_10623_46897# a_10428_46928# a_10933_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X5042 a_5263_45724# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X5043 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5044 VDD a_11823_42460# a_11322_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5045 VSS a_5111_44636# a_8018_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5046 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5047 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5048 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5049 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5050 a_3357_43084# a_4905_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5051 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5052 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5053 a_7903_47542# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5054 VSS a_8667_46634# a_n237_47217# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5056 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5057 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5058 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5059 a_n2472_46090# a_n2293_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5060 VREF a_19237_31679# C0_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X5061 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5062 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5063 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5064 VCM a_5742_30871# C6_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5065 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5066 a_10249_46116# a_9823_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X5067 a_2684_37794# VDAC_Pi a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5068 VSS a_22959_46660# a_21076_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5069 VDD a_10775_45002# a_10180_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5070 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5071 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X5072 a_13467_32519# a_21487_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5073 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5074 a_8696_44636# a_16855_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5075 a_6633_46155# a_5807_45002# a_6419_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X5076 a_n2661_42834# a_8975_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5077 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5078 a_7274_43762# a_6197_43396# a_7112_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5079 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5080 a_10922_42852# a_10835_43094# a_10518_42984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X5081 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5082 VDD a_5807_45002# a_11691_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5083 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5084 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5085 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5086 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5087 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5088 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5089 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5090 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5091 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5092 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5093 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5095 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5096 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5097 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5098 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5099 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5100 VSS RST_Z a_14311_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5101 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5102 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5103 a_18285_46348# a_18834_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5104 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5105 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5107 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5108 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5109 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5110 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5111 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5112 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5113 VSS a_18443_44721# a_18374_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X5114 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5115 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5116 a_18597_46090# a_19431_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5118 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5119 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5120 VSS a_8199_44636# a_10951_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5121 a_7735_45067# a_6709_45028# a_7276_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X5122 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5123 a_1176_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X5124 C8_P_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5125 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5126 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5127 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5128 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X5129 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5130 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5131 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X5132 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5133 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5134 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5135 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5136 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5137 VSS a_n2109_45247# en_comp VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5139 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5140 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5141 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5142 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5143 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5144 a_13348_45260# a_13556_45296# a_13490_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5145 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5146 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5147 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5148 a_n2302_40160# a_n2312_40392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5149 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5150 VSS a_21356_42826# a_n357_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5151 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5153 VDD a_11453_44696# a_22959_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5154 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5155 VSS a_8696_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5156 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5157 VSS a_15037_45618# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5158 a_3878_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5160 a_626_44172# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5161 a_2277_45546# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5162 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5163 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5164 a_18479_45785# a_19268_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X5165 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X5166 a_20273_45572# a_20107_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5167 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5168 VSS a_n443_42852# a_742_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5169 VSS a_n901_43156# a_n967_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5170 a_10555_44260# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X5171 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5172 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5173 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5174 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5175 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5176 a_20820_30879# a_22591_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5178 a_17364_32525# a_22959_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5179 VSS a_13076_44458# a_12883_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5181 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5182 a_685_42968# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5184 a_11633_42558# a_9290_44172# a_11551_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5185 a_13170_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5186 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5188 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5189 a_20731_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5190 VDD a_4791_45118# a_6633_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X5191 a_19700_43370# a_18579_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5192 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5193 a_2382_45260# a_3877_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5194 VDD a_11599_46634# a_20107_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5195 a_16751_45260# a_17023_45118# a_16981_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5196 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5197 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5198 a_11257_43940# a_10807_43548# a_11173_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5199 a_12829_44484# a_12741_44636# a_n2293_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5200 VCM a_6123_31319# C4_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5201 a_5342_30871# a_14456_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5202 VDD a_5937_45572# a_8034_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5203 VSS a_14084_46812# a_14035_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5204 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5205 a_17639_46660# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X5206 a_10809_44734# a_10057_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5207 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5208 VDD a_11823_42460# a_14853_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5209 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5210 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5211 a_20749_43396# a_20974_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5212 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5213 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5214 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5215 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5217 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5218 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5219 a_19511_42282# a_n913_45002# a_21125_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5220 VDD a_11967_42832# a_16243_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5221 a_17517_44484# a_16979_44734# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5222 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5223 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5224 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5225 a_1609_45572# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5226 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5227 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5228 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5229 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5230 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5231 a_20075_46420# a_19900_46494# a_20254_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5232 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5233 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5234 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5235 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5236 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5237 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5238 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5239 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5240 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5241 a_16020_45572# a_15903_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5242 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5243 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5244 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5245 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5246 a_20731_45938# a_20107_45572# a_20623_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5248 VDD a_n3420_39072# a_n2860_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X5249 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5250 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5253 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5254 a_16855_45546# a_16680_45572# a_17034_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5255 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5256 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5257 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5258 VSS a_22731_47423# a_13717_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5259 a_18114_32519# a_22223_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5260 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5261 VSS a_18429_43548# a_16823_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5262 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5263 VSS a_8325_42308# a_8791_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5264 a_17339_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5265 a_n2472_45546# a_n2293_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5266 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5267 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5268 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5269 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5270 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5271 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5272 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5273 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5275 VSS a_768_44030# a_13076_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X5276 VSS a_12861_44030# a_19692_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5277 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5278 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5279 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5280 VDD a_14495_45572# a_n881_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5281 a_18596_45572# a_18479_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5282 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5283 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5284 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5285 a_n2472_45002# a_n2293_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5286 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5287 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5288 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5289 a_3445_43172# a_3357_43084# a_n2293_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5290 a_5326_44056# a_5147_45002# a_5244_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5291 VSS a_22959_42860# a_14097_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5292 VDD a_n881_46662# a_6431_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5293 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5294 a_13003_42852# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5295 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5296 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5299 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5300 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5301 a_3503_45724# a_3775_45552# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5302 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5303 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5304 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5305 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5306 C6_N_btm a_14401_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5307 a_3540_43646# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5309 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5310 a_19929_45028# a_19778_44110# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5311 VDD a_167_45260# a_117_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5312 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5313 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5314 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5315 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5316 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5317 a_3147_46376# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X5318 a_6086_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5319 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5320 a_n1533_46116# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5321 VSS a_n3565_38216# a_n3607_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5322 a_5337_42558# a_5267_42460# a_4905_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X5323 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5324 a_21542_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5325 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5326 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5327 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5328 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5329 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5330 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5331 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5332 a_10216_45572# a_10180_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X5333 a_3626_43646# a_3232_43370# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5334 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5335 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5336 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5337 a_4699_43561# a_3080_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5338 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5339 a_1067_42314# a_1184_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5340 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5342 VDD a_21613_42308# a_22775_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5343 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5344 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5345 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X5346 a_16269_42308# a_15890_42674# a_16197_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X5347 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5348 VDD a_5937_45572# a_6945_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5349 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5350 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5351 a_22545_38993# a_22459_39145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5352 a_21356_42826# a_21381_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5353 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5354 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5355 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5356 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5357 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5358 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5359 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5360 VSS a_19862_44208# a_19808_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5361 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5362 VDD a_1307_43914# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5363 VDD a_5891_43370# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5364 a_20256_43172# a_18494_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X5365 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5366 VREF_GND a_13887_32519# C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5367 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5368 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X5369 a_7927_46660# a_7411_46660# a_7832_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5371 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5372 a_n2472_45546# a_n2293_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5373 VSS C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5374 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5376 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5377 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5378 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5379 a_4649_42852# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5380 a_17668_45572# a_n881_46662# a_17568_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X5381 VSS a_15493_43396# a_19478_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5382 a_16664_43396# a_16547_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5383 VDD a_6511_45714# a_6472_45840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5384 a_6540_46812# a_3877_44458# a_6682_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5385 VDD a_5068_46348# a_4955_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5386 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5387 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5388 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5389 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5390 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5391 a_9159_44484# a_5883_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5392 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5393 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5394 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5396 VSS a_10341_43396# a_22591_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5397 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5398 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5399 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5400 VSS a_17124_42282# a_4958_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5401 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5402 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5403 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5404 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5405 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5406 a_5267_42460# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X5407 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5408 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5409 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5410 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5411 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5412 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5413 a_1138_42852# a_791_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X5414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5415 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5416 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5417 a_n4318_40392# a_n2840_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5418 a_n1644_44306# a_n1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X5419 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5421 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X5422 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5423 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5424 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5425 a_5267_42460# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5426 VDD a_1609_45822# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X5427 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5428 VREF_GND a_17364_32525# C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X5429 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5430 a_2127_44172# a_2675_43914# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5431 a_11787_45002# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X5432 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5433 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5434 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5435 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5436 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5437 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5438 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5439 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5440 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5441 a_n2946_37984# a_n2956_38216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5442 VSS a_19333_46634# a_19123_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5443 a_3316_45546# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X5444 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5445 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5446 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5447 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5448 VSS a_13777_45326# a_13711_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5449 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5450 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5451 a_20712_42282# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5452 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5453 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5454 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5455 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5456 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5457 a_20573_43172# a_20512_43084# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X5458 a_19479_31679# a_22223_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5460 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5462 a_n2293_46634# a_14673_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5463 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5464 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5465 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5466 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5467 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5468 VSS a_526_44458# a_5457_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5469 a_33_46660# a_n133_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5470 VDD a_10903_43370# a_10849_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X5471 VDD a_7754_40130# a_7754_40130# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X5472 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5473 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5474 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5475 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5476 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5477 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5478 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5479 a_8495_42852# a_7871_42858# a_8387_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5480 a_5495_43940# a_5244_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5481 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5482 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5483 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5484 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5485 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5486 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5487 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5488 a_16842_45938# a_15765_45572# a_16680_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5489 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5490 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5491 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5492 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5493 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5494 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5495 VSS a_n961_42308# a_n784_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5496 VDD a_167_45260# a_2521_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5497 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5499 VSS a_13259_45724# a_17303_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5500 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5501 a_22780_40945# COMP_P a_22521_40599# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5502 a_17538_32519# a_22959_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5503 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5504 VDD a_5937_45572# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X5505 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5507 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5508 a_5742_30871# a_10723_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5509 a_9801_43940# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5510 a_21496_47436# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5511 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5512 a_11816_44260# a_11750_44172# a_10729_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5513 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5514 a_2123_42473# a_n784_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5515 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5516 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5517 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5518 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5519 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5520 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5521 a_13565_43940# a_12891_46348# a_13483_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5522 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5523 a_7227_42852# a_n97_42460# a_7309_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5524 VDD a_13747_46662# a_13607_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5525 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5526 a_5257_43370# a_5907_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5527 a_1667_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X5528 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5529 a_n2293_46098# a_5663_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X5530 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5531 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5532 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5533 a_13003_42852# a_12379_42858# a_12895_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5534 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5535 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5536 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5537 a_2711_45572# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5538 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5539 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5540 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5541 a_4883_46098# a_21363_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5542 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5543 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5544 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5545 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X5546 VSS a_16751_45260# a_6171_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X5547 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5548 a_16763_47508# a_16588_47582# a_16942_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5549 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5550 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5551 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5552 a_11750_44172# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5553 VDD a_20835_44721# a_20766_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X5554 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5555 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5556 VSS a_15861_45028# a_17668_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X5557 a_7845_44172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5558 a_15597_42852# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5559 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5560 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5561 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5562 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5563 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5564 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5565 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5568 VSS a_9223_42460# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X5569 VDD a_11967_42832# a_18083_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5570 a_13487_47204# a_13381_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5572 C2_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5573 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5574 a_13297_45572# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X5575 a_n923_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X5576 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5577 VDD a_n3565_38216# a_n3690_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X5578 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5580 C10_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5581 a_6101_43172# a_5891_43370# a_5755_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5582 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5583 a_11901_46660# a_11735_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5584 a_16979_44734# a_14539_43914# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5585 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5586 VSS a_14955_47212# a_10227_46804# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5587 a_18443_44721# a_18248_44752# a_18753_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X5588 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5590 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5592 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5593 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5594 VDD a_18909_45814# a_18799_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X5595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5596 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5597 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5598 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5599 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5600 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5601 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5602 a_1431_46436# a_1138_42852# a_1337_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5603 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5604 VDD a_n4064_37984# a_n2216_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X5605 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5606 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5607 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5608 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5609 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5610 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5611 VDD a_22521_40599# a_22469_40625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5612 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5613 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5616 VDD a_768_44030# a_5326_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5617 a_18443_44721# a_18287_44626# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X5618 VSS a_n4209_39304# a_n4251_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5619 a_n357_42282# a_21356_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5620 a_491_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5622 VSS a_n2288_47178# a_n2312_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5623 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5624 VCM a_1606_42308# C1_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5625 VDD a_20712_42282# a_10193_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5626 VSS a_3483_46348# a_15301_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5627 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X5628 a_n901_46420# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5629 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5630 a_5068_46348# a_5204_45822# a_5210_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5631 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5632 a_14033_45822# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5633 VSS a_6761_42308# a_7227_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5634 VSS a_11599_46634# a_20107_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5635 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5636 w_1575_34946# EN_VIN_BSTR_P VDD w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5638 VDD a_13661_43548# a_15595_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5639 a_9803_42558# a_n97_42460# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5640 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5641 VDD a_10227_46804# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X5642 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5643 a_n1177_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5644 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5645 VREF_GND a_n3420_39616# C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5646 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5647 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5648 a_601_46902# a_383_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X5649 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X5650 a_5024_45822# a_n443_46116# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X5651 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5652 a_17701_42308# a_17531_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5653 VSS a_12861_44030# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X5654 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X5655 a_6598_45938# a_6472_45840# a_6194_45824# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X5656 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5657 a_4808_45572# a_1823_45246# a_4419_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X5658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5659 a_n3607_38304# a_n3674_38216# a_n3690_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X5660 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5661 a_n229_43646# a_n2497_47436# a_n447_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5662 VSS a_6969_46634# a_6903_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5663 a_18214_42558# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X5664 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5667 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5669 VSS a_4883_46098# a_10355_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X5670 VDD a_4646_46812# a_6031_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5671 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5672 a_491_47026# a_n133_46660# a_383_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5673 VDD a_16327_47482# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X5674 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5675 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5676 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5677 VSS a_n1613_43370# a_n1655_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5679 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5680 a_6812_45938# a_6598_45938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X5681 a_8147_43396# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5682 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5683 a_12427_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X5684 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5685 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5686 VDD a_19594_46812# a_19551_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X5687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5688 a_n4318_37592# a_n1736_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5689 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5690 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5691 VSS a_1736_39043# a_1239_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5692 a_1414_42308# a_1067_42314# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X5693 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5694 VSS a_2698_46116# a_2804_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5695 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5696 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5697 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5698 VSS a_5649_42852# a_22223_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5699 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5700 VDD a_13259_45724# a_14797_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X5701 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5702 a_4817_46660# a_4651_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5703 a_n2288_47178# a_n2109_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5704 a_8062_46155# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5705 VDD a_20623_43914# a_20365_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X5706 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5707 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5708 a_13296_44484# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X5709 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5710 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5711 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5712 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5713 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5714 a_11601_46155# a_11309_47204# a_11387_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X5715 a_10210_45822# a_8746_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5716 a_18287_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5717 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5718 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5719 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5720 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5721 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5722 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5723 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5724 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5725 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5726 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5727 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5728 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5729 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5730 VSS a_11189_46129# a_11133_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X5731 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5732 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X5733 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5734 a_6109_44484# a_5518_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5735 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5736 a_6431_45366# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5737 a_14021_43940# a_13483_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5738 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5740 a_17499_43370# a_17324_43396# a_17678_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5741 a_3495_45348# a_3429_45260# a_3316_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X5742 VDD a_1115_44172# a_n2293_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X5743 VDD a_19787_47423# a_19594_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5744 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5745 a_18707_42852# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5746 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5747 a_1208_46090# a_n881_46662# a_1431_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5748 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5749 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5750 a_5431_46482# a_n1151_42308# a_5068_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X5751 a_8667_46634# a_8492_46660# a_8846_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5752 a_19787_47423# START VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5753 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5754 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5755 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5756 a_n2302_39866# a_n2442_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5757 VSS a_n2438_43548# a_2443_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5758 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5759 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5760 a_18797_44260# a_13661_43548# a_18451_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5761 a_19551_46910# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5762 VDD a_10341_43396# a_22591_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5763 a_8697_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X5764 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5765 VDD a_8953_45546# a_8049_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5766 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5767 a_12005_46116# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5768 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5769 VSS a_2123_42473# a_1184_42692# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5770 VSS a_12861_44030# a_18911_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X5771 a_1241_43940# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X5772 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5774 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5775 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5776 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5777 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5778 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5779 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5780 a_16285_47570# a_16241_47178# a_16119_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5781 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5782 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5783 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5784 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5785 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5786 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5787 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5788 VSS a_961_42354# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5789 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X5790 a_10617_44484# a_10440_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5791 a_1423_45028# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5792 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5793 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5794 C7_P_btm a_n4064_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X5795 VDD a_4704_46090# a_1823_45246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5796 a_18479_47436# a_20075_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5797 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5798 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5799 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5800 a_19987_42826# a_10193_42453# a_20573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5801 VDD a_9313_45822# a_11459_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5802 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5803 a_n1809_44850# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5804 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5805 VSS a_3785_47178# a_3815_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5806 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5807 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5808 VDD a_5891_43370# a_8375_44464# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5809 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5810 VSS a_9863_46634# a_2063_45854# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X5811 a_7920_46348# a_n1151_42308# a_8062_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5812 a_19721_31679# a_22959_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5813 a_19808_44306# a_19778_44110# a_19328_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5814 VDD a_10193_42453# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5815 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5816 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5817 VDD a_15559_46634# a_13059_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5818 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5819 VSS a_n2840_43370# a_n4318_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5821 a_15037_43396# a_14205_43396# a_14955_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X5822 VDD a_11189_46129# a_11601_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X5823 a_5263_45724# a_5257_43370# a_5437_45600# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5824 a_12495_44260# a_12429_44172# a_10949_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X5825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5826 a_6452_43396# a_6293_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5827 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5828 VSS a_4915_47217# a_12891_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5829 a_14084_46812# a_13885_46660# a_14226_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5831 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5832 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5833 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5835 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5836 a_19478_44306# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X5837 a_7705_45326# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5838 a_1115_44172# a_1307_43914# a_1241_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X5839 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5840 a_16981_45144# a_16922_45042# a_16886_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X5841 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5842 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5843 a_4223_44672# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5844 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5845 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5846 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5847 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5848 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5850 a_7174_31319# a_20107_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5851 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5852 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5854 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5855 VDD a_10227_46804# a_15051_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5856 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5857 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5858 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5859 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5860 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5861 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5862 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5863 VSS a_8103_44636# a_7640_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X5864 a_15146_44811# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5865 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5866 a_n2833_47464# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X5867 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5868 a_2903_45348# a_n971_45724# a_2809_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5869 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5870 VSS a_3537_45260# a_8103_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5871 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5872 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5873 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5875 VSS a_21137_46414# a_21071_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5876 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5877 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5878 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5879 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5880 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5881 VSS a_1414_42308# a_2889_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5882 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5883 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5884 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5885 VDD a_1848_45724# a_1799_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5886 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5887 VSS a_n13_43084# a_n1853_43023# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5888 a_18479_45785# a_19268_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5889 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5890 VSS a_19279_43940# a_21398_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X5891 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5892 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5893 a_1736_39587# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5894 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5895 VSS a_22485_44484# a_20974_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5896 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5897 VSS a_n3420_37984# a_n2946_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X5898 a_5841_44260# a_5495_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5899 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5900 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5901 a_5275_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5902 C5_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5903 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5904 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5905 a_n2661_45546# a_4093_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5906 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5907 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5908 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5909 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5910 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5911 VSS a_5497_46414# a_5431_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5912 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5913 VDD a_19339_43156# a_19326_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5914 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5915 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5916 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5917 VDD a_6123_31319# a_7963_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5918 a_8137_45348# a_8049_45260# a_n2293_42834# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5919 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5920 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5921 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5923 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5924 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5926 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5927 VDD a_12861_44030# a_17339_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5929 a_10849_43646# a_10807_43548# a_10765_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5930 VSS a_13507_46334# a_18997_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5931 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5933 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5934 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5935 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5936 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5937 a_8560_45348# a_3483_46348# a_8488_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X5938 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5939 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5940 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5941 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5942 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5943 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5944 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5945 a_13249_42308# a_13070_42354# a_13333_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5946 a_6969_46634# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5947 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5948 a_n2216_37984# a_n2810_45572# a_n2302_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X5949 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5950 VSS a_22223_46124# a_20205_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5951 VSS a_n1613_43370# a_n1379_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5952 a_6194_45824# a_6511_45714# a_6469_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X5953 a_n229_43646# a_n97_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5954 a_17613_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5955 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5956 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5957 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5958 VSS a_13747_46662# a_19862_44208# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5959 a_22821_38993# a_22400_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5960 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5961 a_17303_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5962 a_8649_43218# a_8605_42826# a_8483_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5963 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5964 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5965 VSS a_n901_46420# a_n967_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5966 a_15004_44636# a_13556_45296# a_15146_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5967 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5968 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5969 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5970 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5971 a_11186_47026# a_10467_46802# a_10623_46897# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X5972 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X5973 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5974 VSS a_526_44458# a_4169_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5975 a_3353_43940# a_2998_44172# a_2675_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5976 a_n23_45546# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5977 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5978 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5979 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5980 a_18326_43940# a_18079_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5981 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5982 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5983 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5984 a_20922_43172# a_19862_44208# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X5985 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5986 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5987 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5989 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5990 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5991 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5992 C5_P_btm a_5934_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X5993 a_10334_44484# a_10157_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5994 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5995 a_n2017_45002# a_19987_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X5996 VSS a_742_44458# a_1756_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5997 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5998 a_n2956_38216# a_n2472_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5999 VDD a_10193_42453# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6000 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6001 VDD a_8191_45002# a_n2293_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6002 a_13885_46660# a_13607_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6003 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6004 VSS RST_Z a_7754_39964# VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X6005 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6006 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6007 VSS a_4223_44672# a_n2497_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6008 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6009 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6010 a_4699_43561# a_3080_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6011 a_19511_42282# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6012 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6013 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6014 VSS a_19692_46634# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6015 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6016 VDD a_22591_43396# a_14209_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6017 a_n1991_46122# a_n2157_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6018 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6019 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X6020 VDD a_7499_43078# a_8746_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6021 a_n971_45724# a_104_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6023 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6024 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6025 a_20447_31679# a_22959_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6026 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6027 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6028 VDD a_15493_43940# a_22959_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6029 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6030 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6031 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6032 a_n4334_39616# a_n4318_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6033 VDD a_13527_45546# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X6034 a_18147_46436# a_17339_46660# a_17957_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X6035 a_8336_45822# a_8270_45546# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X6036 a_n2956_39304# a_n2840_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6037 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6038 VDD a_584_46384# a_766_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X6039 a_11361_45348# a_10907_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6040 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6041 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6042 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6043 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6044 VDD a_11599_46634# a_11735_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6045 a_19431_45546# a_19256_45572# a_19610_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6046 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6047 VSS a_9290_44172# a_12710_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X6048 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6049 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6050 VDD a_11323_42473# a_10807_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6051 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6052 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6053 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6054 a_2266_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6056 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6057 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6058 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6059 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6060 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6061 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6062 a_2982_43646# a_2479_44172# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6063 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6064 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6065 a_18280_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6066 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6067 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6068 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6069 C1_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X6070 VDD a_8492_46660# a_8667_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6071 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6072 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6073 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6075 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6076 VDD a_11967_42832# a_12379_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6077 VDD a_n1076_46494# a_n901_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6078 a_n4251_38528# a_n4318_38680# a_n4334_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6079 a_4361_42308# a_3823_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6080 VDD a_n971_45724# a_3775_45552# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6081 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6082 VDD a_11599_46634# a_13759_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6083 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6084 VDD a_21811_47423# a_20916_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6085 a_18985_46122# a_18819_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6086 VDD a_5649_42852# a_22223_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6087 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6088 VSS a_5343_44458# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6089 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6090 VSS a_3090_45724# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X6091 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6092 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6094 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6095 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6096 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6097 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6098 a_20528_45572# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6099 a_13487_47204# a_13717_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6100 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6101 VREF_GND a_13678_32519# C2_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X6102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6104 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6105 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6106 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6107 VDD a_20269_44172# a_19319_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6108 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6109 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6110 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6111 a_5807_45002# a_16763_47508# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X6112 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6113 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6114 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6115 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6116 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6117 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6118 VSS a_16327_47482# a_16285_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6119 a_n23_44458# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6120 VDD a_n1059_45260# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6121 a_1847_42826# a_2351_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6122 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6123 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6124 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6125 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6126 VSS a_3503_45724# a_3218_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X6127 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6128 a_19553_46090# a_19335_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6129 VDD a_n2840_45546# a_n2810_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6130 a_15037_45618# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6131 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6132 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6133 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6134 a_14537_43646# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6135 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6136 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6137 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6139 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6140 a_n1699_43638# a_n1917_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6141 VDD a_9313_44734# a_22959_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6142 C6_P_btm a_n3420_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6143 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6144 a_6671_43940# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6145 VSS a_5111_44636# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X6146 a_2124_47436# a_2063_45854# a_2266_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6147 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6148 VSS a_9625_46129# a_9569_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X6149 VDD a_3483_46348# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6150 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6151 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6152 VDD a_19279_43940# a_21398_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X6153 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6155 a_6171_42473# a_5932_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6156 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6157 a_17568_45572# a_8696_44636# a_17478_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X6158 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6162 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6163 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6164 a_18588_44850# a_18374_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X6165 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6166 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6167 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6168 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6169 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6171 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6172 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6173 a_18451_43940# a_18579_44172# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6174 VSS a_5755_42308# a_5932_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6175 a_2959_46660# a_2609_46660# a_2864_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6176 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6178 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6179 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6180 a_21359_45002# a_21513_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6181 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6182 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6183 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6184 a_7_47243# a_n746_45260# a_n452_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6185 a_14493_46090# a_14275_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6186 a_19478_44306# a_15493_43396# a_19478_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X6187 a_7287_43370# a_7112_43396# a_7466_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6188 a_15227_46910# a_3090_45724# a_15009_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6189 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6190 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6191 a_12251_46660# a_11901_46660# a_12156_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6192 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6193 a_8495_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6194 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6195 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6196 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6197 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6199 a_11633_42558# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6200 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6201 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6202 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6203 a_n4251_37440# a_n4318_37592# a_n4334_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6204 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6205 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6206 a_15279_43071# a_5342_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6207 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6208 VDD a_7276_45260# a_7227_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6209 VSS a_2479_44172# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X6210 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6211 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6212 VREF_GND a_14401_32519# C6_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X6213 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6214 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6215 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6216 VDD a_n815_47178# a_n785_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6217 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6218 VDD a_3877_44458# a_3699_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6219 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6220 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6221 a_9313_45822# a_5937_45572# a_9241_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X6222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6223 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6224 a_1239_47204# a_1209_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6225 a_20841_45814# a_20623_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6226 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6227 VDD a_805_46414# a_835_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6228 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6230 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6231 a_961_42354# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6232 a_12379_46436# a_12005_46116# a_n1741_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6233 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6234 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X6235 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6236 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6237 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6238 VDD a_5257_43370# a_3905_42865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6239 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6240 a_n1741_47186# a_12594_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6241 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6242 a_n2956_39768# a_n2840_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6243 VSS a_n473_42460# a_n1761_44111# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6244 a_13163_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X6245 a_10210_45822# a_10586_45546# a_10053_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6246 VDD a_10227_46804# a_9863_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6247 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6248 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6249 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6250 VSS a_4185_45028# a_22959_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6251 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6252 VDD a_n2438_43548# a_n2065_43946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6253 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6254 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6255 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6256 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6257 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6258 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6259 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6260 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6261 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6263 a_5457_43172# a_5111_44636# a_5111_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6264 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6266 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6267 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6268 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6269 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6270 a_10695_43548# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X6271 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6272 VDD a_11787_45002# a_11652_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X6273 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6274 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6275 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6276 a_13059_46348# a_15559_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6277 VDD a_n23_44458# a_7_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6278 a_12891_46348# a_4915_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6279 a_8023_46660# a_7577_46660# a_7927_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6280 VSS a_10057_43914# a_9672_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6281 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6282 a_20637_44484# a_20159_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X6283 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6284 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6285 a_n237_47217# a_8667_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X6286 a_n143_45144# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6287 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6288 a_4520_42826# a_4905_42826# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6289 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6290 VSS RST_Z a_8530_39574# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6291 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6292 VSS a_n971_45724# a_8423_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X6293 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6294 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6295 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6296 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6297 VSS a_3626_43646# a_19647_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6298 a_8697_45822# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X6299 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6300 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6301 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6302 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6303 a_3094_47243# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6304 a_15051_42282# a_15486_42560# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X6305 VDD a_1209_47178# a_1239_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6306 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6307 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6308 VDD a_13661_43548# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X6309 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6310 a_5167_46660# a_4817_46660# a_5072_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6311 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6312 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6313 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6314 VSS a_10835_43094# a_10796_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6315 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6316 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6317 VDD a_20708_46348# a_20411_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6318 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6319 VSS a_16327_47482# a_18005_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X6320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6321 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6322 VSS a_16292_46812# a_15811_47375# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6323 a_9482_43914# a_9838_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6324 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6325 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X6326 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6327 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6328 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6329 a_20623_46660# a_20273_46660# a_20528_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6330 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6331 VDD a_12594_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6332 a_18374_44850# a_18287_44626# a_17970_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X6333 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6334 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6335 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6336 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6337 a_16750_47204# a_15673_47210# a_16588_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6338 a_6545_47178# a_6419_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X6339 VDD a_22223_43396# a_13887_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6340 a_8783_44734# a_8696_44636# a_8701_44490# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6341 a_175_44278# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6342 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6343 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6344 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X6345 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6346 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6347 VDD a_18479_47436# a_20935_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6348 a_3754_38470# a_7754_38470# VSS sky130_fd_pr__res_high_po_0p35 l=18
X6349 VSS a_5907_46634# a_5841_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6350 a_5745_43940# a_5883_43914# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6351 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6352 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6353 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6354 a_1110_47026# a_33_46660# a_948_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6355 a_16434_46987# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6356 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6357 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6358 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6359 a_20974_43370# a_22485_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6360 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6361 a_2998_44172# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6362 a_13381_47204# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6363 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6364 VDD a_4921_42308# a_5755_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6365 a_10991_42826# a_10835_43094# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X6366 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6367 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6368 VDD a_6851_47204# a_7227_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6369 a_3052_44056# a_2998_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X6370 a_n1699_43638# a_n1917_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6372 CAL_N a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6373 a_3177_46902# a_2959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6374 a_9241_44734# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6376 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6377 VSS a_1208_46090# a_472_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6378 a_22365_46825# EN_OFFSET_CAL VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6379 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6380 VSS a_13163_45724# a_11962_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6381 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6382 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6383 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6384 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6385 a_3055_46660# a_2609_46660# a_2959_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6386 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6387 a_19326_42852# a_18249_42858# a_19164_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6388 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6389 a_9885_43646# a_8270_45546# a_9803_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6390 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6391 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6393 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6394 VDD a_18597_46090# a_16375_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6395 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6397 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6398 VSS a_22959_43396# a_17364_32525# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6399 a_19431_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6400 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6401 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6402 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6403 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6405 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X6406 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6407 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6408 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X6409 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6410 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6411 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6412 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6413 VSS a_n1177_44458# a_n1243_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6414 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6415 VSS a_n23_45546# a_n89_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6416 VDD a_12816_46660# a_12991_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6417 a_7499_43940# a_7640_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6418 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6419 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X6420 a_2952_47436# a_n1151_42308# a_3094_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6421 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6422 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6423 a_n452_47436# a_n746_45260# a_n310_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6424 a_4235_43370# a_3935_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X6425 a_5105_45348# a_4558_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6426 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6427 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6428 a_18051_46116# a_765_45546# a_17957_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X6429 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6430 a_n1441_43940# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6431 a_15301_44260# a_15227_44166# a_14955_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6432 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6434 VSS a_n3565_38502# a_n3607_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X6435 a_n746_45260# a_n1177_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6436 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6437 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6438 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6439 a_n2840_43914# a_n2661_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6440 a_6809_43396# a_6765_43638# a_6643_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6441 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6442 VSS a_376_46348# a_171_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6443 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6444 VSS a_8199_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6445 a_7499_43940# a_3090_45724# a_7281_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6446 a_9165_43940# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6447 a_19443_46116# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6448 VSS a_13059_46348# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6449 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6450 a_453_43940# a_175_44278# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6451 a_9885_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6452 a_n3674_39304# a_n2840_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6453 a_2959_46660# a_2443_46660# a_2864_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6454 a_14543_46987# a_13885_46660# a_14084_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6455 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6456 VDD a_413_45260# a_22959_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6457 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6461 a_17969_45144# a_16375_45002# a_17896_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6462 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6463 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6464 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6465 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6466 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6467 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6468 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6469 a_16292_46812# a_n743_46660# a_16434_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6470 a_21188_46660# a_20107_46660# a_20841_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6471 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6472 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6473 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6474 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6475 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6476 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6477 a_4365_46436# a_4185_45028# a_n1925_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6478 a_12251_46660# a_11735_46660# a_12156_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6479 a_n998_44484# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6480 VDD a_n2472_45546# a_n2956_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6481 a_7577_46660# a_7411_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6482 a_10835_43094# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6483 VDD a_3177_46902# a_3067_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6484 a_14976_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6485 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6486 VSS a_13661_43548# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6487 a_12638_46436# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6488 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6489 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6490 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6491 a_12839_46116# a_12891_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6492 VSS a_3090_45724# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6493 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6494 VSS a_22000_46634# a_15227_44166# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6495 VSS a_n863_45724# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6496 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6497 a_14209_32519# a_22591_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6498 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6499 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6500 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6501 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6502 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6503 a_n2012_43396# a_n2129_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6504 VSS a_11823_42460# a_14635_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6505 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6506 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6507 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6508 a_n2661_43922# a_12465_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6509 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6510 VSS a_4520_42826# a_4093_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6511 a_19692_46634# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6512 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6513 a_5013_44260# a_3905_42865# a_5025_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6514 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6515 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6516 VSS C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6517 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6518 a_8018_44260# a_7499_43078# a_7911_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X6519 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6520 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6521 VDD a_11823_42460# a_14358_43442# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X6522 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6523 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6524 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6525 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6526 a_742_44458# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6527 VDD a_10405_44172# a_8016_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X6528 a_20254_46482# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6529 VIN_N EN_VIN_BSTR_N C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X6530 a_167_45260# a_2202_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6532 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6533 VSS a_19332_42282# a_4190_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6534 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6535 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6536 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6537 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6539 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6540 a_20356_42852# a_18184_42460# a_20256_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X6541 a_14840_46494# a_13925_46122# a_14493_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6542 VSS a_1414_42308# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X6543 a_19006_44850# a_18287_44626# a_18443_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6544 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6545 a_9420_43940# a_768_44030# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X6546 VDD a_10903_43370# a_12005_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6547 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6548 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6549 VSS a_13661_43548# a_15685_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6550 VSS a_12861_44030# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6551 C4_P_btm a_6123_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X6552 a_13575_42558# a_n97_42460# a_13657_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6553 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6554 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6555 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6556 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6557 a_8667_46634# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6558 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6559 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6560 VDD a_n971_45724# a_n229_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X6561 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6562 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6563 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6564 a_21335_42336# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6565 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6566 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6567 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6568 VSS a_n3565_37414# a_n3607_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X6569 a_n2946_38778# a_n2956_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6570 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6572 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6573 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6574 VSS a_13351_46090# a_10903_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6576 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6577 a_743_42282# a_12549_44172# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6578 a_14309_45028# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X6579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6580 VSS a_413_45260# a_22959_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6581 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6582 VDD a_3877_44458# a_4185_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6583 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6584 a_13105_45348# a_13017_45260# a_n2661_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6585 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6586 a_8229_43396# a_7499_43078# a_8147_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X6587 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6588 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6590 VSS a_6545_47178# a_6575_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6592 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6593 a_19551_46910# a_19466_46812# a_19333_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6594 a_6945_45028# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6596 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6597 a_18280_46660# a_12549_44172# a_17609_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X6598 VSS a_18285_46348# a_18243_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X6599 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6600 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6601 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6602 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6603 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6604 a_20708_46348# a_20916_46384# a_20850_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6605 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6606 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6607 a_5167_46660# a_4651_46660# a_5072_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6608 VDD a_n1352_44484# a_n1177_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6609 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6610 a_15685_45394# a_15415_45028# a_15595_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X6611 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6613 VDD a_10193_42453# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6614 a_21350_45938# a_20273_45572# a_21188_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6617 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6618 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6619 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6620 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6621 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6622 a_7765_42852# a_7227_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6623 VSS a_526_44458# a_10149_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6624 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6625 a_7639_45394# a_n1151_42308# a_7276_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6627 a_501_45348# a_413_45260# a_375_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6628 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6629 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6630 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6631 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6632 a_16547_43609# a_16414_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X6633 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6635 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6636 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6637 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6638 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6639 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6640 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6641 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6642 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6643 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6644 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6646 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6647 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6648 a_13857_44734# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6649 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6650 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6651 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6652 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6653 a_n2661_46098# a_2107_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6654 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6655 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6656 VSS a_16327_47482# a_18953_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6657 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6659 VSS a_742_44458# a_1568_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6660 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6661 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6662 a_19273_43230# a_18083_42858# a_19164_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6663 a_6123_31319# a_7227_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6664 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6665 a_12293_43646# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6666 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6667 VDD a_2711_45572# a_4099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6668 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6669 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6670 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6671 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6672 C8_N_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6673 a_10306_45572# a_10193_42453# a_10216_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X6674 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6675 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6676 a_8035_47026# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6677 a_18545_45144# a_13259_45724# a_18450_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X6678 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6679 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6680 VDD a_21855_43396# a_13678_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6681 a_16977_43638# a_16759_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6682 a_n1423_46090# a_n1641_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6683 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6684 VDD a_22223_43948# a_14401_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6685 VDD a_6540_46812# a_6491_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6686 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6688 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6689 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6690 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6691 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6692 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6693 VDD a_n863_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6694 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6695 a_n2946_37690# a_n2956_37592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6696 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6697 C10_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X6698 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6699 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6700 a_5111_42852# a_4905_42826# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6701 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6702 VDD a_5263_45724# a_5204_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X6703 a_n467_45028# a_n745_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X6704 VDD a_15095_43370# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X6705 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X6706 VSS a_765_45546# a_1208_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6707 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6708 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X6709 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6710 VDD a_2957_45546# a_2905_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6711 a_8855_44734# a_4791_45118# a_8783_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6712 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6713 a_11963_45334# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X6714 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6715 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6716 a_n2661_44458# a_11453_44696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X6717 VDD a_4915_47217# a_11415_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6718 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6719 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6720 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6721 a_3600_43914# a_3537_45260# a_3820_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6722 a_n1741_47186# a_12005_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6723 a_1848_45724# a_2063_45854# a_1990_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6724 a_21588_30879# a_22223_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6725 a_14537_46482# a_14493_46090# a_14371_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6726 a_16241_44734# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X6727 a_3905_42865# a_5257_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6729 a_10425_46660# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X6730 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6731 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6732 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6733 a_19365_45572# a_18175_45572# a_19256_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6734 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6735 a_21811_47423# SINGLE_ENDED VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6736 VDD a_22959_45572# a_20447_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6737 a_3090_45724# a_18911_45144# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6738 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6739 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6740 a_13777_45326# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6741 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6742 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6743 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6744 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6745 VCM a_5934_30871# C5_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6746 a_n3690_39616# a_n3674_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6747 a_17333_42852# a_16795_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6748 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6749 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6750 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6751 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6752 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6753 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6754 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6755 a_11525_45546# a_11962_45724# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X6756 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6757 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6758 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6759 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6760 a_17595_43084# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X6761 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6762 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6763 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6764 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6766 a_n13_43084# a_n755_45592# a_133_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X6767 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6768 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6769 a_n1838_35608# a_n1386_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6770 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6771 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6772 a_n2840_42282# a_n2661_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6774 a_20193_45348# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6775 a_1756_43548# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6776 a_20719_46660# a_20273_46660# a_20623_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6777 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6778 a_n2302_39072# a_n2312_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6779 VSS a_n1613_43370# a_n1379_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6780 a_n2472_43914# a_n2293_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6781 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6782 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6783 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6784 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6785 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6786 a_14456_42282# a_14635_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6787 VSS a_2711_45572# a_4099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6788 VDD a_20075_46420# a_20062_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6789 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6790 a_4927_45028# a_5147_45002# a_5105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6791 a_21381_43940# a_21115_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6792 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6793 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6794 VSS a_10227_46804# a_10185_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X6795 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6796 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6798 a_4169_42308# a_1823_45246# a_3823_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6799 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6800 a_n3607_38528# a_n3674_38680# a_n3690_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6801 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6802 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6803 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6804 a_4704_46090# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6805 VDD a_20894_47436# a_20843_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6806 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X6807 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6808 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6809 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6810 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6811 VSS a_n913_45002# a_6761_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6812 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6813 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6814 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6815 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6816 VDD a_12465_44636# a_22223_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6817 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6818 VDD a_20193_45348# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6819 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6820 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6821 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6822 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6823 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6824 VDD a_5257_43370# a_3357_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6825 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6826 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X6827 VSS a_14113_42308# a_16522_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X6828 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6829 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6830 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6831 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6832 a_13460_43230# a_12379_42858# a_13113_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6834 a_19240_46482# a_19123_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6835 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6836 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6837 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6838 a_22609_37990# a_22521_39511# CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6839 a_5829_43940# a_5495_43940# a_5745_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6840 VSS C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6841 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6843 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6844 VSS a_21487_43396# a_13467_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6845 a_10227_46804# a_14955_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6846 VDD a_7287_43370# a_7274_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6847 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6848 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6850 a_14955_43940# a_14537_43396# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6852 VDD a_12861_44030# a_18911_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X6853 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6854 a_15953_42852# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6855 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6856 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6857 a_9114_42852# a_8037_42858# a_8952_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6858 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6859 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6860 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6861 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6862 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X6863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6864 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6866 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6867 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6868 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6869 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X6870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6871 VSS a_8199_44636# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X6872 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6873 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6875 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6876 VDD a_15227_44166# a_18285_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6877 a_16375_45002# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6878 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6879 a_15279_43071# a_5342_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6880 a_18780_47178# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6881 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6882 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6883 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6884 a_10193_42453# a_20712_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6885 a_5205_44484# a_5111_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6886 a_19335_46494# a_18985_46122# a_19240_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6887 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6888 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6889 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6890 VSS a_685_42968# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6891 a_4842_47243# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6892 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6893 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6894 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6895 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6896 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6897 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6898 VSS a_22591_45572# a_19963_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6899 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6900 VSS a_11322_45546# a_12016_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X6901 a_20753_42852# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X6902 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6903 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6904 a_509_45572# a_n1099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X6905 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6906 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6907 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6908 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6909 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6910 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6911 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6912 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6913 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6914 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6916 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6917 a_n1991_42858# a_n2157_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6918 a_16789_45572# a_15599_45572# a_16680_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6919 a_20362_44736# a_20640_44752# a_20596_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X6920 a_13622_42852# a_12545_42858# a_13460_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6921 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6922 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6923 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6924 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6925 a_8701_44490# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6926 a_n3607_37440# a_n3674_37592# a_n3690_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6927 VSS a_n746_45260# a_556_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6928 a_15143_45578# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6929 a_10775_45002# a_10951_45334# a_10903_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X6930 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6932 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6933 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6934 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6935 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6936 VDD a_6151_47436# a_14955_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6937 a_15673_47210# a_15507_47210# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6938 a_19120_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X6939 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6940 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6941 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6942 a_20679_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6943 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6944 VDD a_10991_42826# a_10922_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X6945 a_5815_47464# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X6946 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X6947 a_n2956_37592# a_n2472_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6948 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6949 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6950 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6951 a_13667_43396# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X6952 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6953 VSS a_n1920_47178# a_n2312_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6954 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6955 VDD a_n4064_40160# a_n2216_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X6956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6957 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6958 a_5164_46348# a_4927_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6959 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6961 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6962 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6963 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6964 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6965 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6966 a_15940_43402# a_12549_44172# a_15868_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6967 VDD a_4646_46812# a_4651_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6968 a_1427_43646# a_1049_43396# a_1209_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6969 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6970 a_19164_43230# a_18249_42858# a_18817_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6971 a_2982_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X6972 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6973 VDD a_12861_44030# a_21845_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6974 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6975 a_648_43396# a_526_44458# a_548_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X6976 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6977 VDD a_3600_43914# a_3499_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X6978 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6979 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6980 a_16409_43396# a_16243_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6981 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6982 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6983 VSS a_2063_45854# a_11136_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6985 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6986 VSS a_1823_45246# a_2202_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6987 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6988 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6989 VDD a_n3420_39616# a_n2860_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X6990 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6991 a_10903_45394# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X6992 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6993 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6995 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6996 VSS a_n971_45724# a_3775_45552# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6997 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6998 a_18243_46436# a_18189_46348# a_18147_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X6999 a_4700_47436# a_4915_47217# a_4842_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7000 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7001 VDD a_6453_43914# a_n2661_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7002 VSS a_n2438_43548# a_n2433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7003 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7004 VDD a_10053_45546# a_9625_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X7005 VDD a_12861_44030# a_19615_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7006 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7007 VDD a_13113_42826# a_13003_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7008 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7009 VDD a_380_45546# a_n356_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7010 a_11813_46116# a_11387_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X7011 a_2253_43940# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X7012 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7013 a_765_45546# a_17609_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7014 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7015 a_3503_45724# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X7016 VDD a_9625_46129# a_10037_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X7017 VDD a_3699_46348# a_3160_47472# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7018 a_18997_42308# a_18727_42674# a_18907_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7019 a_5755_42852# a_n97_42460# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7020 VDD a_22223_45036# a_18114_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7021 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7023 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7024 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X7025 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7026 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7027 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7028 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7029 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7030 a_12281_43396# a_n913_45002# a_12293_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7031 VDD a_10533_42308# a_10723_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7032 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7033 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7034 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7035 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7036 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7037 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7038 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7039 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7040 VSS a_9863_47436# a_9804_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7041 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7042 VDD a_8791_42308# a_5934_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7043 a_11387_46482# a_11133_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X7044 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7045 VDD a_21005_45260# a_19778_44110# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X7046 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7047 a_8049_45260# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7048 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7049 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7051 VSS a_n3420_38528# a_n2946_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X7052 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7053 VDD a_4646_46812# a_7871_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7054 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7055 a_895_43940# a_644_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7056 C3_P_btm a_n4064_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7057 a_19256_45572# a_18341_45572# a_18909_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7058 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7059 VSS a_2713_42308# a_2903_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7060 a_3067_47026# a_2443_46660# a_2959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7061 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7062 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7063 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7064 a_9863_47436# a_2063_45854# a_10037_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7065 a_15037_45618# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7066 a_10991_42826# a_10796_42968# a_11301_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X7067 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7068 a_3726_37500# CAL_P a_11206_38545# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X7069 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7070 a_2127_44172# a_1307_43914# a_2253_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X7071 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7072 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7073 a_1823_45246# a_4704_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7074 VDD a_n2438_43548# a_n2433_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7075 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7076 a_17678_43396# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7077 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7078 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7079 a_3080_42308# a_2903_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7080 VDD a_10903_43370# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X7081 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7082 a_n452_47436# a_n237_47217# a_n310_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7083 a_18057_42282# a_n1059_45260# a_18310_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7084 VSS a_n452_45724# a_n1853_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X7085 a_n3674_39768# a_n2472_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7087 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7088 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7089 a_8846_46660# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7090 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7091 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7092 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7093 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7094 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7095 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7096 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X7097 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7098 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7099 a_22365_46825# EN_OFFSET_CAL VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7100 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7101 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7102 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7103 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7104 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7105 a_n2472_42282# a_n2293_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7106 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7107 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7108 a_n89_45572# a_n743_46660# a_n452_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7109 VSS a_n2840_45002# a_n2810_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7110 a_15928_47570# a_15811_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7111 a_518_46482# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7112 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7113 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7114 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7115 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X7116 a_15463_44811# a_11691_44458# a_15004_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7117 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7118 a_20556_43646# a_19692_46634# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7119 VSS a_17767_44458# a_17715_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X7120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7121 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7122 a_9061_43230# a_7871_42858# a_8952_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7123 a_14309_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7124 a_16237_45028# a_16375_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7125 a_8791_43396# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7126 VDD a_n4209_38216# a_n4334_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7127 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7128 VDD a_n1423_42826# a_n1533_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7129 a_1568_43370# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7130 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7131 a_22780_39857# a_22465_38105# a_22521_39511# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7132 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7133 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7134 a_13575_42558# a_n97_42460# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7135 a_6667_45809# a_6511_45714# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X7136 a_3754_39964# a_7754_39964# VSS sky130_fd_pr__res_high_po_0p35 l=18
X7137 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7138 a_16115_45572# a_15765_45572# a_16020_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7139 VDD a_18911_45144# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7140 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7141 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7142 VSS a_9290_44172# a_10586_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7143 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7144 VDD a_3499_42826# a_n2293_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7145 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7146 a_2725_42558# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7147 a_18504_43218# a_17333_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7148 a_2253_43940# a_2479_44172# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7149 a_16979_44734# a_14539_43914# a_17061_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7150 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7151 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7153 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7155 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7156 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7158 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7159 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7161 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7162 VSS a_1307_43914# a_3681_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X7163 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7164 VSS a_626_44172# a_648_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X7165 VSS a_n3420_37440# a_n2946_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X7166 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X7167 a_21356_42826# a_21381_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7168 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7169 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7170 a_n310_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X7171 a_5025_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7172 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7173 a_16877_43172# a_16823_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7174 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7175 a_20841_46902# a_20623_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7176 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7177 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7178 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7179 VSS a_6171_45002# a_6125_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7181 VSS a_17595_43084# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X7182 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7183 a_5883_43914# a_8333_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X7184 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7185 a_21137_46414# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7186 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7188 a_20766_44850# a_20640_44752# a_20362_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X7189 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7190 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7191 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7192 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7193 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7194 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7195 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7196 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7197 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7198 a_805_46414# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7199 a_1176_45822# a_997_45618# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X7200 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7201 VDAC_N C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7202 a_21887_42336# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7203 VSS a_11967_42832# a_18083_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7204 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7205 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7206 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7207 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7208 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7209 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7211 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7212 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7213 VDD a_1823_45246# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7214 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7215 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7216 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7217 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7218 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7219 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7220 a_21513_45002# a_21363_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7221 a_8704_45028# a_5937_45572# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X7222 a_3232_43370# a_1823_45246# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7223 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7225 a_22780_40081# en_comp a_22521_40055# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7226 a_13333_42558# a_13291_42460# a_13249_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7227 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7228 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7229 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7230 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7231 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7232 a_13661_43548# a_18780_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7233 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7234 VSS a_n2840_43914# a_n4318_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7235 a_15037_44260# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7236 a_5497_46414# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7237 a_12749_45572# a_12549_44172# a_12649_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X7238 VSS a_22223_45572# a_19479_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7239 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X7240 VDD a_n2438_43548# a_n133_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7241 VDD a_14815_43914# a_n2293_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7242 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7243 VDD a_n984_44318# a_n809_44244# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7244 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7245 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7246 VDD a_22521_39511# a_22469_39537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7247 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7248 a_11530_34132# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7249 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7250 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7251 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7252 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7253 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7254 a_8128_46384# a_7903_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7255 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7256 VDD a_7281_43914# a_7229_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7257 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7258 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7259 VDD a_13507_46334# a_18907_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7260 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7261 VDD a_13904_45546# a_12594_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7262 a_479_46660# a_33_46660# a_383_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7263 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7264 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7266 VSS a_6667_45809# a_6598_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7267 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7268 a_8568_45546# a_8953_45546# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7269 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7270 VREF a_19479_31679# C1_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X7271 VDD a_n881_46662# a_n1021_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7272 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7273 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7275 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7276 a_17767_44458# a_17970_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X7277 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7278 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7280 VSS a_22400_42852# a_22780_40945# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7281 VDD a_n755_45592# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X7282 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7283 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7284 a_10867_43940# a_7499_43078# a_10405_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X7285 VDD a_10723_42308# a_5742_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7286 a_16241_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7287 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7288 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7289 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7290 a_20556_43646# a_20974_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7291 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7292 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7293 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7294 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7295 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X7296 a_4574_45260# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X7297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7299 a_13483_43940# a_13249_42308# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7300 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7301 VDD a_20159_44458# a_19321_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X7302 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7303 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7304 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7305 a_2583_47243# a_584_46384# a_2124_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7306 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7307 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7308 a_22612_30879# a_22959_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7309 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7310 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7311 VDD a_8349_46414# a_8379_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7312 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7313 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7314 a_n2216_40160# a_n2312_40392# a_n2302_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X7315 VSS a_14456_42282# a_5342_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7316 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7317 VSS a_768_44030# a_2711_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7318 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7319 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7321 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7322 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7323 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7324 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7325 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7326 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7327 a_5093_45028# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7328 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7329 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7330 a_11608_46482# a_n1151_42308# a_11387_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7331 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7332 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7333 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7334 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7335 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7336 VDD a_15227_44166# a_15597_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7337 a_19862_44208# a_13747_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7338 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7339 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7340 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7342 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7343 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7344 a_19335_46494# a_18819_46122# a_19240_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7345 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7346 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7347 VSS a_1736_39587# a_1239_39587# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7348 a_n4318_38216# a_n2472_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7349 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7350 a_8953_45546# a_8685_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7351 a_18249_42858# a_18083_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7352 a_12816_46660# a_11735_46660# a_12469_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7353 a_19268_43646# a_13661_43548# a_19177_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X7354 a_20256_42852# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X7355 a_13258_32519# a_19647_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7356 VDD a_16680_45572# a_16855_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7357 VSS a_n447_43370# a_n2129_43609# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7358 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7359 a_20528_45572# a_19466_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7360 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7361 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7362 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7363 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7364 a_11525_45546# a_10586_45546# a_11778_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7365 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7366 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7367 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7368 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7369 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7370 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7371 VDD a_2711_45572# a_20107_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7372 a_16147_45260# a_17478_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7373 a_n2109_45247# a_n2017_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7374 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7375 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7376 a_19963_31679# a_22591_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7377 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7378 a_19610_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7379 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7380 a_5837_43172# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7381 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7382 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7383 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7384 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7385 a_n143_45144# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7386 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7387 a_n310_45572# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7388 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7389 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7390 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7391 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7392 VDD a_22959_47212# a_22612_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7393 a_15015_46420# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7394 a_20596_44850# a_20159_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7395 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7396 VSS a_7227_45028# a_7230_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7397 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7398 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7399 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7400 a_2957_45546# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X7401 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7402 VSS a_14579_43548# a_14537_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7403 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7404 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7405 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X7406 VSS a_5111_44636# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7407 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7408 VDD a_11599_46634# a_15507_47210# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7409 VDD a_6151_47436# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X7410 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7411 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7412 VDD COMP_P a_n1329_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7413 VDD a_20679_44626# a_20640_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7415 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7417 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7418 VSS a_19321_45002# a_20567_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7419 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7420 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7421 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7422 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7423 VSS a_n2472_45002# a_n2956_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7424 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7425 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7426 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7427 a_10903_43370# a_13351_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7428 a_14513_46634# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7429 a_10949_43914# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X7430 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7431 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7432 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7434 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7435 a_10149_43396# a_5111_44636# a_9803_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7436 VSS a_19431_45546# a_19365_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7437 a_13943_43396# a_11823_42460# a_13837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7438 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7440 VSS a_16922_45042# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7441 a_16112_44458# a_14539_43914# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7442 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7443 C8_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X7444 VDD a_4099_45572# a_3483_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7445 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7446 a_6197_43396# a_6031_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7447 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7448 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7449 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X7450 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7451 a_7309_42852# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7452 a_n2840_46634# a_n2661_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7453 a_380_45546# a_n357_42282# a_603_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7454 a_18533_43940# a_18326_43940# a_18451_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7455 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7456 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7457 a_5932_42308# a_5755_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7458 VDD a_n863_45724# a_2448_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7460 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7461 a_16328_43172# a_n97_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7462 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7463 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7464 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7465 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7466 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7467 a_17583_46090# a_17715_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X7468 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7469 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7470 VDD a_n755_45592# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X7471 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7472 VSS a_10991_42826# a_10922_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7473 VDD a_15433_44458# a_15463_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7474 a_n2267_43396# a_n2433_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7475 a_19615_44636# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X7476 a_5732_46660# a_4651_46660# a_5385_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7477 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X7478 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7479 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7480 a_n2840_46090# a_n2661_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7481 VDD a_5129_47502# a_5159_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7482 a_n967_45348# a_n913_45002# a_n955_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7483 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7484 a_19006_44850# a_18248_44752# a_18443_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X7485 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X7486 VDD a_18817_42826# a_18707_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7487 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7488 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7489 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7490 a_15559_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X7491 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7492 a_9803_43646# a_8953_45546# a_9885_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7493 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7494 VDD a_n2840_42282# a_n3674_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7496 VDD a_3232_43370# a_9313_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X7497 a_13460_43230# a_12545_42858# a_13113_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7498 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7499 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7500 a_20362_44736# a_20679_44626# a_20637_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X7501 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7502 a_2713_42308# a_n913_45002# a_2725_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7503 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7504 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7505 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7506 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7507 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7508 a_16241_47178# a_16023_47582# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X7509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7510 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7511 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7512 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7513 a_14955_43396# a_14205_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X7514 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7515 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7516 VSS a_n913_45002# a_10533_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7517 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7518 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7519 a_7466_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7520 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7521 VDD a_6151_47436# a_5907_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7522 a_16697_47582# a_15507_47210# a_16588_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7523 a_n2267_44484# a_n2433_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7524 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7525 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7526 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7527 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7528 a_13693_46688# a_6755_46942# a_13607_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7529 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7530 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7531 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7532 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X7533 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7534 VDD a_19778_44110# a_19741_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7535 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7536 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7538 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7539 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7540 a_2609_46660# a_2443_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7541 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7542 a_5708_44484# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X7543 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7544 VSS a_n2472_43914# a_n3674_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7545 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7546 a_18143_47464# a_18479_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X7547 a_5263_46660# a_4817_46660# a_5167_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7548 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7549 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7550 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7551 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7552 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7553 a_12016_45572# a_11962_45724# a_11525_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X7554 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7556 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7557 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7558 VSS a_18057_42282# a_n356_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X7559 VDD a_21671_42860# a_3422_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7560 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7561 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7562 VDD a_8746_45002# a_8704_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7563 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7564 a_3411_47243# a_3160_47472# a_2952_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7565 a_n2840_46634# a_n2661_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7566 VSS a_7705_45326# a_7639_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7567 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7568 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7569 a_133_43172# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X7570 VDD a_9396_43370# a_5111_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7571 VSS a_167_45260# a_1423_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7572 a_743_42282# a_13661_43548# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7575 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7576 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7577 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7578 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7579 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7580 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7581 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7582 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7583 VDD a_20512_43084# a_19987_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X7584 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7585 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7586 a_1891_43646# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X7587 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7588 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7589 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7590 VSS a_n357_42282# a_17141_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7591 a_n4318_39304# a_n2840_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7593 VIN_P EN_VIN_BSTR_P C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7594 a_14485_44260# a_5807_45002# a_12465_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7596 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7597 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7598 VSS a_n1059_45260# a_8945_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7599 a_11453_44696# a_17719_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X7600 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7601 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7602 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7603 a_10545_42558# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7605 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7606 a_17701_42308# a_17531_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7607 a_8292_43218# a_7765_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7608 a_13657_42558# a_11823_42460# a_13575_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7609 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7610 a_16751_46987# a_5807_45002# a_16292_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7611 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7612 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7613 a_10586_45546# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7614 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7615 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7617 VDD a_3537_45260# a_4223_44672# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7619 VSS a_16855_45546# a_16789_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7620 a_3626_43646# a_1414_42308# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7621 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7622 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7623 a_45_45144# a_n143_45144# a_n37_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7624 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7625 VDD a_20107_42308# a_7174_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7626 a_3815_47204# a_3785_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7627 a_15567_42826# a_15743_43084# a_15953_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7628 VSS a_10341_42308# a_11554_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7629 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7630 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7631 VCM a_5342_30871# C8_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7632 a_n83_35174# VDD EN_VIN_BSTR_P VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X7633 a_6755_46942# a_15015_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7634 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7635 VSS a_4791_45118# a_6640_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X7636 a_2437_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7637 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7638 VDAC_Pi a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X7639 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7640 a_9823_46155# a_9804_47204# a_9823_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7641 a_1990_45899# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X7642 a_15743_43084# a_19339_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X7643 VDD a_5385_46902# a_5275_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7644 a_5129_47502# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7646 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7647 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7648 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7649 VDAC_P C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7650 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7651 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7652 a_9145_43396# a_8791_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7653 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7654 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7655 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7656 VIN_P EN_VIN_BSTR_P C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7657 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7658 VDD a_20841_46902# a_20731_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7659 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7660 a_7276_45260# a_n1151_42308# a_7418_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7661 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7662 VDD a_n785_47204# a_327_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7663 a_8103_44636# a_8375_44464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7664 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7665 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7666 a_4915_47217# a_12991_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X7667 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7670 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7671 VDD a_8199_44636# a_8855_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7672 VDD a_12549_44172# a_21115_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7673 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7674 VDD a_2553_47502# a_2583_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7675 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7676 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7677 a_n327_42558# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X7678 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7679 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7680 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7681 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7682 a_19864_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X7683 a_12800_43218# a_12089_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7684 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7686 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7688 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7689 VSS a_20623_43914# a_20365_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X7690 VSS a_n743_46660# a_16501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X7691 VSS a_22959_45036# a_19721_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7692 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7693 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7694 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7695 a_n4318_38680# a_n2472_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7696 VSS a_11967_42832# a_16243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7697 a_7754_40130# RST_Z VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7698 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7699 a_13483_43940# a_13249_42308# a_13565_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7700 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7701 a_3363_44484# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7702 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7703 a_13249_42558# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7704 a_18504_43218# a_17333_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7705 VDD a_4235_43370# a_n2661_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7706 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7707 a_n39_42308# a_n97_42460# a_n473_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7708 a_10210_45822# a_10180_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X7709 VSS a_11967_42832# a_20512_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7710 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7711 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7712 VSS a_n443_46116# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7713 VSS a_4646_46812# a_7411_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7714 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7715 a_20273_46660# a_20107_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7716 VDD a_11341_43940# a_22223_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7717 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X7718 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7719 a_n2312_38680# a_n2104_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7720 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7721 VDD a_12791_45546# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X7722 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7723 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7724 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7725 a_19237_31679# a_22959_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7726 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7727 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7729 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7730 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7732 VDD a_19328_44172# a_19279_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X7733 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7734 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7735 VDD SMPL_ON_P a_n1605_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7737 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7738 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7739 VSS a_11967_42832# a_12379_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7740 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7741 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7742 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7743 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7744 VDD a_18315_45260# a_18189_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X7745 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7746 VSS a_15227_44166# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7747 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7748 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7749 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7750 a_10951_45334# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7751 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7752 VDD a_2123_42473# a_1184_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7753 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7754 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7755 a_4791_45118# a_4743_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7756 a_21195_42852# a_20922_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X7757 a_4156_43218# a_3905_42865# a_3935_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7758 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7759 a_15227_44166# a_22000_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7760 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7761 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7762 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7763 a_n1899_43946# a_n2065_43946# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7764 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7765 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7766 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7767 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7768 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7769 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7770 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7771 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7772 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7773 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7774 a_n743_46660# a_n1021_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7775 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7776 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7777 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7778 a_n2293_45546# a_2274_45254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7779 a_11633_42308# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7780 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7781 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7782 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7783 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7784 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7785 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7786 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7787 a_20205_31679# a_22223_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7788 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7789 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X7790 a_n2472_46634# a_n2293_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7791 a_2698_46116# a_2521_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7792 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7793 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7794 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7795 VDD a_10193_42453# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7796 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7797 a_22705_37990# a_22521_40055# a_22609_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7798 VDD a_n3565_38502# a_n3690_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7799 a_5342_30871# a_14456_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7800 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7801 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7802 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7803 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7804 VDD a_8325_42308# a_8791_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7805 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7806 a_548_43396# a_n863_45724# a_458_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X7807 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7808 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7809 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7810 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7811 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X7812 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7813 VSS a_1756_43548# a_1467_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X7814 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7815 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7816 VDD a_17517_44484# a_22591_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7817 VSS a_n913_45002# a_19511_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7818 a_288_46660# a_171_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7819 a_15312_46660# a_14976_45028# a_15009_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7820 a_n2472_46090# a_n2293_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7821 VSS a_22959_43948# a_17538_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7822 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7823 C9_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X7824 a_20894_47436# a_20990_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7825 VDD a_n2438_43548# a_n2157_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7826 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7827 VDD a_n4064_38528# a_n2216_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X7828 a_8037_42858# a_7871_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7829 a_n1736_43218# a_n1853_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7830 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7831 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7832 a_13527_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7834 VDD a_n2472_42282# a_n4318_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7835 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7836 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7837 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7839 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7840 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7841 a_n2661_43370# a_11415_45002# a_11361_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7842 VDD a_n2840_42826# a_n3674_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7843 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7844 VSS a_1343_38525# a_2113_38308# VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X7845 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7846 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7847 VDD a_22165_42308# a_22223_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7848 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7850 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7851 VSS a_14180_45002# a_13017_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X7852 a_15681_43442# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7854 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7855 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7856 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7857 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7858 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7859 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7860 a_8488_45348# a_8199_44636# a_8191_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X7861 a_16588_47582# a_15673_47210# a_16241_47178# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7862 a_18220_42308# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7863 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7864 a_n1423_46090# a_n1641_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7866 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X7867 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7868 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7869 a_17609_46634# a_12549_44172# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7871 a_16115_45572# a_15599_45572# a_16020_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7873 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7874 VSS a_19700_43370# a_n97_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7875 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7876 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7877 VSS a_2124_47436# a_1209_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X7878 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7879 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7880 VDD a_6755_46942# a_12741_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7881 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7882 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7883 VSS a_19615_44636# a_18579_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7884 a_15595_45028# a_15415_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7885 a_12545_42858# a_12379_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7886 a_8791_45572# a_7499_43078# a_8697_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7887 a_16942_47570# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7888 a_14853_42852# a_n913_45002# a_14635_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7890 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7891 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7892 VSS a_4958_30871# a_17531_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7893 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7894 a_8333_44056# a_4223_44672# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7895 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7896 a_6511_45714# a_4646_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7897 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7898 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7899 VDD a_10949_43914# a_10867_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X7900 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7901 a_17973_43940# a_17737_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7902 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7903 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7904 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7905 a_18494_42460# a_18907_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X7906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7907 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7908 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7909 a_17061_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7910 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7911 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7913 a_n2472_46634# a_n2293_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7914 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7915 C2_P_btm a_3080_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7916 VSS a_5267_42460# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X7917 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7918 VSS a_n2438_43548# a_n2065_43946# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7919 VDD a_7754_40130# a_3754_38470# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7920 VDD a_n357_42282# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7921 a_9159_45572# a_5937_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7923 a_3483_46348# a_4099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7924 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7925 VDD a_n3565_37414# a_n3690_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7926 a_8238_44734# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X7927 VSS a_17517_44484# a_22591_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7929 VSS a_21613_42308# a_22775_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X7930 VDD a_3381_47502# a_3411_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7931 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7933 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7934 a_10150_46912# a_10467_46802# a_10425_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X7935 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7936 a_n2810_45572# a_n2840_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7937 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7938 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7939 a_13675_47204# a_n1435_47204# a_13569_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X7940 a_22165_42308# a_21887_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X7941 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7942 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7943 VDD a_n4064_37440# a_n2216_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X7944 VSS a_11827_44484# a_22223_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7945 a_5518_44484# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X7946 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7947 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7948 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7949 VDD a_22521_40055# a_22459_39145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7950 a_13678_32519# a_21855_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7951 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7952 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7953 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7954 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7955 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7956 VDD a_8605_42826# a_8495_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7957 a_n2312_40392# a_n2288_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7958 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7959 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7960 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7961 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7962 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7963 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7964 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7965 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7966 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7967 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7968 VDD a_20193_45348# a_21887_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7969 a_13076_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X7970 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X7971 a_18691_45572# a_18341_45572# a_18596_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7972 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X7973 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7974 a_3600_43914# a_1307_43914# a_3992_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X7975 a_4743_43172# a_3537_45260# a_4649_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7976 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7977 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7978 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7979 a_11387_46155# a_11309_47204# a_11387_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7980 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7981 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7982 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7983 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7985 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7986 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7987 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7989 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7990 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7991 a_22609_37990# a_22469_39537# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X7992 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7993 a_11554_42852# a_10835_43094# a_10991_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X7994 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7995 VSS a_9313_44734# a_22959_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7996 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7997 VDD a_2680_45002# a_2274_45254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7998 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7999 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8000 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8001 VSS C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8002 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8003 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8004 VDD a_n1177_43370# a_n1190_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8005 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8006 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X8007 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8009 VDD a_6755_46942# a_13556_45296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8010 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8011 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8012 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8013 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8014 VDD a_n971_45724# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X8015 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8016 a_n785_47204# a_n815_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8017 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8018 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8019 a_n4251_40480# a_n4318_40392# a_n4334_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8020 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8021 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8022 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8023 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8024 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8025 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8026 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X8027 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8028 a_19900_46494# a_18819_46122# a_19553_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8029 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8030 VSS a_n1386_35608# a_n1838_35608# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8031 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8032 a_12561_45572# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X8033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8034 a_10083_42826# a_10518_42984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X8035 a_12359_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8036 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8037 VSS a_10355_46116# a_8199_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8038 a_3422_30871# a_21671_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8039 a_5937_45572# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8040 VDD a_16327_47482# a_17767_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8041 a_21005_45260# a_21101_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X8042 a_12649_45572# a_10903_43370# a_12561_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X8043 VSS a_19321_45002# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8044 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8045 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8046 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8047 a_5111_44636# a_9396_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8048 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8049 a_21297_45572# a_20107_45572# a_21188_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X8050 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8051 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8052 a_12469_46902# a_12251_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8053 a_376_46348# a_584_46384# a_518_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8054 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8056 a_15146_44484# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8057 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8058 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8059 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8060 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8061 VIN_P EN_VIN_BSTR_P C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X8062 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8063 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8064 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8065 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8066 VDD a_n971_45724# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X8067 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X8068 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8069 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8070 a_14180_45002# a_14537_43396# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8071 VDD a_10193_42453# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X8072 a_18681_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X8073 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8074 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8075 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8076 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8077 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8078 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8079 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8080 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8081 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8082 a_17829_46910# a_12549_44172# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X8083 VSS a_15009_46634# a_14180_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X8084 a_2304_45348# a_2274_45254# a_2232_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X8085 a_6598_45938# a_6511_45714# a_6194_45824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X8086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8087 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8088 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8089 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8090 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8091 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8092 a_5745_43940# a_5013_44260# a_5663_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8093 VDD a_10193_42453# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8094 a_5742_30871# a_10723_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8095 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8096 a_19478_44056# a_3090_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X8097 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8098 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8099 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8100 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8101 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8104 a_8192_45572# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X8105 a_10185_46660# a_10150_46912# a_9863_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8106 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8107 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8108 a_10835_43094# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8109 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8110 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8111 a_15890_42674# a_15764_42576# a_15486_42560# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X8112 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8113 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8114 a_n699_43396# a_n1177_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X8115 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8116 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8118 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8119 a_14033_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X8120 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8121 a_6101_44260# a_1307_43914# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8122 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8123 a_7927_46660# a_7577_46660# a_7832_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8124 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8125 a_16721_46634# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8126 a_5826_44734# a_5147_45002# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X8127 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8128 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8129 a_21496_47436# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X8130 VDD a_16763_47508# a_16750_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8131 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8132 VDD a_n746_45260# a_175_44278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8133 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8134 a_2813_43396# a_3232_43370# a_2982_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8135 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8136 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8137 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8138 a_6171_42473# a_5932_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8139 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8140 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8141 VDD a_601_46902# a_491_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8142 VSS a_4646_46812# a_6031_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8143 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8144 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8145 VSS a_13059_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X8146 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8147 VDD a_1123_46634# a_1110_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8148 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8149 a_8292_43218# a_7765_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8150 a_11787_45002# a_11963_45334# a_11915_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X8151 VSS a_584_46384# a_2998_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8152 VDD a_n2472_42826# a_n4318_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8153 a_1667_45002# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X8154 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8155 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8156 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8158 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8159 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8160 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8162 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8163 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8164 a_20731_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8165 a_8062_46482# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8166 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8167 a_n2216_38778# a_n2312_38680# a_n2302_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8168 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8169 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8171 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8172 a_13925_46122# a_13759_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8173 VSS a_11599_46634# a_20107_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8174 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8175 a_5385_46902# a_5167_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8176 VDD a_7499_43078# a_10729_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X8177 a_9803_43646# a_8953_45546# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8178 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8179 VSS a_n2104_46634# a_n2312_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8180 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8181 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8182 a_n1177_44458# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8184 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8185 VDD a_5111_44636# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X8186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8187 VDD a_19256_45572# a_19431_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8188 VDD a_6761_42308# a_7227_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X8189 a_7911_44260# a_7845_44172# a_7542_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X8190 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8191 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8192 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8193 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8194 VDD a_19553_46090# a_19443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8195 a_5205_44484# a_5343_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8196 a_22400_42852# a_22223_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8197 a_12603_44260# a_12549_44172# a_12495_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X8198 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8199 VSS a_18194_35068# a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X8200 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8201 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8202 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8203 a_3638_45822# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X8204 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8205 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8206 a_17324_43396# a_16243_43396# a_16977_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8207 a_5275_47026# a_4651_46660# a_5167_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8208 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8209 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8210 a_19452_47524# a_19386_47436# a_13747_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8211 a_11915_45394# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X8212 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8213 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8214 a_14447_46660# a_n1151_42308# a_14084_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8215 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8216 a_12800_43218# a_12089_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8217 VSS a_n1613_43370# a_n1655_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8218 a_20731_47026# a_20107_46660# a_20623_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8219 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8220 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8221 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8222 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8223 VSS a_20712_42282# a_10193_42453# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8224 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8225 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8226 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8227 VSS a_n443_42852# a_421_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8228 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8229 a_15720_42674# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8230 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8231 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8233 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8234 VDD a_11599_46634# a_15599_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8235 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8236 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8237 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8238 a_n659_45366# a_n746_45260# a_n745_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8239 a_14493_46090# a_14275_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8240 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8241 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8242 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8243 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8244 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X8245 a_n881_46662# a_14495_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8246 a_8685_43396# a_8147_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X8247 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8248 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8249 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8250 C7_P_btm a_n4209_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8252 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8253 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8254 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8255 a_11554_42852# a_10796_42968# a_10991_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X8256 a_765_45546# a_17609_46634# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8257 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X8258 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8259 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8260 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8261 VDD a_15803_42450# a_15764_42576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8262 a_2063_45854# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8263 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8265 a_19386_47436# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X8266 a_8492_46660# a_7411_46660# a_8145_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8267 a_1337_46436# a_1176_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X8268 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8269 VSS a_4419_46090# a_4365_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8270 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8271 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8272 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8273 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8275 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8276 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8277 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8278 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8279 VSS a_6575_47204# a_9067_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X8280 a_n1331_43914# a_n1549_44318# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8281 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8282 VDD a_3537_45260# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8283 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8284 a_20835_44721# a_20640_44752# a_21145_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X8285 VSS a_11189_46129# a_11608_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X8286 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8287 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8288 a_n327_42558# a_n97_42460# a_n473_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X8289 a_8147_43396# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X8290 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8291 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8292 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8293 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8294 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8295 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8296 a_8685_42308# a_8515_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8297 VDD a_17324_43396# a_17499_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8298 a_19431_46494# a_18985_46122# a_19335_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X8299 VDD a_12607_44458# a_n2661_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8300 a_1414_42308# a_1067_42314# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X8301 VDD a_10193_42453# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8302 VDD a_21356_42826# a_n357_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8303 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8304 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8305 a_n2216_37690# a_n2810_45028# a_n2302_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8306 VDD a_4883_46098# a_10355_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8307 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8308 a_16977_43638# a_16759_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8309 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8310 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8312 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8313 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8314 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8315 a_1049_43396# a_458_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8316 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8317 VDD a_n443_42852# a_742_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8318 a_10555_43940# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8319 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8320 VSS a_n237_47217# a_8270_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8321 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8322 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8323 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8324 a_21613_42308# a_21335_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X8325 a_8145_46902# a_7927_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8326 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8327 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8328 VSS a_16019_45002# a_15903_45785# VSS sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X8329 VCM a_5342_30871# C8_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8330 VDD a_n23_45546# a_7_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8331 VDD a_2698_46116# a_2804_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8332 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8333 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8334 a_20935_43940# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8335 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8336 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8337 a_2713_42308# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8338 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8339 VSS C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8340 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8341 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8342 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8343 VDD a_n699_43396# a_4743_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8344 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8345 a_17591_47464# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X8346 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8347 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8348 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8349 a_9223_42460# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8350 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8351 a_12741_44636# a_14537_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8352 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8353 VDD a_20202_43084# a_21335_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8354 a_564_42282# a_743_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8355 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8356 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8357 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8358 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8359 a_2684_37794# a_1736_39587# a_1736_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8360 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8361 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8362 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8363 a_15367_44484# a_13556_45296# a_15004_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8364 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8365 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8366 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8367 VSS a_n452_47436# a_n815_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8368 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8369 VDD a_2063_45854# a_9863_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8370 VSS a_6511_45714# a_6472_45840# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8371 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8372 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8373 a_9223_42460# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X8374 VSS a_19987_42826# a_n2017_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X8375 VSS a_13159_45002# a_13105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8376 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8377 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8378 a_2981_46116# a_2804_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8379 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8380 a_21188_45572# a_20273_45572# a_20841_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8381 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8382 a_20692_30879# a_22959_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8383 a_9028_43914# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X8384 VDD a_17715_44484# a_17737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8385 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8386 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8388 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8389 VSS a_n2840_44458# a_n4318_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8390 VSS a_15004_44636# a_14815_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8391 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8392 a_16759_43396# a_16243_43396# a_16664_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8393 a_4574_45260# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8394 a_17829_46910# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X8395 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8396 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8397 VSS a_n443_46116# a_4880_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X8398 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8400 VDD a_1799_45572# a_1983_46706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X8401 VDD a_21363_45546# a_21350_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8402 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8403 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X8404 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8405 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8406 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8407 a_13259_45724# a_17583_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8408 C1_P_btm a_n4064_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X8409 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8410 VIN_P EN_VIN_BSTR_P C4_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X8411 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8412 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8413 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8414 VSS a_327_44734# a_501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8415 a_6575_47204# a_6545_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8416 VSS a_765_45546# a_380_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X8417 a_104_43370# a_n699_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8418 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8419 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8421 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8423 a_n2293_42282# a_3357_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8424 VDD a_22959_42860# a_14097_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8425 a_3935_42891# a_2382_45260# a_3935_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8426 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8427 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8428 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8429 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8430 VSS a_6171_42473# a_5379_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8431 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8432 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8433 VDD a_n863_45724# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X8434 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8435 VDD a_8145_46902# a_8035_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8436 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8437 a_17141_43172# a_n1059_45260# a_16795_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8438 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8440 VSS a_10193_42453# a_11897_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8441 a_15433_44458# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8442 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8443 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8444 VSS a_4791_45118# a_5066_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8445 VDD a_5691_45260# a_n2109_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X8446 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8447 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8448 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8449 a_15486_42560# a_15803_42450# a_15761_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X8450 a_18753_44484# a_18374_44850# a_18681_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X8451 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8452 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8453 VDD a_1983_46706# a_n2661_46098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8454 a_15227_46910# a_15368_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8455 a_6682_46987# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8456 a_n1079_45724# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8457 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8458 a_12429_44172# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X8459 a_1568_43370# a_1847_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8460 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8462 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8463 VDD a_7227_42308# a_6123_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8464 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8465 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8466 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8467 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8468 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8469 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8470 a_8952_43230# a_8037_42858# a_8605_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8471 a_3457_43396# a_3232_43370# a_3626_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8472 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8473 a_7174_31319# a_20107_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8474 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8475 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8476 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8477 VSS a_167_45260# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8478 a_13490_45067# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8479 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8480 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8481 VSS a_6171_45002# a_11909_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8482 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8483 a_4181_44734# a_3090_45724# a_n2497_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8484 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8485 a_16388_46812# a_17957_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X8486 VDD a_3218_45724# a_3175_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8487 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8488 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8489 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8490 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8491 a_33_46660# a_n133_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8492 a_8283_46482# a_n1151_42308# a_7920_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8493 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8494 VDD a_15279_43071# a_14579_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8495 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8496 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8497 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8498 VDD a_16763_47508# a_5807_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8499 VDD a_310_45028# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8500 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8501 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8502 a_n23_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8503 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8504 a_3935_43218# a_3681_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X8505 VDD a_10903_43370# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X8506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8507 a_n1099_45572# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X8508 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8509 a_14949_46494# a_13759_46122# a_14840_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X8510 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8511 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8512 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8513 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8514 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8515 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8516 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8517 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8518 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8519 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8520 VDD a_n4315_30879# a_n4334_40480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X8521 a_6851_47204# a_6491_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8522 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8523 a_13556_45296# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8524 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8525 VSS a_15227_44166# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X8526 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8527 a_19987_42826# a_18494_42460# a_20356_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X8528 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X8529 a_n2833_47464# a_n2497_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X8530 a_3524_46660# a_2609_46660# a_3177_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8531 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8532 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8533 VSS a_6151_47436# a_6229_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X8534 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8535 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8536 VSS a_22223_47212# a_21588_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8537 a_18533_43940# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8538 a_14205_43396# a_13667_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X8539 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8540 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8541 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8542 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8543 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8544 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8545 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X8546 a_16377_45572# a_16333_45814# a_16211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X8547 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8549 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8550 a_10044_46482# a_n743_46660# a_9823_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8551 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8552 a_19113_45348# a_18911_45144# a_3090_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8553 VSS a_13720_44458# a_12607_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8554 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8556 a_n2860_37984# a_n2956_38216# a_n2946_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8557 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8558 a_5934_30871# a_8791_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8559 a_5837_43396# a_5111_44636# a_5147_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8560 a_2266_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8561 a_10861_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X8562 VSS a_7920_46348# a_7715_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8563 a_14383_46116# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8564 a_2905_42968# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8565 a_2809_45348# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X8566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8568 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8569 a_6540_46812# a_6755_46942# a_6682_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8570 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8571 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8572 a_6709_45028# a_6431_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X8573 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8576 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8577 VSS a_18494_42460# a_20193_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8578 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8579 C7_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X8580 a_n1991_42858# a_n2157_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8581 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8582 a_13249_42308# a_13070_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8583 a_n2442_46660# a_n2472_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8584 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8585 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X8586 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X8587 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8588 a_13348_45260# a_12891_46348# a_13490_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8589 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8590 a_17061_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8591 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8593 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8594 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X8595 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8596 VDD a_18443_44721# a_18374_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X8597 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8598 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8599 VDD a_n3565_39304# a_n3690_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X8600 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8601 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8602 a_1512_43396# a_n443_46116# a_1209_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X8603 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8604 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8605 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8606 VSS a_15803_42450# a_15764_42576# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8607 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8608 VDD a_22591_44484# a_17730_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8609 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8610 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8611 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8613 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X8614 a_11901_46660# a_11735_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8615 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8616 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8617 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8618 a_21076_30879# a_22959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8619 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8620 a_3877_44458# a_3699_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X8621 VDD a_n4064_39072# a_n2216_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X8622 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8623 a_11691_44458# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8625 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8626 a_2813_43396# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X8627 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8628 a_15368_46634# a_15143_45578# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X8629 VSS a_9028_43914# a_8975_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8630 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8631 C8_N_btm a_17538_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8632 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8633 a_5093_45028# a_4558_45348# a_5009_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8634 VSS a_10193_42453# a_13921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8635 a_15597_42852# a_15567_42826# a_15095_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X8636 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8637 VDD a_13059_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8638 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8639 a_3823_42558# a_3065_45002# a_3905_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8640 VDD a_526_44458# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8641 a_2553_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8642 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8643 VSS a_1667_45002# a_n863_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X8644 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8645 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8646 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8647 a_16855_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8648 a_5495_43940# a_5244_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8649 VDD a_21177_47436# a_20990_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X8650 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8651 VDD a_22365_46825# a_20202_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8652 VSS a_19787_47423# a_19594_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8653 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8654 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X8655 a_n1736_46482# a_n1853_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8656 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8657 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8659 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8660 a_5063_47570# a_4915_47217# a_4700_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8662 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8663 a_11322_45546# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8664 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8667 a_19787_47423# START VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8670 VDD a_9127_43156# a_9114_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8671 a_n4251_39616# a_n4318_39768# a_n4334_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8672 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8673 a_3754_39466# a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X8674 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X8675 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8676 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8677 a_10384_47026# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8678 VSS a_11525_45546# a_11189_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8679 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8680 a_10729_43914# a_11750_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8681 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8682 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8684 a_4921_42308# a_n913_45002# a_4933_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8686 VSS a_8568_45546# a_8162_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X8687 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8688 a_20528_46660# a_20411_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8689 VSS a_n23_47502# a_n89_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X8690 a_13657_42558# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8691 VSS a_4223_44672# a_5205_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8692 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8693 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X8694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8695 a_791_42968# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8696 a_13837_43396# a_13259_45724# a_13749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X8697 a_19177_43646# a_17339_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X8698 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8699 a_196_42282# a_375_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8700 a_18005_44484# a_17970_44736# a_17767_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8701 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8702 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8703 a_11309_47204# a_11031_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X8704 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8705 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8706 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8707 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8708 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8709 VSS a_4646_46812# a_7871_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8710 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8711 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8712 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8713 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X8714 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8715 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8716 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8717 a_18691_45572# a_18175_45572# a_18596_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8718 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8719 a_n23_45546# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X8720 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8721 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8722 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8723 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8724 a_9885_42558# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8725 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8726 VSS a_4700_47436# a_3785_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8727 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8729 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8732 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8733 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X8734 a_4361_42308# a_3823_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8735 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8737 VDD a_n2438_43548# a_n2157_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8738 VDD a_n2840_46634# a_n2956_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8739 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8740 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8741 VDD a_13635_43156# a_13622_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8742 a_4817_46660# a_4651_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8744 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8745 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8746 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8747 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8748 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8749 VSS a_1307_43914# a_4156_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X8750 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X8751 a_8415_44056# a_5343_44458# a_8333_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8752 a_n1699_44726# a_n1917_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8753 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8754 a_1525_44260# a_1467_44172# a_1115_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X8755 a_14976_45028# a_14797_45144# a_15060_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X8756 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8757 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8758 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8759 VSS a_15959_42545# a_15890_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X8760 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X8761 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8762 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8763 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X8764 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8766 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8767 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8768 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8769 VDD a_22469_40625# a_22705_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X8770 a_n2312_39304# a_n1920_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X8771 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8772 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8773 VIN_N EN_VIN_BSTR_N C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X8774 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8775 VDD a_1736_39587# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X8776 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8777 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8778 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8779 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8780 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8781 VDD a_n452_44636# a_n2129_44697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X8782 VSS a_21363_45546# a_21297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X8783 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8784 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8785 VDD a_7112_43396# a_7287_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8786 a_19443_46116# a_18819_46122# a_19335_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8787 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8788 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8789 VDD a_5111_44636# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X8790 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8791 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8792 VDD EN_VIN_BSTR_N w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8793 a_310_45028# a_n37_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X8794 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8795 a_17719_45144# a_17613_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8796 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8797 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8798 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8799 VDD a_12563_42308# a_5534_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8800 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8801 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8802 a_17499_43370# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8803 a_n357_42282# a_21356_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8804 VSS a_13747_46662# a_19466_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8805 a_14112_44734# a_768_44030# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X8806 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8807 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8808 VDD a_3483_46348# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8809 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X8810 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X8811 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8812 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X8813 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8814 a_14097_32519# a_22959_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8815 a_8270_45546# a_n237_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8816 a_3094_47570# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8817 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8818 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8819 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8820 VSS a_3232_43370# a_11541_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8821 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8822 VSS C0_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8823 a_8781_46436# a_8199_44636# a_8034_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8824 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8826 a_10533_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8827 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8828 a_20841_46902# a_20623_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8829 a_13527_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8830 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8831 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8832 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8834 a_17896_45144# a_16922_45042# a_17801_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X8835 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8836 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8837 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8838 a_18817_42826# a_18599_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8839 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8840 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8841 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8843 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8844 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8845 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8846 a_104_43370# a_n699_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X8847 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8848 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8850 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8852 a_16211_45572# a_15765_45572# a_16115_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X8853 VSS a_20835_44721# a_20766_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X8854 a_19741_43940# a_19478_44306# a_19328_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8855 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8856 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8857 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8858 VDD a_4223_44672# a_4181_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8859 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8860 VDD a_13747_46662# a_14495_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8861 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8862 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8863 a_2487_47570# a_2063_45854# a_2124_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8864 VSS a_10809_44734# a_22959_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8865 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8866 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8867 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8868 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8869 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8870 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8871 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8873 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8875 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8876 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8877 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8878 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X8879 VSS a_20567_45036# a_12549_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8880 a_18451_43940# a_18579_44172# a_18533_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8881 a_21359_45002# a_21513_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8882 a_13904_45546# a_13249_42308# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8883 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8884 VSS a_13661_43548# a_18587_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8885 a_6547_43396# a_6031_43396# a_6452_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
C0 a_13113_42826# a_12895_43230# 0.209641f
C1 a_3626_43646# a_5934_30871# 0.192998f
C2 a_9290_44172# a_10083_42826# 0.136441f
C3 a_n2661_42282# VDD 0.406474f
C4 a_3483_46348# a_9290_44172# 0.207611f
C5 a_15227_44166# a_13259_45724# 0.916975f
C6 a_16763_47508# VDD 0.392885f
C7 a_n2472_42282# a_n4318_38216# 0.157105f
C8 a_11967_42832# a_3422_30871# 0.139082f
C9 a_16823_43084# VDD 0.159922f
C10 a_6755_46942# a_13556_45296# 0.103107f
C11 a_19321_45002# a_20193_45348# 0.489018f
C12 a_5932_42308# C3_N_btm 0.121156f
C13 a_5742_30871# EN_VIN_BSTR_P 0.645417f
C14 a_12861_44030# a_n743_46660# 0.100542f
C15 a_n971_45724# a_6540_46812# 0.31827f
C16 a_18479_47436# a_19594_46812# 0.108004f
C17 a_19386_47436# a_13747_46662# 0.145228f
C18 a_3754_38470# VDAC_N 0.169096f
C19 a_8530_39574# a_5088_37509# 0.166912f
C20 a_n4064_37440# a_n2302_37690# 0.239588f
C21 a_7754_38470# a_5700_37509# 0.971846f
C22 a_n3420_39072# VDD 1.01442f
C23 a_n2293_43922# COMP_P 0.151768f
C24 a_2274_45254# a_2382_45260# 0.130215f
C25 a_n357_42282# a_5891_43370# 0.304889f
C26 a_15415_45028# VDD 0.191729f
C27 a_12549_44172# a_17639_46660# 0.129285f
C28 a_19279_43940# VDD 0.302681f
C29 a_n743_46660# a_310_45028# 0.143623f
C30 a_12465_44636# a_11823_42460# 0.127538f
C31 a_4185_45028# a_5932_42308# 0.118319f
C32 en_comp a_3080_42308# 1.28517f
C33 a_7112_43396# VDD 0.273193f
C34 a_9290_44172# a_n357_42282# 0.138435f
C35 a_9863_46634# VDD 0.411318f
C36 a_10193_42453# a_9803_42558# 0.20198f
C37 a_18494_42460# a_4190_30871# 0.242908f
C38 a_11136_42852# VDD 0.132515f
C39 a_16763_47508# a_16588_47582# 0.233657f
C40 a_16327_47482# a_10227_46804# 0.630403f
C41 a_4915_47217# a_11415_45002# 0.134061f
C42 a_n971_45724# a_1823_45246# 0.514159f
C43 a_3699_46634# a_3524_46660# 0.233657f
C44 C3_P_btm VREF_GND 0.67174f
C45 C4_P_btm VCM 0.716447f
C46 C10_N_btm VDD 2.40001f
C47 C2_P_btm VREF 0.987884f
C48 C0_P_btm VIN_P 0.529671f
C49 a_2063_45854# a_7499_43078# 0.478913f
C50 a_n2312_40392# a_n2302_40160# 0.151095f
C51 a_9482_43914# a_9672_43914# 0.122568f
C52 a_9801_43940# VDD 0.19512f
C53 a_5937_45572# a_5066_45546# 0.419426f
C54 a_20075_46420# a_19900_46494# 0.233657f
C55 a_20916_46384# VDD 0.302226f
C56 a_22612_30879# C10_N_btm 1.5848f
C57 a_1606_42308# a_6123_31319# 1.43958f
C58 a_742_44458# a_1568_43370# 0.525694f
C59 a_12545_42858# VDD 0.285703f
C60 a_6165_46155# VDD 0.204296f
C61 a_n3420_39072# a_n2946_39072# 0.238708f
C62 a_19332_42282# VDD 0.227361f
C63 a_8696_44636# a_16147_45260# 0.284694f
C64 a_10210_45822# VDD 0.323342f
C65 a_n1613_43370# a_2443_46660# 0.917984f
C66 VDAC_N C0_N_btm 0.324278f
C67 VDAC_P C0_dummy_P_btm 0.284358f
C68 a_n2946_37690# VDD 0.38221f
C69 a_n1838_35608# a_n1386_35608# 0.150796f
C70 a_15415_45028# a_15595_45028# 0.185422f
C71 a_21101_45002# VDD 0.2903f
C72 a_n2661_46098# a_n2157_46122# 0.227082f
C73 a_12545_42858# a_12895_43230# 0.215953f
C74 a_12379_42858# a_13460_43230# 0.102325f
C75 a_n2661_43370# a_n2661_43922# 0.13591f
C76 a_11415_45002# a_10809_44734# 0.140489f
C77 a_n1435_47204# CLK 1.41989f
C78 a_16023_47582# VDD 0.201413f
C79 a_n3674_38680# a_n4318_38216# 2.82961f
C80 a_5342_30871# a_4958_30871# 10.9366f
C81 a_5379_42460# VDD 0.213136f
C82 a_n2293_45546# a_n2293_45010# 0.257189f
C83 a_n863_45724# a_n2661_45010# 0.345234f
C84 a_n443_46116# a_n97_42460# 0.131756f
C85 a_n23_45546# VDD 0.150941f
C86 a_18479_47436# a_19321_45002# 0.262984f
C87 a_18597_46090# a_13747_46662# 0.391702f
C88 a_n443_46116# a_n2661_46098# 0.198865f
C89 a_n3690_39392# VDD 0.363068f
C90 a_7754_38470# a_5088_37509# 0.394117f
C91 a_n1613_43370# a_n1076_43230# 0.224215f
C92 a_10227_46804# a_12379_42858# 0.298444f
C93 a_2711_45572# a_14539_43914# 0.199754f
C94 a_14797_45144# VDD 0.124624f
C95 a_9863_46634# a_10150_46912# 0.233657f
C96 a_13747_46662# a_19123_46287# 0.191545f
C97 a_20766_44850# VDD 0.197657f
C98 a_n743_46660# a_n1099_45572# 0.108295f
C99 a_15227_44166# a_17715_44484# 0.385336f
C100 a_n357_42282# a_16795_42852# 0.180926f
C101 a_3537_45260# a_n97_42460# 0.74108f
C102 a_7287_43370# VDD 0.457521f
C103 a_15227_44166# a_15861_45028# 0.208121f
C104 a_1823_45246# a_2711_45572# 0.262616f
C105 a_8492_46660# VDD 0.273866f
C106 a_18184_42460# a_4190_30871# 0.630738f
C107 a_16327_47482# a_17591_47464# 0.339529f
C108 a_11599_46634# a_18597_46090# 0.191253f
C109 a_n97_42460# a_1049_43396# 0.195034f
C110 a_13507_46334# a_15743_43084# 0.158635f
C111 a_13747_46662# a_6755_46942# 0.316914f
C112 C4_P_btm VREF_GND 0.671882f
C113 C5_P_btm VCM 0.719982f
C114 C9_N_btm VDD 0.345685f
C115 C3_P_btm VREF 0.984942f
C116 C1_P_btm VIN_P 0.39234f
C117 a_13556_45296# a_11691_44458# 0.399095f
C118 a_n23_44458# VDD 0.169093f
C119 a_n2438_43548# a_526_44458# 0.107408f
C120 a_13747_46662# a_8049_45260# 0.208778f
C121 a_16388_46812# a_765_45546# 0.164902f
C122 a_n881_46662# a_13259_45724# 0.507296f
C123 a_3877_44458# a_2324_44458# 0.153319f
C124 a_6151_47436# a_6598_45938# 0.173467f
C125 a_n2312_40392# a_n4064_40160# 0.103899f
C126 a_12281_43396# a_12563_42308# 0.173003f
C127 a_10440_44484# a_10617_44484# 0.134298f
C128 a_8199_44636# a_5066_45546# 0.178583f
C129 a_1414_42308# a_453_43940# 0.248504f
C130 a_644_44056# a_895_43940# 0.106452f
C131 a_12089_42308# VDD 0.807892f
C132 a_n4318_37592# a_n3420_37984# 0.404896f
C133 a_n3674_38216# a_n4064_37984# 0.65176f
C134 a_5497_46414# VDD 0.200657f
C135 a_n3565_39304# a_n4064_39072# 0.344587f
C136 a_5891_43370# a_9127_43156# 0.457718f
C137 a_18907_42674# VDD 0.148872f
C138 a_11599_46634# a_6755_46942# 0.321942f
C139 a_n1613_43370# a_n2661_46098# 1.40554f
C140 VDAC_N C0_dummy_N_btm 0.287929f
C141 VDAC_P C0_P_btm 0.322595f
C142 a_n3420_37440# VDD 2.26579f
C143 a_n357_42282# a_3422_30871# 0.122733f
C144 a_n2293_46098# a_n97_42460# 0.333817f
C145 a_21005_45260# VDD 0.184261f
C146 a_15009_46634# a_3090_45724# 0.154981f
C147 a_n2497_47436# a_n755_45592# 0.45034f
C148 a_11599_46634# a_8049_45260# 0.14064f
C149 a_3626_43646# a_6123_31319# 0.109715f
C150 a_2982_43646# a_5934_30871# 0.178f
C151 a_12545_42858# a_13113_42826# 0.178024f
C152 a_n2661_43370# a_n2661_42834# 0.306215f
C153 a_4646_46812# a_6511_45714# 0.421269f
C154 a_n881_46662# a_17478_45572# 0.11503f
C155 a_16327_47482# VDD 2.81451f
C156 a_n2661_42834# a_2998_44172# 0.790177f
C157 a_14539_43914# a_15682_43940# 0.161926f
C158 a_22400_42852# a_22465_38105# 0.199207f
C159 a_19321_45002# a_19113_45348# 0.147788f
C160 a_12594_46348# a_11962_45724# 0.177228f
C161 a_10903_43370# a_11823_42460# 1.16382f
C162 a_n967_45348# a_n961_42308# 0.174237f
C163 a_n2017_45002# a_n1630_35242# 0.111641f
C164 a_5267_42460# VDD 0.170631f
C165 a_7499_43078# a_8696_44636# 0.155392f
C166 a_n356_45724# VDD 0.719282f
C167 a_n2956_37592# a_n4315_30879# 0.107228f
C168 a_18597_46090# a_13661_43548# 0.266647f
C169 a_n3565_39304# VDD 0.888861f
C170 a_n3565_39590# VREF 0.417978f
C171 a_n4209_39590# VCM 0.179761f
C172 a_3754_38470# a_5700_37509# 0.124176f
C173 a_7754_38470# a_4338_37500# 0.208284f
C174 a_8530_39574# a_3726_37500# 1.35509f
C175 a_n1613_43370# a_n901_43156# 0.281398f
C176 a_2711_45572# a_16112_44458# 0.183744f
C177 a_13661_43548# a_743_42282# 0.132115f
C178 a_8953_45002# CLK 0.310391f
C179 a_14537_43396# VDD 0.779752f
C180 a_2063_45854# a_10809_44734# 0.169005f
C181 a_7411_46660# a_6755_46942# 0.265786f
C182 a_3232_43370# a_3363_44484# 0.103472f
C183 a_21101_45002# a_21359_45002# 0.22264f
C184 a_20835_44721# VDD 0.198384f
C185 a_4190_30871# a_17303_42282# 0.279034f
C186 a_6547_43396# VDD 0.219105f
C187 a_15227_44166# a_8696_44636# 0.203885f
C188 a_16327_47482# a_11827_44484# 0.107078f
C189 a_5257_43370# a_3357_43084# 0.894879f
C190 a_8667_46634# VDD 0.39254f
C191 a_9290_44172# a_10951_45334# 0.136064f
C192 a_n1613_43370# a_n984_44318# 0.245331f
C193 a_3483_46348# a_1423_45028# 0.110369f
C194 a_2063_45854# a_n881_46662# 0.612456f
C195 a_16327_47482# a_16588_47582# 0.276601f
C196 a_21381_43940# a_2982_43646# 0.236232f
C197 a_10809_44734# a_n2661_42834# 0.14417f
C198 a_20273_45572# a_3357_43084# 0.358383f
C199 a_20731_45938# VDD 0.142103f
C200 C5_P_btm VREF_GND 0.676559f
C201 C6_P_btm VCM 0.877162f
C202 C8_N_btm VDD 0.19922f
C203 C4_P_btm VREF 0.98728f
C204 C2_P_btm VIN_P 0.502408f
C205 a_n2661_42282# a_5379_42460# 0.121051f
C206 a_9482_43914# a_11691_44458# 0.616964f
C207 a_n356_44636# VDD 1.17667f
C208 a_16388_46812# a_17339_46660# 0.24887f
C209 a_12891_46348# a_12638_46436# 0.13727f
C210 a_6151_47436# a_6667_45809# 0.1609f
C211 a_1307_43914# a_3499_42826# 0.532672f
C212 a_5883_43914# a_n2661_42834# 0.106812f
C213 a_2982_43646# CAL_N 0.181412f
C214 a_9165_43940# VDD 0.192035f
C215 a_11453_44696# a_6171_45002# 1.39146f
C216 a_20843_47204# VDD 0.188032f
C217 a_21588_30879# C9_N_btm 0.786375f
C218 a_19321_45002# START 0.10793f
C219 a_3823_42558# a_3905_42558# 0.171361f
C220 a_12379_42858# VDD 0.484153f
C221 a_584_46384# a_2998_44172# 0.181241f
C222 a_n1613_43370# a_n2661_43922# 0.113996f
C223 a_5204_45822# VDD 0.359177f
C224 a_2063_45854# a_n443_46116# 0.177177f
C225 a_n3690_39392# a_n3420_39072# 0.414961f
C226 a_n3565_39304# a_n2946_39072# 0.410957f
C227 a_1736_39587# a_1736_39043# 1.92825f
C228 a_n4334_39392# a_n4064_39072# 0.410653f
C229 a_n4209_39304# a_n2302_39072# 0.407162f
C230 a_18727_42674# VDD 0.181095f
C231 a_8697_45822# VDD 0.189893f
C232 VDAC_P C1_P_btm 0.560533f
C233 a_n3690_37440# VDD 0.363068f
C234 a_n1761_44111# a_n473_42460# 0.110251f
C235 a_2982_43646# a_5649_42852# 0.205161f
C236 a_20567_45036# VDD 0.237324f
C237 a_12379_42858# a_12895_43230# 0.109156f
C238 a_18479_45785# a_15493_43396# 0.235084f
C239 a_413_45260# a_2127_44172# 0.104737f
C240 a_4223_44672# a_5343_44458# 0.229803f
C241 a_n699_43396# a_4743_44484# 0.235328f
C242 a_4646_46812# a_6472_45840# 0.129446f
C243 a_n881_46662# a_15861_45028# 0.153795f
C244 a_16241_47178# VDD 0.208959f
C245 a_17517_44484# a_22591_44484# 0.196232f
C246 a_2324_44458# a_9049_44484# 0.102942f
C247 a_16721_46634# VDD 0.186443f
C248 a_15493_43396# a_14021_43940# 0.139192f
C249 a_3823_42558# VDD 0.170296f
C250 a_3503_45724# VDD 0.129733f
C251 en_comp a_22465_38105# 0.533581f
C252 a_12465_44636# a_768_44030# 0.120859f
C253 a_10227_46804# a_19321_45002# 0.111029f
C254 a_18780_47178# a_13661_43548# 0.153988f
C255 a_n3420_37440# a_n4064_37440# 8.19012f
C256 a_3754_38470# a_5088_37509# 0.632585f
C257 a_7754_38470# a_3726_37500# 0.124796f
C258 VDAC_Ni a_6886_37412# 0.178275f
C259 a_n4334_39392# VDD 0.385989f
C260 a_19319_43548# a_19268_43646# 0.17076f
C261 a_6293_42852# a_6452_43396# 0.157972f
C262 a_7287_43370# a_7112_43396# 0.234322f
C263 a_8696_44636# a_n2661_43370# 0.674122f
C264 a_n1613_43370# a_n1641_43230# 0.152896f
C265 a_10227_46804# a_10922_42852# 0.159426f
C266 a_14180_45002# VDD 0.151315f
C267 a_n2293_42834# a_5343_44458# 0.165923f
C268 a_20679_44626# VDD 0.439119f
C269 a_768_44030# a_2711_45572# 0.529995f
C270 a_22959_46660# a_21076_30879# 0.165603f
C271 a_4190_30871# a_4958_30871# 11.510201f
C272 a_n699_43396# a_1414_42308# 0.104607f
C273 a_n913_45002# a_4905_42826# 0.101072f
C274 a_6765_43638# VDD 0.218204f
C275 a_5066_45546# a_8034_45724# 0.242476f
C276 a_7927_46660# VDD 0.187888f
C277 a_11551_42558# a_11633_42558# 0.171361f
C278 a_10057_43914# a_10695_43548# 0.148476f
C279 a_n357_42282# a_20712_42282# 0.173926f
C280 a_3090_45724# a_4223_44672# 0.269823f
C281 a_8199_44636# a_9482_43914# 0.276776f
C282 a_n1613_43370# a_n809_44244# 0.291484f
C283 a_9290_44172# a_10775_45002# 0.215292f
C284 a_584_46384# a_n881_46662# 0.286501f
C285 a_16327_47482# a_16763_47508# 0.338544f
C286 a_22465_38105# a_22469_39537# 0.576946f
C287 a_16327_47482# a_16823_43084# 0.535969f
C288 a_3090_45724# a_15493_43940# 0.255251f
C289 a_20107_45572# a_3357_43084# 0.308463f
C290 a_526_44458# a_5891_43370# 1.12739f
C291 a_10227_46804# a_13059_46348# 0.656528f
C292 a_2063_45854# a_n2293_46098# 0.994164f
C293 a_5807_45002# a_6755_46942# 1.47519f
C294 a_2609_46660# a_3524_46660# 0.118759f
C295 C7_P_btm VCM 1.58335f
C296 C6_P_btm VREF_GND 0.836236f
C297 C7_N_btm VDD 0.121904f
C298 C5_P_btm VREF 0.987144f
C299 C9_N_btm C10_N_btm 37.815998f
C300 C3_P_btm VIN_P 0.455045f
C301 a_3232_43370# a_n2661_44458# 0.468391f
C302 a_5807_45002# a_8049_45260# 1.37423f
C303 a_6151_47436# a_6511_45714# 0.3215f
C304 a_n2312_40392# a_n4315_30879# 0.389397f
C305 a_n4318_38680# a_n3674_38680# 3.04229f
C306 a_18184_42460# a_18579_44172# 0.161593f
C307 a_n755_45592# a_743_42282# 0.160592f
C308 a_9290_44172# a_526_44458# 0.200352f
C309 a_18985_46122# a_19900_46494# 0.118759f
C310 a_11453_44696# a_3232_43370# 0.132496f
C311 a_19594_46812# VDD 0.349555f
C312 a_1467_44172# a_1414_42308# 0.335735f
C313 a_1115_44172# a_453_43940# 0.150214f
C314 a_10341_42308# VDD 0.931019f
C315 a_10809_44734# a_8696_44636# 0.117876f
C316 a_16327_47482# a_19279_43940# 0.446333f
C317 a_n1613_43370# a_n2661_42834# 0.112184f
C318 a_5164_46348# VDD 0.717083f
C319 a_584_46384# a_n443_46116# 0.496286f
C320 a_n3565_39304# a_n3420_39072# 0.241179f
C321 a_n4209_39304# a_n4064_39072# 0.19711f
C322 a_18057_42282# VDD 0.130308f
C323 a_n1613_43370# a_n1352_43396# 0.244933f
C324 a_n755_45592# a_626_44172# 0.100613f
C325 a_10193_42453# a_n913_45002# 0.562004f
C326 VDAC_P C2_P_btm 1.03235f
C327 a_n3565_37414# VDD 0.783539f
C328 a_3626_43646# a_4361_42308# 5.20633f
C329 a_18494_42460# VDD 0.73193f
C330 a_n2661_46098# a_n2840_46090# 0.170439f
C331 a_n2293_46634# a_3483_46348# 0.157275f
C332 a_12089_42308# a_12545_42858# 0.261463f
C333 a_2982_43646# a_6123_31319# 0.163265f
C334 a_n97_42460# a_13575_42558# 0.179828f
C335 a_3499_42826# VDD 0.333472f
C336 a_n881_46662# a_8696_44636# 0.178516f
C337 a_584_46384# a_3537_45260# 0.108506f
C338 a_15673_47210# VDD 0.569224f
C339 a_22400_42852# COMP_P 0.614467f
C340 a_n2840_42282# a_n3674_38680# 0.154001f
C341 a_17517_44484# a_22485_44484# 0.110643f
C342 a_n356_44636# a_n2661_42282# 2.54767f
C343 a_13661_43548# a_11691_44458# 0.263889f
C344 a_3090_45724# a_413_45260# 0.135828f
C345 a_n1613_43370# a_n1352_44484# 0.232498f
C346 a_10903_43370# a_11962_45724# 0.357882f
C347 a_16388_46812# VDD 0.797417f
C348 a_n2017_45002# a_n3674_37592# 0.241068f
C349 a_2479_44172# a_n97_42460# 0.196935f
C350 a_3318_42354# VDD 0.203036f
C351 a_5934_30871# C5_P_btm 0.139996f
C352 a_584_46384# a_1049_43396# 0.148494f
C353 a_3316_45546# VDD 0.428912f
C354 a_n3420_37440# a_n2946_37690# 0.236674f
C355 a_3754_38470# a_4338_37500# 0.473597f
C356 a_n4209_39590# VREF 0.860047f
C357 a_n4209_39304# VDD 0.984278f
C358 a_n1613_43370# a_n1423_42826# 0.15981f
C359 a_10227_46804# a_10991_42826# 0.152133f
C360 a_13661_43548# a_4190_30871# 0.147163f
C361 a_3483_46348# a_9672_43914# 0.125466f
C362 a_13777_45326# VDD 0.145151f
C363 a_10193_42453# a_18451_43940# 0.20167f
C364 a_4185_45028# a_4190_30871# 0.16524f
C365 a_21005_45260# a_21101_45002# 0.419086f
C366 a_20640_44752# VDD 0.246486f
C367 a_12549_44172# a_2711_45572# 2.05236f
C368 a_15227_44166# a_2324_44458# 0.190521f
C369 a_6197_43396# VDD 0.408793f
C370 a_8145_46902# VDD 0.199702f
C371 a_7499_43078# a_9803_42558# 0.158876f
C372 a_n1613_43370# a_n1549_44318# 0.16289f
C373 a_5066_45546# VDD 1.34058f
C374 a_15673_47210# a_16588_47582# 0.125324f
C375 a_15507_47210# a_10227_46804# 0.23187f
C376 a_16327_47482# a_16023_47582# 0.159305f
C377 a_21188_45572# VDD 0.288663f
C378 a_11599_46634# a_765_45546# 0.332797f
C379 a_2443_46660# a_3524_46660# 0.102325f
C380 a_3177_46902# a_2959_46660# 0.209641f
C381 C7_P_btm VREF_GND 1.61142f
C382 C8_P_btm VCM 2.61094f
C383 C6_N_btm VDD 0.210613f
C384 C6_P_btm VREF 1.41944f
C385 C8_N_btm C10_N_btm 0.878696f
C386 C4_P_btm VIN_P 0.50261f
C387 a_18597_46090# a_n357_42282# 0.250702f
C388 a_5257_43370# a_5937_45572# 0.262028f
C389 a_n3674_39304# a_n3674_38680# 0.17962f
C390 a_19778_44110# a_18579_44172# 0.268475f
C391 a_19553_46090# a_19335_46494# 0.209641f
C392 a_18819_46122# a_19900_46494# 0.102355f
C393 a_19321_45002# VDD 1.01574f
C394 a_5267_42460# a_5379_42460# 0.156424f
C395 a_1115_44172# a_1414_42308# 0.134389f
C396 a_n913_45002# a_2075_43172# 0.175893f
C397 a_10922_42852# VDD 0.216186f
C398 a_n356_45724# a_n23_45546# 0.360492f
C399 a_n2661_45546# a_2711_45572# 0.359276f
C400 a_21076_30879# a_413_45260# 0.141502f
C401 a_16327_47482# a_20766_44850# 0.17113f
C402 a_n755_45592# a_1609_45822# 0.12055f
C403 a_n1741_47186# a_9313_45822# 0.102019f
C404 a_n3565_39304# a_n3690_39392# 0.247167f
C405 a_5891_43370# a_8037_42858# 0.12253f
C406 a_17531_42308# VDD 0.262303f
C407 a_n1613_43370# a_n1177_43370# 0.325171f
C408 a_n357_42282# a_626_44172# 0.551369f
C409 a_10193_42453# a_n1059_45260# 0.440111f
C410 VDAC_P C3_P_btm 1.99006f
C411 a_n4334_37440# VDD 0.385859f
C412 en_comp a_n2661_43370# 0.164814f
C413 a_18184_42460# VDD 2.05053f
C414 a_n2312_39304# a_n2956_39304# 6.38528f
C415 a_12379_42858# a_12545_42858# 0.810394f
C416 a_4223_44672# a_n699_43396# 0.217586f
C417 a_413_45260# a_1414_42308# 0.12534f
C418 a_3483_46348# a_8953_45546# 0.133493f
C419 a_15811_47375# VDD 0.979053f
C420 a_11459_47204# DATA[5] 0.370451f
C421 a_n1059_45260# a_16137_43396# 0.438785f
C422 a_20679_44626# a_19279_43940# 0.279785f
C423 a_20835_44721# a_20766_44850# 0.209641f
C424 a_10193_42453# a_19987_42826# 0.164153f
C425 a_5807_45002# a_11691_44458# 0.117249f
C426 a_n1613_43370# a_n1177_44458# 0.332209f
C427 a_13059_46348# VDD 0.955445f
C428 a_18057_42282# a_18214_42558# 0.18824f
C429 a_15493_43940# a_22959_43948# 0.182001f
C430 en_comp COMP_P 1.92051f
C431 a_2903_42308# VDD 0.22017f
C432 a_6123_31319# C4_P_btm 0.132906f
C433 a_3218_45724# VDD 0.133843f
C434 a_10227_46804# a_13747_46662# 0.16398f
C435 a_n3565_37414# a_n4064_37440# 0.230258f
C436 a_3754_38470# a_3726_37500# 0.554457f
C437 VDAC_Ni a_5088_37509# 1.70462f
C438 a_1343_38525# VDD 3.25389f
C439 a_13556_45296# VDD 0.569056f
C440 a_8667_46634# a_8492_46660# 0.233657f
C441 a_n3674_39304# a_n4318_38680# 2.92578f
C442 a_10193_42453# a_18326_43940# 0.130866f
C443 a_20362_44736# VDD 0.275577f
C444 a_12741_44636# a_22959_46660# 0.17409f
C445 a_20820_30879# a_21076_30879# 8.6867f
C446 a_n2293_42282# a_n3674_38216# 0.111055f
C447 a_6293_42852# VDD 0.401011f
C448 a_7577_46660# VDD 0.249866f
C449 a_1606_42308# a_7174_31319# 2.41314f
C450 a_10057_43914# a_9145_43396# 0.121499f
C451 a_8016_46348# a_9482_43914# 0.293982f
C452 a_7227_45028# a_7230_45938# 0.170618f
C453 a_n1613_43370# a_n1331_43914# 0.16678f
C454 a_13059_46348# a_11827_44484# 0.495367f
C455 a_8270_45546# a_8975_43940# 0.207334f
C456 a_16241_47178# a_16023_47582# 0.209641f
C457 a_11599_46634# a_10227_46804# 0.60865f
C458 a_2684_37794# VDAC_Pi 0.133177f
C459 a_22465_38105# a_22545_38993# 0.253407f
C460 a_21363_45546# VDD 0.36538f
C461 a_11599_46634# a_17339_46660# 0.131185f
C462 a_2609_46660# a_2959_46660# 0.216095f
C463 C8_P_btm VREF_GND 2.58605f
C464 C9_P_btm VCM 6.06251f
C465 C5_N_btm VDD 0.267489f
C466 C7_P_btm VREF 1.818f
C467 C7_N_btm C10_N_btm 0.680974f
C468 C8_N_btm C9_N_btm 29.256199f
C469 C5_P_btm VIN_P 0.502041f
C470 a_413_45260# a_n699_43396# 0.100762f
C471 a_4791_45118# a_7227_45028# 0.288276f
C472 a_6151_47436# a_6194_45824# 0.227219f
C473 a_18494_42460# a_19279_43940# 0.137363f
C474 a_n356_44636# a_n23_44458# 0.220577f
C475 a_7499_43940# VDD 0.193884f
C476 a_n1613_43370# a_n967_45348# 0.213625f
C477 a_18985_46122# a_19335_46494# 0.210876f
C478 a_1606_42308# a_5932_42308# 0.111585f
C479 a_1115_44172# a_1467_44172# 0.115277f
C480 a_n913_45002# a_1847_42826# 0.294312f
C481 a_175_44278# a_453_43940# 0.112594f
C482 a_n3674_38216# a_n3565_38216# 0.128699f
C483 a_10991_42826# VDD 0.201891f
C484 a_16327_47482# a_20835_44721# 0.157393f
C485 a_n755_45592# a_n443_42852# 0.469263f
C486 a_4704_46090# VDD 0.225404f
C487 a_3160_47472# a_n1151_42308# 0.357683f
C488 a_2905_45572# a_3381_47502# 0.208262f
C489 a_5891_43370# a_7765_42852# 0.168516f
C490 a_17303_42282# VDD 0.379254f
C491 a_n1613_43370# a_n1917_43396# 0.153085f
C492 a_n755_45592# a_375_42282# 0.366231f
C493 a_2747_46873# a_2864_46660# 0.174836f
C494 a_11599_46634# a_10467_46802# 0.261176f
C495 a_12861_44030# a_6755_46942# 0.376009f
C496 VDAC_P C4_P_btm 3.9276f
C497 a_n4209_37414# VDD 0.817347f
C498 a_8530_39574# RST_Z 0.431385f
C499 a_2982_43646# a_4361_42308# 0.545077f
C500 a_19778_44110# VDD 0.469922f
C501 a_12549_44172# a_10903_43370# 0.792848f
C502 a_n2438_43548# a_1138_42852# 0.646257f
C503 a_12861_44030# a_8049_45260# 0.109405f
C504 a_12379_42858# a_12089_42308# 0.16885f
C505 a_3483_46348# a_5937_45572# 0.767636f
C506 a_n1151_42308# a_413_45260# 0.135643f
C507 SMPL_ON_N a_21589_35634# 0.399184f
C508 a_15507_47210# VDD 0.441662f
C509 a_n2017_45002# a_16137_43396# 0.63011f
C510 a_20640_44752# a_19279_43940# 0.22152f
C511 a_19615_44636# a_18579_44172# 0.158449f
C512 a_5111_44636# a_9803_43646# 0.118936f
C513 a_n1613_43370# a_n1917_44484# 0.153277f
C514 a_9290_44172# a_11823_42460# 0.864145f
C515 a_15227_46910# VDD 0.229766f
C516 a_18727_42674# a_18907_42674# 0.185422f
C517 a_2713_42308# VDD 0.208275f
C518 a_526_44458# a_1423_45028# 0.133656f
C519 a_4185_45028# a_22959_45036# 0.17601f
C520 a_584_46384# a_458_43396# 0.196763f
C521 a_2957_45546# VDD 0.192471f
C522 a_n4064_40160# VCM 0.121302f
C523 a_n4334_37440# a_n4064_37440# 0.448688f
C524 a_n3690_37440# a_n3420_37440# 0.431074f
C525 a_n3565_37414# a_n2946_37690# 0.407439f
C526 a_n4209_37414# a_n2302_37690# 0.407594f
C527 VDAC_Ni a_4338_37500# 0.640521f
C528 a_7754_38636# a_5088_37509# 0.288061f
C529 a_n4209_39590# VIN_P 0.105382f
C530 a_14021_43940# a_22959_43396# 0.191956f
C531 a_6197_43396# a_7112_43396# 0.118423f
C532 a_n1613_43370# a_n1853_43023# 0.423772f
C533 a_10227_46804# a_10835_43094# 0.295543f
C534 a_413_45260# a_327_44734# 0.195096f
C535 a_9482_43914# VDD 1.75061f
C536 a_13661_43548# a_17339_46660# 0.599051f
C537 a_5807_45002# a_765_45546# 0.103324f
C538 a_5649_42852# a_5111_42852# 0.110096f
C539 a_15743_43084# a_15567_42826# 0.215954f
C540 a_1823_45246# a_4361_42308# 0.11884f
C541 a_20159_44458# VDD 0.345429f
C542 a_6031_43396# VDD 0.47547f
C543 a_12861_44030# a_20193_45348# 0.680394f
C544 a_13661_43548# a_1307_43914# 0.396211f
C545 a_n2661_46634# a_13017_45260# 0.123713f
C546 a_7715_46873# VDD 0.414019f
C547 a_13661_43548# a_18579_44172# 0.229269f
C548 a_15507_47210# a_16588_47582# 0.102325f
C549 a_14955_47212# a_10227_46804# 0.175517f
C550 a_15673_47210# a_16023_47582# 0.228897f
C551 a_16241_47178# a_16327_47482# 0.185907f
C552 a_22465_38105# a_22521_39511# 0.902378f
C553 a_n4318_40392# a_n4315_30879# 0.151169f
C554 a_20623_45572# VDD 0.200978f
C555 a_12861_44030# a_18285_46348# 0.247326f
C556 a_2443_46660# a_2959_46660# 0.110816f
C557 a_2609_46660# a_3177_46902# 0.17072f
C558 C9_P_btm VREF_GND 5.18245f
C559 C10_P_btm VCM 10.3108f
C560 C4_N_btm VDD 0.265463f
C561 C8_P_btm VREF 3.6701f
C562 C6_N_btm C10_N_btm 0.421276f
C563 C7_N_btm C9_N_btm 0.227839f
C564 C6_P_btm VIN_P 0.391898f
C565 a_n1809_44850# VDD 0.132538f
C566 a_3090_45724# a_11415_45002# 0.16525f
C567 a_6151_47436# a_5907_45546# 0.274247f
C568 a_12089_42308# a_12800_43218# 0.15794f
C569 a_7499_43078# a_10695_43548# 0.124597f
C570 a_18184_42460# a_19279_43940# 0.132218f
C571 a_6671_43940# VDD 0.227011f
C572 a_18985_46122# a_19553_46090# 0.16939f
C573 a_18819_46122# a_19335_46494# 0.108964f
C574 a_13747_46662# VDD 3.70214f
C575 a_n699_43396# a_104_43370# 0.21575f
C576 a_10796_42968# VDD 0.270235f
C577 a_16327_47482# a_20679_44626# 0.318301f
C578 a_10227_46804# a_11967_42832# 0.461417f
C579 a_12465_44636# a_14673_44172# 0.101564f
C580 a_10586_45546# a_11962_45724# 0.137051f
C581 a_n357_42282# a_n443_42852# 0.763015f
C582 a_4419_46090# VDD 0.664887f
C583 a_n2661_42282# a_6293_42852# 0.16527f
C584 a_14539_43914# a_17595_43084# 0.141972f
C585 a_4958_30871# VDD 1.06745f
C586 a_n1613_43370# a_n1699_43638# 0.160308f
C587 a_2711_45572# a_6171_45002# 0.457554f
C588 a_n357_42282# a_375_42282# 0.142311f
C589 a_17339_46660# a_11967_42832# 0.493072f
C590 VDAC_P C5_P_btm 7.72471f
C591 a_8530_39574# VDD 0.346613f
C592 a_14180_45002# a_14537_43396# 0.143922f
C593 a_18911_45144# VDD 0.218047f
C594 a_12891_46348# a_10903_43370# 0.132903f
C595 a_n13_43084# a_133_42852# 0.171361f
C596 a_3483_46348# a_8199_44636# 1.81719f
C597 a_3090_45724# a_13259_45724# 0.261789f
C598 a_2107_46812# a_9049_44484# 0.240008f
C599 a_3160_47472# a_413_45260# 0.208121f
C600 a_n1435_47204# a_3357_43084# 1.08491f
C601 a_5164_46348# a_5497_46414# 0.203417f
C602 a_11599_46634# VDD 5.64965f
C603 a_20679_44626# a_20835_44721# 0.105995f
C604 a_20640_44752# a_20766_44850# 0.17072f
C605 a_13249_42308# a_5534_30871# 0.215947f
C606 a_11967_42832# a_18579_44172# 0.158329f
C607 a_12465_44636# a_12607_44458# 0.186652f
C608 a_n1613_43370# a_n1699_44726# 0.166123f
C609 a_10903_43370# a_11322_45546# 0.313957f
C610 a_n2293_43922# a_12281_43396# 0.147288f
C611 a_1414_42308# a_n97_42460# 0.196768f
C612 a_n784_42308# VCM 0.195503f
C613 a_1848_45724# VDD 0.100884f
C614 a_10227_46804# a_5807_45002# 0.262866f
C615 a_n4064_40160# VREF_GND 0.493568f
C616 a_n4209_37414# a_n4064_37440# 0.265895f
C617 a_n3565_37414# a_n3420_37440# 0.307576f
C618 VDAC_Ni a_3726_37500# 1.5261f
C619 a_18494_42460# a_18907_42674# 0.11494f
C620 a_6765_43638# a_6547_43396# 0.209641f
C621 a_n1613_43370# a_n2157_42858# 0.303592f
C622 a_10227_46804# a_10518_42984# 0.225803f
C623 a_4791_45118# a_2324_44458# 0.19212f
C624 a_3232_43370# a_9313_44734# 0.11426f
C625 a_19615_44636# VDD 0.203841f
C626 a_n881_46662# a_6511_45714# 0.149116f
C627 a_20820_30879# a_12741_44636# 0.103478f
C628 a_n2442_46660# a_n2302_39866# 0.161638f
C629 a_3080_42308# VCM 0.148824f
C630 a_12861_44030# a_11691_44458# 0.196929f
C631 a_3090_45724# a_17478_45572# 0.128299f
C632 a_7411_46660# VDD 0.41059f
C633 a_11323_42473# a_5742_30871# 0.198522f
C634 a_16922_45042# a_743_42282# 0.120316f
C635 a_n1613_43370# a_n1761_44111# 0.148121f
C636 a_167_45260# a_1423_45028# 0.123079f
C637 a_n237_47217# a_8128_46384# 0.113499f
C638 a_15673_47210# a_16327_47482# 0.206019f
C639 a_n4064_37984# a_n2302_37984# 0.250408f
C640 a_20841_45814# VDD 0.209907f
C641 C10_P_btm VREF_GND 10.3207f
C642 C3_N_btm VDD 0.26836f
C643 C9_P_btm VREF 7.369471f
C644 C5_N_btm C10_N_btm 0.285351f
C645 C6_N_btm C9_N_btm 0.169882f
C646 C7_N_btm C8_N_btm 23.7884f
C647 C7_P_btm VIN_P 1.52449f
C648 a_n2293_46634# a_526_44458# 0.579444f
C649 a_8975_43940# a_9313_44734# 0.391938f
C650 a_5829_43940# VDD 0.156797f
C651 a_765_45546# a_n357_42282# 0.209746f
C652 a_2324_44458# a_6945_45028# 0.183081f
C653 a_13661_43548# VDD 3.93017f
C654 a_20202_43084# a_21335_42336# 0.227943f
C655 a_n1059_45260# a_791_42968# 0.122941f
C656 a_n699_43396# a_n97_42460# 0.152094f
C657 a_10835_43094# VDD 0.43308f
C658 a_310_45028# a_n443_42852# 0.376934f
C659 a_4185_45028# VDD 1.65665f
C660 a_2905_45572# a_3160_47472# 0.54473f
C661 a_n237_47217# a_6151_47436# 0.360224f
C662 a_n4209_39304# a_n3565_39304# 6.82668f
C663 a_5891_43370# a_7227_42852# 0.129383f
C664 a_n863_45724# a_1423_45028# 0.113534f
C665 a_7499_43078# a_n913_45002# 0.548687f
C666 a_6151_47436# a_8270_45546# 0.142873f
C667 VDAC_P C6_P_btm 15.441001f
C668 a_7754_38470# VDD 0.302129f
C669 SMPL_ON_P a_n1630_35242# 6.11548f
C670 a_n2497_47436# a_n863_45724# 0.337007f
C671 a_16327_47482# a_21188_45572# 0.227468f
C672 a_584_46384# a_2382_45260# 0.185451f
C673 a_2905_45572# a_413_45260# 0.124898f
C674 a_5164_46348# a_5204_45822# 0.132894f
C675 a_14955_47212# VDD 0.301751f
C676 a_14311_47204# RST_Z 0.184572f
C677 a_20640_44752# a_20835_44721# 0.20669f
C678 a_13661_43548# a_11827_44484# 0.120515f
C679 a_11341_43940# a_15493_43940# 0.216602f
C680 a_3422_30871# a_2982_43646# 0.140944f
C681 a_1467_44172# a_n97_42460# 0.190191f
C682 a_12549_44172# a_12429_44172# 0.137881f
C683 a_3090_45724# a_n2661_42834# 0.164804f
C684 a_526_44458# a_626_44172# 0.180416f
C685 a_997_45618# VDD 0.12359f
C686 a_16327_47482# a_19321_45002# 0.925259f
C687 a_13507_46334# a_12549_44172# 0.363125f
C688 a_n971_45724# a_4646_46812# 0.303249f
C689 a_n3565_37414# a_n3690_37440# 0.247968f
C690 a_n4315_30879# VCM 0.473529f
C691 a_1736_39587# VDD 3.14139f
C692 a_6197_43396# a_6547_43396# 0.216095f
C693 a_6031_43396# a_7112_43396# 0.101963f
C694 a_10227_46804# a_10083_42826# 0.292997f
C695 a_13159_45002# VDD 0.321035f
C696 a_7577_46660# a_8492_46660# 0.118423f
C697 a_16922_45042# a_20193_45348# 0.328274f
C698 a_11967_42832# VDD 2.67441f
C699 a_3090_45724# a_17715_44484# 0.108364f
C700 a_n881_46662# a_6472_45840# 0.179318f
C701 a_n2442_46660# a_n4064_39616# 0.224005f
C702 a_n2293_42282# a_n2472_42282# 0.163758f
C703 a_3090_45724# a_15861_45028# 0.125763f
C704 a_13661_43548# a_15595_45028# 0.214904f
C705 a_16327_47482# a_18184_42460# 0.168018f
C706 a_5257_43370# VDD 0.922495f
C707 a_10723_42308# a_5742_30871# 0.185564f
C708 a_2711_45572# a_10193_42453# 0.218272f
C709 a_n1613_43370# a_n2065_43946# 0.30437f
C710 a_1337_46116# VDD 0.20087f
C711 a_12861_44030# a_18143_47464# 0.394543f
C712 a_15507_47210# a_16023_47582# 0.109156f
C713 a_15673_47210# a_16241_47178# 0.183195f
C714 a_22465_38105# a_22459_39145# 0.98555f
C715 a_20273_45572# VDD 0.571099f
C716 a_11453_44696# a_15227_44166# 0.979188f
C717 a_2443_46660# a_2609_46660# 0.579196f
C718 a_12861_44030# a_765_45546# 0.190301f
C719 C2_N_btm VDD 0.268945f
C720 C10_P_btm VREF 14.773f
C721 C5_N_btm C9_N_btm 0.153949f
C722 C4_N_btm C10_N_btm 0.348092f
C723 C6_N_btm C8_N_btm 0.170091f
C724 C8_P_btm VIN_P 0.907642f
C725 a_18989_43940# VDD 0.342796f
C726 a_10227_46804# a_n357_42282# 0.103631f
C727 a_16388_46812# a_16721_46634# 0.222024f
C728 a_10057_43914# a_9313_44734# 0.139382f
C729 a_5745_43940# VDD 0.144352f
C730 a_5204_45822# a_5066_45546# 0.402457f
C731 a_n881_46662# a_n745_45366# 0.152998f
C732 a_18819_46122# a_18985_46122# 0.749955f
C733 a_5807_45002# VDD 1.75047f
C734 a_n1059_45260# a_685_42968# 0.103646f
C735 a_10518_42984# VDD 0.273357f
C736 a_10586_45546# a_11525_45546# 0.115475f
C737 a_584_46384# a_453_43940# 0.125447f
C738 a_16327_47482# a_20362_44736# 0.213851f
C739 a_13059_46348# a_14537_43396# 0.30244f
C740 a_3699_46348# VDD 0.208984f
C741 a_n2810_45572# a_n3565_38502# 0.409424f
C742 a_2952_47436# a_3160_47472# 0.192116f
C743 a_n971_45724# a_6545_47178# 0.295443f
C744 a_n4209_39304# a_n4334_39392# 0.253307f
C745 a_14021_43940# a_20974_43370# 0.893848f
C746 a_5891_43370# a_5755_42852# 0.160849f
C747 a_7499_43078# a_n1059_45260# 0.277353f
C748 a_12741_44636# a_n2293_43922# 0.114756f
C749 a_n1613_43370# a_n2129_43609# 0.44294f
C750 a_2324_44458# a_6298_44484# 0.315008f
C751 a_15143_45578# VDD 0.12071f
C752 VDAC_P C7_P_btm 30.8442f
C753 a_3754_38470# RST_Z 0.203816f
C754 a_2982_43646# a_21487_43396# 0.169809f
C755 a_3626_43646# a_743_42282# 0.147999f
C756 a_13556_45296# a_14537_43396# 0.590856f
C757 a_18315_45260# VDD 0.12623f
C758 a_768_44030# a_9290_44172# 0.189655f
C759 a_n97_42460# a_5742_30871# 0.259664f
C760 a_16327_47482# a_21363_45546# 0.276554f
C761 a_n881_46662# a_15765_45572# 0.58719f
C762 a_n1151_42308# a_n467_45028# 0.406349f
C763 a_5068_46348# a_5204_45822# 0.20685f
C764 a_14311_47204# VDD 0.241476f
C765 a_5891_43370# a_7845_44172# 0.119969f
C766 a_20640_44752# a_20679_44626# 0.582607f
C767 a_n2293_42834# a_n97_42460# 0.17628f
C768 a_16867_43762# VDD 0.132317f
C769 a_17364_32525# EN_VIN_BSTR_N 0.959329f
C770 a_19321_45002# a_20567_45036# 0.205038f
C771 a_11341_43940# a_22223_43948# 0.175191f
C772 a_5932_42308# C3_P_btm 0.121156f
C773 a_n755_45592# VDD 2.41485f
C774 a_n971_45724# a_3877_44458# 0.927248f
C775 a_n4209_37414# a_n3420_37440# 0.245806f
C776 a_n4315_30879# VREF_GND 0.168163f
C777 a_1239_39587# VDD 0.530104f
C778 a_6197_43396# a_6765_43638# 0.17072f
C779 a_4185_45028# a_n2661_42282# 0.833759f
C780 a_13017_45260# VDD 0.263701f
C781 a_8145_46902# a_7927_46660# 0.209641f
C782 a_n2661_43370# a_n2661_44458# 1.0558f
C783 a_16922_45042# a_11691_44458# 0.428229f
C784 a_19778_44110# a_21005_45260# 0.135527f
C785 a_22591_46660# a_20820_30879# 0.166885f
C786 a_11415_45002# a_12741_44636# 1.07921f
C787 a_n2293_46634# a_n863_45724# 0.157683f
C788 a_n1151_42308# a_n452_44636# 0.238824f
C789 a_167_45260# a_2277_45546# 0.214157f
C790 a_13661_43548# a_15415_45028# 0.133591f
C791 a_16922_45042# a_4190_30871# 0.353708f
C792 a_8199_44636# a_10951_45334# 0.237774f
C793 a_10903_43370# a_3232_43370# 0.114259f
C794 a_n1741_47186# a_12891_46348# 0.107238f
C795 a_12861_44030# a_10227_46804# 0.291378f
C796 a_15507_47210# a_16327_47482# 0.425757f
C797 a_22465_38105# a_22521_40055# 0.214039f
C798 a_20107_45572# VDD 0.458237f
C799 a_12861_44030# a_17339_46660# 1.25428f
C800 C9_P_btm VIN_P 1.82823f
C801 C1_N_btm VDD 0.264503f
C802 C6_N_btm C7_N_btm 20.5296f
C803 C5_N_btm C8_N_btm 0.148944f
C804 C3_N_btm C10_N_btm 0.208539f
C805 C4_N_btm C9_N_btm 0.1579f
C806 a_15743_43084# a_4190_30871# 0.290729f
C807 a_16751_45260# a_17023_45118# 0.13675f
C808 a_18374_44850# VDD 0.203584f
C809 a_5257_43370# a_6419_46155# 0.186651f
C810 a_n699_43396# a_n2661_42834# 0.131393f
C811 a_12741_44636# a_13259_45724# 0.113445f
C812 a_16131_47204# VDD 0.142103f
C813 a_n784_42308# a_5934_30871# 0.142087f
C814 a_n4318_38216# a_n4209_38216# 0.135236f
C815 a_10083_42826# VDD 0.461256f
C816 a_10586_45546# a_11322_45546# 0.220166f
C817 a_16327_47482# a_20159_44458# 0.270426f
C818 a_12861_44030# a_18579_44172# 0.221909f
C819 a_584_46384# a_1414_42308# 0.321387f
C820 a_3483_46348# VDD 2.29096f
C821 a_2063_45854# a_n1151_42308# 0.425035f
C822 a_n971_45724# a_6151_47436# 0.29974f
C823 a_2952_47436# a_2905_45572# 0.318161f
C824 a_n2661_42834# a_n4318_38680# 0.102282f
C825 a_18579_44172# a_19700_43370# 0.175511f
C826 a_4958_30871# C9_N_btm 0.209166f
C827 a_n1613_43370# a_n2433_43396# 0.299968f
C828 a_2324_44458# a_5518_44484# 0.112753f
C829 a_14495_45572# VDD 0.238674f
C830 a_n881_46662# a_2107_46812# 0.138703f
C831 a_19321_45002# a_19594_46812# 0.267862f
C832 VDAC_P C8_P_btm 61.723297f
C833 a_3754_38470# VDD 2.52245f
C834 a_n356_44636# a_17303_42282# 0.10316f
C835 a_n97_42460# a_n13_43084# 0.13246f
C836 a_17719_45144# VDD 0.1297f
C837 a_12991_46634# a_12816_46660# 0.233657f
C838 a_11453_44696# a_10809_44734# 0.274367f
C839 a_n2497_47436# a_n2293_45546# 0.307373f
C840 a_3080_42308# a_5934_30871# 1.27306f
C841 a_n755_45592# a_8147_43396# 0.134231f
C842 a_16327_47482# a_20623_45572# 0.168593f
C843 a_n1435_47204# a_2437_43646# 0.191468f
C844 a_n971_45724# a_5111_44636# 0.381443f
C845 a_5068_46348# a_5164_46348# 0.31819f
C846 a_9067_47204# DATA[4] 0.354356f
C847 a_13487_47204# VDD 0.273369f
C848 a_12861_44030# RST_Z 0.290405f
C849 a_20362_44736# a_20679_44626# 0.102355f
C850 a_n2661_43370# a_n2840_43370# 0.172532f
C851 a_n1613_43370# a_n2433_44484# 0.29864f
C852 a_10903_43370# a_10193_42453# 0.402091f
C853 a_13259_45724# a_16375_45002# 0.60955f
C854 a_526_44458# a_n443_42852# 2.06448f
C855 a_14513_46634# VDD 0.223375f
C856 a_2351_42308# VDD 0.188239f
C857 a_n357_42282# VDD 1.90108f
C858 a_16327_47482# a_13747_46662# 0.128159f
C859 a_16763_47508# a_5807_45002# 0.127783f
C860 a_n4315_30879# VREF 1.73216f
C861 a_18184_42460# a_18057_42282# 0.19301f
C862 a_6031_43396# a_6547_43396# 0.105995f
C863 a_n143_45144# a_n37_45144# 0.13675f
C864 a_n913_45002# a_3537_45260# 0.148413f
C865 a_11963_45334# VDD 0.229584f
C866 a_7577_46660# a_7927_46660# 0.206455f
C867 a_7411_46660# a_8492_46660# 0.102325f
C868 a_18184_42460# a_18494_42460# 1.31047f
C869 a_7229_43940# a_7640_43914# 0.177622f
C870 a_18588_44850# VDD 0.132317f
C871 a_20202_43084# a_12741_44636# 0.22243f
C872 a_11823_42460# a_743_42282# 0.147603f
C873 a_4185_45028# a_5379_42460# 0.189676f
C874 a_18287_44626# a_18579_44172# 0.107662f
C875 a_22165_42308# a_21887_42336# 0.110763f
C876 a_167_45260# a_1609_45822# 0.141505f
C877 a_13661_43548# a_14797_45144# 0.116989f
C878 a_18189_46348# a_16375_45002# 0.165328f
C879 a_584_46384# a_n699_43396# 0.632931f
C880 a_16922_45042# a_21259_43561# 0.108631f
C881 a_11599_46634# a_16327_47482# 0.526398f
C882 a_15811_47375# a_15673_47210# 0.281607f
C883 a_n3420_37984# a_n4064_37984# 8.18485f
C884 a_11341_43940# a_10341_43396# 0.289072f
C885 a_n2497_47436# a_1138_42852# 0.144386f
C886 C10_P_btm VIN_P 3.66034f
C887 C0_N_btm VDD 1.02806f
C888 C5_N_btm C7_N_btm 0.15419f
C889 C2_N_btm C10_N_btm 0.215144f
C890 C3_N_btm C9_N_btm 0.138859f
C891 C4_N_btm C8_N_btm 0.149948f
C892 a_2982_43646# a_5342_30871# 0.178973f
C893 a_16751_45260# a_16922_45042# 0.12103f
C894 SMPL_ON_N COMP_P 2.13516f
C895 a_18443_44721# VDD 0.193515f
C896 a_5257_43370# a_6165_46155# 0.11382f
C897 a_3626_43646# a_19647_42308# 0.170024f
C898 a_10341_42308# a_11554_42852# 0.170124f
C899 a_n1613_43370# a_n913_45002# 0.686014f
C900 a_765_45546# a_380_45546# 0.141908f
C901 a_n881_46662# a_n1059_45260# 0.121542f
C902 a_8952_43230# VDD 0.273404f
C903 a_3218_45724# a_3316_45546# 0.162813f
C904 a_n863_45724# a_1609_45822# 0.117311f
C905 a_10586_45546# a_10490_45724# 0.235237f
C906 a_3147_46376# VDD 0.341038f
C907 a_18597_46090# a_2982_43646# 0.239147f
C908 a_19692_46634# a_20512_43084# 0.387138f
C909 a_2324_44458# a_5343_44458# 0.255488f
C910 a_13249_42308# VDD 0.653917f
C911 a_2747_46873# a_2609_46660# 0.347674f
C912 VDAC_P C9_P_btm 0.123386p
C913 a_n356_44636# a_4958_30871# 0.46356f
C914 a_13556_45296# a_13777_45326# 0.101558f
C915 a_n2293_46634# a_1823_45246# 0.230429f
C916 a_n2293_42834# a_n2661_42834# 0.202366f
C917 a_742_44458# a_949_44458# 0.185221f
C918 a_n1441_43940# VDD 0.142719f
C919 a_16327_47482# a_20841_45814# 0.161808f
C920 a_n881_46662# a_15599_45572# 0.601034f
C921 a_4791_45118# a_n913_45002# 0.254334f
C922 a_6575_47204# DATA[4] 0.15718f
C923 a_12861_44030# VDD 3.56689f
C924 a_13717_47436# RST_Z 4.51263f
C925 a_20362_44736# a_20640_44752# 0.118759f
C926 a_19700_43370# VDD 0.28578f
C927 a_3483_46348# a_10907_45822# 0.140023f
C928 a_n2956_38680# a_n2946_38778# 0.14863f
C929 a_14180_46812# VDD 0.755623f
C930 a_2123_42473# VDD 0.1936f
C931 a_310_45028# VDD 0.360949f
C932 a_16327_47482# a_13661_43548# 0.132061f
C933 a_n4209_37414# a_n3565_37414# 6.90997f
C934 a_n97_42460# a_10341_43396# 0.917198f
C935 a_6293_42852# a_6197_43396# 0.213423f
C936 a_n1059_45260# a_3537_45260# 0.162323f
C937 a_11787_45002# VDD 0.153399f
C938 a_7577_46660# a_8145_46902# 0.170059f
C939 a_n901_43156# a_n1076_43230# 0.234322f
C940 a_n1853_43023# a_n1736_43218# 0.183149f
C941 a_3090_45724# a_2324_44458# 0.684819f
C942 a_n881_46662# a_5263_45724# 0.180025f
C943 a_11415_45002# a_22591_46660# 0.172844f
C944 a_167_45260# a_n443_42852# 0.246952f
C945 a_12861_44030# a_11827_44484# 0.466435f
C946 a_13661_43548# a_14537_43396# 0.505634f
C947 a_n743_46660# a_6171_45002# 0.140224f
C948 a_10533_42308# a_10723_42308# 0.23663f
C949 a_n2293_43922# a_n97_42460# 0.136247f
C950 a_8495_42852# VDD 0.132018f
C951 a_12549_44172# a_3422_30871# 0.148646f
C952 a_8270_45546# a_5883_43914# 0.20967f
C953 a_8199_44636# a_8953_45002# 0.12099f
C954 a_5937_45572# a_8191_45002# 0.180306f
C955 a_n237_47217# a_n881_46662# 0.958566f
C956 a_15507_47210# a_15673_47210# 0.81159f
C957 a_n3420_37984# a_n2946_37984# 0.238664f
C958 a_21363_45546# a_21188_45572# 0.233657f
C959 a_19864_35138# VIN_N 0.367112f
C960 C4_N_btm C7_N_btm 0.148546f
C961 C5_N_btm C6_N_btm 18.2841f
C962 C1_N_btm C10_N_btm 0.204172f
C963 C2_N_btm C9_N_btm 0.144261f
C964 C3_N_btm C8_N_btm 0.13616f
C965 EN_VIN_BSTR_N VCM 0.927905f
C966 a_17339_46660# a_15743_43084# 0.450316f
C967 a_18287_44626# VDD 0.389383f
C968 a_n971_45724# a_7499_43078# 0.857375f
C969 a_3626_43646# a_19511_42282# 0.182478f
C970 a_n1613_43370# a_n1059_45260# 0.202724f
C971 a_8270_45546# a_8162_45546# 0.170838f
C972 a_n784_42308# a_6123_31319# 0.144274f
C973 a_9127_43156# VDD 0.468721f
C974 a_16327_47482# a_11967_42832# 0.241578f
C975 a_13059_46348# a_13556_45296# 0.274813f
C976 a_n863_45724# a_n443_42852# 0.556081f
C977 a_584_46384# a_1115_44172# 0.174981f
C978 a_2804_46116# VDD 0.159351f
C979 a_n237_47217# a_n443_46116# 0.110841f
C980 a_17124_42282# VDD 0.28176f
C981 a_n2293_45546# a_626_44172# 0.150062f
C982 a_4185_45028# a_n356_44636# 1.54308f
C983 a_n863_45724# a_375_42282# 0.451905f
C984 a_13904_45546# VDD 0.135068f
C985 a_n1613_43370# a_948_46660# 0.281392f
C986 a_2747_46873# a_2443_46660# 0.129886f
C987 a_22609_38406# a_22609_37990# 0.32625f
C988 VDAC_P C10_P_btm 0.24639p
C989 VDAC_Ni VDD 0.288547f
C990 a_3422_30871# a_n1630_35242# 0.828871f
C991 a_9482_43914# a_13777_45326# 0.206086f
C992 a_3626_43646# a_4921_42308# 0.431551f
C993 a_3080_42308# a_6123_31319# 1.45722f
C994 a_10991_42826# a_10922_42852# 0.209641f
C995 a_10796_42968# a_10341_42308# 0.65943f
C996 a_11691_44458# a_16979_44734# 0.12231f
C997 a_n1151_42308# a_n967_45348# 0.170453f
C998 a_584_46384# a_413_45260# 0.164383f
C999 a_13717_47436# VDD 0.314317f
C1000 a_n1435_47204# RST_Z 0.179508f
C1001 a_7640_43914# a_7542_44172# 0.20977f
C1002 a_11823_42460# a_5534_30871# 0.511874f
C1003 a_19268_43646# VDD 0.237793f
C1004 a_19321_45002# a_19778_44110# 0.568668f
C1005 a_12741_44636# a_8696_44636# 2.20704f
C1006 a_16327_47482# a_18989_43940# 0.100946f
C1007 a_n2956_38680# a_n3420_38528# 0.233147f
C1008 a_14035_46660# VDD 0.363878f
C1009 a_13483_43940# a_14021_43940# 0.109097f
C1010 a_1755_42282# VDD 0.215277f
C1011 a_1606_42308# RST_Z 1.44945f
C1012 a_526_44458# a_1307_43914# 0.467539f
C1013 a_n1099_45572# VDD 0.89411f
C1014 a_16327_47482# a_5807_45002# 0.451783f
C1015 a_n4315_30879# VIN_P 0.187185f
C1016 a_n4209_37414# a_n4334_37440# 0.253282f
C1017 a_n2302_39866# VDD 0.361509f
C1018 a_6031_43396# a_6197_43396# 0.581047f
C1019 a_n913_45002# a_3065_45002# 0.225034f
C1020 a_10951_45334# VDD 0.226705f
C1021 a_9313_45822# a_5937_45572# 0.137696f
C1022 a_7411_46660# a_7927_46660# 0.105839f
C1023 a_19778_44110# a_18184_42460# 0.119002f
C1024 a_13259_45724# a_n97_42460# 0.182889f
C1025 a_765_45546# a_167_45260# 0.276049f
C1026 a_n2956_39768# a_n2946_39866# 0.14868f
C1027 a_n2442_46660# a_n3565_39590# 0.134948f
C1028 a_1823_45246# a_1609_45822# 0.35471f
C1029 a_8199_44636# a_8191_45002# 0.234072f
C1030 a_n443_42852# a_11823_42460# 0.356965f
C1031 a_n1925_42282# VDD 0.728242f
C1032 a_n746_45260# a_n881_46662# 0.190303f
C1033 a_15507_47210# a_15811_47375# 0.170975f
C1034 a_22465_38105# a_22521_40599# 0.132396f
C1035 a_n3565_38216# a_n4064_37984# 0.342209f
C1036 a_11967_42832# a_12379_42858# 0.492977f
C1037 a_11599_46634# a_16388_46812# 0.24092f
C1038 C3_N_btm C7_N_btm 0.136068f
C1039 C4_N_btm C6_N_btm 0.145942f
C1040 C0_N_btm C10_N_btm 0.251079f
C1041 C1_N_btm C9_N_btm 0.133953f
C1042 C2_N_btm C8_N_btm 0.14124f
C1043 EN_VIN_BSTR_N VREF_GND 0.85739f
C1044 a_18248_44752# VDD 0.251171f
C1045 a_3737_43940# VDD 0.18423f
C1046 a_11415_45002# a_13259_45724# 0.505354f
C1047 a_15227_44166# a_2711_45572# 0.113396f
C1048 a_2713_42308# a_2903_42308# 0.23738f
C1049 a_5111_44636# a_5649_42852# 0.121004f
C1050 a_8387_43230# VDD 0.200672f
C1051 a_13059_46348# a_9482_43914# 0.448068f
C1052 a_n2293_45546# a_1609_45822# 0.159696f
C1053 a_10586_45546# a_10193_42453# 0.380236f
C1054 a_12861_44030# a_19279_43940# 0.152657f
C1055 a_2698_46116# VDD 0.195879f
C1056 a_n237_47217# a_4791_45118# 0.10712f
C1057 a_13527_45546# VDD 0.1902f
C1058 a_n1613_43370# a_1123_46634# 0.358475f
C1059 a_768_44030# a_n2293_46634# 0.26984f
C1060 CAL_P a_22609_37990# 0.205305f
C1061 a_2982_43646# a_4190_30871# 0.3223f
C1062 a_5205_44484# a_1423_45028# 0.821456f
C1063 a_9482_43914# a_13556_45296# 0.726155f
C1064 a_18114_32519# EN_VIN_BSTR_N 0.187697f
C1065 a_16922_45042# VDD 1.54713f
C1066 a_11901_46660# a_12816_46660# 0.125324f
C1067 SMPL_ON_P a_n4315_30879# 3.70932f
C1068 a_10835_43094# a_10341_42308# 0.541777f
C1069 a_10796_42968# a_10922_42852# 0.170059f
C1070 a_11691_44458# a_14539_43914# 0.268287f
C1071 a_16327_47482# a_20107_45572# 0.674639f
C1072 a_n2661_46634# a_11823_42460# 0.331717f
C1073 a_n743_46660# a_10193_42453# 0.25279f
C1074 a_n1435_47204# VDD 0.267875f
C1075 a_20159_44458# a_20362_44736# 0.233657f
C1076 a_11967_42832# a_20679_44626# 0.863531f
C1077 a_15743_43084# VDD 0.572249f
C1078 a_13747_46662# a_18184_42460# 0.123281f
C1079 a_16327_47482# a_18374_44850# 0.16003f
C1080 a_11189_46129# a_10193_42453# 0.123385f
C1081 a_13885_46660# VDD 0.499249f
C1082 a_4958_30871# a_17531_42308# 0.192941f
C1083 a_20935_43940# a_21115_43940# 0.185422f
C1084 a_1606_42308# VDD 0.631207f
C1085 a_380_45546# VDD 0.154763f
C1086 a_n913_45002# a_21613_42308# 0.259761f
C1087 a_n4064_39616# VDD 1.6861f
C1088 a_6031_43396# a_6293_42852# 0.163953f
C1089 a_12549_44172# a_20556_43646# 0.125209f
C1090 a_n755_45592# a_n356_44636# 2.42652f
C1091 a_10775_45002# VDD 0.148349f
C1092 a_7715_46873# a_7577_46660# 0.205227f
C1093 a_13747_46662# a_13059_46348# 0.273684f
C1094 a_5807_45002# a_16721_46634# 0.112018f
C1095 a_3232_43370# a_5891_43370# 0.137859f
C1096 a_n2956_39768# a_n3420_39616# 0.233256f
C1097 a_10193_42453# a_4361_42308# 0.274131f
C1098 a_3539_42460# VDD 0.363092f
C1099 a_768_44030# a_626_44172# 0.186913f
C1100 a_1823_45246# a_n443_42852# 0.125287f
C1101 COMP_P a_22469_40625# 0.120018f
C1102 a_5937_45572# a_6709_45028# 0.629301f
C1103 a_526_44458# VDD 2.35177f
C1104 a_n971_45724# a_n881_46662# 0.236696f
C1105 a_n746_45260# a_n1613_43370# 0.146842f
C1106 a_2553_47502# a_2747_46873# 0.14563f
C1107 a_11599_46634# a_15811_47375# 0.107881f
C1108 a_2684_37794# a_2113_38308# 0.468006f
C1109 a_n4209_38216# a_n2302_37984# 0.407312f
C1110 a_n3565_38216# a_n2946_37984# 0.411006f
C1111 a_n3690_38304# a_n3420_37984# 0.414894f
C1112 a_n4334_38304# a_n4064_37984# 0.410244f
C1113 a_n2293_43922# a_n2293_42282# 0.19201f
C1114 a_3090_45724# a_15493_43396# 0.134629f
C1115 a_2711_45572# a_n2661_43370# 0.112998f
C1116 a_13507_46334# a_19692_46634# 0.823157f
C1117 a_11599_46634# a_13059_46348# 0.371555f
C1118 C0_P_btm VDD 1.02806f
C1119 C2_N_btm C7_N_btm 0.139982f
C1120 C3_N_btm C6_N_btm 0.134599f
C1121 C4_N_btm C5_N_btm 15.915401f
C1122 C0_dummy_N_btm C10_N_btm 0.63636f
C1123 C0_N_btm C9_N_btm 0.14782f
C1124 C1_N_btm C8_N_btm 0.131002f
C1125 a_n2661_42282# a_1755_42282# 0.145244f
C1126 a_17970_44736# VDD 0.27753f
C1127 a_15227_44166# a_22000_46634# 0.154332f
C1128 a_4915_47217# a_2711_45572# 0.265557f
C1129 a_16327_47482# a_n357_42282# 0.49929f
C1130 a_5883_43914# a_9313_44734# 0.124999f
C1131 a_14401_32519# EN_VIN_BSTR_N 0.772414f
C1132 a_11823_42460# a_13291_42460# 0.257506f
C1133 a_n809_44244# a_n984_44318# 0.234322f
C1134 a_8605_42826# VDD 0.204898f
C1135 a_n1151_42308# a_n1761_44111# 0.642214f
C1136 a_n755_45592# a_3503_45724# 0.163919f
C1137 a_1823_45246# a_2437_43646# 0.324477f
C1138 a_2521_46116# VDD 0.163553f
C1139 a_n971_45724# a_n443_46116# 0.129009f
C1140 a_16104_42674# VDD 0.134357f
C1141 a_2324_44458# a_4223_44672# 0.56408f
C1142 a_n2293_45546# a_375_42282# 0.104283f
C1143 a_9290_44172# a_8975_43940# 0.114958f
C1144 a_13163_45724# VDD 0.322298f
C1145 a_n1613_43370# a_383_46660# 0.182504f
C1146 a_9804_47204# a_n743_46660# 0.295465f
C1147 en_comp a_n2293_42834# 0.103485f
C1148 a_13348_45260# a_13556_45296# 0.189446f
C1149 a_n1925_42282# a_n2661_42282# 2.27741f
C1150 a_12469_46902# a_12251_46660# 0.209641f
C1151 a_10796_42968# a_10991_42826# 0.206455f
C1152 a_n971_45724# a_3537_45260# 0.266743f
C1153 a_13381_47204# VDD 0.130765f
C1154 a_7227_47204# DATA[3] 0.357377f
C1155 a_11967_42832# a_20640_44752# 0.588649f
C1156 a_18783_43370# VDD 0.289099f
C1157 a_13747_46662# a_19778_44110# 0.670692f
C1158 a_10903_43370# a_7499_43078# 0.888628f
C1159 a_16327_47482# a_18443_44721# 0.1665f
C1160 a_9290_44172# a_10193_42453# 1.23123f
C1161 a_n2956_38680# a_n3565_38502# 0.302523f
C1162 a_4958_30871# a_17303_42282# 0.168656f
C1163 a_19862_44208# a_15493_43940# 0.534481f
C1164 a_2324_44458# a_n2293_42834# 0.168086f
C1165 a_768_44030# a_9028_43914# 0.113848f
C1166 a_584_46384# a_n97_42460# 0.526796f
C1167 a_n452_45724# VDD 0.112977f
C1168 a_12465_44636# a_n881_46662# 0.813228f
C1169 a_584_46384# a_n2661_46098# 0.17431f
C1170 a_n2946_39866# VDD 0.393552f
C1171 a_12549_44172# a_743_42282# 0.119701f
C1172 a_n357_42282# a_n356_44636# 0.308599f
C1173 a_8953_45002# VDD 1.24336f
C1174 a_5807_45002# a_16388_46812# 0.235518f
C1175 a_13661_43548# a_13059_46348# 0.267127f
C1176 a_7411_46660# a_7577_46660# 0.634781f
C1177 a_n2472_42826# a_n4318_38680# 0.158196f
C1178 a_n1991_42858# a_n1076_43230# 0.123255f
C1179 a_n1853_43023# a_n13_43084# 0.109925f
C1180 a_16547_43609# a_16414_43172# 0.143695f
C1181 a_n2293_46634# a_n2661_45546# 0.85166f
C1182 a_10227_46804# a_11823_42460# 0.428745f
C1183 a_n881_46662# a_2711_45572# 0.170524f
C1184 a_n2661_42834# a_n2661_43922# 0.841361f
C1185 a_3626_43646# VDD 0.340378f
C1186 a_17715_44484# a_13259_45724# 0.391904f
C1187 a_1138_42852# a_n443_42852# 0.14758f
C1188 a_15368_46634# a_15599_45572# 0.100853f
C1189 a_13661_43548# a_13556_45296# 0.559682f
C1190 a_5275_47026# VDD 0.135766f
C1191 COMP_P a_22521_40599# 0.204681f
C1192 a_5937_45572# a_7229_43940# 0.126047f
C1193 a_19321_45002# a_11967_42832# 0.266816f
C1194 a_13259_45724# a_15861_45028# 0.16873f
C1195 a_2981_46116# VDD 0.111597f
C1196 a_11599_46634# a_15507_47210# 0.267808f
C1197 a_12861_44030# a_16327_47482# 0.120085f
C1198 a_n971_45724# a_n1613_43370# 0.6298f
C1199 a_n3565_38216# a_n3420_37984# 0.238595f
C1200 a_n4209_38216# a_n4064_37984# 0.19304f
C1201 a_3090_45724# a_19328_44172# 0.153704f
C1202 a_15227_44166# a_14955_43940# 0.134177f
C1203 a_20273_45572# a_21188_45572# 0.125324f
C1204 a_12549_44172# a_6755_46942# 0.553062f
C1205 a_4883_46098# a_15227_44166# 0.176028f
C1206 a_n971_45724# a_n2293_46098# 0.110318f
C1207 EN_VIN_BSTR_N VIN_N 1.41696f
C1208 C1_P_btm VDD 0.264503f
C1209 C1_N_btm C7_N_btm 0.129707f
C1210 C2_N_btm C6_N_btm 0.138423f
C1211 C0_dummy_N_btm C9_N_btm 0.11363f
C1212 C0_N_btm C8_N_btm 0.148433f
C1213 C3_N_btm C5_N_btm 0.136119f
C1214 EN_VIN_BSTR_P VCM 0.929333f
C1215 a_17767_44458# VDD 0.348803f
C1216 a_7499_43078# a_8685_43396# 0.153217f
C1217 a_10057_43914# a_5891_43370# 0.197199f
C1218 a_n755_45592# a_3318_42354# 0.152654f
C1219 a_8037_42858# VDD 0.344922f
C1220 a_310_45028# a_n356_45724# 0.12349f
C1221 a_167_45260# VDD 1.41955f
C1222 a_584_46384# a_2553_47502# 0.100103f
C1223 a_n3420_39616# a_n4064_39072# 6.32746f
C1224 a_1736_39587# a_1343_38525# 0.289453f
C1225 a_12791_45546# VDD 0.205486f
C1226 a_n1613_43370# a_601_46902# 0.178721f
C1227 a_5807_45002# a_19321_45002# 0.376188f
C1228 w_11334_34010# a_n1630_35242# 3.10971f
C1229 a_13348_45260# a_9482_43914# 0.352976f
C1230 a_13017_45260# a_13777_45326# 0.195607f
C1231 a_526_44458# a_n2661_42282# 0.191497f
C1232 a_11901_46660# a_12251_46660# 0.219633f
C1233 a_11735_46660# a_12816_46660# 0.102325f
C1234 a_10835_43094# a_10991_42826# 0.105839f
C1235 a_11691_44458# a_15004_44636# 0.221929f
C1236 a_n971_45724# a_3429_45260# 0.171338f
C1237 a_n2109_47186# a_5691_45260# 0.113268f
C1238 a_11459_47204# VDD 0.34771f
C1239 a_6851_47204# DATA[3] 0.146601f
C1240 a_4185_45028# a_17303_42282# 0.235259f
C1241 a_6109_44484# a_6453_43914# 0.165572f
C1242 a_18525_43370# VDD 0.263553f
C1243 a_12549_44172# a_20193_45348# 0.587618f
C1244 a_16327_47482# a_18287_44626# 0.552724f
C1245 a_11415_45002# a_8696_44636# 0.10924f
C1246 a_20692_30879# a_20447_31679# 9.02991f
C1247 a_n863_45724# VDD 1.89058f
C1248 a_11599_46634# a_13747_46662# 0.25325f
C1249 a_584_46384# a_1799_45572# 0.179456f
C1250 a_n3420_39616# VDD 0.568506f
C1251 a_8191_45002# VDD 0.39677f
C1252 a_n971_45724# a_6945_45028# 0.247957f
C1253 a_5807_45002# a_13059_46348# 0.1145f
C1254 a_7411_46660# a_7715_46873# 0.162909f
C1255 a_n1423_42826# a_n1641_43230# 0.209641f
C1256 a_1307_43914# a_14539_43914# 0.131617f
C1257 a_22365_46825# a_20202_43084# 0.115624f
C1258 a_n2956_39768# a_n3565_39590# 0.302561f
C1259 a_3540_43646# VDD 0.209044f
C1260 a_13661_43548# a_9482_43914# 0.127225f
C1261 a_17583_46090# a_13259_45724# 0.191869f
C1262 a_n2293_46098# a_2711_45572# 0.530463f
C1263 a_13059_46348# a_15143_45578# 0.262261f
C1264 a_n2293_42834# a_n2472_42826# 0.199703f
C1265 a_7309_42852# VDD 0.177437f
C1266 a_13259_45724# a_8696_44636# 0.259609f
C1267 a_n3565_38216# a_n3690_38304# 0.247167f
C1268 a_20107_45572# a_21188_45572# 0.102355f
C1269 a_20841_45814# a_20623_45572# 0.209641f
C1270 a_11453_44696# a_3090_45724# 0.232756f
C1271 a_11530_34132# VIN_N 1.547f
C1272 C2_P_btm VDD 0.268945f
C1273 C0_N_btm C7_N_btm 0.142187f
C1274 C0_dummy_N_btm C8_N_btm 0.236317f
C1275 C1_N_btm C6_N_btm 0.128559f
C1276 C3_N_btm C4_N_btm 7.90108f
C1277 C2_N_btm C5_N_btm 0.138678f
C1278 EN_VIN_BSTR_P VREF_GND 0.85739f
C1279 a_10193_42453# a_3422_30871# 0.404849f
C1280 a_8696_44636# a_n2661_43922# 0.257466f
C1281 a_16979_44734# VDD 0.256327f
C1282 a_4791_45118# a_2711_45572# 0.160646f
C1283 a_743_42282# a_564_42282# 0.169821f
C1284 a_18479_45785# a_19319_43548# 0.102555f
C1285 a_2455_43940# VDD 0.144352f
C1286 a_768_44030# a_2437_43646# 0.137571f
C1287 a_10903_43370# a_10809_44734# 0.353301f
C1288 a_7765_42852# VDD 0.333322f
C1289 a_17715_44484# a_15861_45028# 0.184272f
C1290 a_2202_46116# VDD 0.20904f
C1291 a_584_46384# a_2063_45854# 0.406382f
C1292 a_8696_44636# a_17478_45572# 0.185985f
C1293 a_2324_44458# a_949_44458# 0.323116f
C1294 a_11823_42460# VDD 4.44574f
C1295 a_n1613_43370# a_33_46660# 0.599895f
C1296 a_22469_39537# a_22609_37990# 0.490939f
C1297 a_15095_43370# a_14955_43396# 0.130374f
C1298 a_n97_42460# a_n1853_43023# 0.151542f
C1299 a_3090_45724# a_9145_43396# 0.189557f
C1300 w_1575_34946# a_n1630_35242# 3.10971f
C1301 a_3232_43370# a_1423_45028# 0.396815f
C1302 a_11901_46660# a_12469_46902# 0.175891f
C1303 a_10835_43094# a_10796_42968# 0.671797f
C1304 a_n2293_45010# a_895_43940# 0.283316f
C1305 a_n971_45724# a_3065_45002# 0.220337f
C1306 a_6151_47436# DATA[5] 0.19492f
C1307 a_9313_45822# VDD 0.5747f
C1308 a_4185_45028# a_4958_30871# 0.121495f
C1309 a_n913_45002# a_12281_43396# 0.28203f
C1310 a_13259_45724# a_22400_42852# 0.34531f
C1311 a_18429_43548# VDD 0.163446f
C1312 a_n2956_38680# a_n4209_38502# 0.235751f
C1313 a_15493_43396# a_15493_43940# 0.188034f
C1314 a_20205_31679# a_20447_31679# 9.01329f
C1315 a_n1079_45724# VDD 0.172275f
C1316 a_4883_46098# a_n881_46662# 0.193691f
C1317 a_7754_38470# a_8530_39574# 0.143675f
C1318 a_n3690_39616# VDD 0.358567f
C1319 a_12549_44172# a_4190_30871# 0.270972f
C1320 a_7705_45326# VDD 0.211554f
C1321 a_n1991_42858# a_n1641_43230# 0.229804f
C1322 a_n2840_42826# a_n3674_39304# 0.16082f
C1323 a_n2157_42858# a_n1076_43230# 0.102325f
C1324 a_16137_43396# a_16414_43172# 0.179708f
C1325 a_5111_44636# a_5891_43370# 0.702087f
C1326 a_1423_45028# a_8975_43940# 0.331942f
C1327 en_comp a_n2293_43922# 0.412872f
C1328 a_765_45546# a_1176_45822# 0.241847f
C1329 a_13059_46348# a_3483_46348# 0.319214f
C1330 a_2982_43646# VDD 1.40372f
C1331 a_n784_42308# a_7174_31319# 1.93626f
C1332 a_5837_42852# VDD 0.1774f
C1333 a_3483_46348# a_13556_45296# 0.375978f
C1334 a_1138_42852# a_1307_43914# 0.123153f
C1335 a_5937_45572# a_5205_44484# 0.481405f
C1336 a_4646_46812# a_7640_43914# 0.183308f
C1337 a_n2293_46634# a_14673_44172# 0.100552f
C1338 a_n1177_43370# a_n1352_43396# 0.233657f
C1339 a_n2129_43609# a_n2012_43396# 0.183186f
C1340 a_20273_45572# a_20623_45572# 0.219856f
C1341 a_16327_47482# a_15743_43084# 1.21037f
C1342 a_n357_42282# a_18184_42460# 0.106442f
C1343 a_13507_46334# a_15227_44166# 0.235687f
C1344 a_12861_44030# a_16388_46812# 0.11634f
C1345 C3_P_btm VDD 0.26836f
C1346 C0_dummy_N_btm C7_N_btm 0.120543f
C1347 C0_N_btm C6_N_btm 0.140033f
C1348 C1_N_btm C5_N_btm 0.128021f
C1349 C2_N_btm C4_N_btm 7.19288f
C1350 a_11967_42832# a_4958_30871# 0.239255f
C1351 a_14539_43914# VDD 0.873589f
C1352 a_19692_46634# a_20411_46873# 0.215749f
C1353 a_3080_42308# a_7174_31319# 0.22305f
C1354 a_2253_43940# VDD 0.156797f
C1355 a_17583_46090# a_17715_44484# 0.22771f
C1356 a_n1613_43370# a_n2661_45010# 0.223356f
C1357 a_n784_42308# a_5932_42308# 0.151611f
C1358 a_n755_45592# a_2713_42308# 0.243663f
C1359 a_n1899_43946# a_n984_44318# 0.118759f
C1360 a_7871_42858# VDD 0.395222f
C1361 a_n2661_45546# a_n443_42852# 0.141363f
C1362 a_1823_45246# VDD 1.7584f
C1363 a_n3420_39616# a_n3420_39072# 0.115485f
C1364 a_8696_44636# a_15861_45028# 0.26484f
C1365 a_19692_46634# a_3422_30871# 0.208985f
C1366 a_12427_45724# VDD 0.33808f
C1367 a_8128_46384# a_n1925_46634# 0.21095f
C1368 a_n1613_43370# a_171_46873# 0.11335f
C1369 a_5807_45002# a_13747_46662# 0.103485f
C1370 a_14205_43396# a_14955_43396# 0.157423f
C1371 a_13159_45002# a_13348_45260# 0.105274f
C1372 a_14309_45028# VDD 0.189806f
C1373 a_11735_46660# a_12251_46660# 0.105995f
C1374 a_3080_42308# a_5932_42308# 14.0282f
C1375 a_10518_42984# a_10796_42968# 0.118759f
C1376 a_n1177_44458# a_n1352_44484# 0.233657f
C1377 a_n3674_39768# VDD 0.398971f
C1378 a_n971_45724# a_2680_45002# 0.108251f
C1379 a_n1151_42308# a_n913_45002# 0.395136f
C1380 a_4915_47217# CLK 0.198293f
C1381 a_11031_47542# VDD 0.214104f
C1382 a_6545_47178# DATA[3] 0.178561f
C1383 a_3232_43370# a_3457_43396# 0.131408f
C1384 a_17324_43396# VDD 0.274722f
C1385 a_16327_47482# a_17970_44736# 0.219775f
C1386 a_n2438_43548# a_n2661_43370# 0.147387f
C1387 a_4646_46812# a_1423_45028# 0.415897f
C1388 a_12891_46348# a_11691_44458# 0.141379f
C1389 a_20365_43914# a_20623_43914# 0.22264f
C1390 a_10193_42453# a_20712_42282# 0.157661f
C1391 a_1184_42692# VDD 0.813074f
C1392 a_13259_45724# en_comp 0.19355f
C1393 a_n2293_45546# VDD 2.06545f
C1394 a_11599_46634# a_5807_45002# 0.303048f
C1395 a_12861_44030# a_19321_45002# 0.10527f
C1396 a_7754_40130# a_11206_38545# 0.736866f
C1397 a_n3565_39590# VDD 1.26658f
C1398 a_n356_44636# a_1606_42308# 0.282657f
C1399 a_3357_43084# a_3232_43370# 0.118744f
C1400 a_6709_45028# VDD 0.390566f
C1401 a_12549_44172# a_765_45546# 0.118284f
C1402 a_n1991_42858# a_n1423_42826# 0.186387f
C1403 a_15227_44166# a_17701_42308# 0.172697f
C1404 en_comp a_n2661_43922# 0.237031f
C1405 a_7499_43078# a_11750_44172# 0.195997f
C1406 a_765_45546# a_1208_46090# 0.134766f
C1407 a_n2956_39768# a_n4209_39590# 0.334714f
C1408 a_22959_42860# a_14097_32519# 0.166017f
C1409 a_2896_43646# VDD 0.208317f
C1410 a_13059_46348# a_13249_42308# 0.306398f
C1411 a_12861_44030# a_18184_42460# 0.266953f
C1412 a_768_44030# a_1307_43914# 1.13357f
C1413 a_5732_46660# VDD 0.277366f
C1414 a_5193_42852# VDD 0.187605f
C1415 a_3483_46348# a_9482_43914# 0.130172f
C1416 a_5937_45572# a_6431_45366# 0.129839f
C1417 a_13661_43548# a_11967_42832# 0.165876f
C1418 a_4791_45118# a_4883_46098# 0.135093f
C1419 a_12861_44030# a_15811_47375# 0.144648f
C1420 a_11967_42832# a_10835_43094# 0.263495f
C1421 a_20107_45572# a_20623_45572# 0.103168f
C1422 a_20273_45572# a_20841_45814# 0.175891f
C1423 a_526_44458# a_n356_44636# 0.142971f
C1424 a_18799_45938# VDD 0.132317f
C1425 a_12861_44030# a_13059_46348# 0.504219f
C1426 C4_P_btm VDD 0.265463f
C1427 C0_dummy_N_btm C6_N_btm 0.120464f
C1428 C2_N_btm C3_N_btm 5.64696f
C1429 C0_N_btm C5_N_btm 0.138736f
C1430 C1_N_btm C4_N_btm 0.128692f
C1431 a_18429_43548# a_16823_43084# 0.130506f
C1432 a_16112_44458# VDD 0.182397f
C1433 a_19692_46634# a_20107_46660# 0.126737f
C1434 a_1443_43940# VDD 0.144342f
C1435 a_n1331_43914# a_n1549_44318# 0.209641f
C1436 a_n3674_38216# a_n3420_38528# 0.152701f
C1437 a_7227_42852# VDD 0.254613f
C1438 a_n452_45724# a_n356_45724# 0.318161f
C1439 a_1138_42852# VDD 0.397518f
C1440 a_2124_47436# a_584_46384# 0.220021f
C1441 a_n1741_47186# a_4915_47217# 0.128899f
C1442 a_11962_45724# VDD 0.210594f
C1443 a_n1613_43370# a_n133_46660# 0.347805f
C1444 a_22469_39537# a_22609_38406# 0.198764f
C1445 a_n4318_39304# a_n3674_39304# 2.9537f
C1446 a_7499_43078# a_5891_43370# 1.00892f
C1447 a_n2438_43548# a_n2157_46122# 0.270054f
C1448 a_11813_46116# a_11901_46660# 0.211542f
C1449 a_13507_46334# a_10809_44734# 0.603934f
C1450 a_10518_42984# a_10835_43094# 0.102355f
C1451 a_n4318_39768# VDD 0.469044f
C1452 a_11599_46634# a_20107_45572# 0.246047f
C1453 a_3483_46348# a_4419_46090# 0.218073f
C1454 a_13747_46662# a_14495_45572# 0.288916f
C1455 a_n1151_42308# a_n1059_45260# 0.16984f
C1456 a_9863_47436# VDD 0.207794f
C1457 a_526_44458# a_3823_42558# 0.183187f
C1458 a_375_42282# a_n1557_42282# 0.450989f
C1459 a_10193_42453# a_5342_30871# 0.151919f
C1460 a_17499_43370# VDD 0.453381f
C1461 a_16327_47482# a_17767_44458# 0.269619f
C1462 a_9290_44172# a_7499_43078# 0.597117f
C1463 a_1576_42282# VDD 0.26017f
C1464 a_20205_31679# a_19963_31679# 9.023429f
C1465 a_n2956_38216# VDD 0.484692f
C1466 a_10227_46804# a_12549_44172# 0.360691f
C1467 a_n4334_39616# VDD 0.385881f
C1468 a_7754_40130# VDAC_P 0.334598f
C1469 VDAC_Pi a_6886_37412# 0.259481f
C1470 a_5937_45572# a_6453_43914# 0.144397f
C1471 a_7229_43940# VDD 0.821851f
C1472 a_11453_44696# a_12741_44636# 1.02327f
C1473 a_n1741_47186# a_10809_44734# 0.332771f
C1474 a_n2157_42858# a_n1641_43230# 0.110532f
C1475 a_16922_45042# a_18494_42460# 0.242236f
C1476 a_7499_43078# a_10807_43548# 0.119721f
C1477 a_18315_45260# a_18587_45118# 0.13675f
C1478 a_10193_42453# a_743_42282# 1.1645f
C1479 a_3357_43084# a_3080_42308# 0.233522f
C1480 a_12861_44030# a_19778_44110# 0.113118f
C1481 a_12549_44172# a_1307_43914# 1.82879f
C1482 a_5907_46634# VDD 0.341121f
C1483 a_4649_42852# VDD 0.194775f
C1484 a_5937_45572# a_6171_45002# 0.206948f
C1485 a_12549_44172# a_18579_44172# 0.154956f
C1486 a_n1741_47186# a_n881_46662# 0.179671f
C1487 a_n4209_38216# a_n3565_38216# 6.80743f
C1488 a_n2293_46634# a_4646_46812# 0.135642f
C1489 a_5807_45002# a_5257_43370# 0.683815f
C1490 C5_P_btm VDD 0.267489f
C1491 EN_VIN_BSTR_P VIN_P 1.41696f
C1492 C0_N_btm C4_N_btm 0.138884f
C1493 C0_dummy_N_btm C5_N_btm 0.11443f
C1494 C1_N_btm C3_N_btm 7.40325f
C1495 a_16137_43396# a_743_42282# 0.183525f
C1496 a_413_45260# a_n2661_44458# 0.69469f
C1497 a_19692_46634# a_20556_43646# 0.118928f
C1498 a_n2312_38680# a_n2956_38680# 6.25577f
C1499 a_11453_44696# a_16375_45002# 0.104273f
C1500 a_11691_44458# a_14673_44172# 0.371587f
C1501 a_1241_43940# VDD 0.162129f
C1502 a_768_44030# VDD 1.53454f
C1503 a_n1899_43946# a_n1549_44318# 0.218775f
C1504 a_n2065_43946# a_n984_44318# 0.102325f
C1505 a_5755_42852# VDD 0.179985f
C1506 a_n755_45592# a_997_45618# 0.133124f
C1507 a_1176_45822# VDD 0.781481f
C1508 a_n237_47217# a_n1151_42308# 0.63407f
C1509 a_1239_39587# a_1736_39587# 0.105143f
C1510 a_n2293_46634# a_14021_43940# 0.202404f
C1511 a_11652_45724# VDD 0.155048f
C1512 a_n881_46662# a_n743_46660# 0.527182f
C1513 a_n1613_43370# a_n2438_43548# 1.04064f
C1514 VDAC_N EN_VIN_BSTR_N 0.341021f
C1515 a_22521_39511# a_22609_37990# 0.333805f
C1516 a_13017_45260# a_13159_45002# 0.160415f
C1517 a_n2438_43548# a_n2293_46098# 0.409291f
C1518 a_11735_46660# a_11901_46660# 0.579036f
C1519 a_13661_43548# a_3483_46348# 0.381471f
C1520 a_3539_42460# a_3318_42354# 0.161793f
C1521 a_n2293_45010# a_453_43940# 0.181603f
C1522 a_413_45260# a_19237_31679# 0.119197f
C1523 a_13259_45724# a_13667_43396# 0.160676f
C1524 a_7845_44172# VDD 0.11772f
C1525 a_3483_46348# a_4185_45028# 0.430982f
C1526 a_13747_46662# a_13249_42308# 0.134714f
C1527 a_4915_47217# DATA[5] 0.121371f
C1528 a_9067_47204# VDD 0.47483f
C1529 a_n2293_43922# a_n2472_43914# 0.189122f
C1530 a_8975_43940# a_9028_43914# 0.184602f
C1531 a_10057_43914# a_9672_43914# 0.143523f
C1532 a_11823_42460# a_12089_42308# 0.335983f
C1533 a_16759_43396# VDD 0.191873f
C1534 a_5937_45572# a_8746_45002# 0.121678f
C1535 a_19321_45002# a_16922_45042# 0.493823f
C1536 a_526_44458# a_3316_45546# 0.128261f
C1537 a_768_44030# a_11827_44484# 0.831344f
C1538 a_17124_42282# a_17303_42282# 0.172579f
C1539 a_20269_44172# a_20365_43914# 0.419086f
C1540 a_1067_42314# VDD 0.128996f
C1541 a_9290_44172# a_n2661_43370# 0.185465f
C1542 a_3090_45724# a_9313_44734# 2.43867f
C1543 a_11525_45546# a_11682_45822# 0.18824f
C1544 a_n2472_45546# VDD 0.290266f
C1545 a_12861_44030# a_13747_46662# 0.139424f
C1546 a_n443_46116# a_n743_46660# 0.532861f
C1547 a_n4209_39590# VDD 2.06918f
C1548 VDAC_Pi a_5700_37509# 2.20213f
C1549 a_7754_40130# a_8912_37509# 1.81084f
C1550 a_10193_42453# a_20193_45348# 0.305022f
C1551 a_n863_45724# a_n356_44636# 0.301674f
C1552 a_5937_45572# a_5663_43940# 0.177912f
C1553 a_4646_46812# a_6755_46942# 0.362783f
C1554 a_3877_44458# a_6969_46634# 0.101189f
C1555 a_n1853_43023# a_n1991_42858# 0.237526f
C1556 a_7499_43078# a_10949_43914# 0.152939f
C1557 a_17517_44484# VDD 2.99662f
C1558 a_22223_42860# a_22400_42852# 0.154104f
C1559 a_18989_43940# a_19006_44850# 0.168452f
C1560 a_12861_44030# a_18911_45144# 0.169f
C1561 a_5167_46660# VDD 0.203378f
C1562 a_9803_42558# a_9885_42558# 0.171361f
C1563 a_n784_42308# a_13258_32519# 0.140549f
C1564 a_18184_42460# a_15743_43084# 0.182123f
C1565 a_5937_45572# a_3232_43370# 0.662525f
C1566 a_8199_44636# a_6171_45002# 0.163434f
C1567 a_12861_44030# a_11599_46634# 0.169929f
C1568 a_n4209_38216# a_n4334_38304# 0.253307f
C1569 a_n2267_43396# a_n1352_43396# 0.124988f
C1570 a_n2129_43609# a_n447_43370# 0.119518f
C1571 a_3483_46348# a_11967_42832# 0.264293f
C1572 a_20107_45572# a_20273_45572# 0.667378f
C1573 a_19256_45572# VDD 0.27151f
C1574 a_1983_46706# a_n2661_46098# 0.147223f
C1575 C6_P_btm VDD 0.210613f
C1576 a_n923_35174# VIN_P 1.547f
C1577 C0_N_btm C3_N_btm 0.409996f
C1578 C1_N_btm C2_N_btm 5.0586f
C1579 C0_dummy_N_btm C4_N_btm 0.113746f
C1580 a_19692_46634# a_743_42282# 0.150479f
C1581 a_3232_43370# a_11691_44458# 0.251483f
C1582 a_13720_44458# VDD 0.202097f
C1583 a_n2312_38680# a_n2956_39304# 5.96956f
C1584 a_5883_43914# a_5891_43370# 0.216958f
C1585 SMPL_ON_N a_413_45260# 0.199669f
C1586 a_9290_44172# a_10809_44734# 0.239594f
C1587 a_3090_45724# a_2711_45572# 0.555348f
C1588 a_12549_44172# VDD 3.08339f
C1589 a_n1899_43946# a_n1331_43914# 0.171939f
C1590 a_n4318_38216# a_n3420_38528# 0.31769f
C1591 a_5111_42852# VDD 0.178652f
C1592 a_n3674_38680# a_n4064_38528# 0.557806f
C1593 a_1208_46090# VDD 0.178097f
C1594 a_n746_45260# a_n1151_42308# 0.116939f
C1595 a_n2109_47186# a_4915_47217# 0.352259f
C1596 a_22959_43948# a_17538_32519# 0.168682f
C1597 a_16855_45546# a_8696_44636# 0.112262f
C1598 a_11525_45546# VDD 0.133093f
C1599 a_n1613_43370# a_n743_46660# 0.521102f
C1600 a_n881_46662# a_n1021_46688# 0.15991f
C1601 VDAC_P EN_VIN_BSTR_P 0.339793f
C1602 a_14358_43442# a_14205_43396# 0.163543f
C1603 a_9803_43646# a_10341_43396# 0.11445f
C1604 a_14579_43548# a_15095_43370# 0.109081f
C1605 a_n357_42282# a_11967_42832# 0.153035f
C1606 a_6171_45002# a_16751_45260# 0.104212f
C1607 a_n2017_45002# a_n2293_42834# 0.28698f
C1608 a_n743_46660# a_n2293_46098# 0.213418f
C1609 a_11735_46660# a_11813_46116# 0.162547f
C1610 a_13507_46334# a_6945_45028# 0.187229f
C1611 a_10083_42826# a_10518_42984# 0.234322f
C1612 a_413_45260# a_22959_44484# 0.202222f
C1613 a_n2267_44484# a_n1352_44484# 0.118759f
C1614 a_7542_44172# VDD 0.412456f
C1615 a_n746_45260# a_327_44734# 0.256943f
C1616 a_13661_43548# a_13249_42308# 0.486588f
C1617 a_6575_47204# VDD 1.32036f
C1618 a_20193_45348# a_14021_43940# 0.118757f
C1619 a_10193_42453# a_5534_30871# 0.136243f
C1620 a_16977_43638# VDD 0.206333f
C1621 a_4190_30871# C10_P_btm 0.446355f
C1622 a_8199_44636# a_8746_45002# 0.680077f
C1623 a_12549_44172# a_11827_44484# 1.40268f
C1624 a_17124_42282# a_4958_30871# 0.20224f
C1625 en_comp a_22400_42852# 0.730145f
C1626 a_n1630_35242# VDD 3.16282f
C1627 a_n2661_45546# VDD 0.733118f
C1628 a_12861_44030# a_13661_43548# 0.8566f
C1629 VDAC_Pi a_5088_37509# 0.391059f
C1630 a_7754_40130# VDAC_N 0.434929f
C1631 a_n745_45366# a_n467_45028# 0.110406f
C1632 a_3357_43084# a_5111_44636# 0.318002f
C1633 a_5205_44484# VDD 0.508148f
C1634 a_3877_44458# a_6755_46942# 0.388535f
C1635 a_n1741_47186# a_6945_45028# 2.51584f
C1636 a_n2157_42858# a_n1991_42858# 0.905962f
C1637 a_10227_46804# a_15890_42674# 0.159412f
C1638 a_3537_45260# a_5891_43370# 0.359819f
C1639 a_7499_43078# a_10729_43914# 0.23002f
C1640 a_14537_43396# a_14539_43914# 0.135541f
C1641 a_17061_44734# VDD 0.17647f
C1642 a_3422_30871# EN_VIN_BSTR_N 0.182769f
C1643 a_n2442_46660# a_n4315_30879# 0.361271f
C1644 a_5534_30871# a_n784_42308# 9.92256f
C1645 a_n913_45002# a_n97_42460# 0.109647f
C1646 a_10193_42453# a_4190_30871# 0.305842f
C1647 a_1427_43646# VDD 0.19291f
C1648 a_n2293_46634# a_5111_44636# 0.130609f
C1649 a_n971_45724# a_n699_43396# 0.139047f
C1650 a_5385_46902# VDD 0.203316f
C1651 a_n356_44636# a_2982_43646# 0.434193f
C1652 a_1307_43914# a_3935_42891# 0.318189f
C1653 a_3483_46348# a_13017_45260# 0.51131f
C1654 a_8199_44636# a_3232_43370# 0.32342f
C1655 a_n1533_46116# VDD 0.143145f
C1656 a_n1699_43638# a_n1917_43396# 0.209641f
C1657 a_4791_45118# a_4361_42308# 0.111224f
C1658 a_16327_47482# a_17324_43396# 0.216094f
C1659 a_19431_45546# VDD 0.342308f
C1660 a_13507_46334# a_15559_46634# 0.216791f
C1661 C7_P_btm VDD 0.121904f
C1662 C0_N_btm C2_N_btm 0.698973f
C1663 a_16137_43396# a_4190_30871# 0.113768f
C1664 a_n913_45002# a_742_44458# 0.302053f
C1665 a_19692_46634# a_20301_43646# 0.110092f
C1666 a_13076_44458# VDD 0.180665f
C1667 a_2063_45854# a_6472_45840# 0.545607f
C1668 a_4646_46812# a_5937_45572# 0.105447f
C1669 a_22165_42308# a_22223_42860# 0.171681f
C1670 a_2324_44458# a_15682_46116# 0.343876f
C1671 a_12891_46348# VDD 1.01428f
C1672 a_n2065_43946# a_n1549_44318# 0.110816f
C1673 a_4520_42826# VDD 0.142755f
C1674 a_12861_44030# a_11967_42832# 0.209245f
C1675 a_n357_42282# a_n755_45592# 0.664842f
C1676 a_805_46414# VDD 0.154663f
C1677 a_21076_30879# VREF 0.417978f
C1678 a_n971_45724# a_n1151_42308# 0.682801f
C1679 a_1209_47178# a_584_46384# 0.104123f
C1680 a_n2661_42834# a_n2840_42826# 0.174935f
C1681 a_n913_45002# a_10533_42308# 0.246621f
C1682 a_5742_30871# VCM 0.211981f
C1683 a_16855_45546# a_16680_45572# 0.233657f
C1684 a_15903_45785# a_16020_45572# 0.157972f
C1685 a_n2810_45028# a_n3565_38216# 0.349341f
C1686 a_11322_45546# VDD 0.370908f
C1687 a_n881_46662# a_n1925_46634# 0.467945f
C1688 a_6151_47436# a_6755_46942# 0.361724f
C1689 a_22521_39511# a_22609_38406# 0.23688f
C1690 a_22459_39145# a_22609_37990# 0.172129f
C1691 a_9803_43646# a_9885_43646# 0.171361f
C1692 a_3422_30871# COMP_P 0.208163f
C1693 a_3357_43084# a_3905_42865# 0.125186f
C1694 a_n1699_44726# a_n1917_44484# 0.209641f
C1695 a_7281_43914# VDD 0.198809f
C1696 a_n1925_46634# a_8162_45546# 0.104508f
C1697 a_n2661_46634# a_10193_42453# 0.351509f
C1698 a_5807_45002# a_13249_42308# 0.725941f
C1699 a_7903_47542# VDD 0.202868f
C1700 a_n2661_43922# a_n2840_43914# 0.171265f
C1701 a_18479_45785# a_4190_30871# 0.123942f
C1702 a_16409_43396# VDD 0.250832f
C1703 a_8199_44636# a_10193_42453# 0.236934f
C1704 a_8049_45260# a_20205_31679# 0.301209f
C1705 a_12359_47026# VDD 0.142103f
C1706 a_10193_42453# a_19511_42282# 0.133376f
C1707 a_564_42282# VDD 0.293756f
C1708 a_13259_45724# a_n913_45002# 0.142601f
C1709 a_n2810_45572# VDD 0.557886f
C1710 a_12861_44030# a_5807_45002# 0.214011f
C1711 a_7754_39964# a_5088_37509# 0.392826f
C1712 VDAC_Pi a_4338_37500# 1.92369f
C1713 a_5343_44458# a_7963_42308# 0.108654f
C1714 a_13661_43548# a_19268_43646# 0.136251f
C1715 a_6431_45366# VDD 0.203167f
C1716 a_11453_44696# a_11415_45002# 0.123733f
C1717 a_n2157_42858# a_n1853_43023# 0.290902f
C1718 a_10227_46804# a_15959_42545# 0.152289f
C1719 a_3537_45260# a_8375_44464# 0.10437f
C1720 a_7499_43078# a_10405_44172# 0.132405f
C1721 a_1423_45028# a_9838_44484# 0.254741f
C1722 a_16241_44734# VDD 0.189894f
C1723 a_3422_30871# a_11530_34132# 0.127528f
C1724 a_10227_46804# a_8746_45002# 0.117547f
C1725 a_1823_45246# a_3823_42558# 0.137565f
C1726 a_18287_44626# a_11967_42832# 0.789765f
C1727 a_n1059_45260# a_n97_42460# 0.869353f
C1728 a_n1557_42282# VDD 0.355513f
C1729 a_1823_45246# a_3503_45724# 0.295715f
C1730 a_4817_46660# VDD 0.370615f
C1731 a_1307_43914# a_3681_42891# 0.236785f
C1732 a_22400_42852# a_22821_38993# 0.136515f
C1733 a_6511_45714# a_7227_45028# 0.213161f
C1734 a_6667_45809# a_6598_45938# 0.209641f
C1735 a_8953_45546# a_5111_44636# 0.181796f
C1736 a_n2433_43396# a_n1352_43396# 0.102325f
C1737 a_n2267_43396# a_n1917_43396# 0.227165f
C1738 a_16327_47482# a_17499_43370# 0.34052f
C1739 a_18691_45572# VDD 0.191893f
C1740 C8_P_btm VDD 0.19922f
C1741 a_n1386_35608# VIN_P 0.367112f
C1742 C0_N_btm C1_N_btm 10.8764f
C1743 C0_dummy_N_btm C2_N_btm 6.66125f
C1744 a_413_45260# a_19721_31679# 0.116395f
C1745 a_12883_44458# VDD 0.263743f
C1746 a_19333_46634# a_19123_46287# 0.113955f
C1747 a_11453_44696# a_13259_45724# 0.251534f
C1748 a_n2661_44458# a_n2661_43922# 6.64988f
C1749 a_18287_44626# a_18989_43940# 0.193279f
C1750 a_18443_44721# a_18374_44850# 0.209641f
C1751 a_1307_43914# a_5663_43940# 0.11718f
C1752 a_4185_45028# a_n1925_42282# 0.638728f
C1753 a_11309_47204# VDD 0.358104f
C1754 a_n1761_44111# a_n1899_43946# 0.737653f
C1755 a_20202_43084# a_n913_45002# 0.322116f
C1756 a_472_46348# VDD 0.706547f
C1757 a_n2109_47186# a_4791_45118# 0.34446f
C1758 a_1239_47204# a_1431_47204# 0.219138f
C1759 a_375_42282# a_196_42282# 0.165785f
C1760 a_15890_42674# VDD 0.203548f
C1761 a_5742_30871# VREF_GND 0.191352f
C1762 a_1138_42852# a_n356_44636# 0.29814f
C1763 a_8199_44636# a_10057_43914# 0.113262f
C1764 a_n2956_37592# a_n4209_38216# 0.104159f
C1765 a_10490_45724# VDD 0.162001f
C1766 a_n1613_43370# a_n1925_46634# 0.33524f
C1767 a_22521_40055# a_22609_37990# 0.234448f
C1768 a_14579_43548# a_14358_43442# 0.142377f
C1769 a_3090_45724# a_8685_43396# 2.11639f
C1770 a_3232_43370# a_1307_43914# 0.14252f
C1771 a_11453_44696# a_18189_46348# 0.534507f
C1772 a_13259_45724# a_9145_43396# 0.155949f
C1773 a_n2433_44484# a_n1352_44484# 0.102355f
C1774 a_n2267_44484# a_n1917_44484# 0.212549f
C1775 a_6453_43914# VDD 0.194953f
C1776 a_n2293_46634# a_7499_43078# 0.14773f
C1777 a_n971_45724# a_413_45260# 0.937818f
C1778 a_3147_46376# a_3483_46348# 0.207919f
C1779 a_7227_47204# VDD 0.430714f
C1780 a_5342_30871# a_14113_42308# 0.203397f
C1781 a_16547_43609# VDD 0.31275f
C1782 a_8199_44636# a_10180_45724# 0.216999f
C1783 a_19692_46634# a_2437_43646# 0.293918f
C1784 a_3483_46348# a_13249_42308# 0.338396f
C1785 a_n3674_37592# VDD 0.357168f
C1786 a_13259_45724# a_n1059_45260# 0.390886f
C1787 a_n2840_45546# VDD 0.302566f
C1788 a_2063_45854# a_2107_46812# 0.214026f
C1789 a_7754_38636# a_7754_38470# 0.296258f
C1790 VDAC_Pi a_3726_37500# 1.17174f
C1791 a_n2302_40160# VDD 0.428934f
C1792 a_n1059_45260# a_n467_45028# 0.229142f
C1793 a_6171_45002# VDD 0.441339f
C1794 a_12465_44636# a_12741_44636# 0.914049f
C1795 a_2711_45572# a_15493_43940# 0.128282f
C1796 a_10227_46804# a_15803_42450# 0.296174f
C1797 a_n2017_45002# a_n2293_43922# 0.654835f
C1798 a_14673_44172# VDD 0.381917f
C1799 w_11334_34010# a_18194_35068# 0.796644f
C1800 a_18248_44752# a_11967_42832# 0.500539f
C1801 a_n2017_45002# a_n97_42460# 0.169401f
C1802 a_13059_46348# a_11823_42460# 0.256727f
C1803 a_4955_46873# VDD 0.467566f
C1804 a_13259_45724# a_15599_45572# 0.205417f
C1805 a_6472_45840# a_7227_45028# 0.208286f
C1806 a_12861_44030# a_13487_47204# 0.127147f
C1807 a_n2267_43396# a_n1699_43638# 0.179796f
C1808 a_16327_47482# a_16759_43396# 0.152273f
C1809 a_18909_45814# VDD 0.205795f
C1810 a_18597_46090# a_15227_44166# 0.150202f
C1811 C9_P_btm VDD 0.345685f
C1812 C0_dummy_N_btm C1_N_btm 1.2494f
C1813 a_10193_42453# a_18579_44172# 0.12582f
C1814 a_12607_44458# VDD 0.188171f
C1815 a_14180_46812# a_14513_46634# 0.253235f
C1816 a_18248_44752# a_18989_43940# 0.207562f
C1817 a_5111_44636# a_8333_44056# 0.280148f
C1818 a_11827_44484# a_14673_44172# 0.150125f
C1819 a_8103_44636# a_8375_44464# 0.13675f
C1820 a_4185_45028# a_526_44458# 0.162857f
C1821 a_12465_44636# a_413_45260# 0.28925f
C1822 a_n755_45592# a_1755_42282# 1.52791f
C1823 a_n2065_43946# a_n1899_43946# 0.614122f
C1824 a_3681_42891# VDD 0.223661f
C1825 a_n1099_45572# a_n755_45592# 0.193775f
C1826 a_310_45028# a_n357_42282# 0.113929f
C1827 a_n746_45260# a_175_44278# 0.159759f
C1828 a_376_46348# VDD 0.116284f
C1829 a_n971_45724# a_2905_45572# 0.118495f
C1830 a_n3565_39590# a_n4209_39304# 5.4667f
C1831 a_11967_42832# a_15743_43084# 0.180938f
C1832 a_15959_42545# VDD 0.19373f
C1833 a_n443_42852# a_5111_44636# 0.584506f
C1834 a_15903_45785# a_15861_45028# 0.232345f
C1835 a_8746_45002# VDD 0.970181f
C1836 a_22459_39145# a_22609_38406# 0.12318f
C1837 a_11787_45002# a_11963_45334# 0.185422f
C1838 a_6755_46942# a_15227_44166# 0.288173f
C1839 a_3357_43084# a_2998_44172# 0.119142f
C1840 a_n2267_44484# a_n1699_44726# 0.172319f
C1841 a_20202_43084# a_19987_42826# 0.177726f
C1842 a_5663_43940# VDD 0.133666f
C1843 a_16327_47482# a_19256_45572# 0.235006f
C1844 a_n1151_42308# a_n2661_45010# 0.155007f
C1845 a_6851_47204# VDD 0.287724f
C1846 a_16243_43396# VDD 0.39865f
C1847 a_8016_46348# a_10193_42453# 0.125497f
C1848 a_n2293_46634# a_n2661_43370# 2.59564f
C1849 a_3483_46348# a_13904_45546# 0.125708f
C1850 a_8953_45546# a_7499_43078# 0.108436f
C1851 a_5937_45572# a_9049_44484# 0.311862f
C1852 a_n327_42558# VDD 0.198414f
C1853 a_10490_45724# a_10907_45822# 0.229517f
C1854 a_n971_45724# a_104_43370# 0.156156f
C1855 a_n237_47217# a_1799_45572# 0.417887f
C1856 a_6151_47436# a_n2661_46634# 0.140541f
C1857 a_16327_47482# a_12549_44172# 0.123271f
C1858 VDAC_Ni a_3754_38470# 0.911632f
C1859 a_n4064_40160# VDD 2.37253f
C1860 a_3232_43370# VDD 2.96597f
C1861 a_3422_30871# EN_VIN_BSTR_P 0.182769f
C1862 SMPL_ON_P a_n1838_35608# 0.399535f
C1863 w_11334_34010# EN_VIN_BSTR_N 3.99277f
C1864 a_4905_42826# VDD 0.439034f
C1865 a_167_45260# a_1848_45724# 0.359783f
C1866 a_4651_46660# VDD 0.457722f
C1867 a_5934_30871# a_5742_30871# 16.7261f
C1868 a_6453_43914# a_n2661_42282# 0.122766f
C1869 a_n3674_37592# a_n4064_37440# 0.651412f
C1870 a_6472_45840# a_6598_45938# 0.178024f
C1871 a_6511_45714# a_6667_45809# 0.113977f
C1872 a_n1151_42308# a_4883_46098# 0.407909f
C1873 a_n2497_47436# a_n1613_43370# 0.402561f
C1874 a_n2433_43396# a_n1917_43396# 0.108815f
C1875 a_16327_47482# a_16977_43638# 0.15941f
C1876 a_18341_45572# VDD 0.2432f
C1877 a_6151_47436# a_765_45546# 0.191559f
C1878 a_10227_46804# a_19692_46634# 0.239326f
C1879 a_12861_44030# a_14180_46812# 0.238709f
C1880 C10_P_btm VDD 2.40001f
C1881 C0_dummy_N_btm C0_N_btm 7.61701f
C1882 a_10341_43396# a_22591_43396# 0.172197f
C1883 a_n2661_42282# a_n3674_37592# 0.12829f
C1884 a_4791_45118# a_5932_42308# 0.212275f
C1885 a_8975_43940# VDD 0.257588f
C1886 a_2982_43646# a_17303_42282# 0.139588f
C1887 a_8103_44636# a_7640_43914# 0.101633f
C1888 a_18287_44626# a_18443_44721# 0.10279f
C1889 a_18248_44752# a_18374_44850# 0.170059f
C1890 a_1307_43914# a_5013_44260# 0.358053f
C1891 a_3483_46348# a_n1925_42282# 0.536704f
C1892 a_4791_45118# a_1423_45028# 0.721318f
C1893 a_n755_45592# a_1606_42308# 0.104938f
C1894 a_n2065_43946# a_n1761_44111# 0.617556f
C1895 a_n3674_38680# a_n3565_38502# 0.128677f
C1896 a_2905_42968# VDD 0.142081f
C1897 a_20820_30879# VREF 0.195875f
C1898 a_n1076_46494# VDD 0.294742f
C1899 a_1209_47178# a_1239_47204# 0.264529f
C1900 a_n237_47217# a_2063_45854# 0.947844f
C1901 a_22223_43948# a_14401_32519# 0.157135f
C1902 a_15803_42450# VDD 0.448709f
C1903 a_15765_45572# a_16680_45572# 0.118759f
C1904 a_10193_42453# VDD 2.18892f
C1905 a_4915_47217# a_6755_46942# 0.260675f
C1906 a_22521_40055# a_22609_38406# 0.1922f
C1907 a_22469_40625# a_22609_37990# 0.130478f
C1908 a_9145_43396# a_15095_43370# 0.213415f
C1909 a_8696_44636# a_n2661_44458# 1.37553f
C1910 a_8128_46384# a_8349_46414# 0.101217f
C1911 a_9127_43156# a_8952_43230# 0.234322f
C1912 a_n2433_44484# a_n1917_44484# 0.113784f
C1913 a_5495_43940# VDD 0.173477f
C1914 a_1823_45246# a_4704_46090# 0.164557f
C1915 a_11453_44696# a_8696_44636# 2.67247f
C1916 a_16327_47482# a_19431_45546# 0.344862f
C1917 a_13747_46662# a_11823_42460# 0.521845f
C1918 a_6491_46660# VDD 0.436756f
C1919 a_n1059_45260# a_15095_43370# 0.108103f
C1920 a_9290_44172# a_13070_42354# 0.140007f
C1921 a_16137_43396# VDD 0.483673f
C1922 a_12549_44172# a_20567_45036# 0.176249f
C1923 a_8016_46348# a_10180_45724# 0.259851f
C1924 a_8953_45546# a_8568_45546# 0.136365f
C1925 a_9313_44734# a_10341_43396# 0.175125f
C1926 a_14955_43940# a_15493_43940# 0.110232f
C1927 a_n784_42308# VDD 0.597561f
C1928 a_13904_45546# a_13249_42308# 0.13587f
C1929 a_n971_45724# a_n97_42460# 0.581616f
C1930 a_15811_47375# a_15928_47570# 0.161235f
C1931 a_n4334_40480# VDD 0.390668f
C1932 a_10193_42453# a_11827_44484# 0.121679f
C1933 a_n913_45002# a_n967_45348# 1.00127f
C1934 a_n2810_45028# a_n2956_37592# 6.13705f
C1935 a_5691_45260# VDD 0.205518f
C1936 a_n1151_42308# a_11387_46155# 0.195225f
C1937 a_2711_45572# a_11341_43940# 1.54309f
C1938 a_16922_45042# a_17719_45144# 0.22253f
C1939 a_10227_46804# a_15486_42560# 0.227612f
C1940 w_11334_34010# a_11530_34132# 37.743603f
C1941 a_n443_42852# a_685_42968# 0.104532f
C1942 a_3080_42308# VDD 0.849483f
C1943 a_n2293_46634# a_3537_45260# 0.155982f
C1944 a_4646_46812# VDD 2.53408f
C1945 a_1307_43914# a_1847_42826# 0.428505f
C1946 a_9313_44734# a_n97_42460# 1.76217f
C1947 a_6472_45840# a_6667_45809# 0.215953f
C1948 a_n443_42852# a_7499_43078# 0.375366f
C1949 a_15227_44166# a_11691_44458# 0.443265f
C1950 a_13717_47436# a_12861_44030# 0.319645f
C1951 a_n1435_47204# a_13487_47204# 0.135076f
C1952 a_n3420_38528# a_n4064_37984# 7.35343f
C1953 a_n2129_43609# a_n2267_43396# 0.230013f
C1954 a_18479_45785# VDD 0.536075f
C1955 a_12861_44030# a_14035_46660# 0.153051f
C1956 a_18479_47436# a_15227_44166# 0.199537f
C1957 a_21589_35634# VDD 0.525446f
C1958 a_10057_43914# VDD 0.399284f
C1959 a_18834_46812# a_18285_46348# 0.144972f
C1960 a_13885_46660# a_14513_46634# 0.101344f
C1961 a_21195_42852# a_21671_42860# 0.177876f
C1962 a_2982_43646# a_4958_30871# 0.136637f
C1963 a_5343_44458# a_5891_43370# 1.06553f
C1964 a_18248_44752# a_18443_44721# 0.206455f
C1965 a_n443_42852# a_15781_43660# 0.22553f
C1966 a_14021_43940# VDD 1.60583f
C1967 a_15015_46420# a_14840_46494# 0.233657f
C1968 a_3483_46348# a_526_44458# 0.134907f
C1969 a_n1613_43370# a_3357_43084# 0.228593f
C1970 a_9804_47204# VDD 0.410522f
C1971 a_1606_42308# a_2351_42308# 0.191324f
C1972 a_n1099_45572# a_310_45028# 0.333219f
C1973 a_n2293_46098# a_3357_43084# 0.16657f
C1974 a_n901_46420# VDD 0.518805f
C1975 a_21076_30879# EN_OFFSET_CAL 0.2809f
C1976 a_n237_47217# a_584_46384# 0.645142f
C1977 a_n971_45724# a_2553_47502# 0.23907f
C1978 a_15764_42576# VDD 0.258303f
C1979 a_8953_45546# a_5883_43914# 0.262126f
C1980 a_16333_45814# a_16115_45572# 0.209641f
C1981 a_n443_46116# a_2813_43396# 0.124521f
C1982 en_comp a_1177_38525# 0.205977f
C1983 a_10180_45724# VDD 0.336512f
C1984 a_n1613_43370# a_n2293_46634# 0.103089f
C1985 a_22545_38993# a_22821_38993# 0.235701f
C1986 a_22521_39511# a_22469_39537# 1.02751f
C1987 a_7754_39632# VDD 0.205733f
C1988 a_9145_43396# a_14205_43396# 0.13322f
C1989 a_5111_44636# a_1307_43914# 0.114933f
C1990 a_2711_45572# a_n97_42460# 0.137121f
C1991 a_n2129_44697# a_n2267_44484# 0.698671f
C1992 a_5013_44260# VDD 0.198233f
C1993 a_4791_45118# a_3357_43084# 0.144996f
C1994 a_1823_45246# a_4419_46090# 0.340207f
C1995 a_16327_47482# a_18691_45572# 0.162157f
C1996 a_13661_43548# a_11823_42460# 0.116839f
C1997 a_6545_47178# VDD 0.386368f
C1998 a_17517_44484# a_20640_44752# 0.54753f
C1999 a_5111_44636# a_9396_43370# 0.203348f
C2000 a_15227_44166# a_2437_43646# 0.167451f
C2001 a_12549_44172# a_18494_42460# 0.331306f
C2002 a_8199_44636# a_7499_43078# 0.859274f
C2003 a_526_44458# a_n357_42282# 0.220537f
C2004 a_19692_46634# VDD 2.53528f
C2005 a_15493_43396# a_19478_44306# 0.154347f
C2006 a_196_42282# VDD 0.291844f
C2007 a_3090_45724# a_5891_43370# 0.166094f
C2008 a_n971_45724# a_n447_43370# 0.113797f
C2009 a_5937_45572# a_n2661_43370# 0.202031f
C2010 a_20692_30879# VDD 0.499615f
C2011 a_584_46384# a_1123_46634# 0.370049f
C2012 a_n4315_30879# VDD 4.0486f
C2013 a_14401_32519# a_10341_43396# 0.133035f
C2014 a_16147_45260# a_1307_43914# 0.150161f
C2015 a_4927_45028# VDD 0.159822f
C2016 a_12465_44636# a_11415_45002# 0.375509f
C2017 a_n1151_42308# a_11133_46155# 0.162011f
C2018 a_1423_45028# a_6298_44484# 0.103777f
C2019 a_13556_45296# a_15004_44636# 0.127354f
C2020 a_16922_45042# a_17613_45144# 0.10967f
C2021 a_10227_46804# a_15051_42282# 0.361922f
C2022 a_12861_44030# a_13527_45546# 0.274077f
C2023 a_3090_45724# a_9290_44172# 0.196232f
C2024 a_4699_43561# VDD 0.262218f
C2025 a_768_44030# a_13556_45296# 0.267809f
C2026 a_167_45260# a_n755_45592# 1.02724f
C2027 a_12861_44030# a_16922_45042# 0.120012f
C2028 a_11415_45002# a_2711_45572# 0.337384f
C2029 a_3877_44458# VDD 0.786903f
C2030 a_6123_31319# a_5742_30871# 0.106954f
C2031 a_22400_42852# a_22459_39145# 0.242947f
C2032 a_19321_45002# a_17517_44484# 0.264473f
C2033 a_3483_46348# a_8953_45002# 0.121322f
C2034 a_6472_45840# a_6511_45714# 0.781352f
C2035 a_13381_47204# a_13487_47204# 0.152045f
C2036 a_2112_39137# a_2113_38308# 0.479143f
C2037 a_n2433_43396# a_n2267_43396# 0.756435f
C2038 a_18175_45572# VDD 0.38478f
C2039 a_19864_35138# VDD 0.332629f
C2040 C3_P_btm C3_N_btm 2.90968f
C2041 a_6293_42852# a_5755_42852# 0.114235f
C2042 a_11823_42460# a_11967_42832# 0.573139f
C2043 a_4185_45028# a_2982_43646# 0.243496f
C2044 a_10440_44484# VDD 0.159539f
C2045 a_13885_46660# a_14180_46812# 0.150851f
C2046 a_17609_46634# a_18285_46348# 0.115413f
C2047 a_14209_32519# a_14097_32519# 10.7606f
C2048 a_18248_44752# a_18287_44626# 0.633819f
C2049 a_1307_43914# a_3905_42865# 0.224019f
C2050 a_3147_46376# a_526_44458# 0.352f
C2051 a_8128_46384# VDD 0.403575f
C2052 a_1847_42826# VDD 0.527555f
C2053 a_12465_44636# a_n2661_43922# 0.17969f
C2054 a_n863_45724# a_n755_45592# 1.76733f
C2055 a_13259_45724# a_2711_45572# 1.26722f
C2056 a_13661_43548# a_14539_43914# 0.193767f
C2057 a_n1641_46494# VDD 0.226065f
C2058 a_n1741_47186# a_n1151_42308# 2.98024f
C2059 a_n2109_47186# a_3785_47178# 0.190973f
C2060 a_n971_45724# a_2063_45854# 0.164981f
C2061 a_n746_45260# a_584_46384# 0.491308f
C2062 a_n2661_42282# a_3080_42308# 0.161683f
C2063 a_20512_43084# a_10341_43396# 0.758407f
C2064 a_15486_42560# VDD 0.275297f
C2065 a_5937_45572# a_5883_43914# 0.454323f
C2066 a_10809_44734# a_11691_44458# 0.354084f
C2067 a_15765_45572# a_16115_45572# 0.20669f
C2068 a_15599_45572# a_16680_45572# 0.102355f
C2069 a_2324_44458# a_n2661_44458# 0.134417f
C2070 a_10053_45546# VDD 0.150582f
C2071 a_12549_44172# a_19321_45002# 0.238866f
C2072 a_22521_39511# a_22821_38993# 0.112629f
C2073 a_19862_44208# a_20922_43172# 0.164553f
C2074 a_8128_46384# a_7920_46348# 0.197919f
C2075 a_n881_46662# a_5937_45572# 0.195456f
C2076 a_n97_42460# a_5934_30871# 0.221607f
C2077 a_n2433_44484# a_n2267_44484# 0.730194f
C2078 a_5244_44056# VDD 0.146618f
C2079 a_16327_47482# a_18909_45814# 0.16767f
C2080 a_4915_47217# a_2437_43646# 0.114772f
C2081 a_2698_46116# a_2804_46116# 0.313533f
C2082 a_6151_47436# VDD 4.39915f
C2083 a_4007_47204# DATA[2] 0.337596f
C2084 a_5342_30871# a_14456_42282# 0.160195f
C2085 a_5883_43914# a_8333_44056# 0.152643f
C2086 a_n913_45002# a_14579_43548# 0.239851f
C2087 a_n971_45724# a_n2661_42834# 0.165951f
C2088 a_n2438_43548# a_n2293_42834# 0.138621f
C2089 a_8199_44636# a_8568_45546# 0.141772f
C2090 a_19466_46812# VDD 0.664497f
C2091 a_19328_44172# a_19478_44306# 0.188181f
C2092 a_n473_42460# VDD 0.27195f
C2093 a_11823_42460# a_15143_45578# 0.120787f
C2094 a_8199_44636# a_n2661_43370# 0.126664f
C2095 a_20205_31679# VDD 0.737305f
C2096 a_n1151_42308# a_n743_46660# 0.195953f
C2097 a_n4209_39304# C7_P_btm 0.184297f
C2098 a_3357_43084# a_3065_45002# 0.316449f
C2099 a_16147_45260# a_16019_45002# 0.186254f
C2100 a_5111_44636# VDD 1.28013f
C2101 a_12549_44172# a_13059_46348# 0.808395f
C2102 a_13507_46334# a_12741_44636# 0.137731f
C2103 a_n1151_42308# a_11189_46129# 0.12414f
C2104 a_13556_45296# a_13720_44458# 0.212774f
C2105 a_9482_43914# a_15004_44636# 0.34299f
C2106 a_10227_46804# a_14113_42308# 0.627404f
C2107 a_9290_44172# a_12281_43396# 0.36475f
C2108 a_22612_30879# a_20205_31679# 0.111294f
C2109 a_14539_43914# a_11967_42832# 0.512158f
C2110 a_4235_43370# VDD 0.229422f
C2111 a_n4318_38680# a_n4209_38502# 0.105064f
C2112 a_768_44030# a_9482_43914# 0.77718f
C2113 a_167_45260# a_n357_42282# 0.148401f
C2114 a_n2293_46634# a_3065_45002# 0.102991f
C2115 a_8685_42308# a_9223_42460# 0.166964f
C2116 a_22400_42852# a_22521_40055# 0.681186f
C2117 a_6194_45824# a_6511_45714# 0.102325f
C2118 a_10809_44734# a_2437_43646# 0.13907f
C2119 a_n2956_38680# VDD 0.871805f
C2120 a_n1435_47204# a_13717_47436# 0.196889f
C2121 a_n3420_38528# a_n3420_37984# 0.113087f
C2122 a_n2433_43396# a_n2129_43609# 0.283605f
C2123 a_7499_43078# a_1307_43914# 0.109806f
C2124 a_16327_47482# a_16243_43396# 0.295263f
C2125 en_comp a_22459_39145# 0.415926f
C2126 a_16147_45260# VDD 0.197706f
C2127 a_4915_47217# a_765_45546# 0.169406f
C2128 a_171_46873# a_n2661_46098# 0.168482f
C2129 a_19120_35138# VDD 0.318963f
C2130 a_n2661_45010# a_742_44458# 0.694478f
C2131 a_10334_44484# VDD 0.19332f
C2132 a_2063_45854# a_2711_45572# 0.185507f
C2133 a_13885_46660# a_14035_46660# 0.25868f
C2134 a_17609_46634# a_17829_46910# 0.111805f
C2135 a_n443_46116# a_n443_42852# 0.145452f
C2136 a_15227_44166# a_17339_46660# 0.524034f
C2137 a_17970_44736# a_18287_44626# 0.102355f
C2138 a_1307_43914# a_3600_43914# 0.153686f
C2139 a_5343_44458# a_7640_43914# 0.152634f
C2140 a_1606_42308# a_1755_42282# 0.278431f
C2141 a_791_42968# VDD 0.128737f
C2142 a_n1079_45724# a_n755_45592# 0.109544f
C2143 a_n863_45724# a_n357_42282# 0.172013f
C2144 a_380_45546# a_n1099_45572# 0.148825f
C2145 a_12741_44636# EN_OFFSET_CAL 0.230064f
C2146 a_n1423_46090# VDD 0.227012f
C2147 a_n971_45724# a_584_46384# 0.152617f
C2148 a_n4064_39616# a_n2302_39866# 0.239588f
C2149 a_n2293_43922# a_5649_42852# 1.78418f
C2150 a_15051_42282# VDD 0.461307f
C2151 a_n443_42852# a_3537_45260# 0.567413f
C2152 a_15765_45572# a_16333_45814# 0.17072f
C2153 a_3483_46348# a_16979_44734# 0.173123f
C2154 a_9049_44484# VDD 0.680993f
C2155 a_768_44030# a_13747_46662# 0.434325f
C2156 VDAC_Pi VDD 0.591846f
C2157 a_22521_39511# a_22545_38993# 0.27533f
C2158 a_22459_39145# a_22469_39537# 0.351623f
C2159 a_7754_39964# RST_Z 0.843939f
C2160 a_8685_43396# a_10341_43396# 2.41562f
C2161 a_10775_45002# a_10951_45334# 0.185422f
C2162 a_17715_44484# a_17737_43940# 0.289085f
C2163 a_n1613_43370# a_5937_45572# 0.117604f
C2164 a_8037_42858# a_8952_43230# 0.118759f
C2165 a_4905_42826# a_5267_42460# 0.146764f
C2166 a_n755_45592# a_2982_43646# 0.221452f
C2167 a_n2433_44484# a_n2129_44697# 0.130072f
C2168 a_n1059_45260# a_n1761_44111# 0.535535f
C2169 a_3905_42865# VDD 0.788273f
C2170 a_n443_46116# a_2437_43646# 0.410719f
C2171 a_765_45546# a_10809_44734# 2.52248f
C2172 a_5815_47464# VDD 0.399354f
C2173 a_n1059_45260# a_14579_43548# 0.250544f
C2174 a_9290_44172# a_11551_42558# 0.123803f
C2175 a_1307_43914# a_1756_43548# 0.267667f
C2176 a_12549_44172# a_19778_44110# 0.294084f
C2177 a_3483_46348# a_11823_42460# 0.377948f
C2178 a_8199_44636# a_8162_45546# 0.119979f
C2179 a_19333_46634# VDD 0.199048f
C2180 a_7542_44172# a_7499_43940# 0.157633f
C2181 a_n961_42308# VDD 0.24416f
C2182 a_8162_45546# a_8192_45572# 0.134163f
C2183 a_n1151_42308# a_n1021_46688# 0.105326f
C2184 a_n443_46116# a_n2661_46634# 0.121882f
C2185 a_22465_38105# VDD 1.3089f
C2186 a_n2661_45010# a_n467_45028# 0.227953f
C2187 a_5147_45002# VDD 0.574918f
C2188 a_413_45260# EN_OFFSET_CAL 0.114452f
C2189 a_12891_46348# a_13059_46348# 0.372745f
C2190 a_4791_45118# a_5937_45572# 0.151145f
C2191 a_n881_46662# a_765_45546# 0.333008f
C2192 a_n1151_42308# a_9290_44172# 0.10853f
C2193 a_20916_46384# a_19692_46634# 0.117693f
C2194 a_n2661_45010# a_n2661_43922# 0.111071f
C2195 a_9482_43914# a_13720_44458# 0.188323f
C2196 a_1423_45028# a_5343_44458# 0.128331f
C2197 a_16327_47482# a_10193_42453# 0.163668f
C2198 a_12861_44030# a_12791_45546# 0.248928f
C2199 a_22000_46634# a_20202_43084# 0.154237f
C2200 w_1575_34946# EN_VIN_BSTR_P 3.99222f
C2201 a_4093_43548# VDD 0.216874f
C2202 a_10903_43370# a_13259_45724# 0.600111f
C2203 a_12891_46348# a_13556_45296# 0.29495f
C2204 a_526_44458# a_n1925_42282# 0.213917f
C2205 a_1823_45246# a_n755_45592# 0.390511f
C2206 a_8685_42308# a_8791_42308# 0.147376f
C2207 a_n3674_37592# a_n3565_37414# 0.129086f
C2208 a_n784_42308# a_n3420_37440# 0.140549f
C2209 a_6194_45824# a_6472_45840# 0.118423f
C2210 a_8199_44636# a_3537_45260# 0.199536f
C2211 a_n2956_39304# VDD 0.455981f
C2212 a_9313_44734# a_22959_42860# 0.174475f
C2213 a_3090_45724# a_10729_43914# 0.135702f
C2214 a_11823_42460# a_11963_45334# 0.110904f
C2215 a_20202_43084# a_20512_43084# 0.130366f
C2216 en_comp a_22521_40055# 0.260972f
C2217 a_n443_46116# a_765_45546# 0.297346f
C2218 a_n2438_43548# a_2443_46660# 0.237765f
C2219 a_18194_35068# VDD 2.17116f
C2220 C0_P_btm C0_dummy_P_btm 7.61701f
C2221 a_n2956_37592# a_n4318_40392# 2.71462f
C2222 a_10157_44484# VDD 0.174233f
C2223 a_17609_46634# a_765_45546# 0.256159f
C2224 a_20922_43172# a_21195_42852# 0.119168f
C2225 a_13887_32519# a_14097_32519# 10.5943f
C2226 a_17970_44736# a_18248_44752# 0.117156f
C2227 a_1307_43914# a_2998_44172# 0.233292f
C2228 a_13259_45724# a_5649_42852# 1.92021f
C2229 a_5343_44458# a_6109_44484# 0.285594f
C2230 a_13925_46122# a_14840_46494# 0.118759f
C2231 a_2804_46116# a_2981_46116# 0.134298f
C2232 a_5937_45572# a_6945_45028# 0.22046f
C2233 a_n2438_43548# a_949_44458# 1.62911f
C2234 a_3090_45724# a_1423_45028# 0.450367f
C2235 a_20820_30879# EN_OFFSET_CAL 0.107181f
C2236 a_n1991_46122# VDD 0.581018f
C2237 a_n2109_47186# a_n1151_42308# 0.235661f
C2238 a_n785_47204# a_327_47204# 0.237391f
C2239 a_n971_45724# a_2124_47436# 0.352461f
C2240 a_n237_47217# a_1239_47204# 0.203126f
C2241 a_2479_44172# a_2813_43396# 0.115852f
C2242 a_14113_42308# VDD 0.365578f
C2243 a_8199_44636# a_8701_44490# 0.25266f
C2244 a_15599_45572# a_16115_45572# 0.105995f
C2245 a_3483_46348# a_14539_43914# 1.24006f
C2246 a_7499_43078# VDD 1.87959f
C2247 a_n2497_47436# a_3090_45724# 0.16041f
C2248 a_n1613_43370# a_n2661_46634# 0.279652f
C2249 a_768_44030# a_13661_43548# 0.175469f
C2250 CAL_N a_22609_38406# 0.204621f
C2251 a_7754_39964# VDD 0.848281f
C2252 a_20202_43084# a_21381_43940# 0.108097f
C2253 a_10193_42453# a_n356_44636# 2.49128f
C2254 a_10227_46804# a_10809_44734# 0.17883f
C2255 a_18479_47436# a_6945_45028# 0.348097f
C2256 a_8605_42826# a_8387_43230# 0.209641f
C2257 a_3626_43646# a_1755_42282# 0.119352f
C2258 a_n97_42460# a_6123_31319# 0.182488f
C2259 a_n2293_42834# a_5891_43370# 0.669411f
C2260 a_3600_43914# VDD 0.22716f
C2261 a_16327_47482# a_18479_45785# 0.841261f
C2262 a_n971_45724# a_n967_45348# 0.581053f
C2263 a_2521_46116# a_2698_46116# 0.159555f
C2264 a_5129_47502# VDD 0.20906f
C2265 a_3785_47178# DATA[2] 0.119025f
C2266 a_9290_44172# a_5742_30871# 0.118117f
C2267 a_1307_43914# a_1568_43370# 0.182552f
C2268 a_15781_43660# VDD 0.196099f
C2269 a_15227_44166# VDD 2.69945f
C2270 a_n2956_39304# a_n2946_39072# 0.150476f
C2271 a_n1329_42308# VDD 0.237697f
C2272 a_13163_45724# a_13527_45546# 0.124682f
C2273 a_13507_46334# a_11341_43940# 0.162723f
C2274 a_10053_45546# a_10210_45822# 0.18824f
C2275 a_11823_42460# a_13249_42308# 0.360411f
C2276 a_n1151_42308# a_n1925_46634# 0.105874f
C2277 a_10227_46804# a_n881_46662# 0.146883f
C2278 a_7754_38968# a_3754_38470# 0.209356f
C2279 a_20447_31679# a_413_45260# 0.226658f
C2280 a_7499_43078# a_11827_44484# 0.104754f
C2281 a_3357_43084# a_2382_45260# 0.219664f
C2282 a_n2109_45247# en_comp 0.108653f
C2283 a_4558_45348# VDD 0.25277f
C2284 a_4791_45118# a_8199_44636# 0.14611f
C2285 a_4883_46098# a_20202_43084# 0.135688f
C2286 a_n1613_43370# a_765_45546# 0.205521f
C2287 a_2063_45854# a_10903_43370# 0.277624f
C2288 a_9482_43914# a_13076_44458# 0.103066f
C2289 a_1307_43914# a_5883_43914# 0.289388f
C2290 a_526_44458# a_3539_42460# 0.213772f
C2291 a_20273_46660# a_12741_44636# 0.540506f
C2292 a_12861_44030# a_11823_42460# 1.2465f
C2293 w_1575_34946# a_n923_35174# 37.7438f
C2294 a_1756_43548# VDD 0.138878f
C2295 a_1176_45822# a_997_45618# 0.140567f
C2296 a_12891_46348# a_9482_43914# 0.314487f
C2297 a_8325_42308# a_8791_42308# 0.173196f
C2298 a_22400_42852# a_22469_40625# 0.954861f
C2299 a_n2438_43548# a_n2293_43922# 0.575621f
C2300 a_6945_45028# a_2437_43646# 2.26888f
C2301 a_12549_44172# a_19615_44636# 0.157395f
C2302 a_22959_46124# VDD 0.309939f
C2303 a_2063_45854# a_4883_46098# 0.116597f
C2304 a_n4064_40160# a_n3565_37414# 4.29714f
C2305 a_3090_45724# a_10405_44172# 0.126512f
C2306 a_11823_42460# a_11787_45002# 0.217891f
C2307 a_10903_43370# a_n2661_42834# 0.269313f
C2308 a_20193_45348# a_21613_42308# 0.137559f
C2309 a_2107_46812# a_1983_46706# 0.212212f
C2310 a_n2438_43548# a_n2661_46098# 0.391488f
C2311 C1_P_btm C0_dummy_P_btm 1.2494f
C2312 EN_VIN_BSTR_N VDD 1.13406f
C2313 a_18783_43370# a_15743_43084# 0.303966f
C2314 a_4791_45118# a_4921_42308# 0.172224f
C2315 a_9838_44484# VDD 0.242131f
C2316 a_3232_43370# a_3499_42826# 0.339727f
C2317 a_7499_43078# a_8147_43396# 0.227361f
C2318 a_13759_46122# a_14840_46494# 0.102325f
C2319 a_14493_46090# a_14275_46494# 0.209641f
C2320 a_n443_46116# a_1307_43914# 0.442637f
C2321 a_n881_46662# RST_Z 0.351994f
C2322 a_14635_42282# a_14456_42282# 0.172313f
C2323 a_n2438_43548# a_742_44458# 0.171623f
C2324 a_n863_45724# a_n1099_45572# 0.172847f
C2325 a_8034_45724# a_8162_45546# 0.14162f
C2326 a_13661_43548# a_13720_44458# 0.122691f
C2327 a_n1853_46287# VDD 0.645231f
C2328 a_n237_47217# a_1209_47178# 0.206644f
C2329 a_n23_47502# a_327_47204# 0.140943f
C2330 a_5111_44636# a_5379_42460# 0.118194f
C2331 a_15493_43940# a_19319_43548# 0.36082f
C2332 a_13657_42558# VDD 0.195727f
C2333 a_8199_44636# a_8103_44636# 0.256009f
C2334 a_15903_45785# a_15765_45572# 0.205788f
C2335 a_13059_46348# a_14673_44172# 0.108306f
C2336 a_8568_45546# VDD 0.182812f
C2337 a_6151_47436# a_8492_46660# 0.302615f
C2338 a_12549_44172# a_13661_43548# 0.149087f
C2339 CAL_N CAL_P 5.91728f
C2340 a_22521_40055# a_22821_38993# 0.131339f
C2341 a_22459_39145# a_22545_38993# 0.121283f
C2342 a_8685_43396# a_14955_43396# 0.111211f
C2343 a_3537_45260# a_1307_43914# 0.290878f
C2344 a_n2661_43370# VDD 1.53673f
C2345 a_8037_42858# a_8387_43230# 0.225358f
C2346 a_7871_42858# a_8952_43230# 0.102355f
C2347 a_13556_45296# a_14673_44172# 0.137701f
C2348 a_n2293_45010# a_n1899_43946# 0.18948f
C2349 a_2998_44172# VDD 0.362233f
C2350 a_16327_47482# a_18175_45572# 0.346603f
C2351 a_765_45546# a_6945_45028# 4.99804f
C2352 a_4915_47217# VDD 3.43172f
C2353 a_17517_44484# a_11967_42832# 0.342031f
C2354 a_5111_44636# a_7287_43370# 0.104641f
C2355 a_15681_43442# VDD 0.159054f
C2356 a_3090_45724# a_3357_43084# 0.546562f
C2357 a_18834_46812# VDD 0.116625f
C2358 a_n2956_39304# a_n3420_39072# 0.208204f
C2359 COMP_P VDD 3.48893f
C2360 a_11599_46634# a_12891_46348# 0.150715f
C2361 a_11453_44696# a_22959_47212# 0.182671f
C2362 a_3754_38802# VDAC_Ni 0.301032f
C2363 a_4574_45260# VDD 0.122256f
C2364 a_13507_46334# a_11415_45002# 0.160889f
C2365 a_n2293_46634# a_3090_45724# 1.2853f
C2366 a_10807_43548# a_11323_42473# 0.109765f
C2367 a_768_44030# a_n755_45592# 0.202175f
C2368 w_1575_34946# a_n1532_35090# 0.796778f
C2369 a_n357_42282# a_7227_42852# 0.185359f
C2370 a_1568_43370# VDD 0.433732f
C2371 a_1138_42852# a_n357_42282# 0.325445f
C2372 a_n2497_47436# a_n699_43396# 0.355158f
C2373 a_8325_42308# a_8685_42308# 0.141819f
C2374 a_18494_42460# a_16137_43396# 0.115144f
C2375 a_22400_42852# a_22521_40599# 0.133947f
C2376 a_5907_45546# a_6194_45824# 0.233657f
C2377 a_n2293_46098# a_1307_43914# 0.107603f
C2378 a_12549_44172# a_11967_42832# 0.193926f
C2379 a_10809_44734# VDD 2.67671f
C2380 a_20193_45348# a_21887_42336# 0.169001f
C2381 a_16327_47482# a_19466_46812# 0.203994f
C2382 a_n743_46660# a_n2661_46098# 0.414618f
C2383 a_n2438_43548# a_1799_45572# 0.137623f
C2384 C2_P_btm C0_dummy_P_btm 6.66125f
C2385 C1_P_btm C0_P_btm 10.8764f
C2386 a_11530_34132# VDD 0.362839f
C2387 a_5883_43914# VDD 0.859221f
C2388 a_4955_46873# a_4704_46090# 0.109136f
C2389 a_17767_44458# a_17970_44736# 0.233657f
C2390 a_1307_43914# a_2675_43914# 0.453622f
C2391 a_626_44172# a_453_43940# 0.163589f
C2392 a_13925_46122# a_14275_46494# 0.20669f
C2393 a_n881_46662# VDD 2.6692f
C2394 a_1184_42692# a_2123_42473# 0.107417f
C2395 a_n863_45724# a_1606_42308# 0.20593f
C2396 a_15227_44166# a_15415_45028# 0.222342f
C2397 a_n1079_45724# a_n1099_45572# 0.15766f
C2398 a_n2293_45546# a_310_45028# 0.113595f
C2399 a_n2157_46122# VDD 0.42567f
C2400 a_11415_45002# EN_OFFSET_CAL 0.14622f
C2401 a_n2497_47436# a_n1151_42308# 0.156942f
C2402 a_n2109_47186# a_2905_45572# 0.124881f
C2403 a_n3420_39616# a_n4064_39616# 6.66063f
C2404 a_n913_45002# a_8325_42308# 0.233489f
C2405 a_15599_45572# a_15765_45572# 0.576512f
C2406 a_8162_45546# VDD 0.266272f
C2407 a_6151_47436# a_8667_46634# 0.357581f
C2408 a_12549_44172# a_5807_45002# 0.675558f
C2409 a_11206_38545# CAL_P 0.234643f
C2410 a_22469_40625# a_22469_39537# 0.604831f
C2411 a_7754_40130# VDD 13.6809f
C2412 a_n97_42460# a_4361_42308# 0.15989f
C2413 a_10227_46804# a_6945_45028# 0.220094f
C2414 a_768_44030# a_3483_46348# 0.281593f
C2415 a_8037_42858# a_8605_42826# 0.178024f
C2416 a_9482_43914# a_14673_44172# 0.42967f
C2417 a_n2293_45010# a_n1761_44111# 0.148418f
C2418 a_2889_44172# VDD 0.1447f
C2419 a_3090_45724# a_8049_45260# 1.23904f
C2420 a_167_45260# a_2521_46116# 0.328009f
C2421 a_n443_46116# VDD 3.87014f
C2422 a_2063_45854# CLK 0.271193f
C2423 a_2324_44458# a_2711_45572# 0.804101f
C2424 a_526_44458# a_n863_45724# 0.801581f
C2425 a_11453_44696# a_n2661_44458# 0.174607f
C2426 a_17609_46634# VDD 0.501057f
C2427 a_5742_30871# a_7174_31319# 0.34728f
C2428 a_n4318_37592# VDD 0.919667f
C2429 a_n2293_46634# a_1414_42308# 0.260739f
C2430 a_19443_46116# VDD 0.132317f
C2431 a_13487_47204# a_768_44030# 0.371206f
C2432 a_n1059_45260# a_n913_45002# 1.19505f
C2433 a_10193_42453# a_18184_42460# 0.216199f
C2434 a_4646_46812# a_6197_43396# 0.601282f
C2435 a_n2472_45002# en_comp 0.117861f
C2436 a_3537_45260# VDD 3.9063f
C2437 a_20916_46384# a_15227_44166# 0.681561f
C2438 a_13507_46334# a_20202_43084# 0.205796f
C2439 a_19594_46812# a_19692_46634# 0.134424f
C2440 a_9482_43914# a_12607_44458# 0.151452f
C2441 a_9290_44172# a_10341_43396# 0.157042f
C2442 a_768_44030# a_n357_42282# 0.175577f
C2443 a_20107_46660# a_12741_44636# 0.527863f
C2444 a_12861_44030# a_11962_45724# 0.184706f
C2445 a_n357_42282# a_5755_42852# 0.179701f
C2446 a_13259_45724# a_17701_42308# 0.137488f
C2447 a_1049_43396# VDD 0.196328f
C2448 a_n746_45260# a_n2129_44697# 0.17701f
C2449 a_5932_42308# a_5742_30871# 1.14154f
C2450 a_5891_43370# a_n97_42460# 0.957548f
C2451 a_22223_46124# VDD 0.300745f
C2452 a_n2840_43370# a_n4318_39304# 0.158695f
C2453 a_9290_44172# a_n2293_43922# 0.369185f
C2454 C2_P_btm C0_P_btm 0.698973f
C2455 a_n83_35174# VDD 0.313947f
C2456 EN_VIN_BSTR_N C10_N_btm 0.320569f
C2457 a_18525_43370# a_18783_43370# 0.22264f
C2458 a_9290_44172# a_n97_42460# 0.351467f
C2459 a_8701_44490# VDD 0.164475f
C2460 a_21588_30879# a_10809_44734# 0.110956f
C2461 a_1307_43914# a_895_43940# 0.754684f
C2462 a_11691_44458# a_15433_44458# 0.110923f
C2463 a_13759_46122# a_14275_46494# 0.105995f
C2464 a_13925_46122# a_14493_46090# 0.17072f
C2465 a_19321_45002# a_18479_45785# 0.114441f
C2466 a_n1613_43370# VDD 4.75085f
C2467 a_n1533_42852# VDD 0.142813f
C2468 a_n2661_45546# a_n755_45592# 0.14317f
C2469 a_n2293_46098# VDD 1.7963f
C2470 a_n3420_39616# a_n2946_39866# 0.236674f
C2471 a_4958_30871# C9_P_btm 0.209166f
C2472 a_15599_45572# a_15903_45785# 0.161702f
C2473 a_1609_45822# a_2274_45254# 0.11737f
C2474 a_6151_47436# a_7927_46660# 0.182356f
C2475 a_22521_40055# a_22521_39511# 0.457858f
C2476 a_22521_40599# a_22469_39537# 0.380006f
C2477 a_3232_43370# a_9482_43914# 0.129525f
C2478 a_413_45260# a_1423_45028# 0.194002f
C2479 a_2324_44458# a_15682_43940# 0.321744f
C2480 a_12549_44172# a_3483_46348# 0.185475f
C2481 a_7871_42858# a_8387_43230# 0.106107f
C2482 a_3080_42308# a_2903_42308# 0.154008f
C2483 a_2675_43914# VDD 0.200923f
C2484 a_n746_45260# a_n745_45366# 0.119822f
C2485 a_4791_45118# VDD 3.05095f
C2486 a_5534_30871# a_12563_42308# 0.179331f
C2487 a_5883_43914# a_n2661_42282# 0.107496f
C2488 a_19466_46812# a_20528_45572# 0.157758f
C2489 a_16292_46812# VDD 0.123916f
C2490 a_n2956_39304# a_n3565_39304# 0.307358f
C2491 a_18326_43940# a_18451_43940# 0.145292f
C2492 a_n1736_42282# VDD 0.227152f
C2493 a_n971_45724# a_n2129_43609# 0.173854f
C2494 a_2063_45854# a_n743_46660# 1.58762f
C2495 a_12861_44030# a_768_44030# 0.260776f
C2496 SMPL_ON_N a_11453_44696# 0.147722f
C2497 a_n4064_39072# EN_VIN_BSTR_P 0.959329f
C2498 a_7754_38968# a_7754_38636# 0.296258f
C2499 a_3540_43646# a_3626_43646# 0.100706f
C2500 a_n2017_45002# a_n913_45002# 0.275686f
C2501 a_n2661_45010# en_comp 0.10363f
C2502 a_n2472_45002# a_n2956_37592# 0.152938f
C2503 a_3429_45260# VDD 0.142923f
C2504 a_2063_45854# a_11189_46129# 0.294233f
C2505 a_19594_46812# a_19466_46812# 0.100902f
C2506 a_22959_43396# a_17364_32525# 0.156288f
C2507 a_1423_45028# a_2779_44458# 0.246285f
C2508 a_9482_43914# a_8975_43940# 0.186623f
C2509 a_20202_43084# a_4361_42308# 0.472299f
C2510 a_13259_45724# a_17595_43084# 0.118887f
C2511 a_1209_43370# VDD 0.191694f
C2512 a_167_45260# a_n863_45724# 0.424358f
C2513 a_12891_46348# a_13017_45260# 0.210934f
C2514 a_3483_46348# a_n2661_45546# 0.163728f
C2515 a_9290_44172# a_13259_45724# 0.272297f
C2516 a_3090_45724# a_11691_44458# 0.245063f
C2517 a_13661_43548# a_14673_44172# 0.36897f
C2518 a_6945_45028# VDD 1.30257f
C2519 a_16327_47482# a_15227_44166# 0.239667f
C2520 C4_P_btm C0_dummy_P_btm 0.113746f
C2521 C2_P_btm C1_P_btm 5.0586f
C2522 C3_P_btm C0_P_btm 0.409996f
C2523 EN_VIN_BSTR_P VDD 0.917313f
C2524 EN_VIN_BSTR_N C9_N_btm 0.226529f
C2525 a_n97_42460# a_16795_42852# 0.126591f
C2526 a_1823_45246# a_3539_42460# 0.678673f
C2527 a_n3674_39768# a_n4064_39616# 0.464693f
C2528 a_8103_44636# VDD 0.124028f
C2529 a_1307_43914# a_2479_44172# 0.300587f
C2530 a_3537_45260# a_n2661_42282# 0.105917f
C2531 a_3090_45724# a_n443_42852# 0.269331f
C2532 a_19123_46287# a_19240_46482# 0.157972f
C2533 a_1823_45246# a_526_44458# 1.93329f
C2534 a_13747_46662# a_18341_45572# 0.554429f
C2535 a_1576_42282# a_1755_42282# 0.168925f
C2536 a_1184_42692# a_1606_42308# 0.125247f
C2537 a_13291_42460# a_13070_42354# 0.155164f
C2538 a_22959_44484# a_19237_31679# 0.155744f
C2539 a_15227_44166# a_14537_43396# 0.105881f
C2540 a_n2472_46090# VDD 0.224658f
C2541 a_22365_46825# EN_OFFSET_CAL 0.195393f
C2542 a_n746_45260# a_n785_47204# 0.198992f
C2543 a_n3565_39590# a_n4064_39616# 0.231239f
C2544 a_11967_42832# a_16547_43609# 0.176385f
C2545 a_19862_44208# a_21381_43940# 0.113704f
C2546 a_14456_42282# VDD 0.265543f
C2547 a_6812_45938# VDD 0.132317f
C2548 a_n1151_42308# a_6755_46942# 0.142929f
C2549 a_6151_47436# a_8145_46902# 0.178565f
C2550 a_327_44734# a_626_44172# 0.120093f
C2551 a_7765_42852# a_8037_42858# 0.309282f
C2552 a_n2840_44458# a_n2661_44458# 0.179135f
C2553 a_n755_45592# a_n1557_42282# 0.199254f
C2554 a_895_43940# VDD 0.318652f
C2555 a_2202_46116# a_167_45260# 0.159883f
C2556 a_11599_46634# a_18341_45572# 0.588263f
C2557 a_3483_46348# a_11322_45546# 0.554731f
C2558 a_15559_46634# VDD 0.301657f
C2559 a_5663_43940# a_5829_43940# 0.143754f
C2560 a_10729_43914# a_11341_43940# 0.243062f
C2561 a_10193_42453# a_4958_30871# 0.108497f
C2562 a_n3674_38216# VDD 0.309006f
C2563 a_584_46384# a_n743_46660# 0.42078f
C2564 a_12861_44030# a_12549_44172# 1.20253f
C2565 a_22775_42308# VDD 0.426018f
C2566 a_2982_43646# a_3626_43646# 6.553431f
C2567 a_n2017_45002# a_n1059_45260# 6.27837f
C2568 a_3357_43084# a_413_45260# 7.24598f
C2569 a_4646_46812# a_6031_43396# 0.849684f
C2570 a_n2293_46098# a_n2661_42282# 0.182071f
C2571 a_n2661_45010# a_n2956_37592# 0.163638f
C2572 a_3065_45002# VDD 0.501045f
C2573 a_18597_46090# a_12741_44636# 0.267775f
C2574 a_768_44030# a_14035_46660# 0.270355f
C2575 a_n1151_42308# a_8953_45546# 0.120628f
C2576 a_4791_45118# a_6419_46155# 0.371259f
C2577 a_2063_45854# a_9290_44172# 0.655982f
C2578 a_19321_45002# a_19466_46812# 0.130025f
C2579 a_20202_43084# a_13467_32519# 0.333168f
C2580 a_9482_43914# a_10057_43914# 0.401746f
C2581 a_11599_46634# a_10193_42453# 0.100544f
C2582 a_458_43396# VDD 0.431902f
C2583 a_10903_43370# a_12839_46116# 0.115226f
C2584 a_n2497_47436# a_949_44458# 0.127971f
C2585 a_n2293_46634# a_413_45260# 0.497204f
C2586 a_5807_45002# a_6171_45002# 0.193427f
C2587 a_3067_47026# VDD 0.132018f
C2588 a_n2017_45002# a_19987_42826# 0.142839f
C2589 a_3090_45724# a_19113_45348# 0.128103f
C2590 a_21137_46414# VDD 0.219745f
C2591 a_9313_45822# a_11459_47204# 0.210847f
C2592 a_n3565_38502# a_n4209_38216# 5.84657f
C2593 a_n1613_43370# a_7112_43396# 0.245085f
C2594 a_10227_46804# a_14976_45028# 0.536884f
C2595 a_1123_46634# a_948_46660# 0.234322f
C2596 C5_P_btm C0_dummy_P_btm 0.11443f
C2597 C3_P_btm C1_P_btm 7.40325f
C2598 C4_P_btm C0_P_btm 0.138884f
C2599 a_n923_35174# VDD 0.340432f
C2600 a_18429_43548# a_18525_43370# 0.419086f
C2601 a_n443_42852# a_1414_42308# 0.193113f
C2602 a_n2661_45010# a_n2267_44484# 0.260289f
C2603 a_13507_46334# a_22400_42852# 0.235269f
C2604 a_6298_44484# VDD 1.21616f
C2605 a_768_44030# a_n1925_42282# 0.145535f
C2606 a_n443_46116# a_n23_45546# 0.118272f
C2607 a_18597_46090# a_16375_45002# 0.105669f
C2608 a_6755_46942# a_12741_44636# 0.131965f
C2609 a_1307_43914# a_2127_44172# 0.127867f
C2610 a_13759_46122# a_13925_46122# 0.576786f
C2611 a_1576_42282# a_1606_42308# 0.176925f
C2612 a_n2840_46090# VDD 0.295278f
C2613 a_n971_45724# a_n785_47204# 0.385455f
C2614 a_n746_45260# a_n23_47502# 0.148631f
C2615 a_n3690_39616# a_n3420_39616# 0.431154f
C2616 a_n3565_39590# a_n2946_39866# 0.406088f
C2617 a_n4334_39616# a_n4064_39616# 0.4504f
C2618 a_n4209_39590# a_n2302_39866# 0.406459f
C2619 a_11967_42832# a_16243_43396# 0.269605f
C2620 a_13575_42558# VDD 0.182133f
C2621 a_8049_45260# a_n2293_42834# 0.224469f
C2622 a_6151_47436# a_7577_46660# 0.578207f
C2623 a_n237_47217# a_8270_45546# 0.552109f
C2624 a_22521_40055# a_22459_39145# 0.129251f
C2625 a_22469_40625# a_22521_39511# 0.65678f
C2626 a_n2293_43922# a_5932_42308# 0.178011f
C2627 a_17538_32519# a_17364_32525# 9.64512f
C2628 a_13259_45724# a_3422_30871# 0.587088f
C2629 a_2382_45260# a_1307_43914# 0.53878f
C2630 a_6755_46942# a_13607_46688# 0.129798f
C2631 a_7871_42858# a_8037_42858# 0.772842f
C2632 a_n2840_44458# a_n4318_40392# 0.161548f
C2633 a_n357_42282# a_n1557_42282# 0.384406f
C2634 a_2479_44172# VDD 0.431428f
C2635 a_12891_46348# a_13249_42308# 0.166217f
C2636 a_1823_45246# a_167_45260# 0.155648f
C2637 a_n971_45724# a_n913_45002# 0.101346f
C2638 a_n746_45260# a_n1059_45260# 0.138039f
C2639 a_19123_46287# a_18985_46122# 0.215692f
C2640 a_13661_43548# a_10193_42453# 0.211481f
C2641 a_4007_47204# VDD 0.41212f
C2642 a_7499_43078# a_10341_42308# 0.42152f
C2643 a_3537_45260# a_7287_43370# 0.400907f
C2644 a_20193_45348# a_15493_43940# 0.10893f
C2645 a_3483_46348# a_10490_45724# 0.207668f
C2646 a_4185_45028# a_10193_42453# 3.16135f
C2647 a_15368_46634# VDD 0.324877f
C2648 a_n2956_39304# a_n4209_39304# 0.328727f
C2649 a_15764_42576# a_4958_30871# 0.413236f
C2650 a_18079_43940# a_18326_43940# 0.152347f
C2651 a_n2104_42282# VDD 0.280329f
C2652 a_11962_45724# a_13163_45724# 0.113317f
C2653 a_8049_45260# a_413_45260# 0.140877f
C2654 a_12427_45724# a_12791_45546# 0.124682f
C2655 a_22731_47423# SMPL_ON_N 0.194951f
C2656 a_16327_47482# a_n881_46662# 0.195459f
C2657 a_n3420_39072# EN_VIN_BSTR_P 0.772414f
C2658 a_21613_42308# VDD 0.273985f
C2659 a_n443_42852# a_n699_43396# 0.333516f
C2660 a_5257_43370# a_4905_42826# 0.254437f
C2661 a_2680_45002# VDD 0.145087f
C2662 a_4646_46812# a_7411_46660# 0.266058f
C2663 a_n1151_42308# a_5937_45572# 0.11638f
C2664 a_4791_45118# a_6165_46155# 0.291653f
C2665 a_375_42282# a_n699_43396# 0.127058f
C2666 a_18248_44752# a_17517_44484# 0.561898f
C2667 a_n229_43646# VDD 0.278436f
C2668 a_1823_45246# a_n863_45724# 0.207189f
C2669 a_n2497_47436# a_742_44458# 0.153038f
C2670 a_167_45260# a_n2293_45546# 0.681309f
C2671 a_n2438_43548# en_comp 0.915368f
C2672 a_8515_42308# a_8685_42308# 0.108744f
C2673 a_5934_30871# a_8791_42308# 0.223675f
C2674 a_3600_43914# a_3499_42826# 0.125876f
C2675 a_19466_46812# a_19778_44110# 0.116901f
C2676 a_2063_45854# a_10949_43914# 0.129837f
C2677 a_3483_46348# a_6171_45002# 0.153232f
C2678 a_20202_43084# a_3422_30871# 0.527141f
C2679 a_n1613_43370# a_7287_43370# 0.337957f
C2680 a_10227_46804# a_3090_45724# 0.320681f
C2681 a_171_46873# a_288_46660# 0.159893f
C2682 C6_P_btm C0_dummy_P_btm 0.120464f
C2683 C3_P_btm C2_P_btm 5.64696f
C2684 C5_P_btm C0_P_btm 0.138736f
C2685 C4_P_btm C1_P_btm 0.128692f
C2686 a_n1532_35090# VDD 2.19114f
C2687 EN_VIN_BSTR_N C7_N_btm 0.115875f
C2688 a_16547_43609# a_16664_43396# 0.161376f
C2689 a_11967_42832# a_15803_42450# 0.258862f
C2690 a_21381_43940# a_21195_42852# 0.238789f
C2691 a_n2661_45010# a_n2129_44697# 0.18531f
C2692 a_10193_42453# a_11967_42832# 0.752992f
C2693 a_4791_45118# a_5379_42460# 0.197725f
C2694 a_5518_44484# VDD 0.40715f
C2695 a_768_44030# a_526_44458# 0.341438f
C2696 a_n443_46116# a_n356_45724# 0.113738f
C2697 a_14539_43914# a_16979_44734# 0.132799f
C2698 a_626_44172# a_644_44056# 0.126386f
C2699 a_n863_45724# a_1184_42692# 0.563857f
C2700 a_n357_42282# a_n3674_37592# 0.327427f
C2701 a_n2293_45546# a_n863_45724# 0.17075f
C2702 a_3090_45724# a_1307_43914# 2.66267f
C2703 a_n746_45260# a_n237_47217# 0.285294f
C2704 a_n971_45724# a_n23_47502# 0.225828f
C2705 a_n2109_47186# a_584_46384# 0.352889f
C2706 a_n3565_39590# a_n3420_39616# 0.281955f
C2707 a_n4209_39590# a_n4064_39616# 0.269818f
C2708 a_11967_42832# a_16137_43396# 0.300696f
C2709 a_13070_42354# VDD 0.18656f
C2710 a_n2293_46634# a_11341_43940# 0.487839f
C2711 a_3090_45724# a_18579_44172# 0.16932f
C2712 a_13661_43548# a_14021_43940# 0.103152f
C2713 a_6491_46660# a_5257_43370# 0.1719f
C2714 a_22521_40599# a_22521_39511# 0.365591f
C2715 a_n2438_43548# a_n2157_42858# 0.266513f
C2716 a_13507_46334# a_22165_42308# 0.126777f
C2717 a_18597_46090# a_18819_46122# 0.230891f
C2718 a_7871_42858# a_7765_42852# 0.379881f
C2719 a_2127_44172# VDD 0.138239f
C2720 a_n971_45724# a_n1059_45260# 0.322275f
C2721 a_11599_46634# a_18175_45572# 0.844188f
C2722 a_19123_46287# a_18819_46122# 0.172712f
C2723 a_1138_42852# a_167_45260# 0.250282f
C2724 a_1823_45246# a_2202_46116# 0.25354f
C2725 a_3815_47204# VDD 0.260661f
C2726 a_4223_44672# a_8333_44056# 0.122173f
C2727 a_5111_44636# a_6031_43396# 0.207345f
C2728 a_3483_46348# a_8746_45002# 0.605995f
C2729 a_n1925_42282# a_n2661_45546# 0.181908f
C2730 a_12549_44172# a_16922_45042# 0.803336f
C2731 a_14976_45028# VDD 0.484864f
C2732 a_n4318_38216# VDD 0.538766f
C2733 a_12741_44636# a_11691_44458# 0.81445f
C2734 a_12427_45724# a_11823_42460# 0.17307f
C2735 a_11962_45724# a_12791_45546# 0.124167f
C2736 a_n2497_47436# a_n447_43370# 0.192476f
C2737 a_18051_46116# VDD 0.189782f
C2738 a_n1151_42308# a_n2661_46634# 0.832521f
C2739 a_21887_42336# VDD 0.210392f
C2740 a_n2109_45247# a_n2017_45002# 0.193269f
C2741 a_n2840_45002# a_n2810_45028# 0.161831f
C2742 a_n2293_46634# a_10341_43396# 2.04894f
C2743 a_2382_45260# VDD 1.6285f
C2744 a_19321_45002# a_15227_44166# 0.145462f
C2745 a_n1151_42308# a_8199_44636# 0.161616f
C2746 a_13747_46662# a_19466_46812# 0.869986f
C2747 a_n443_42852# a_15493_43940# 0.301211f
C2748 a_15433_44458# VDD 0.201121f
C2749 a_18114_32519# a_19237_31679# 8.86333f
C2750 a_3357_43084# a_n97_42460# 0.113127f
C2751 a_3080_42308# C2_N_btm 0.108823f
C2752 a_1138_42852# a_n863_45724# 0.135594f
C2753 a_2324_44458# a_10586_45546# 0.436403f
C2754 a_5807_45002# a_5691_45260# 0.19412f
C2755 a_3524_46660# VDD 0.278519f
C2756 a_8515_42308# a_8325_42308# 0.134955f
C2757 a_5934_30871# a_8685_42308# 0.186981f
C2758 a_3483_46348# a_3232_43370# 0.220803f
C2759 a_19900_46494# VDD 0.279179f
C2760 a_n2293_46634# a_n97_42460# 0.108602f
C2761 a_n1613_43370# a_6547_43396# 0.154311f
C2762 a_n443_42852# a_n2293_42834# 1.60683f
C2763 a_n2438_43548# a_n2267_43396# 0.120634f
C2764 a_n1151_42308# a_765_45546# 1.7705f
C2765 a_11599_46634# a_19466_46812# 0.453656f
C2766 C7_P_btm C0_dummy_P_btm 0.120543f
C2767 C6_P_btm C0_P_btm 0.140033f
C2768 C5_P_btm C1_P_btm 0.128021f
C2769 C4_P_btm C2_P_btm 7.19288f
C2770 a_n1386_35608# VDD 0.360375f
C2771 EN_VIN_BSTR_N C6_N_btm 0.118916f
C2772 a_21381_43940# a_21356_42826# 0.196864f
C2773 a_n2661_45010# a_n2433_44484# 0.217176f
C2774 a_4791_45118# a_5267_42460# 0.138738f
C2775 a_5343_44458# VDD 0.49245f
C2776 a_20916_46384# a_21137_46414# 0.118131f
C2777 a_3877_44458# a_4185_45028# 0.338483f
C2778 a_19339_43156# a_19164_43230# 0.233657f
C2779 a_7227_42852# a_7309_42852# 0.171361f
C2780 a_526_44458# a_5111_42852# 0.265994f
C2781 a_1307_43914# a_1414_42308# 0.147738f
C2782 a_5807_45002# a_18479_45785# 0.174313f
C2783 a_1184_42692# a_961_42354# 0.100246f
C2784 a_n755_45592# a_n784_42308# 0.711298f
C2785 a_n2438_43548# a_n2267_44484# 0.120608f
C2786 a_n815_47178# a_n785_47204# 0.123817f
C2787 a_n971_45724# a_n237_47217# 0.134971f
C2788 a_n3565_39590# a_n3690_39616# 0.246863f
C2789 a_n913_45002# a_5934_30871# 0.126791f
C2790 a_12563_42308# VDD 0.254292f
C2791 a_n971_45724# a_8270_45546# 0.251101f
C2792 a_6151_47436# a_7411_46660# 0.330209f
C2793 a_22469_40625# a_22459_39145# 0.245891f
C2794 a_14401_32519# a_17364_32525# 7.51978f
C2795 a_n97_42460# a_743_42282# 0.107736f
C2796 a_413_45260# a_375_42282# 0.112554f
C2797 a_16327_47482# a_6945_45028# 0.111399f
C2798 a_n1741_47186# a_12839_46116# 0.113988f
C2799 a_7227_42852# a_7765_42852# 0.118623f
C2800 a_n755_45592# a_3080_42308# 0.237742f
C2801 a_453_43940# VDD 0.225569f
C2802 a_12549_44172# a_13163_45724# 0.172293f
C2803 a_3785_47178# VDD 0.387755f
C2804 a_20193_45348# a_11341_43940# 0.21261f
C2805 a_3483_46348# a_10193_42453# 0.359034f
C2806 a_3090_45724# VDD 2.05725f
C2807 a_17973_43940# a_18079_43940# 0.419086f
C2808 a_17730_32519# a_17538_32519# 9.37324f
C2809 a_n2472_42282# VDD 0.278905f
C2810 a_n2438_43548# a_n2065_43946# 0.265458f
C2811 a_11962_45724# a_11823_42460# 0.177935f
C2812 a_13381_47204# a_12549_44172# 0.135267f
C2813 a_21335_42336# VDD 0.199586f
C2814 a_2896_43646# a_2982_43646# 0.100706f
C2815 a_2437_43646# a_413_45260# 0.20387f
C2816 a_2274_45254# VDD 0.256655f
C2817 a_3877_44458# a_5257_43370# 0.142219f
C2818 a_22591_43396# a_14209_32519# 0.158752f
C2819 a_9482_43914# a_10157_44484# 0.321004f
C2820 a_14815_43914# VDD 0.307386f
C2821 a_n443_42852# a_n13_43084# 0.13203f
C2822 a_1823_45246# a_n2293_45546# 0.234971f
C2823 a_3699_46634# VDD 0.347281f
C2824 a_5934_30871# a_8325_42308# 0.173576f
C2825 a_n357_42282# a_10193_42453# 0.634772f
C2826 a_20075_46420# VDD 0.347847f
C2827 a_n1151_42308# a_10227_46804# 0.458569f
C2828 a_6151_47436# a_14955_47212# 0.192081f
C2829 SMPL_ON_P a_n2312_40392# 4.89949f
C2830 a_n4064_38528# a_n2302_38778# 0.239588f
C2831 a_n1613_43370# a_6765_43638# 0.164755f
C2832 a_33_46660# a_948_46660# 0.117156f
C2833 C8_P_btm C0_dummy_P_btm 0.236317f
C2834 C6_P_btm C1_P_btm 0.128559f
C2835 C7_P_btm C0_P_btm 0.142187f
C2836 C4_P_btm C3_P_btm 7.90108f
C2837 C5_P_btm C2_P_btm 0.138678f
C2838 a_n1838_35608# VDD 0.523851f
C2839 EN_VIN_BSTR_N C5_N_btm 0.115337f
C2840 a_16409_43396# a_15743_43084# 0.586918f
C2841 a_4743_44484# VDD 0.266843f
C2842 a_n3674_39768# a_n3565_39590# 0.128683f
C2843 a_n881_46662# a_5066_45546# 0.801045f
C2844 a_20916_46384# a_20708_46348# 0.189941f
C2845 a_16112_44458# a_14539_43914# 0.13299f
C2846 a_526_44458# a_4520_42826# 0.247914f
C2847 a_n357_42282# a_16137_43396# 1.09442f
C2848 a_1307_43914# a_1467_44172# 0.228571f
C2849 a_4915_47217# a_13556_45296# 0.146395f
C2850 a_11415_45002# a_8049_45260# 0.426371f
C2851 a_22591_44484# a_17730_32519# 0.156987f
C2852 a_n863_45724# a_1067_42314# 0.289393f
C2853 a_11415_45002# a_19479_31679# 0.224531f
C2854 a_21076_30879# VDD 1.17389f
C2855 a_n971_45724# a_n746_45260# 0.393354f
C2856 a_n4209_39590# a_n3420_39616# 0.234699f
C2857 a_20269_44172# a_19319_43548# 0.12985f
C2858 a_11633_42558# VDD 0.193501f
C2859 a_n443_42852# a_n37_45144# 0.137227f
C2860 a_4883_46098# a_2107_46812# 2.95673f
C2861 a_22521_40599# a_22459_39145# 1.41583f
C2862 a_7229_43940# a_7705_45326# 0.203098f
C2863 a_n443_46116# a_5066_45546# 0.130975f
C2864 a_17730_32519# VREF_GND 0.241027f
C2865 a_1414_42308# VDD 0.657887f
C2866 a_18285_46348# a_17957_46116# 0.12677f
C2867 a_3381_47502# VDD 0.197761f
C2868 a_3537_45260# a_6197_43396# 0.337459f
C2869 a_12281_43396# VDD 0.341026f
C2870 a_5257_43370# a_5111_44636# 0.22597f
C2871 a_8049_45260# a_13259_45724# 0.895805f
C2872 a_19466_46812# a_20273_45572# 0.328586f
C2873 a_15009_46634# VDD 0.205396f
C2874 a_n1059_45260# a_16245_42852# 0.130348f
C2875 a_n3674_38680# VDD 0.503323f
C2876 a_n784_42308# C0_N_btm 0.281635f
C2877 a_20512_43084# a_19987_42826# 0.11919f
C2878 a_1667_45002# VDD 0.315476f
C2879 a_10227_46804# a_12741_44636# 0.188309f
C2880 a_n881_46662# a_13059_46348# 0.642888f
C2881 a_n1151_42308# a_8016_46348# 0.580516f
C2882 a_4791_45118# a_5164_46348# 0.42219f
C2883 a_5807_45002# a_19466_46812# 0.178376f
C2884 VREF_GND VCM 2.79113f
C2885 a_15095_43370# a_15567_42826# 0.167909f
C2886 a_9482_43914# a_9838_44484# 0.175591f
C2887 a_526_44458# a_n1557_42282# 0.31675f
C2888 a_20202_43084# a_743_42282# 0.135735f
C2889 a_n443_42852# a_11341_43940# 0.51832f
C2890 a_1307_43914# a_4223_44672# 0.747516f
C2891 a_18114_32519# a_17730_32519# 9.1497f
C2892 a_16979_44734# a_17517_44484# 0.109784f
C2893 a_17538_32519# VREF_GND 0.117023f
C2894 a_5807_45002# a_5111_44636# 0.204193f
C2895 a_2959_46660# VDD 0.19762f
C2896 a_n4318_39768# a_n3674_39768# 3.06574f
C2897 a_3357_43084# a_n2293_42282# 0.146926f
C2898 a_18579_44172# a_15493_43940# 0.377126f
C2899 a_2711_45572# a_4099_45572# 0.176427f
C2900 a_19335_46494# VDD 0.198512f
C2901 a_6151_47436# a_14311_47204# 0.136645f
C2902 a_n1920_47178# a_n2312_39304# 0.157528f
C2903 a_n2293_43922# a_5534_30871# 0.271171f
C2904 a_n2438_43548# a_n2433_43396# 0.415301f
C2905 a_11599_46634# a_15227_44166# 0.101252f
C2906 a_601_46902# a_383_46660# 0.209641f
C2907 C9_P_btm C0_dummy_P_btm 0.11363f
C2908 C6_P_btm C2_P_btm 0.138423f
C2909 C7_P_btm C1_P_btm 0.129707f
C2910 C8_P_btm C0_P_btm 0.148433f
C2911 C5_P_btm C3_P_btm 0.136119f
C2912 EN_VIN_BSTR_N C4_N_btm 0.116925f
C2913 a_n97_42460# a_5534_30871# 0.109695f
C2914 a_17499_43370# a_17324_43396# 0.234322f
C2915 a_18114_32519# VCM 0.121302f
C2916 a_n699_43396# VDD 0.922998f
C2917 a_16292_46812# a_16388_46812# 0.318472f
C2918 a_5755_42852# a_5837_42852# 0.171361f
C2919 a_n443_42852# a_10341_43396# 0.23026f
C2920 a_1307_43914# a_1115_44172# 0.115939f
C2921 a_22959_43948# VDD 0.297936f
C2922 a_4915_47217# a_9482_43914# 0.269756f
C2923 a_n2293_46098# a_5066_45546# 0.140248f
C2924 SMPL_ON_N VIN_N 0.587565f
C2925 a_n784_42308# a_2123_42473# 0.216332f
C2926 a_1067_42314# a_961_42354# 0.13675f
C2927 a_n4318_38680# VDD 0.417422f
C2928 a_n2438_43548# a_n2433_44484# 0.421822f
C2929 a_14976_45028# a_14797_45144# 0.137651f
C2930 a_22959_46660# VDD 0.299681f
C2931 a_n452_47436# a_n746_45260# 0.187792f
C2932 a_3065_45002# a_3823_42558# 0.198186f
C2933 a_n913_45002# a_6123_31319# 0.21316f
C2934 a_11551_42558# VDD 0.192086f
C2935 a_3316_45546# a_3429_45260# 0.142842f
C2936 a_584_46384# a_3457_43396# 0.120485f
C2937 a_16375_45002# a_1307_43914# 0.101951f
C2938 a_n443_42852# a_n143_45144# 0.104427f
C2939 a_5257_43370# a_3905_42865# 0.106385f
C2940 a_2063_45854# a_6755_46942# 0.131005f
C2941 a_5891_43370# a_9223_42460# 0.13879f
C2942 a_n97_42460# a_4190_30871# 0.140814f
C2943 a_8685_43396# a_9145_43396# 0.201058f
C2944 a_14401_32519# a_14209_32519# 10.7535f
C2945 a_7229_43940# a_6709_45028# 0.136786f
C2946 a_768_44030# a_1823_45246# 0.287407f
C2947 a_4791_45118# a_5066_45546# 0.238282f
C2948 a_21588_30879# a_21076_30879# 8.21286f
C2949 en_comp a_3422_30871# 0.357746f
C2950 a_n443_42852# a_n97_42460# 0.822111f
C2951 a_1467_44172# VDD 0.391994f
C2952 a_12549_44172# a_11823_42460# 0.624462f
C2953 a_n971_45724# a_n2293_45010# 0.549225f
C2954 a_18285_46348# a_18189_46348# 0.118603f
C2955 a_n1151_42308# VDD 2.57238f
C2956 a_20202_43084# a_13258_32519# 0.685083f
C2957 a_5257_43370# a_5147_45002# 0.836149f
C2958 a_19466_46812# a_20107_45572# 0.283769f
C2959 a_17737_43940# a_17973_43940# 0.22264f
C2960 a_n2840_42282# VDD 0.294987f
C2961 a_20202_43084# a_20193_45348# 0.116706f
C2962 a_584_46384# a_n2293_46634# 0.374996f
C2963 a_12465_44636# a_22223_47212# 0.175138f
C2964 a_4915_47217# a_13747_46662# 0.710704f
C2965 a_n4064_39616# C9_P_btm 0.215899f
C2966 a_7754_39964# a_7754_38470# 0.241119f
C2967 a_3754_39134# a_3754_38802# 0.296258f
C2968 a_n443_42852# a_742_44458# 0.168627f
C2969 a_413_45260# RST_Z 0.199496f
C2970 a_327_44734# VDD 0.667364f
C2971 a_13661_43548# a_15227_44166# 0.805606f
C2972 a_5907_46634# a_5732_46660# 0.233657f
C2973 VREF VCM 45.073803f
C2974 a_15095_43370# a_5342_30871# 0.238762f
C2975 a_9290_44172# a_13667_43396# 0.136018f
C2976 a_1307_43914# a_2779_44458# 0.332183f
C2977 a_13857_44734# VDD 0.18416f
C2978 a_1847_42826# a_2351_42308# 0.120686f
C2979 a_n443_42852# a_n901_43156# 0.367747f
C2980 a_2437_43646# a_n97_42460# 0.201806f
C2981 a_16979_44734# a_17061_44734# 0.171361f
C2982 a_n3674_39304# a_n4064_39072# 0.539144f
C2983 a_n1809_43762# VDD 0.142403f
C2984 a_3177_46902# VDD 0.200982f
C2985 a_n2017_45002# a_18249_42858# 0.545311f
C2986 a_n1059_45260# a_17333_42852# 0.270324f
C2987 a_133_42852# VDD 0.184203f
C2988 a_n4318_37592# a_n4209_37414# 0.105251f
C2989 a_3483_46348# a_5111_44636# 0.340106f
C2990 a_19553_46090# VDD 0.204238f
C2991 a_n237_47217# a_4883_46098# 0.181672f
C2992 en_comp a_7174_31319# 5.65154f
C2993 a_13259_45724# a_11691_44458# 0.337184f
C2994 a_4883_46098# a_8270_45546# 0.278829f
C2995 a_10227_46804# a_12816_46660# 0.253017f
C2996 a_n2438_43548# a_2107_46812# 0.111283f
C2997 a_n133_46660# a_948_46660# 0.102355f
C2998 a_33_46660# a_383_46660# 0.20669f
C2999 C10_P_btm C0_dummy_P_btm 0.63636f
C3000 C6_P_btm C3_P_btm 0.134599f
C3001 C7_P_btm C2_P_btm 0.139982f
C3002 C5_P_btm C4_P_btm 15.915401f
C3003 C9_P_btm C0_P_btm 0.14782f
C3004 C8_P_btm C1_P_btm 0.131002f
C3005 EN_VIN_BSTR_N C3_N_btm 0.100325f
C3006 a_16243_43396# a_15743_43084# 0.600668f
C3007 a_18114_32519# VREF_GND 0.493553f
C3008 a_4223_44672# VDD 2.99073f
C3009 a_n971_45724# a_2711_45572# 0.214535f
C3010 a_18249_42858# a_19164_43230# 0.118759f
C3011 a_13259_45724# a_4190_30871# 0.271537f
C3012 a_15493_43940# VDD 1.4617f
C3013 a_584_46384# a_626_44172# 0.450256f
C3014 a_1067_42314# a_1184_42692# 0.147283f
C3015 a_n357_42282# a_n473_42460# 0.179066f
C3016 a_22485_44484# a_22591_44484# 0.15878f
C3017 a_n3674_39304# VDD 0.587205f
C3018 a_n3674_38680# a_n3420_39072# 0.172947f
C3019 a_12549_44172# a_14539_43914# 0.110516f
C3020 a_n2438_43548# a_n2661_44458# 0.136664f
C3021 a_n2472_45546# a_n2293_45546# 0.171197f
C3022 a_12741_44636# VDD 0.988199f
C3023 a_n2109_47186# a_1209_47178# 0.226908f
C3024 a_n452_47436# a_n971_45724# 0.330438f
C3025 a_n4209_39590# a_n3565_39590# 6.15218f
C3026 a_n4064_40160# a_n4064_39616# 5.80394f
C3027 a_3065_45002# a_3318_42354# 0.146272f
C3028 en_comp a_5932_42308# 0.233106f
C3029 a_9313_44734# a_13887_32519# 0.191376f
C3030 a_5742_30871# VDD 0.556959f
C3031 a_5934_30871# VCM 0.121361f
C3032 a_3316_45546# a_3065_45002# 0.141454f
C3033 a_15227_44166# a_11967_42832# 0.132673f
C3034 a_n881_46662# a_13747_46662# 0.550574f
C3035 a_n2302_37984# VDD 0.350854f
C3036 a_3726_37500# CAL_P 0.102027f
C3037 a_7276_45260# a_6709_45028# 0.215102f
C3038 a_n2293_42834# VDD 0.853754f
C3039 a_6755_46942# a_11901_46660# 0.587021f
C3040 a_16327_47482# a_19900_46494# 0.216811f
C3041 a_n2661_46634# a_11415_45002# 0.494836f
C3042 a_1115_44172# VDD 0.165092f
C3043 a_12549_44172# a_12427_45724# 0.152925f
C3044 a_765_45546# a_17957_46116# 0.133328f
C3045 a_1176_45822# a_1138_42852# 0.41217f
C3046 a_n746_45260# a_n2661_45010# 0.400342f
C3047 a_3160_47472# VDD 0.256092f
C3048 a_n1925_42282# a_n784_42308# 0.235613f
C3049 a_18479_45785# a_19268_43646# 0.12682f
C3050 a_3483_46348# a_9049_44484# 0.117501f
C3051 a_13607_46688# VDD 0.209568f
C3052 a_22485_44484# a_20974_43370# 0.101193f
C3053 a_526_44458# a_3232_43370# 0.461444f
C3054 a_11322_45546# a_11823_42460# 0.133185f
C3055 a_12741_44636# a_11827_44484# 0.305294f
C3056 a_2324_44458# a_1423_45028# 0.154419f
C3057 a_18479_47436# a_20935_43940# 0.207572f
C3058 a_16375_45002# VDD 1.14948f
C3059 a_11599_46634# a_n881_46662# 0.100714f
C3060 a_11459_47204# a_11309_47204# 0.183357f
C3061 a_n746_45260# a_171_46873# 0.120194f
C3062 VDAC_Pi a_3754_38470# 0.389564f
C3063 a_3422_30871# a_21671_42860# 0.199876f
C3064 a_n2472_45002# a_n2293_45010# 0.177252f
C3065 a_413_45260# VDD 1.203f
C3066 a_n2497_47436# a_2324_44458# 0.796031f
C3067 a_13661_43548# a_18834_46812# 0.1407f
C3068 a_n443_46116# a_4419_46090# 0.20069f
C3069 VREF VREF_GND 45.064804f
C3070 VIN_N VCM 1.7189f
C3071 a_15095_43370# a_15279_43071# 0.105784f
C3072 a_n97_42460# a_13291_42460# 0.419357f
C3073 a_526_44458# a_4905_42826# 0.202895f
C3074 a_n1925_42282# a_3080_42308# 0.897997f
C3075 a_1307_43914# a_11341_43940# 2.31482f
C3076 a_n4318_38680# a_n3420_39072# 0.310238f
C3077 a_1823_45246# a_n2661_45546# 0.181403f
C3078 a_22612_30879# a_413_45260# 0.11791f
C3079 a_2609_46660# VDD 0.312974f
C3080 a_n2017_45002# a_17333_42852# 0.314084f
C3081 a_3483_46348# a_5147_45002# 0.363215f
C3082 a_n755_45592# a_7499_43078# 0.157526f
C3083 a_15227_44166# a_18315_45260# 0.272047f
C3084 a_18985_46122# VDD 0.253642f
C3085 a_6151_47436# a_12861_44030# 0.39397f
C3086 a_n3420_38528# a_n4064_38528# 8.203589f
C3087 a_14401_32519# a_20974_43370# 0.118041f
C3088 a_10807_43548# a_10695_43548# 0.159782f
C3089 a_8746_45002# a_8953_45002# 0.257529f
C3090 a_n1613_43370# a_6031_43396# 0.308901f
C3091 a_10227_46804# a_10341_43396# 0.188948f
C3092 a_2324_44458# a_6109_44484# 0.101116f
C3093 a_16327_47482# a_3090_45724# 1.00134f
C3094 a_10227_46804# a_12991_46634# 0.349162f
C3095 a_n743_46660# a_2107_46812# 0.72755f
C3096 a_33_46660# a_601_46902# 0.17072f
C3097 C6_P_btm C4_P_btm 0.145942f
C3098 C7_P_btm C3_P_btm 0.136068f
C3099 C10_P_btm C0_P_btm 0.251079f
C3100 C9_P_btm C1_P_btm 0.133953f
C3101 C8_P_btm C2_P_btm 0.14124f
C3102 EN_VIN_BSTR_N C2_N_btm 0.118072f
C3103 a_n2661_42282# a_n2840_42282# 0.173771f
C3104 a_2779_44458# VDD 0.38604f
C3105 a_n4318_39768# a_n4209_39590# 0.105246f
C3106 a_15559_46634# a_13059_46348# 0.167936f
C3107 a_18817_42826# a_18599_43230# 0.209641f
C3108 a_5111_42852# a_5193_42852# 0.171361f
C3109 a_22223_43948# VDD 0.254313f
C3110 a_10903_43370# a_13351_46090# 0.181897f
C3111 a_n784_42308# a_1606_42308# 15.027599f
C3112 a_n913_45002# a_4361_42308# 0.250497f
C3113 a_n13_43084# VDD 0.260551f
C3114 a_n2472_45546# a_n2956_38216# 0.157892f
C3115 a_3090_45724# a_14537_43396# 0.530123f
C3116 a_20202_43084# a_2437_43646# 0.129143f
C3117 a_20820_30879# VDD 0.719502f
C3118 a_n4209_39590# a_n4334_39616# 0.25243f
C3119 a_15493_43396# a_19319_43548# 0.120111f
C3120 a_n913_45002# a_6761_42308# 0.350952f
C3121 a_11323_42473# VDD 0.205172f
C3122 a_10227_46804# a_n97_42460# 0.18445f
C3123 a_n4064_37984# VDD 1.70621f
C3124 a_22521_40599# a_22469_40625# 1.99151f
C3125 a_7276_45260# a_7229_43940# 0.322065f
C3126 a_16327_47482# a_20075_46420# 0.270434f
C3127 a_1799_45572# a_765_45546# 0.225248f
C3128 a_3080_42308# a_1606_42308# 4.87174f
C3129 a_644_44056# VDD 0.147321f
C3130 a_2063_45854# a_2437_43646# 0.392331f
C3131 a_1431_47204# DATA[1] 0.334099f
C3132 a_2905_45572# VDD 1.22598f
C3133 a_16922_45042# a_14021_43940# 0.11663f
C3134 a_1307_43914# a_n97_42460# 0.23336f
C3135 a_3232_43370# a_3626_43646# 0.204337f
C3136 a_7499_43078# a_10083_42826# 0.375624f
C3137 a_3483_46348# a_7499_43078# 0.207714f
C3138 a_12816_46660# VDD 0.293798f
C3139 a_20753_42852# VDD 0.193909f
C3140 a_n784_42308# C0_P_btm 0.281635f
C3141 a_n2497_47436# a_n2267_43396# 0.222725f
C3142 a_2063_45854# a_n2661_46634# 1.75382f
C3143 a_4915_47217# a_5807_45002# 0.766023f
C3144 a_7754_40130# a_7754_38470# 0.111791f
C3145 a_7754_39300# a_7754_38968# 0.296258f
C3146 a_3422_30871# a_21195_42852# 0.289298f
C3147 a_n2661_45010# a_n2293_45010# 0.400159f
C3148 a_n37_45144# VDD 0.138f
C3149 a_10227_46804# a_11415_45002# 0.139042f
C3150 a_4955_46873# a_5072_46660# 0.17431f
C3151 VIN_N VREF_GND 16.4969f
C3152 VIN_P VCM 1.7189f
C3153 a_12281_43396# a_12089_42308# 0.210903f
C3154 a_22223_43396# a_13887_32519# 0.154411f
C3155 a_1307_43914# a_742_44458# 0.355379f
C3156 a_n913_45002# a_5891_43370# 0.255618f
C3157 a_13213_44734# VDD 0.184239f
C3158 a_15227_44166# a_3483_46348# 0.595533f
C3159 a_6755_46942# a_15682_46116# 0.116442f
C3160 a_104_43370# VDD 0.252393f
C3161 a_n2438_43548# a_n2017_45002# 0.29197f
C3162 a_2443_46660# VDD 0.413663f
C3163 a_5934_30871# a_8515_42308# 0.222946f
C3164 a_2324_44458# a_3357_43084# 0.216574f
C3165 a_9290_44172# a_n913_45002# 0.632534f
C3166 a_n357_42282# a_7499_43078# 0.259858f
C3167 a_15227_44166# a_17719_45144# 0.187414f
C3168 a_4185_45028# a_3537_45260# 1.06643f
C3169 a_18819_46122# VDD 0.453432f
C3170 a_6151_47436# a_13717_47436# 0.17202f
C3171 a_n2288_47178# a_n2312_40392# 0.153632f
C3172 a_n3420_38528# a_n2946_38778# 0.236674f
C3173 a_11823_42460# a_6171_45002# 0.123118f
C3174 a_16223_45938# VDD 0.132317f
C3175 a_10227_46804# a_12251_46660# 0.188053f
C3176 a_n133_46660# a_383_46660# 0.105995f
C3177 a_n881_46662# a_5257_43370# 0.447042f
C3178 a_2063_45854# a_765_45546# 1.71006f
C3179 C6_P_btm C5_P_btm 18.2841f
C3180 C7_P_btm C4_P_btm 0.148546f
C3181 C10_P_btm C1_P_btm 0.204172f
C3182 C9_P_btm C2_P_btm 0.144261f
C3183 C8_P_btm C3_P_btm 0.13616f
C3184 EN_VIN_BSTR_N C1_N_btm 0.110046f
C3185 a_16409_43396# a_17324_43396# 0.118759f
C3186 a_949_44458# VDD 1.2275f
C3187 a_584_46384# a_n443_42852# 1.36389f
C3188 a_10227_46804# a_13259_45724# 0.335001f
C3189 a_15368_46634# a_13059_46348# 0.101997f
C3190 a_18249_42858# a_18599_43230# 0.210876f
C3191 a_18083_42858# a_19164_43230# 0.101963f
C3192 a_7765_42852# a_8292_43218# 0.157652f
C3193 a_526_44458# a_2075_43172# 0.227071f
C3194 a_10193_42453# a_3626_43646# 0.13905f
C3195 a_11341_43940# VDD 1.23655f
C3196 a_10903_43370# a_12594_46348# 0.169312f
C3197 a_584_46384# a_375_42282# 0.480677f
C3198 COMP_P a_1239_39587# 0.388733f
C3199 a_n1076_43230# VDD 0.292942f
C3200 a_768_44030# a_13720_44458# 0.178939f
C3201 a_n2661_45546# a_n2956_38216# 0.15505f
C3202 a_20202_43084# a_21513_45002# 0.13666f
C3203 a_22591_46660# VDD 0.251892f
C3204 a_21076_30879# C8_N_btm 0.384801f
C3205 a_n2109_47186# a_n785_47204# 0.43597f
C3206 a_n815_47178# a_n452_47436# 0.107449f
C3207 a_18451_43940# a_18533_43940# 0.171361f
C3208 a_10723_42308# VDD 0.223902f
C3209 a_6123_31319# VCM 0.144585f
C3210 a_12549_44172# a_768_44030# 0.490163f
C3211 a_n881_46662# a_5807_45002# 0.243322f
C3212 a_n2946_37984# VDD 0.38275f
C3213 a_20974_43370# a_5649_42852# 0.186094f
C3214 a_6431_45366# a_6709_45028# 0.112564f
C3215 a_8696_44636# a_11691_44458# 0.141053f
C3216 a_6755_46942# a_11735_46660# 0.61229f
C3217 a_n881_46662# a_3699_46348# 0.203393f
C3218 a_16327_47482# a_19335_46494# 0.155998f
C3219 a_175_44278# VDD 0.20887f
C3220 a_17339_46660# a_18189_46348# 0.170772f
C3221 a_765_45546# a_17715_44484# 0.117636f
C3222 a_584_46384# a_2437_43646# 0.302508f
C3223 a_1208_46090# a_1176_45822# 0.141891f
C3224 a_12089_42308# a_11551_42558# 0.109508f
C3225 a_11827_44484# a_11341_43940# 0.231114f
C3226 a_n356_44636# a_1414_42308# 0.179164f
C3227 a_10341_43396# VDD 0.401264f
C3228 a_10903_43370# a_2711_45572# 0.213719f
C3229 a_3483_46348# a_8568_45546# 0.137016f
C3230 a_n1151_42308# a_n23_44458# 0.101137f
C3231 a_12991_46634# VDD 0.357655f
C3232 a_9313_44734# a_8685_43396# 0.124273f
C3233 a_10490_45724# a_12427_45724# 0.108721f
C3234 a_18597_46090# a_19862_44208# 0.536021f
C3235 a_3483_46348# a_n2661_43370# 0.953959f
C3236 a_11322_45546# a_11962_45724# 0.270736f
C3237 a_11525_45546# a_11652_45724# 0.138143f
C3238 a_n2497_47436# a_n2129_43609# 0.216536f
C3239 a_n237_47217# a_n743_46660# 0.192378f
C3240 a_11031_47542# a_11309_47204# 0.110775f
C3241 a_n3565_39590# C8_P_btm 0.384801f
C3242 VDAC_Pi VDAC_Ni 3.18068f
C3243 a_4699_43561# a_3539_42460# 0.109444f
C3244 a_n743_46660# a_8270_45546# 0.274248f
C3245 a_11453_44696# a_20273_46660# 0.545219f
C3246 a_4817_46660# a_5732_46660# 0.118759f
C3247 VIN_N VREF 0.775904f
C3248 VIN_P VREF_GND 16.4969f
C3249 a_n1925_42282# a_4235_43370# 0.199349f
C3250 a_327_44734# a_n23_44458# 0.141544f
C3251 a_n1059_45260# a_5891_43370# 0.186322f
C3252 a_9290_44172# a_9145_43396# 0.103991f
C3253 a_n2293_43922# VDD 0.735248f
C3254 a_6755_46942# a_2324_44458# 0.155169f
C3255 a_n863_45724# a_2905_42968# 0.269475f
C3256 a_14539_43914# a_14673_44172# 0.205935f
C3257 a_n97_42460# VDD 3.61113f
C3258 a_n2661_46098# VDD 0.979859f
C3259 a_7542_44172# a_7845_44172# 0.137004f
C3260 a_n2017_45002# a_17701_42308# 0.132871f
C3261 a_17957_46116# VDD 0.138777f
C3262 a_6575_47204# a_9067_47204# 0.210614f
C3263 a_2063_45854# a_10227_46804# 0.186188f
C3264 a_n2497_47436# a_n2312_40392# 0.194574f
C3265 a_n3565_38502# a_n4064_38528# 0.228245f
C3266 a_10807_43548# a_9145_43396# 0.290878f
C3267 a_10180_45724# a_8953_45002# 0.107499f
C3268 a_12861_44030# a_15227_44166# 0.810382f
C3269 a_10227_46804# a_12469_46902# 0.181535f
C3270 a_n1925_46634# a_2107_46812# 1.12874f
C3271 a_171_46873# a_33_46660# 0.207108f
C3272 C7_P_btm C5_P_btm 0.15419f
C3273 C10_P_btm C2_P_btm 0.215144f
C3274 C9_P_btm C3_P_btm 0.138859f
C3275 C8_P_btm C4_P_btm 0.149948f
C3276 VDAC_P VCM 10.716001f
C3277 EN_VIN_BSTR_N C0_N_btm 0.12803f
C3278 a_16977_43638# a_16759_43396# 0.209641f
C3279 a_742_44458# VDD 1.3845f
C3280 a_n443_46116# a_n755_45592# 0.651643f
C3281 a_14976_45028# a_13059_46348# 0.209989f
C3282 a_18249_42858# a_18817_42826# 0.16939f
C3283 a_n443_42852# a_14205_43396# 0.118229f
C3284 a_526_44458# a_1847_42826# 0.154735f
C3285 a_7229_43940# a_7281_43914# 0.164835f
C3286 a_21115_43940# VDD 0.145936f
C3287 a_10903_43370# a_12005_46116# 0.277468f
C3288 a_n863_45724# a_n784_42308# 0.358682f
C3289 a_n901_43156# VDD 0.475947f
C3290 a_n1630_35242# a_n4209_39590# 0.12484f
C3291 a_768_44030# a_13076_44458# 0.132449f
C3292 a_n2810_45572# a_n2956_38216# 6.20057f
C3293 a_8199_44636# a_8696_44636# 0.265919f
C3294 a_11415_45002# VDD 1.84504f
C3295 a_20193_45348# a_22165_42308# 0.252856f
C3296 a_10533_42308# VDD 0.216201f
C3297 a_12891_46348# a_768_44030# 0.193145f
C3298 a_4791_45118# a_5257_43370# 0.36404f
C3299 a_n3420_37984# VDD 0.930532f
C3300 a_n881_46662# a_3483_46348# 0.5947f
C3301 a_16327_47482# a_19553_46090# 0.172776f
C3302 a_13507_46334# a_13351_46090# 0.214666f
C3303 a_1307_43914# a_n2661_42834# 3.43601f
C3304 a_13556_45296# a_15433_44458# 0.1084f
C3305 a_n913_45002# a_3422_30871# 0.145467f
C3306 a_n984_44318# VDD 0.281427f
C3307 a_n881_46662# a_14495_45572# 0.170589f
C3308 a_2553_47502# VDD 0.150286f
C3309 a_3232_43370# a_2982_43646# 0.416054f
C3310 a_9885_43646# VDD 0.190473f
C3311 a_12251_46660# VDD 0.195617f
C3312 a_526_44458# a_5111_44636# 0.338508f
C3313 a_11415_45002# a_11827_44484# 0.169126f
C3314 a_10490_45724# a_11962_45724# 0.114064f
C3315 a_10193_42453# a_11823_42460# 0.235429f
C3316 a_n2497_47436# a_n2433_43396# 0.173242f
C3317 a_11322_45546# a_11652_45724# 0.26844f
C3318 a_13259_45724# VDD 2.41738f
C3319 a_13487_47204# a_n881_46662# 0.108977f
C3320 a_4791_45118# a_5807_45002# 0.129041f
C3321 a_7754_39964# VDAC_Ni 0.207118f
C3322 a_7754_40130# a_3754_38470# 0.191861f
C3323 a_8696_44636# a_16751_45260# 0.265287f
C3324 a_n467_45028# VDD 0.385804f
C3325 a_13747_46662# a_15368_46634# 0.110984f
C3326 a_5807_45002# a_16292_46812# 0.202526f
C3327 a_n1151_42308# a_5204_45822# 0.487224f
C3328 a_5385_46902# a_5167_46660# 0.209641f
C3329 a_19321_45002# a_3090_45724# 0.163821f
C3330 a_n2661_46634# a_11813_46116# 0.162517f
C3331 VIN_P VREF 0.775904f
C3332 a_5649_42852# a_22223_43396# 0.165664f
C3333 a_14579_43548# a_15279_43071# 0.108607f
C3334 a_13678_32519# a_13887_32519# 10.751599f
C3335 a_n2661_43922# VDD 0.611934f
C3336 a_4915_47217# a_13249_42308# 0.161597f
C3337 a_8270_45546# a_9290_44172# 0.433963f
C3338 a_n443_42852# a_n1853_43023# 0.141267f
C3339 a_n3674_39304# a_n3565_39304# 0.128699f
C3340 a_n447_43370# VDD 0.204801f
C3341 a_3080_42308# C2_P_btm 0.108823f
C3342 a_1799_45572# VDD 0.381212f
C3343 a_n1059_45260# a_16795_42852# 0.182174f
C3344 a_1823_45246# a_3232_43370# 0.344002f
C3345 a_3483_46348# a_3537_45260# 0.605469f
C3346 a_18189_46348# VDD 0.211855f
C3347 a_1343_38525# a_2113_38308# 0.325474f
C3348 a_n4334_38528# a_n4064_38528# 0.449049f
C3349 a_n3690_38528# a_n3420_38528# 0.431104f
C3350 a_n3565_38502# a_n2946_38778# 0.406164f
C3351 a_n4209_38502# a_n2302_38778# 0.406492f
C3352 a_20512_43084# a_5649_42852# 0.141324f
C3353 a_19431_45546# a_19256_45572# 0.233657f
C3354 a_12861_44030# a_15681_43442# 0.137136f
C3355 a_10227_46804# a_15095_43370# 0.264777f
C3356 a_17478_45572# VDD 0.411207f
C3357 a_11599_46634# a_15368_46634# 0.320705f
C3358 a_n133_46660# a_33_46660# 0.580914f
C3359 C7_P_btm C6_P_btm 20.5296f
C3360 C8_P_btm C5_P_btm 0.148944f
C3361 C10_P_btm C3_P_btm 0.208539f
C3362 C9_P_btm C4_P_btm 0.1579f
C3363 VDAC_P VREF_GND 0.327446f
C3364 a_22609_38406# VDD 0.317066f
C3365 CAL_P RST_Z 0.551895f
C3366 a_16409_43396# a_16759_43396# 0.20669f
C3367 a_16243_43396# a_17324_43396# 0.102355f
C3368 a_1823_45246# a_4905_42826# 0.110836f
C3369 a_4646_46812# a_7765_42852# 0.122773f
C3370 a_n3674_39768# a_n4064_40160# 0.139482f
C3371 a_n452_44636# VDD 0.112149f
C3372 a_3090_45724# a_13059_46348# 0.167043f
C3373 a_n443_46116# a_n357_42282# 0.153614f
C3374 a_18083_42858# a_18599_43230# 0.113784f
C3375 a_10193_42453# a_2982_43646# 0.231527f
C3376 a_11827_44484# a_n2661_43922# 0.32722f
C3377 a_20935_43940# VDD 0.184334f
C3378 a_5937_45572# a_2324_44458# 0.407894f
C3379 a_584_46384# a_1307_43914# 0.314947f
C3380 a_3090_45724# a_3218_45724# 0.100752f
C3381 a_12465_44636# CLK 0.795478f
C3382 a_2747_46873# VDD 0.626468f
C3383 a_n2293_43922# a_n2661_42282# 0.133253f
C3384 a_n1641_43230# VDD 0.203991f
C3385 a_13507_46334# a_9313_44734# 0.145766f
C3386 a_20202_43084# VDD 0.987622f
C3387 a_n2109_47186# a_n237_47217# 0.730469f
C3388 a_n1741_47186# a_n971_45724# 0.157081f
C3389 a_n913_45002# a_5932_42308# 0.220872f
C3390 a_n357_42282# a_3537_45260# 0.200175f
C3391 a_12891_46348# a_12549_44172# 0.309821f
C3392 a_n2312_39304# a_n2442_46660# 0.15211f
C3393 a_n3690_38304# VDD 0.363068f
C3394 a_n356_44636# a_5742_30871# 0.120133f
C3395 a_n97_42460# a_16823_43084# 0.205258f
C3396 a_10193_42453# a_14539_43914# 0.278963f
C3397 a_526_44458# a_3905_42865# 0.321601f
C3398 a_5837_45028# VDD 0.191549f
C3399 a_10249_46116# a_11186_47026# 0.172467f
C3400 a_12861_44030# a_10809_44734# 0.156561f
C3401 a_9482_43914# a_15433_44458# 0.20244f
C3402 a_13556_45296# a_14815_43914# 0.378519f
C3403 a_n809_44244# VDD 0.47719f
C3404 a_472_46348# a_1176_45822# 0.146555f
C3405 a_2063_45854# VDD 3.60498f
C3406 a_8953_45546# a_9223_42460# 0.166987f
C3407 a_14955_43396# VDD 0.401358f
C3408 a_12469_46902# VDD 0.203316f
C3409 a_14113_42308# a_16522_42674# 0.183181f
C3410 a_3600_43914# a_3737_43940# 0.126609f
C3411 a_18479_47436# a_19862_44208# 0.138185f
C3412 a_14383_46116# VDD 0.132317f
C3413 a_n971_45724# a_n743_46660# 0.122713f
C3414 a_9313_45822# a_9804_47204# 0.171044f
C3415 a_12861_44030# a_n881_46662# 0.135351f
C3416 a_n3420_37984# a_n4064_37440# 7.43287f
C3417 a_n2840_45002# a_n2661_45010# 0.189331f
C3418 a_4651_46660# a_5732_46660# 0.102355f
C3419 a_n1925_46634# a_8270_45546# 0.109762f
C3420 a_n1151_42308# a_5164_46348# 0.110485f
C3421 a_n1741_47186# a_12594_46348# 0.150956f
C3422 a_4817_46660# a_5167_46660# 0.218775f
C3423 a_526_44458# a_4093_43548# 0.107158f
C3424 a_1423_45028# a_n2661_44458# 0.164701f
C3425 a_n2661_42834# VDD 1.00348f
C3426 a_6755_46942# a_15015_46420# 0.133517f
C3427 a_n863_45724# a_1847_42826# 0.216819f
C3428 a_n1352_43396# VDD 0.288329f
C3429 a_n2497_47436# a_n2661_44458# 0.138848f
C3430 a_6123_31319# a_5934_30871# 15.8951f
C3431 a_n2293_42282# VDD 0.464485f
C3432 a_15227_44166# a_16922_45042# 0.533576f
C3433 a_17715_44484# VDD 0.526119f
C3434 a_1736_39043# a_2684_37794# 0.193802f
C3435 a_n4209_38502# a_n4064_38528# 0.265711f
C3436 a_n3565_38502# a_n3420_38528# 0.278952f
C3437 a_10227_46804# a_14205_43396# 0.422372f
C3438 a_15861_45028# VDD 0.690795f
C3439 a_12861_44030# a_17609_46634# 0.183853f
C3440 a_n2438_43548# a_33_46660# 0.588568f
C3441 a_n133_46660# a_171_46873# 0.163873f
C3442 C9_P_btm C5_P_btm 0.153949f
C3443 C10_P_btm C4_P_btm 0.348092f
C3444 C8_P_btm C6_P_btm 0.170091f
C3445 VDAC_N VCM 10.717099f
C3446 CAL_P VDD 22.4716f
C3447 VDAC_P VREF 0.254986f
C3448 a_16409_43396# a_16977_43638# 0.17072f
C3449 a_15227_44166# a_15743_43084# 0.513622f
C3450 a_4646_46812# a_7871_42858# 0.26422f
C3451 a_n4318_39768# a_n4064_40160# 0.293052f
C3452 a_n1352_44484# VDD 0.276725f
C3453 a_17333_42852# a_18249_42858# 0.311255f
C3454 a_20623_43914# VDD 0.258478f
C3455 a_8199_44636# a_2324_44458# 0.412215f
C3456 a_3090_45724# a_2957_45546# 0.167712f
C3457 a_564_42282# a_n1630_35242# 0.156633f
C3458 a_n1423_42826# VDD 0.211036f
C3459 a_12891_46348# a_13076_44458# 0.182315f
C3460 a_768_44030# a_12607_44458# 0.215512f
C3461 a_10586_45546# a_2711_45572# 0.295169f
C3462 a_526_44458# a_7499_43078# 0.2203f
C3463 a_22365_46825# VDD 0.193587f
C3464 a_n2109_47186# a_n746_45260# 0.295988f
C3465 a_9885_42558# VDD 0.18767f
C3466 a_n2312_40392# a_n2442_46660# 5.91846f
C3467 a_n3565_38216# VDD 0.901259f
C3468 a_n2293_43922# a_5379_42460# 0.4571f
C3469 a_20974_43370# a_4361_42308# 0.122936f
C3470 a_3232_43370# a_7229_43940# 0.180766f
C3471 a_n1613_43370# a_8952_43230# 0.213002f
C3472 a_5093_45028# VDD 0.168437f
C3473 a_n1151_42308# a_5066_45546# 0.5423f
C3474 a_16327_47482# a_18819_46122# 0.324239f
C3475 a_n1557_42282# a_n1630_35242# 0.865968f
C3476 a_14579_43548# a_14635_42282# 0.124652f
C3477 a_n1549_44318# VDD 0.200608f
C3478 a_n743_46660# a_2711_45572# 0.525746f
C3479 a_584_46384# VDD 2.50905f
C3480 a_327_47204# DATA[0] 0.353891f
C3481 a_15095_43370# VDD 0.169652f
C3482 a_11901_46660# VDD 0.57548f
C3483 a_14097_32519# VDD 0.284675f
C3484 a_12741_44636# a_18494_42460# 0.114105f
C3485 a_21496_47436# a_4883_46098# 0.257837f
C3486 a_n4209_39590# C9_P_btm 0.786375f
C3487 a_3877_44458# a_6540_46812# 0.244975f
C3488 a_13507_46334# a_22000_46634# 0.183978f
C3489 a_n1741_47186# a_12005_46116# 0.174477f
C3490 a_13661_43548# a_14976_45028# 0.162789f
C3491 a_13747_46662# a_3090_45724# 0.139869f
C3492 a_4817_46660# a_5385_46902# 0.170485f
C3493 a_13678_32519# a_5649_42852# 0.506367f
C3494 a_2063_45854# a_10907_45822# 0.22153f
C3495 a_21363_46634# a_21188_46660# 0.233657f
C3496 a_n863_45724# a_791_42968# 0.338631f
C3497 a_n1177_43370# VDD 0.354704f
C3498 a_768_44030# a_3232_43370# 0.224083f
C3499 a_15368_46634# a_15143_45578# 0.105334f
C3500 a_n2438_43548# a_n2661_45010# 0.220364f
C3501 a_6123_31319# a_7963_42308# 0.192155f
C3502 a_n913_45002# a_5342_30871# 0.122483f
C3503 a_22959_42860# VDD 0.30747f
C3504 a_3090_45724# a_18911_45144# 0.190188f
C3505 a_13507_46334# a_20512_43084# 0.497215f
C3506 a_17583_46090# VDD 0.23578f
C3507 a_n3565_38502# a_n3690_38528# 0.246863f
C3508 a_n2293_43922# a_12089_42308# 0.183316f
C3509 a_16327_47482# a_10341_43396# 0.159266f
C3510 a_9290_44172# a_9313_44734# 0.140741f
C3511 a_8696_44636# VDD 1.12228f
C3512 a_4915_47217# a_13885_46660# 0.179458f
C3513 a_10227_46804# a_11735_46660# 0.54163f
C3514 a_11599_46634# a_3090_45724# 0.133107f
C3515 C10_P_btm C5_P_btm 0.285351f
C3516 C9_P_btm C6_P_btm 0.169882f
C3517 C8_P_btm C7_P_btm 23.7884f
C3518 VDAC_N VREF_GND 0.327524f
C3519 a_16243_43396# a_16759_43396# 0.106647f
C3520 a_n1177_44458# VDD 0.347966f
C3521 a_2107_46812# a_9625_46129# 0.184645f
C3522 a_3877_44458# a_1823_45246# 0.231164f
C3523 a_n443_46116# a_n1099_45572# 0.368941f
C3524 a_18083_42858# a_18249_42858# 0.699797f
C3525 a_12883_44458# a_13076_44458# 0.142643f
C3526 a_12607_44458# a_13720_44458# 0.122704f
C3527 a_20365_43914# VDD 0.261299f
C3528 a_18597_46090# a_n913_45002# 0.126328f
C3529 a_n2312_40392# CLK_DATA 0.213071f
C3530 COMP_P a_1606_42308# 2.6775f
C3531 a_n913_45002# a_743_42282# 0.25834f
C3532 a_n1991_42858# VDD 0.575656f
C3533 a_n2840_45546# a_n2661_45546# 0.175179f
C3534 a_768_44030# a_8975_43940# 0.124155f
C3535 a_20820_30879# C7_N_btm 0.184297f
C3536 a_n2109_47186# a_n971_45724# 1.21934f
C3537 SMPL_ON_P a_n1605_47204# 0.194856f
C3538 a_5742_30871# C6_N_btm 0.170624f
C3539 a_16327_47482# a_n97_42460# 0.113034f
C3540 a_3316_45546# a_413_45260# 0.110075f
C3541 a_7227_45028# VDD 0.501104f
C3542 a_n2312_39304# a_n2661_46634# 0.105298f
C3543 a_2063_45854# a_9863_46634# 0.10786f
C3544 a_n4334_38304# VDD 0.385989f
C3545 a_n2661_42282# a_n2293_42282# 1.04835f
C3546 a_n1613_43370# a_9127_43156# 0.267842f
C3547 a_10903_43370# a_12429_44172# 0.116356f
C3548 a_5009_45028# VDD 0.151712f
C3549 a_12861_44030# a_6945_45028# 0.108969f
C3550 a_19321_45002# a_12741_44636# 0.113088f
C3551 a_20916_46384# a_20202_43084# 0.181561f
C3552 a_n1331_43914# VDD 0.203823f
C3553 a_3422_30871# VCM 1.12142f
C3554 a_472_46348# a_805_46414# 0.360492f
C3555 a_n2497_47436# a_n2017_45002# 0.125552f
C3556 a_n2312_38680# a_n2302_38778# 0.161815f
C3557 a_n785_47204# DATA[0] 0.598846f
C3558 SMPL_ON_P VIN_P 0.587766f
C3559 a_8953_45546# a_8685_42308# 0.250058f
C3560 a_7499_43078# a_8037_42858# 0.160087f
C3561 a_14205_43396# VDD 0.311811f
C3562 a_4646_46812# a_7229_43940# 0.104864f
C3563 a_11813_46116# VDD 0.434656f
C3564 a_11823_42460# a_15051_42282# 0.367924f
C3565 a_22400_42852# VDD 0.829052f
C3566 a_10193_42453# a_11652_45724# 0.197229f
C3567 a_10490_45724# a_11322_45546# 0.246478f
C3568 a_2324_44458# a_1307_43914# 0.129761f
C3569 a_13507_46334# a_4883_46098# 4.09671f
C3570 a_n971_45724# a_n1925_46634# 0.163523f
C3571 a_9863_47436# a_9804_47204# 0.109361f
C3572 a_n3420_37984# a_n3420_37440# 0.132162f
C3573 a_13507_46334# a_5649_42852# 0.136078f
C3574 a_n2293_46634# a_9145_43396# 0.238561f
C3575 a_n967_45348# VDD 0.556063f
C3576 en_comp RST_Z 4.34313f
C3577 a_4651_46660# a_5167_46660# 0.102946f
C3578 a_16327_47482# a_11415_45002# 0.94171f
C3579 a_13661_43548# a_3090_45724# 0.177565f
C3580 a_526_44458# a_1568_43370# 0.220609f
C3581 a_9313_45822# a_9049_44484# 0.119007f
C3582 a_3090_45724# a_4185_45028# 0.770164f
C3583 a_n1917_43396# VDD 0.204644f
C3584 a_6755_46942# a_15903_45785# 0.192397f
C3585 a_10903_43370# a_10586_45546# 0.238199f
C3586 a_n356_44636# a_n97_42460# 1.46232f
C3587 a_22223_42860# VDD 0.250812f
C3588 a_15682_46116# VDD 1.25004f
C3589 a_1736_39587# a_2113_38308# 0.100626f
C3590 a_n4209_38502# a_n3420_38528# 0.230544f
C3591 a_18479_45785# a_18596_45572# 0.183223f
C3592 a_18341_45572# a_19256_45572# 0.116691f
C3593 a_10227_46804# a_14579_43548# 0.118896f
C3594 a_16680_45572# VDD 0.275078f
C3595 a_n2438_43548# a_n133_46660# 0.848709f
C3596 VDAC_P VIN_P 0.252066f
C3597 C10_P_btm C6_P_btm 0.421276f
C3598 C9_P_btm C7_P_btm 0.227839f
C3599 VDAC_N VREF 0.254986f
C3600 a_4905_42826# a_5111_42852# 0.105155f
C3601 a_16547_43609# a_16409_43396# 0.206231f
C3602 a_n913_45002# a_20193_45348# 0.224918f
C3603 a_19963_31679# a_19721_31679# 9.01086f
C3604 a_n1917_44484# VDD 0.186988f
C3605 a_16327_47482# a_13259_45724# 0.584328f
C3606 a_18083_42858# a_17333_42852# 0.284837f
C3607 a_742_44458# a_n356_44636# 0.207503f
C3608 a_12607_44458# a_13076_44458# 0.200168f
C3609 a_20269_44172# VDD 0.169009f
C3610 a_11189_46129# a_10903_43370# 0.151119f
C3611 a_22315_44484# a_22485_44484# 0.109468f
C3612 a_n1059_45260# a_743_42282# 0.198704f
C3613 a_n1853_43023# VDD 0.370563f
C3614 a_n2840_45546# a_n2810_45572# 0.162234f
C3615 a_5932_42308# VCM 0.146001f
C3616 a_3090_45724# a_11967_42832# 0.12811f
C3617 a_2107_46812# a_9028_43914# 0.110155f
C3618 a_6598_45938# VDD 0.204705f
C3619 a_n2312_39304# a_n2956_39768# 5.91067f
C3620 a_4883_46098# a_n743_46660# 5.6639f
C3621 a_n4209_38216# VDD 0.833976f
C3622 VDAC_P a_11206_38545# 0.101449f
C3623 a_21381_43940# a_4361_42308# 0.195418f
C3624 a_3232_43370# a_5205_44484# 0.217288f
C3625 a_n1613_43370# a_8387_43230# 0.163582f
C3626 a_10903_43370# a_11750_44172# 0.135933f
C3627 a_2809_45028# VDD 0.189682f
C3628 a_n443_46116# a_526_44458# 0.366438f
C3629 a_10227_46804# a_14840_46494# 0.275527f
C3630 a_2711_45572# a_19319_43548# 0.225335f
C3631 a_19479_31679# a_19237_31679# 9.049419f
C3632 a_n1899_43946# VDD 0.475205f
C3633 a_3422_30871# VREF_GND 0.10463f
C3634 a_12549_44172# a_10193_42453# 0.116594f
C3635 a_1431_47204# VDD 0.423871f
C3636 a_n2312_38680# a_n4064_38528# 0.22404f
C3637 a_n237_47217# DATA[1] 0.139838f
C3638 a_3537_45260# a_3539_42460# 0.264936f
C3639 a_14358_43442# VDD 0.170277f
C3640 a_11735_46660# VDD 0.407307f
C3641 a_11823_42460# a_14113_42308# 0.103699f
C3642 a_526_44458# a_3537_45260# 0.938783f
C3643 a_15227_44166# a_16979_44734# 0.181002f
C3644 a_13507_46334# a_21496_47436# 0.167302f
C3645 a_3754_39466# a_3754_39134# 0.296258f
C3646 a_n755_45592# a_5343_44458# 0.349527f
C3647 a_1823_45246# a_3905_42865# 0.218008f
C3648 en_comp VDD 4.26539f
C3649 a_11453_44696# a_18285_46348# 0.236771f
C3650 a_16327_47482# a_20202_43084# 0.475502f
C3651 a_4955_46873# a_4817_46660# 0.318259f
C3652 a_21855_43396# a_13678_32519# 0.17881f
C3653 a_526_44458# a_1049_43396# 0.121121f
C3654 a_10617_44484# VDD 0.141193f
C3655 a_20411_46873# a_20528_46660# 0.170785f
C3656 a_n2312_39304# a_n2302_39072# 0.130454f
C3657 a_16795_42852# a_16877_42852# 0.171361f
C3658 a_n1699_43638# VDD 0.210236f
C3659 a_7227_42308# a_6123_31319# 0.189956f
C3660 a_n913_45002# a_5534_30871# 0.274894f
C3661 a_22165_42308# VDD 0.336187f
C3662 a_12741_44636# a_9482_43914# 0.101234f
C3663 a_8953_45546# a_n1059_45260# 0.318691f
C3664 a_2324_44458# VDD 2.73366f
C3665 a_n1151_42308# a_11599_46634# 0.116147f
C3666 a_18909_45814# a_18691_45572# 0.209641f
C3667 a_16855_45546# VDD 0.339227f
C3668 a_n743_46660# a_n133_46660# 0.205551f
C3669 VDAC_N VIN_N 0.253278f
C3670 C10_P_btm C7_P_btm 0.680974f
C3671 C9_P_btm C8_P_btm 29.256199f
C3672 a_22469_39537# VDD 0.356405f
C3673 a_4905_42826# a_4520_42826# 0.147708f
C3674 a_16243_43396# a_16409_43396# 0.575934f
C3675 a_1823_45246# a_4093_43548# 0.17443f
C3676 a_n1699_44726# VDD 0.198612f
C3677 a_n443_46116# a_n452_45724# 0.188857f
C3678 a_n237_47217# a_2277_45546# 0.104529f
C3679 a_n1613_43370# a_526_44458# 0.826565f
C3680 a_n452_44636# a_n356_44636# 0.318214f
C3681 a_12607_44458# a_12883_44458# 0.11453f
C3682 a_n443_42852# a_9803_43646# 0.102893f
C3683 a_19862_44208# VDD 0.588967f
C3684 a_12549_44172# a_18479_45785# 0.105486f
C3685 a_9290_44172# a_10903_43370# 0.340316f
C3686 a_11189_46129# a_11387_46155# 0.320331f
C3687 a_n2017_45002# a_743_42282# 7.84646f
C3688 a_n2157_42858# VDD 0.424058f
C3689 a_n1741_47186# SMPL_ON_P 0.178214f
C3690 a_n2497_47436# a_n971_45724# 0.229429f
C3691 a_n2109_47186# a_n815_47178# 0.160027f
C3692 a_n4315_30879# a_n4209_39590# 4.31257f
C3693 a_9803_42558# VDD 0.253745f
C3694 a_12549_44172# a_14021_43940# 0.150377f
C3695 a_n443_42852# a_n913_45002# 0.796158f
C3696 a_6667_45809# VDD 0.195842f
C3697 a_8912_37509# a_11206_38545# 1.26605f
C3698 a_n1613_43370# a_8605_42826# 0.159791f
C3699 a_10903_43370# a_10807_43548# 0.193971f
C3700 a_n237_47217# a_8049_45260# 0.109887f
C3701 a_n881_46662# a_167_45260# 0.108232f
C3702 a_10227_46804# a_15015_46420# 0.287571f
C3703 a_n863_45724# a_1568_43370# 0.202455f
C3704 a_n2661_45546# a_3080_42308# 0.155045f
C3705 a_1138_42852# a_791_42968# 0.100783f
C3706 a_1423_45028# a_9313_44734# 0.241551f
C3707 a_n1761_44111# VDD 0.620042f
C3708 a_8270_45546# a_8049_45260# 0.321896f
C3709 a_376_46348# a_472_46348# 0.318161f
C3710 a_n2497_47436# a_n2293_45010# 0.233882f
C3711 a_16388_46812# a_17957_46116# 0.140894f
C3712 a_1239_47204# VDD 0.278979f
C3713 a_8199_44636# a_8685_42308# 0.114007f
C3714 a_7499_43078# a_7871_42858# 0.146369f
C3715 a_14579_43548# VDD 0.278225f
C3716 a_n2956_38680# a_n2956_38216# 0.10753f
C3717 a_5937_45572# a_5907_45546# 0.104991f
C3718 a_15959_42545# a_15890_42674# 0.209641f
C3719 a_13249_42308# a_13070_42354# 0.141799f
C3720 a_n913_45002# a_14635_42282# 0.332583f
C3721 a_5891_43370# a_8685_43396# 0.145735f
C3722 a_768_44030# a_5244_44056# 0.167173f
C3723 a_8746_45002# a_10490_45724# 0.116339f
C3724 a_15227_44166# a_14539_43914# 0.520312f
C3725 a_12839_46116# VDD 0.347766f
C3726 a_10586_45546# CLK 0.125859f
C3727 a_n2956_37592# VDD 1.25966f
C3728 a_2063_45854# a_5204_45822# 0.174206f
C3729 a_12549_44172# a_19692_46634# 0.491923f
C3730 a_11599_46634# a_12741_44636# 0.183316f
C3731 a_4651_46660# a_4817_46660# 0.57393f
C3732 a_n443_46116# a_167_45260# 0.794635f
C3733 a_13747_46662# a_13607_46688# 0.168294f
C3734 a_9290_44172# a_8685_43396# 0.207262f
C3735 a_20273_46660# a_21188_46660# 0.118759f
C3736 a_8270_45546# a_8953_45546# 1.06716f
C3737 a_n2267_43396# VDD 0.570924f
C3738 a_2107_46812# a_2437_43646# 0.185914f
C3739 a_768_44030# a_5111_44636# 0.154519f
C3740 a_491_47026# VDD 0.132552f
C3741 a_6761_42308# a_6123_31319# 0.187371f
C3742 a_21671_42860# VDD 0.229963f
C3743 a_5342_30871# VCM 0.325566f
C3744 a_14840_46494# VDD 0.275785f
C3745 a_6851_47204# a_7227_47204# 0.241208f
C3746 a_6545_47178# a_6575_47204# 0.11927f
C3747 a_4915_47217# a_9313_45822# 0.366722f
C3748 a_n4209_38502# a_n3565_38502# 6.84323f
C3749 a_n913_45002# a_19511_42282# 0.120073f
C3750 a_n356_44636# a_n2293_42282# 1.10197f
C3751 a_18175_45572# a_19256_45572# 0.102355f
C3752 a_18341_45572# a_18691_45572# 0.206455f
C3753 a_8270_45546# a_9028_43914# 0.233359f
C3754 a_16115_45572# VDD 0.194492f
C3755 a_n743_46660# a_n2438_43548# 0.426835f
C3756 C10_P_btm C8_P_btm 0.878696f
C3757 a_22821_38993# VDD 0.431879f
C3758 EN_VIN_BSTR_P C0_P_btm 0.12803f
C3759 a_16243_43396# a_16547_43609# 0.165289f
C3760 a_n2267_44484# VDD 0.289888f
C3761 a_11599_46634# a_16375_45002# 0.407484f
C3762 a_n237_47217# a_1609_45822# 0.141985f
C3763 a_2905_45572# a_2957_45546# 0.137248f
C3764 en_comp a_n2661_42282# 0.103098f
C3765 a_n443_42852# a_9145_43396# 2.32123f
C3766 a_19478_44306# VDD 0.127794f
C3767 a_11189_46129# a_11133_46155# 0.203074f
C3768 a_11453_44696# a_2437_43646# 0.189184f
C3769 a_n2312_39304# VDD 0.587668f
C3770 a_n1059_45260# a_4190_30871# 0.133926f
C3771 a_3422_30871# a_20512_43084# 0.125955f
C3772 a_n2472_42826# VDD 0.229608f
C3773 a_n1630_35242# a_n4315_30879# 0.129428f
C3774 a_10809_44734# a_11823_42460# 0.215753f
C3775 a_n4064_40160# a_n2302_40160# 0.249627f
C3776 a_n913_45002# a_4921_42308# 0.169235f
C3777 a_9223_42460# VDD 0.205797f
C3778 a_13661_43548# a_15493_43940# 1.28948f
C3779 a_n443_42852# a_n1059_45260# 0.130036f
C3780 a_6511_45714# VDD 0.405279f
C3781 a_n971_45724# a_6969_46634# 0.235123f
C3782 VDAC_N a_11206_38545# 0.15219f
C3783 a_8912_37509# VDAC_P 3.15325f
C3784 a_10903_43370# a_10949_43914# 0.451961f
C3785 a_3232_43370# a_6171_45002# 0.314056f
C3786 a_11599_46634# a_18985_46122# 0.570252f
C3787 a_10227_46804# a_14275_46494# 0.18614f
C3788 a_13661_43548# a_12741_44636# 0.13948f
C3789 a_4883_46098# a_10355_46116# 0.23167f
C3790 a_n2065_43946# VDD 0.4213f
C3791 a_n971_45724# a_3357_43084# 0.565799f
C3792 a_1209_47178# VDD 0.38145f
C3793 a_3065_45002# a_3539_42460# 0.300764f
C3794 a_n1925_42282# a_n2104_42282# 0.166917f
C3795 a_7499_43078# a_7227_42852# 0.126148f
C3796 a_13667_43396# VDD 0.402378f
C3797 a_584_46384# a_n356_44636# 0.268036f
C3798 a_10768_47026# VDD 0.132317f
C3799 a_5934_30871# a_7174_31319# 0.473128f
C3800 a_20202_43084# a_18494_42460# 0.166633f
C3801 a_1823_45246# a_n2661_43370# 0.112095f
C3802 a_526_44458# a_3065_45002# 0.138202f
C3803 a_n1151_42308# a_5807_45002# 1.52318f
C3804 a_6151_47436# a_12549_44172# 0.214024f
C3805 a_6575_47204# a_8128_46384# 0.105633f
C3806 a_9313_45822# a_n881_46662# 1.00227f
C3807 a_21177_47436# a_13507_46334# 0.329096f
C3808 a_7754_39632# a_7754_39300# 0.296258f
C3809 a_n755_45592# a_n699_43396# 0.185444f
C3810 a_n2810_45028# VDD 0.526631f
C3811 a_4646_46812# a_4817_46660# 0.588038f
C3812 a_4651_46660# a_4955_46873# 0.140348f
C3813 a_4361_42308# a_21855_43396# 0.167446f
C3814 a_13467_32519# a_13678_32519# 10.9526f
C3815 a_6171_45002# a_8975_43940# 0.175346f
C3816 a_3422_30871# CAL_N 0.236929f
C3817 a_13059_46348# a_11415_45002# 0.225168f
C3818 a_20841_46902# a_20623_46660# 0.209641f
C3819 a_8270_45546# a_5937_45572# 0.29626f
C3820 a_n2661_43370# a_n3674_39768# 0.144159f
C3821 a_n2129_43609# VDD 0.400674f
C3822 a_768_44030# a_5147_45002# 0.191082f
C3823 a_6761_42308# a_7227_42308# 0.173849f
C3824 a_5932_42308# a_5934_30871# 1.37963f
C3825 a_11967_42832# a_15493_43940# 0.299734f
C3826 a_5111_44636# a_5111_42852# 0.148196f
C3827 a_21195_42852# VDD 0.285496f
C3828 a_4185_45028# a_413_45260# 0.191095f
C3829 a_11415_45002# a_13556_45296# 0.16025f
C3830 a_3503_45724# a_3775_45552# 0.13675f
C3831 a_15015_46420# VDD 0.337162f
C3832 a_9290_44172# CLK 0.151406f
C3833 a_4915_47217# a_11031_47542# 0.125943f
C3834 a_n4209_38502# a_n4334_38528# 0.25243f
C3835 a_3422_30871# a_5649_42852# 0.291966f
C3836 a_10193_42453# a_6171_45002# 0.411891f
C3837 a_8746_45002# a_3232_43370# 0.439467f
C3838 a_18341_45572# a_18909_45814# 0.170692f
C3839 a_n2293_45546# a_n2661_43370# 0.131199f
C3840 a_16333_45814# VDD 0.201203f
C3841 a_n2810_45028# a_n2302_37690# 0.162246f
C3842 a_12861_44030# a_3090_45724# 0.496275f
C3843 C10_P_btm C9_P_btm 37.815998f
C3844 a_22545_38993# VDD 0.536989f
C3845 EN_VIN_BSTR_P C1_P_btm 0.110046f
C3846 a_16137_43396# a_16547_43609# 0.151161f
C3847 a_19479_31679# a_19721_31679# 9.039419f
C3848 a_n2129_44697# VDD 1.4165f
C3849 a_16795_42852# a_17333_42852# 0.108694f
C3850 a_15493_43396# VDD 2.34659f
C3851 a_12465_44636# a_3357_43084# 1.30897f
C3852 a_13059_46348# a_13259_45724# 0.812126f
C3853 a_10227_46804# a_n913_45002# 0.344574f
C3854 a_n2312_40392# VDD 0.947797f
C3855 a_n784_42308# a_n3674_37592# 0.254719f
C3856 a_n2840_42826# VDD 0.302305f
C3857 a_n1920_47178# a_n1741_47186# 0.173125f
C3858 a_8791_42308# VDD 0.226318f
C3859 a_n443_46116# a_2982_43646# 0.140614f
C3860 a_6472_45840# VDD 0.257073f
C3861 a_n971_45724# a_6755_46942# 0.185154f
C3862 a_2684_37794# VDD 0.286898f
C3863 VDAC_N VDAC_P 4.74149f
C3864 a_n913_45002# a_1307_43914# 0.298747f
C3865 a_5111_44636# a_5205_44484# 0.200189f
C3866 a_11599_46634# a_18819_46122# 0.314824f
C3867 a_10227_46804# a_14493_46090# 0.202633f
C3868 a_n881_46662# a_1823_45246# 0.155149f
C3869 a_n2472_43914# VDD 0.236691f
C3870 a_768_44030# a_7499_43078# 0.101779f
C3871 a_16327_47482# a_16680_45572# 0.223571f
C3872 a_n2497_47436# a_n2661_45010# 0.281004f
C3873 a_327_47204# VDD 0.367528f
C3874 a_n971_45724# DATA[0] 0.213213f
C3875 a_3065_45002# a_3626_43646# 0.480498f
C3876 a_10695_43548# VDD 0.201247f
C3877 a_15803_42450# a_15959_42545# 0.110532f
C3878 a_15764_42576# a_15890_42674# 0.181217f
C3879 a_2711_45572# a_20107_42308# 0.164316f
C3880 a_18707_42852# VDD 0.132317f
C3881 a_10193_42453# a_8746_45002# 0.11003f
C3882 a_20202_43084# a_18184_42460# 0.299795f
C3883 a_768_44030# a_3600_43914# 0.182408f
C3884 a_526_44458# a_2680_45002# 0.119733f
C3885 a_6151_47436# a_12891_46348# 0.169139f
C3886 a_7903_47542# a_8128_46384# 0.109077f
C3887 a_11031_47542# a_n881_46662# 0.183988f
C3888 a_n4064_40160# C10_P_btm 0.460005f
C3889 a_2113_38308# VDAC_Ni 0.315941f
C3890 a_n745_45366# VDD 0.20887f
C3891 a_3160_47472# a_3699_46348# 0.109505f
C3892 a_n443_46116# a_1823_45246# 0.217935f
C3893 a_7499_43078# a_7845_44172# 0.112307f
C3894 a_3232_43370# a_8975_43940# 0.620589f
C3895 a_20273_46660# a_20623_46660# 0.20669f
C3896 a_20107_46660# a_21188_46660# 0.102355f
C3897 a_8270_45546# a_8199_44636# 0.95539f
C3898 a_5649_42852# a_5932_42308# 0.126438f
C3899 a_17333_42852# a_18504_43218# 0.157683f
C3900 a_n2433_43396# VDD 0.416276f
C3901 a_9290_44172# a_10586_45546# 0.264957f
C3902 a_1983_46706# VDD 0.119964f
C3903 a_18579_44172# a_18451_43940# 0.147572f
C3904 a_5495_43940# a_5663_43940# 0.227135f
C3905 a_13259_45724# a_17303_42282# 0.460497f
C3906 a_21356_42826# VDD 0.225688f
C3907 a_11415_45002# a_9482_43914# 0.309633f
C3908 a_1823_45246# a_3537_45260# 0.482502f
C3909 a_14275_46494# VDD 0.196859f
C3910 a_6491_46660# a_6851_47204# 0.132946f
C3911 a_3422_30871# a_13678_32519# 0.452533f
C3912 a_18175_45572# a_18691_45572# 0.105995f
C3913 a_n2956_37592# a_n2946_37690# 0.148852f
C3914 a_15765_45572# VDD 0.249471f
C3915 a_n2810_45028# a_n4064_37440# 0.22413f
C3916 a_n237_47217# a_765_45546# 0.1364f
C3917 a_n1925_46634# a_n2438_43548# 0.166008f
C3918 a_n1021_46688# a_n743_46660# 0.11001f
C3919 a_22521_39511# VDD 0.910209f
C3920 EN_VIN_BSTR_P C2_P_btm 0.118072f
C3921 a_16137_43396# a_16243_43396# 0.182209f
C3922 a_19479_31679# a_18114_32519# 0.182316f
C3923 a_n2433_44484# VDD 0.40658f
C3924 a_15009_46634# a_14180_46812# 0.123843f
C3925 a_n746_45260# a_n443_42852# 0.136813f
C3926 a_17595_43084# a_17701_42308# 0.141211f
C3927 a_19328_44172# VDD 0.263964f
C3928 a_n746_45260# a_375_42282# 0.41439f
C3929 a_9290_44172# a_11189_46129# 0.199578f
C3930 a_6755_46942# a_2711_45572# 0.612305f
C3931 a_22959_47212# VDD 0.245964f
C3932 a_196_42282# a_n3674_37592# 0.1528f
C3933 a_14537_43396# a_14358_43442# 0.1418f
C3934 a_4190_30871# VCM 1.23535f
C3935 a_8049_45260# a_2711_45572# 2.31131f
C3936 a_n2109_47186# a_n1741_47186# 0.18579f
C3937 a_n4334_40480# a_n4064_40160# 0.43652f
C3938 a_n4315_30879# a_n2302_40160# 0.407166f
C3939 a_8685_42308# VDD 0.286875f
C3940 a_13259_45724# a_9482_43914# 0.321549f
C3941 a_19321_45002# a_20623_43914# 0.294126f
C3942 a_15227_44166# a_17517_44484# 0.104904f
C3943 a_13661_43548# a_11341_43940# 0.15891f
C3944 a_6194_45824# VDD 0.274689f
C3945 a_22959_47212# a_22612_30879# 0.156518f
C3946 a_1177_38525# VDD 0.373535f
C3947 VDAC_N a_8912_37509# 3.43288f
C3948 a_n1613_43370# a_7871_42858# 0.659491f
C3949 a_5691_45260# a_3232_43370# 0.123939f
C3950 a_n881_46662# a_1138_42852# 0.148785f
C3951 a_10227_46804# a_13925_46122# 0.635045f
C3952 a_n863_45724# a_458_43396# 0.122956f
C3953 a_n2661_45546# a_4093_43548# 0.343267f
C3954 a_9290_44172# a_4361_42308# 0.1126f
C3955 a_n2840_43914# VDD 0.304745f
C3956 a_n2293_46098# a_1823_45246# 0.107882f
C3957 a_3090_45724# a_n1925_42282# 0.157861f
C3958 a_16327_47482# a_16855_45546# 0.305145f
C3959 a_n785_47204# VDD 0.452945f
C3960 a_n2312_38680# a_n3565_38502# 0.134976f
C3961 a_2382_45260# a_3539_42460# 0.110439f
C3962 a_9803_43646# VDD 0.261557f
C3963 a_4646_46812# a_3232_43370# 0.305673f
C3964 a_n2956_38680# a_n2810_45572# 5.73878f
C3965 a_6123_31319# a_7174_31319# 13.9919f
C3966 a_15764_42576# a_15959_42545# 0.21686f
C3967 a_10949_43914# a_12429_44172# 0.156922f
C3968 a_20193_45348# a_13887_32519# 0.277027f
C3969 a_n1630_35242# a_18194_35068# 0.465356f
C3970 a_10180_45724# a_8746_45002# 0.304016f
C3971 a_16327_47482# a_19862_44208# 0.209324f
C3972 a_768_44030# a_2998_44172# 0.571981f
C3973 a_2324_44458# a_14537_43396# 0.341957f
C3974 a_4915_47217# a_768_44030# 0.187438f
C3975 a_9863_47436# a_n881_46662# 0.164043f
C3976 a_20990_47178# a_21177_47436# 0.159555f
C3977 a_15903_45785# a_16019_45002# 0.139976f
C3978 a_n913_45002# VDD 9.190901f
C3979 a_3160_47472# a_3483_46348# 0.154179f
C3980 a_4646_46812# a_4651_46660# 0.844575f
C3981 a_12549_44172# a_15227_44166# 0.354423f
C3982 a_13467_32519# a_4361_42308# 0.121732f
C3983 a_3422_30871# VDAC_P 0.476038f
C3984 a_20273_46660# a_20841_46902# 0.17072f
C3985 a_10193_42453# a_16137_43396# 0.329316f
C3986 a_n755_45592# a_n13_43084# 0.113444f
C3987 a_n4318_39304# VDD 0.643395f
C3988 a_2107_46812# VDD 0.350275f
C3989 a_5932_42308# a_6123_31319# 1.49414f
C3990 a_20922_43172# VDD 0.192467f
C3991 a_3090_45724# a_16922_45042# 0.206138f
C3992 a_14493_46090# VDD 0.203567f
C3993 a_6545_47178# a_6851_47204# 0.134581f
C3994 a_16375_45002# a_17719_45144# 0.201099f
C3995 a_9290_44172# a_5891_43370# 0.302383f
C3996 a_18479_45785# a_18341_45572# 0.21997f
C3997 a_n357_42282# a_n2293_42834# 4.06139f
C3998 a_n2956_37592# a_n3420_37440# 0.233174f
C3999 a_15903_45785# VDD 0.291109f
C4000 a_n1613_43370# a_5732_46660# 0.268372f
C4001 a_n1925_46634# a_n743_46660# 0.193773f
C4002 EN_VIN_BSTR_P C3_P_btm 0.100325f
C4003 a_n2661_44458# VDD 1.06317f
C4004 a_14084_46812# a_14180_46812# 0.318161f
C4005 a_n971_45724# a_n443_42852# 0.329303f
C4006 a_2905_45572# a_n755_45592# 0.168143f
C4007 a_11599_46634# a_13259_45724# 0.249721f
C4008 a_18451_43940# VDD 0.172318f
C4009 a_11453_44696# VDD 3.75355f
C4010 SMPL_ON_N RST_Z 2.43362f
C4011 a_20193_45348# a_14401_32519# 0.175398f
C4012 a_4190_30871# VREF_GND 0.105109f
C4013 a_17364_32525# VDD 0.511443f
C4014 a_n2497_47436# SMPL_ON_P 0.131317f
C4015 a_n4315_30879# a_n4064_40160# 0.363059f
C4016 a_8325_42308# VDD 0.313956f
C4017 a_5907_45546# VDD 0.390381f
C4018 a_2063_45854# a_7715_46873# 0.178294f
C4019 a_6886_37412# a_8912_37509# 0.339465f
C4020 a_20974_43370# a_4190_30871# 0.214288f
C4021 a_9290_44172# a_10807_43548# 0.364112f
C4022 a_13661_43548# a_11415_45002# 0.107787f
C4023 a_13747_46662# a_20202_43084# 0.308003f
C4024 a_4883_46098# a_9625_46129# 0.164961f
C4025 a_11599_46634# a_18189_46348# 0.101491f
C4026 a_10227_46804# a_13759_46122# 0.920747f
C4027 a_3080_42308# a_n784_42308# 0.170007f
C4028 a_19237_31679# VDD 0.746512f
C4029 a_n971_45724# a_2437_43646# 0.204278f
C4030 a_n901_46420# a_n1076_46494# 0.234322f
C4031 a_16327_47482# a_16115_45572# 0.163022f
C4032 a_n23_47502# VDD 0.152616f
C4033 a_n1059_45260# a_8791_43396# 0.196029f
C4034 a_8953_45546# a_5934_30871# 0.113715f
C4035 a_9145_43396# VDD 2.43736f
C4036 a_12465_44636# a_11691_44458# 0.15589f
C4037 a_n2438_43548# a_1423_45028# 0.242599f
C4038 a_11453_44696# a_11827_44484# 0.170003f
C4039 a_15764_42576# a_15803_42450# 0.901878f
C4040 a_11967_42832# a_n97_42460# 0.489711f
C4041 a_12861_44030# a_15493_43940# 0.370814f
C4042 a_10180_45724# a_10193_42453# 0.145672f
C4043 a_n443_46116# a_768_44030# 0.177051f
C4044 a_4915_47217# a_12549_44172# 0.316329f
C4045 a_n971_45724# a_n2661_46634# 0.190714f
C4046 a_n2497_47436# a_n2438_43548# 0.206216f
C4047 a_n3565_38216# a_n4209_37414# 5.88577f
C4048 a_n4315_30879# C10_P_btm 1.5848f
C4049 a_3905_42865# a_3935_42891# 0.240349f
C4050 a_n2293_46634# a_8685_43396# 0.335608f
C4051 a_5257_43370# a_n97_42460# 0.167676f
C4052 a_22959_45572# a_20447_31679# 0.154273f
C4053 a_n1059_45260# VDD 4.75361f
C4054 a_3160_47472# a_3147_46376# 0.208295f
C4055 a_n971_45724# a_8199_44636# 0.247183f
C4056 a_12861_44030# a_12741_44636# 0.366155f
C4057 a_20107_46660# a_20623_46660# 0.105914f
C4058 a_13661_43548# a_13259_45724# 0.250875f
C4059 a_n2312_39304# a_n3565_39304# 0.104981f
C4060 a_n357_42282# a_n13_43084# 0.194173f
C4061 a_20193_45348# a_20512_43084# 0.160912f
C4062 a_n2840_43370# VDD 0.246858f
C4063 a_768_44030# a_3537_45260# 0.341201f
C4064 a_10903_43370# a_8049_45260# 0.114138f
C4065 a_4185_45028# a_13259_45724# 0.194989f
C4066 a_948_46660# VDD 0.278482f
C4067 a_19279_43940# a_19328_44172# 0.120319f
C4068 a_5013_44260# a_5495_43940# 0.251039f
C4069 a_19987_42826# VDD 0.588466f
C4070 a_11415_45002# a_13159_45002# 0.141106f
C4071 a_1823_45246# a_3065_45002# 0.607468f
C4072 a_13925_46122# VDD 0.251868f
C4073 a_2063_45854# a_11599_46634# 0.19861f
C4074 a_4915_47217# a_6575_47204# 0.849579f
C4075 a_6545_47178# a_6491_46660# 0.181574f
C4076 a_18184_42460# a_22400_42852# 0.16156f
C4077 a_13258_32519# VIN_N 0.143165f
C4078 a_n2661_45546# a_n2661_43370# 0.145941f
C4079 a_18175_45572# a_18341_45572# 0.577068f
C4080 a_15599_45572# VDD 0.390565f
C4081 a_n971_45724# a_765_45546# 0.140618f
C4082 a_n1613_43370# a_5907_46634# 0.338694f
C4083 a_22459_39145# VDD 0.682253f
C4084 EN_VIN_BSTR_P C4_P_btm 0.116925f
C4085 a_14401_32519# a_5534_30871# 0.339008f
C4086 a_n4318_40392# VDD 0.573389f
C4087 a_4883_46098# a_8049_45260# 0.469963f
C4088 a_n743_46660# a_9823_46155# 0.196587f
C4089 a_12549_44172# a_10809_44734# 2.27272f
C4090 a_18326_43940# VDD 0.129408f
C4091 a_12465_44636# a_2437_43646# 0.18195f
C4092 SMPL_ON_N VDD 0.503419f
C4093 a_n473_42460# a_n327_42558# 0.171361f
C4094 COMP_P a_n1630_35242# 2.45645f
C4095 a_22959_43396# VDD 0.303237f
C4096 a_n4315_30879# a_n4334_40480# 0.253307f
C4097 a_14955_43940# a_15037_43940# 0.171361f
C4098 a_15227_44166# a_16241_44734# 0.105126f
C4099 a_n863_45724# a_2382_45260# 0.119625f
C4100 a_5263_45724# VDD 0.202719f
C4101 a_n881_46662# a_12549_44172# 0.225257f
C4102 SMPL_ON_N a_22612_30879# 5.16049f
C4103 a_5088_37509# VDAC_P 1.15441f
C4104 a_5700_37509# a_8912_37509# 15.051701f
C4105 a_14401_32519# a_4190_30871# 0.10855f
C4106 a_5111_44636# a_3232_43370# 0.134191f
C4107 a_9290_44172# a_10949_43914# 0.113864f
C4108 a_13259_45724# a_11967_42832# 0.141918f
C4109 a_n755_45592# a_n97_42460# 1.02989f
C4110 a_22959_45036# a_19721_31679# 0.156264f
C4111 a_22959_44484# VDD 0.303517f
C4112 a_16327_47482# a_16333_45814# 0.168559f
C4113 a_n237_47217# VDD 4.05131f
C4114 a_10341_42308# a_9803_42558# 0.108853f
C4115 a_5111_44636# a_4905_42826# 0.128918f
C4116 a_5883_43914# a_7542_44172# 0.187537f
C4117 a_8270_45546# VDD 1.26092f
C4118 a_15486_42560# a_15803_42450# 0.102355f
C4119 a_10729_43914# a_11750_44172# 0.144893f
C4120 a_2711_45572# a_19511_42282# 0.234026f
C4121 a_4915_47217# a_12891_46348# 0.156543f
C4122 a_6575_47204# a_n881_46662# 0.708623f
C4123 a_20894_47436# a_20990_47178# 0.313533f
C4124 a_3905_42865# a_3681_42891# 0.101054f
C4125 a_4699_43561# a_3080_42308# 0.223965f
C4126 a_19692_46634# a_14021_43940# 0.775991f
C4127 a_n2017_45002# VDD 3.8321f
C4128 a_3357_43084# CLK 2.63944f
C4129 a_12549_44172# a_17609_46634# 0.487224f
C4130 a_3422_30871# VDAC_N 0.480069f
C4131 a_20411_46873# a_20273_46660# 0.219954f
C4132 a_1123_46634# VDD 0.469393f
C4133 a_3537_45260# a_5111_42852# 0.123919f
C4134 a_n913_45002# a_12545_42858# 0.548984f
C4135 a_5244_44056# a_5495_43940# 0.107037f
C4136 a_19164_43230# VDD 0.278643f
C4137 a_11415_45002# a_13017_45260# 0.100288f
C4138 a_13759_46122# VDD 0.399995f
C4139 a_6151_47436# a_6491_46660# 0.31912f
C4140 a_3422_30871# a_13467_32519# 0.421402f
C4141 a_18175_45572# a_18479_45785# 0.280208f
C4142 a_526_44458# a_n699_43396# 0.285f
C4143 a_13259_45724# a_18315_45260# 0.144632f
C4144 a_9049_44484# a_3232_43370# 0.17048f
C4145 a_n2956_37592# a_n3565_37414# 0.304738f
C4146 a_n2293_46634# a_n2438_43548# 0.807205f
C4147 a_n1613_43370# a_5167_46660# 0.177362f
C4148 a_n1151_42308# a_13885_46660# 0.333314f
C4149 a_19864_35138# a_21589_35634# 0.150796f
C4150 a_22521_40055# VDD 1.04757f
C4151 EN_VIN_BSTR_P C5_P_btm 0.115337f
C4152 a_n2840_44458# VDD 0.247948f
C4153 a_14084_46812# a_13885_46660# 0.237373f
C4154 a_n443_46116# a_n2661_45546# 0.136593f
C4155 a_n743_46660# a_9569_46155# 0.104962f
C4156 a_12891_46348# a_10809_44734# 0.102888f
C4157 a_10903_43370# a_5534_30871# 0.134296f
C4158 a_18079_43940# VDD 0.162408f
C4159 a_13717_47436# a_413_45260# 4.36729f
C4160 a_22731_47423# VDD 0.196667f
C4161 a_21811_47423# SINGLE_ENDED 0.215228f
C4162 a_n4318_37592# a_n1630_35242# 0.847279f
C4163 a_n1059_45260# a_16823_43084# 0.318918f
C4164 a_3422_30871# a_22315_44484# 0.19914f
C4165 a_14209_32519# VDD 0.284433f
C4166 a_10809_44734# a_11322_45546# 0.22629f
C4167 a_10227_46804# a_9313_44734# 0.875947f
C4168 a_n2288_47178# a_n2109_47186# 0.177673f
C4169 a_n913_45002# a_5379_42460# 0.179494f
C4170 a_3905_42865# a_4905_42826# 0.404829f
C4171 a_310_45028# a_n37_45144# 0.112458f
C4172 a_10193_42453# a_16147_45260# 0.193225f
C4173 a_18189_46348# a_18315_45260# 0.101775f
C4174 a_15227_44166# a_14673_44172# 0.357896f
C4175 a_n755_45592# a_n467_45028# 0.26002f
C4176 a_n863_45724# a_2274_45254# 0.17549f
C4177 a_n2661_45546# a_3537_45260# 0.780422f
C4178 a_n2956_37592# a_n4209_39304# 0.102982f
C4179 a_4099_45572# VDD 0.296272f
C4180 a_2063_45854# a_5257_43370# 0.426517f
C4181 SMPL_ON_N a_21588_30879# 0.119129f
C4182 a_6151_47436# a_4646_46812# 0.153739f
C4183 a_5700_37509# VDAC_N 1.09421f
C4184 a_5088_37509# a_8912_37509# 16.1906f
C4185 a_3726_37500# a_11206_38545# 0.11542f
C4186 a_n2302_38778# VDD 0.35162f
C4187 a_5111_44636# a_5691_45260# 0.130044f
C4188 a_5147_45002# a_3232_43370# 0.253159f
C4189 a_5649_42852# a_5534_30871# 0.234793f
C4190 a_1847_42826# a_2075_43172# 0.103349f
C4191 a_n1557_42282# COMP_P 0.123881f
C4192 a_n357_42282# a_n97_42460# 0.900712f
C4193 a_1423_45028# a_5891_43370# 0.301629f
C4194 a_17730_32519# VDD 0.289738f
C4195 a_n746_45260# VDD 1.41433f
C4196 a_2382_45260# a_2982_43646# 0.468592f
C4197 a_8199_44636# a_5934_30871# 0.159294f
C4198 a_10903_43370# a_n443_42852# 0.176275f
C4199 a_15486_42560# a_15764_42576# 0.118759f
C4200 a_10729_43914# a_10807_43548# 0.238591f
C4201 a_2127_44172# a_2253_43940# 0.143754f
C4202 a_10053_45546# a_10180_45724# 0.144403f
C4203 a_12741_44636# a_16922_45042# 0.139755f
C4204 a_7499_43078# a_8746_45002# 0.153858f
C4205 a_7903_47542# a_n881_46662# 0.178742f
C4206 VDAC_Pi a_3754_39466# 0.308867f
C4207 a_15493_43940# a_15743_43084# 0.206331f
C4208 a_2437_43646# a_n2661_45010# 0.15182f
C4209 a_n2109_45247# VDD 0.266396f
C4210 VDD VCM 1.51164f
C4211 a_21487_43396# a_13467_32519# 0.152042f
C4212 a_4190_30871# a_5649_42852# 0.434284f
C4213 a_20107_46660# a_20273_46660# 0.608339f
C4214 a_10227_46804# a_2711_45572# 0.130695f
C4215 a_n2312_39304# a_n4209_39304# 0.19527f
C4216 a_17538_32519# VDD 0.352239f
C4217 a_n881_46662# a_6431_45366# 0.177591f
C4218 a_n2293_46098# a_n2661_45546# 3.03243f
C4219 a_768_44030# a_3065_45002# 0.288972f
C4220 a_n1613_43370# a_5205_44484# 0.551795f
C4221 a_3483_46348# a_13259_45724# 0.230226f
C4222 a_383_46660# VDD 0.198466f
C4223 a_22612_30879# VCM 0.473529f
C4224 a_1606_42308# a_5742_30871# 3.46204f
C4225 a_19339_43156# VDD 0.338297f
C4226 a_1823_45246# a_2382_45260# 0.801932f
C4227 a_13351_46090# VDD 0.238036f
C4228 a_6151_47436# a_6545_47178# 0.39775f
C4229 a_2711_45572# a_1307_43914# 0.187968f
C4230 a_16375_45002# a_16922_45042# 0.170835f
C4231 a_7499_43078# a_3232_43370# 0.318423f
C4232 a_n2810_45028# a_n3565_37414# 0.135518f
C4233 a_n1613_43370# a_5385_46902# 0.182522f
C4234 a_11599_46634# a_11813_46116# 0.106062f
C4235 EN_VIN_BSTR_P C6_P_btm 0.118916f
C4236 a_n863_45724# a_1414_42308# 0.711805f
C4237 a_6171_45002# a_n2661_43370# 2.37006f
C4238 a_n755_45592# a_n809_44244# 0.404418f
C4239 a_2711_45572# a_18579_44172# 0.170319f
C4240 a_13059_46348# a_14579_43548# 0.171744f
C4241 a_19721_31679# VDD 0.521328f
C4242 a_13607_46688# a_13885_46660# 0.11044f
C4243 a_n2661_46634# a_10903_43370# 0.663878f
C4244 a_n743_46660# a_9625_46129# 0.206271f
C4245 a_n443_42852# a_8685_43396# 0.281116f
C4246 a_17973_43940# VDD 0.265874f
C4247 a_4883_46098# a_2437_43646# 0.458866f
C4248 a_16327_47482# a_n913_45002# 0.137194f
C4249 a_4883_46098# SINGLE_ENDED 0.1664f
C4250 a_22223_47212# VDD 0.236555f
C4251 a_n961_42308# a_n784_42308# 0.154417f
C4252 a_5891_43370# a_10405_44172# 0.15894f
C4253 a_22591_43396# VDD 0.280354f
C4254 a_20731_47026# VDD 0.132317f
C4255 a_n2497_47436# a_n2109_47186# 0.197671f
C4256 a_13483_43940# a_13565_43940# 0.171361f
C4257 a_526_44458# a_n2293_42834# 1.7774f
C4258 a_n863_45724# a_1667_45002# 0.20954f
C4259 a_3175_45822# VDD 0.193907f
C4260 a_5700_37509# a_6886_37412# 0.13762f
C4261 a_5088_37509# VDAC_N 0.420254f
C4262 a_4338_37500# a_8912_37509# 0.331796f
C4263 a_n4064_38528# VDD 1.69517f
C4264 a_n97_42460# a_19700_43370# 0.154491f
C4265 a_7499_43078# a_8975_43940# 0.519621f
C4266 a_5111_44636# a_4927_45028# 0.134309f
C4267 a_4883_46098# a_8199_44636# 0.242f
C4268 a_11599_46634# a_15682_46116# 1.8289f
C4269 a_22223_45036# a_18114_32519# 0.15655f
C4270 a_22591_44484# VDD 0.223346f
C4271 a_n1991_46122# a_n1076_46494# 0.124988f
C4272 a_n971_45724# VDD 4.911799f
C4273 SMPL_ON_P CLK_DATA 0.200962f
C4274 a_19778_44110# a_19862_44208# 0.213467f
C4275 a_n755_45592# a_n2293_42282# 0.208531f
C4276 a_13507_46334# a_20193_45348# 0.253904f
C4277 a_14113_42308# a_15803_42450# 0.289859f
C4278 a_10729_43914# a_10949_43914# 0.418928f
C4279 a_10809_44734# a_6171_45002# 0.244599f
C4280 a_526_44458# a_413_45260# 0.103799f
C4281 a_7499_43078# a_10193_42453# 0.298293f
C4282 a_1049_43396# a_n1557_42282# 0.211757f
C4283 a_n863_45724# a_n699_43396# 0.23135f
C4284 a_n2293_45010# VDD 1.885f
C4285 a_2063_45854# a_3483_46348# 0.164542f
C4286 VDD VREF_GND 0.482759f
C4287 a_3422_30871# a_7174_31319# 2.22059f
C4288 a_743_42282# a_4361_42308# 7.66647f
C4289 a_n913_45002# a_n356_44636# 0.640597f
C4290 a_9313_44734# VDD 0.389068f
C4291 a_20107_46660# a_20411_46873# 0.316529f
C4292 a_n743_46660# a_8049_45260# 2.07544f
C4293 a_5649_42852# a_4921_42308# 0.133152f
C4294 a_10903_43370# a_13291_42460# 0.135558f
C4295 a_4185_45028# a_22400_42852# 0.105692f
C4296 a_20974_43370# VDD 0.550101f
C4297 a_15227_44166# a_10193_42453# 0.205591f
C4298 a_601_46902# VDD 0.204253f
C4299 a_22612_30879# VREF_GND 0.168163f
C4300 a_21588_30879# VCM 0.179761f
C4301 a_3905_42865# a_5013_44260# 0.182997f
C4302 a_18599_43230# VDD 0.197104f
C4303 a_13259_45724# a_13249_42308# 0.358931f
C4304 a_167_45260# a_327_44734# 0.199136f
C4305 a_n755_45592# a_3775_45552# 0.100709f
C4306 a_n2293_46634# a_5891_43370# 0.105307f
C4307 a_1823_45246# a_2274_45254# 0.255985f
C4308 a_12594_46348# VDD 1.03351f
C4309 a_4915_47217# a_6851_47204# 0.172567f
C4310 a_16147_45260# a_18175_45572# 0.108647f
C4311 a_n2956_37592# a_n4209_37414# 0.145558f
C4312 a_n1613_43370# a_4817_46660# 0.330391f
C4313 a_n2104_46634# a_n1925_46634# 0.167849f
C4314 a_11599_46634# a_11735_46660# 0.268769f
C4315 EN_VIN_BSTR_P C7_P_btm 0.115875f
C4316 a_22469_40625# VDD 0.564837f
C4317 a_18114_32519# VDD 0.550312f
C4318 a_n2293_46634# a_9290_44172# 0.102393f
C4319 a_12861_44030# a_13259_45724# 0.435853f
C4320 a_3626_43646# a_5742_30871# 0.168508f
C4321 a_10334_44484# a_10440_44484# 0.313533f
C4322 a_5147_45002# a_5013_44260# 0.189328f
C4323 a_17737_43940# VDD 0.285511f
C4324 a_4646_46812# a_7499_43078# 0.158236f
C4325 a_16327_47482# a_n1059_45260# 0.235708f
C4326 a_12465_44636# VDD 0.773277f
C4327 a_n4318_37592# a_n3674_37592# 3.06402f
C4328 a_n3674_38216# a_n1630_35242# 0.333493f
C4329 a_14537_43396# a_9145_43396# 0.129182f
C4330 a_13887_32519# VDD 0.424101f
C4331 a_8515_42308# VDD 0.194691f
C4332 a_n863_45724# a_327_44734# 0.353745f
C4333 a_n971_45724# a_8147_43396# 0.116186f
C4334 a_13747_46662# a_19862_44208# 0.15289f
C4335 a_2711_45572# VDD 1.22011f
C4336 a_22223_47212# a_21588_30879# 0.164932f
C4337 a_n443_46116# a_4955_46873# 0.126551f
C4338 a_5088_37509# a_6886_37412# 0.136505f
C4339 a_3726_37500# a_8912_37509# 0.267651f
C4340 a_n2946_38778# VDD 0.383009f
C4341 a_7499_43078# a_10057_43914# 0.262644f
C4342 a_5147_45002# a_4927_45028# 0.168157f
C4343 a_n357_42282# a_n2661_42834# 0.239713f
C4344 a_2905_45572# a_526_44458# 0.142766f
C4345 a_11599_46634# a_2324_44458# 0.428445f
C4346 a_n1557_42282# a_n1736_42282# 0.170341f
C4347 a_1423_45028# a_7640_43914# 0.105665f
C4348 a_9290_44172# a_743_42282# 0.117511f
C4349 a_22485_44484# VDD 0.258874f
C4350 a_n2109_47186# a_3357_43084# 0.170493f
C4351 a_16327_47482# a_15599_45572# 0.331892f
C4352 a_n1423_46090# a_n1641_46494# 0.209641f
C4353 a_5883_43914# a_5663_43940# 0.153361f
C4354 a_12465_44636# a_11827_44484# 0.785011f
C4355 a_15051_42282# a_15486_42560# 0.234322f
C4356 a_14113_42308# a_15764_42576# 0.229529f
C4357 a_5932_42308# a_7174_31319# 13.0265f
C4358 a_11823_42460# a_11551_42558# 0.138126f
C4359 a_16877_42852# VDD 0.192454f
C4360 a_10809_44734# a_3232_43370# 0.158726f
C4361 a_10227_46804# a_4883_46098# 0.200137f
C4362 a_7754_39964# a_7754_39632# 0.296522f
C4363 a_1209_43370# a_n1557_42282# 0.113851f
C4364 a_22591_45572# a_19963_31679# 0.161955f
C4365 a_13507_46334# a_4190_30871# 0.186424f
C4366 a_n1925_42282# a_n2293_43922# 2.06056f
C4367 a_n2472_45002# VDD 0.217954f
C4368 a_2437_43646# CLK 0.101524f
C4369 a_10227_46804# a_21188_46660# 0.22222f
C4370 C10_N_btm VCM 10.3108f
C4371 VDD VREF 4.8299f
C4372 a_7229_43940# a_5343_44458# 0.196399f
C4373 a_3232_43370# a_5883_43914# 0.337937f
C4374 a_n3674_39304# a_n3420_39616# 0.152699f
C4375 a_14401_32519# VDD 0.562673f
C4376 a_33_46660# VDD 0.272723f
C4377 a_22612_30879# VREF 1.73216f
C4378 a_18817_42826# VDD 0.204624f
C4379 a_167_45260# a_413_45260# 0.120357f
C4380 a_1823_45246# a_1667_45002# 0.24808f
C4381 a_8199_44636# CLK 0.231904f
C4382 a_12005_46116# VDD 0.518463f
C4383 a_4915_47217# a_6491_46660# 0.19739f
C4384 a_5815_47464# a_6151_47436# 0.235454f
C4385 a_1343_38525# a_2684_37794# 0.224374f
C4386 a_n3420_39072# a_n4064_38528# 7.47287f
C4387 a_1736_39043# a_2112_39137# 0.554188f
C4388 a_n1059_45260# a_18727_42674# 0.20226f
C4389 a_n863_45724# a_n2293_42834# 0.107229f
C4390 a_10809_44734# a_8975_43940# 0.169586f
C4391 a_8953_45546# a_5891_43370# 0.321625f
C4392 a_10227_46804# a_8685_43396# 0.227547f
C4393 a_4883_46098# a_9396_43370# 0.172323f
C4394 a_14033_45822# VDD 0.195067f
C4395 a_n2661_46634# a_n2438_43548# 0.493975f
C4396 a_n2104_46634# a_n2312_38680# 0.154937f
C4397 a_22521_40599# VDD 0.804442f
C4398 a_10341_43396# a_15743_43084# 0.464206f
C4399 a_1414_42308# a_1184_42692# 0.115223f
C4400 a_584_46384# a_n357_42282# 0.107436f
C4401 a_15227_44166# a_19692_46634# 0.116169f
C4402 a_19333_46634# a_19466_46812# 0.167526f
C4403 a_13661_43548# a_2324_44458# 0.307974f
C4404 a_5883_43914# a_8975_43940# 0.50976f
C4405 a_5147_45002# a_5244_44056# 0.122327f
C4406 a_15682_43940# VDD 1.22657f
C4407 a_13507_46334# a_2437_43646# 0.117533f
C4408 a_n2497_47436# a_1423_45028# 1.36987f
C4409 a_16327_47482# a_n2017_45002# 0.209709f
C4410 a_8953_45546# a_9290_44172# 0.373944f
C4411 a_13507_46334# SINGLE_ENDED 0.111959f
C4412 a_21811_47423# VDD 0.201359f
C4413 COMP_P a_n784_42308# 0.10915f
C4414 a_22223_43396# VDD 0.279195f
C4415 a_20411_46873# a_3357_43084# 0.157199f
C4416 a_22000_46634# VDD 0.257047f
C4417 a_5934_30871# VDD 0.431204f
C4418 a_n863_45724# a_413_45260# 0.140312f
C4419 a_n237_47217# a_8667_46634# 0.171086f
C4420 a_4338_37500# a_6886_37412# 1.95816f
C4421 a_5088_37509# a_5700_37509# 1.48771f
C4422 a_n3420_38528# VDD 0.522772f
C4423 a_n97_42460# a_15743_43084# 0.205305f
C4424 a_3537_45260# a_3232_43370# 0.530258f
C4425 a_16327_47482# a_19164_43230# 0.292734f
C4426 a_5147_45002# a_5111_44636# 0.562127f
C4427 a_4558_45348# a_4927_45028# 0.123258f
C4428 a_9290_44172# a_9028_43914# 0.169653f
C4429 a_4883_46098# a_8016_46348# 0.289691f
C4430 a_3080_42308# COMP_P 4.43551f
C4431 a_n4318_39304# a_n4209_39304# 0.135369f
C4432 a_20512_43084# VDD 0.317257f
C4433 a_17730_32519# C9_N_btm 0.215899f
C4434 a_n743_46660# a_n443_42852# 0.378464f
C4435 a_n1991_46122# a_n1641_46494# 0.219633f
C4436 a_n2157_46122# a_n1076_46494# 0.102355f
C4437 a_n1741_47186# a_2437_43646# 4.86702f
C4438 a_n815_47178# VDD 0.380339f
C4439 a_13467_32519# a_13258_32519# 11.0084f
C4440 a_5343_44458# a_7845_44172# 0.103601f
C4441 a_3537_45260# a_4905_42826# 0.339989f
C4442 a_22959_46124# a_20692_30879# 0.155635f
C4443 a_5204_45822# a_5263_45724# 0.109078f
C4444 a_n1630_35242# a_n1532_35090# 0.462421f
C4445 a_16245_42852# VDD 0.205729f
C4446 a_8049_45260# a_22959_45572# 0.176374f
C4447 a_768_44030# a_453_43940# 0.110708f
C4448 a_n1741_47186# a_n2661_46634# 0.22396f
C4449 a_4093_43548# a_4235_43370# 0.515101f
C4450 a_n2293_46098# a_5663_43940# 0.142661f
C4451 a_n2661_45010# VDD 0.842431f
C4452 a_n1925_46634# a_6755_46942# 0.12389f
C4453 a_768_44030# a_3090_45724# 0.115303f
C4454 a_10227_46804# a_21363_46634# 0.273017f
C4455 VDD VIN_N 1.46155f
C4456 C9_N_btm VCM 6.06251f
C4457 C10_N_btm VREF_GND 10.3207f
C4458 a_526_44458# a_n97_42460# 0.277959f
C4459 a_5205_44484# a_5518_44484# 0.135771f
C4460 a_21381_43940# VDD 0.344882f
C4461 a_n2956_39304# a_n2956_38680# 0.163045f
C4462 a_22612_30879# VIN_N 0.19035f
C4463 a_171_46873# VDD 0.539781f
C4464 a_21588_30879# VREF 0.860047f
C4465 a_6171_42473# a_5932_42308# 0.224949f
C4466 a_18249_42858# VDD 0.250132f
C4467 a_167_45260# a_n37_45144# 0.277898f
C4468 a_10903_43370# VDD 2.60588f
C4469 a_1343_38525# a_1177_38525# 0.238422f
C4470 a_n1059_45260# a_18057_42282# 0.141112f
C4471 a_526_44458# a_742_44458# 0.54618f
C4472 a_7499_43078# a_5111_44636# 0.753731f
C4473 a_13259_45724# a_16922_45042# 0.401687f
C4474 a_n1741_47186# a_765_45546# 0.536367f
C4475 a_n2293_46634# a_n2312_38680# 0.131017f
C4476 a_n1613_43370# a_4651_46660# 0.686447f
C4477 EN_VIN_BSTR_P C9_P_btm 0.226529f
C4478 a_18194_35068# a_19120_35138# 0.558402f
C4479 EN_VIN_BSTR_N a_19864_35138# 0.573134f
C4480 a_11206_38545# RST_Z 0.382319f
C4481 CAL_N VDD 26.069302f
C4482 a_n1059_45260# a_18494_42460# 0.187733f
C4483 a_18114_32519# C10_N_btm 0.460005f
C4484 a_15227_44166# a_19466_46812# 0.310201f
C4485 a_5807_45002# a_2324_44458# 0.232399f
C4486 a_2982_43646# a_5742_30871# 0.196805f
C4487 a_10157_44484# a_10334_44484# 0.159555f
C4488 a_9290_44172# a_5534_30871# 0.472376f
C4489 a_14955_43940# VDD 0.253201f
C4490 a_n1151_42308# a_6709_45028# 0.286957f
C4491 a_n1853_46287# a_n1736_46482# 0.170096f
C4492 a_4791_45118# a_3232_43370# 0.268929f
C4493 a_9625_46129# a_9823_46155# 0.321686f
C4494 a_10227_46804# CLK 0.207445f
C4495 a_4883_46098# VDD 1.12729f
C4496 a_14539_43914# a_15493_43940# 0.625897f
C4497 a_5649_42852# VDD 0.438443f
C4498 w_11334_34010# a_3422_30871# 1.91172f
C4499 a_21188_46660# VDD 0.284105f
C4500 a_20107_42308# a_7174_31319# 0.175129f
C4501 a_n2833_47464# a_n2497_47436# 0.217831f
C4502 a_7963_42308# VDD 0.266057f
C4503 a_4791_45118# a_4905_42826# 0.516502f
C4504 a_3726_37500# a_6886_37412# 0.702909f
C4505 a_4338_37500# a_5700_37509# 2.69237f
C4506 a_n3690_38528# VDD 0.363159f
C4507 a_16327_47482# a_19339_43156# 0.346029f
C4508 a_n443_42852# a_5891_43370# 0.175668f
C4509 a_n1613_43370# a_n1076_46494# 0.232314f
C4510 a_n743_46660# a_765_45546# 0.148721f
C4511 a_685_42968# a_791_42968# 0.13675f
C4512 a_n1991_46122# a_n1423_46090# 0.175891f
C4513 a_n1605_47204# VDD 0.20224f
C4514 a_n2293_42282# a_1755_42282# 0.875855f
C4515 a_8685_43396# VDD 0.261626f
C4516 a_9290_44172# a_n443_42852# 0.483812f
C4517 a_n746_45260# a_n356_44636# 0.418585f
C4518 a_15227_44166# a_16147_45260# 0.282941f
C4519 a_4646_46812# a_3537_45260# 0.361823f
C4520 a_8049_45260# a_19963_31679# 0.2062f
C4521 a_10227_46804# a_13507_46334# 0.120657f
C4522 a_n2497_47436# a_n2293_46634# 0.174929f
C4523 a_n4064_40160# EN_VIN_BSTR_P 0.187697f
C4524 a_n97_42460# a_3626_43646# 0.394673f
C4525 a_3357_43084# a_22591_45572# 0.181818f
C4526 a_13661_43548# a_13667_43396# 0.168674f
C4527 a_19479_31679# a_19963_31679# 0.104687f
C4528 a_526_44458# a_n2661_43922# 0.154533f
C4529 a_n2840_45002# VDD 0.289706f
C4530 a_10227_46804# a_20623_46660# 0.156341f
C4531 a_n443_46116# a_n901_46420# 0.367344f
C4532 VDD VIN_P 1.47957f
C4533 C8_N_btm VCM 2.61094f
C4534 C9_N_btm VREF_GND 5.18245f
C4535 C10_N_btm VREF 14.773f
C4536 a_3422_30871# a_13258_32519# 0.410904f
C4537 a_n443_42852# a_10807_43548# 0.173997f
C4538 a_5205_44484# a_5343_44458# 0.129692f
C4539 a_10249_46116# a_10355_46116# 0.182836f
C4540 a_4361_42308# a_4921_42308# 0.472085f
C4541 a_n1925_42282# a_n2293_42282# 0.234055f
C4542 a_19741_43940# VDD 0.153579f
C4543 a_n133_46660# VDD 0.483405f
C4544 a_21588_30879# VIN_N 0.106594f
C4545 a_5755_42308# a_5932_42308# 0.196877f
C4546 a_17333_42852# VDD 0.525529f
C4547 a_13259_45724# a_13163_45724# 0.166368f
C4548 a_4915_47217# a_6151_47436# 0.783303f
C4549 a_n3420_39072# a_n3420_38528# 0.127439f
C4550 a_n913_45002# a_17303_42282# 1.81467f
C4551 a_8199_44636# a_5891_43370# 0.399007f
C4552 a_3090_45724# a_7542_44172# 0.137368f
C4553 a_n1613_43370# a_4646_46812# 1.38979f
C4554 a_n881_46662# a_3877_44458# 0.142507f
C4555 EN_VIN_BSTR_P C10_P_btm 0.320569f
C4556 EN_VIN_BSTR_N a_19120_35138# 0.652984f
C4557 a_11530_34132# a_19864_35138# 0.201937f
C4558 VDAC_P RST_Z 0.158793f
C4559 a_11206_38545# VDD 8.87267f
C4560 a_1414_42308# a_1067_42314# 0.100434f
C4561 a_1568_43370# a_1847_42826# 0.153113f
C4562 a_n863_45724# a_175_44278# 0.113317f
C4563 a_n1059_45260# a_18184_42460# 0.52106f
C4564 a_10227_46804# a_10586_45546# 0.306536f
C4565 a_n2129_44697# a_n2012_44484# 0.172424f
C4566 a_13483_43940# VDD 0.219591f
C4567 a_9625_46129# a_9569_46155# 0.204034f
C4568 a_n2497_47436# a_626_44172# 0.249352f
C4569 a_3090_45724# a_n2661_45546# 0.561435f
C4570 a_8199_44636# a_9290_44172# 0.516297f
C4571 a_3483_46348# a_2324_44458# 0.668551f
C4572 a_13747_46662# a_15765_45572# 0.5661f
C4573 a_21496_47436# VDD 0.198362f
C4574 a_13678_32519# VDD 0.454512f
C4575 w_1575_34946# a_3422_30871# 1.88476f
C4576 a_768_44030# a_n699_43396# 1.37533f
C4577 a_16327_47482# a_9313_44734# 0.169217f
C4578 a_10903_43370# a_10907_45822# 0.199567f
C4579 a_21363_46634# VDD 0.357368f
C4580 a_n913_45002# a_2713_42308# 0.291963f
C4581 a_18184_42460# a_19987_42826# 0.208392f
C4582 a_6123_31319# VDD 0.532709f
C4583 a_13661_43548# a_15493_43396# 0.491785f
C4584 a_n881_46662# a_8128_46384# 0.206292f
C4585 a_21811_47423# a_20916_46384# 0.109084f
C4586 a_4791_45118# a_4646_46812# 0.485113f
C4587 a_10227_46804# a_n743_46660# 0.134234f
C4588 a_4338_37500# a_5088_37509# 0.896828f
C4589 a_3726_37500# a_5700_37509# 0.574743f
C4590 a_n3565_38502# VDD 0.762011f
C4591 a_19319_43548# a_4190_30871# 0.188868f
C4592 a_16327_47482# a_18599_43230# 0.182696f
C4593 a_15861_45028# a_16922_45042# 0.259169f
C4594 a_3537_45260# a_4927_45028# 0.216859f
C4595 a_584_46384# a_n1925_42282# 0.194054f
C4596 a_n1613_43370# a_n901_46420# 0.406381f
C4597 a_n237_47217# a_5066_45546# 1.48406f
C4598 a_n863_45724# a_n97_42460# 0.581863f
C4599 a_8270_45546# a_5066_45546# 0.189476f
C4600 a_n2157_46122# a_n1641_46494# 0.105995f
C4601 SMPL_ON_P VDD 0.614138f
C4602 a_n2293_42282# a_1606_42308# 0.192228f
C4603 a_2107_46812# a_9482_43914# 0.109711f
C4604 a_3877_44458# a_3537_45260# 0.12249f
C4605 a_8035_47026# VDD 0.132317f
C4606 a_15597_42852# VDD 0.239357f
C4607 a_6151_47436# a_n881_46662# 1.58776f
C4608 a_n863_45724# a_742_44458# 0.629795f
C4609 a_10227_46804# a_20841_46902# 0.164019f
C4610 a_18479_47436# a_20411_46873# 0.192791f
C4611 C10_N_btm VIN_N 3.66034f
C4612 VDD CLK 0.49309f
C4613 C9_N_btm VREF 7.369471f
C4614 C8_N_btm VREF_GND 2.58605f
C4615 C7_N_btm VCM 1.58335f
C4616 a_3232_43370# a_6298_44484# 0.256727f
C4617 a_n357_42282# a_19862_44208# 0.138067f
C4618 a_5111_44636# a_5883_43914# 0.281106f
C4619 a_16327_47482# a_2711_45572# 0.101699f
C4620 a_n2293_46634# a_3357_43084# 0.963711f
C4621 a_n2438_43548# VDD 3.40589f
C4622 a_n913_45002# a_10796_42968# 0.545674f
C4623 a_18083_42858# VDD 0.408512f
C4624 a_11133_46155# VDD 0.176249f
C4625 a_4791_45118# a_6545_47178# 0.112353f
C4626 a_1736_39587# a_2684_37794# 0.565517f
C4627 a_3422_30871# a_4190_30871# 12.909901f
C4628 a_2711_45572# a_14537_43396# 0.249285f
C4629 a_3090_45724# a_7281_43914# 0.170855f
C4630 a_n1613_43370# a_3877_44458# 1.43013f
C4631 a_n2109_47186# a_765_45546# 0.126431f
C4632 a_n2661_46634# a_n1925_46634# 4.75867f
C4633 a_11530_34132# a_19120_35138# 0.480251f
C4634 EN_VIN_BSTR_N a_18194_35068# 0.340036f
C4635 VDAC_P VDD 5.19214f
C4636 a_7229_43940# a_n2293_42834# 0.148023f
C4637 a_11823_42460# a_n2293_43922# 0.494696f
C4638 a_n2017_45002# a_18184_42460# 0.205351f
C4639 a_n743_46660# a_8016_46348# 0.155955f
C4640 a_11823_42460# a_n97_42460# 0.324041f
C4641 a_12429_44172# VDD 0.169047f
C4642 a_18597_46090# a_3357_43084# 0.160577f
C4643 a_8199_44636# a_10355_46116# 0.176325f
C4644 a_13507_46334# VDD 1.4135f
C4645 a_21855_43396# VDD 0.289066f
C4646 a_768_44030# a_4223_44672# 0.136643f
C4647 a_10227_46804# a_5891_43370# 0.2393f
C4648 a_20623_46660# VDD 0.194217f
C4649 a_7227_42308# VDD 0.296912f
C4650 a_4883_46098# a_20916_46384# 0.471396f
C4651 a_3726_37500# a_5088_37509# 0.189392f
C4652 a_n4334_38528# VDD 0.385889f
C4653 a_16327_47482# a_18817_42826# 0.215236f
C4654 a_8696_44636# a_16922_45042# 0.10244f
C4655 a_n863_45724# a_n2661_43922# 0.115404f
C4656 a_3537_45260# a_5111_44636# 1.36722f
C4657 a_10227_46804# a_9290_44172# 0.918064f
C4658 a_584_46384# a_526_44458# 0.458472f
C4659 a_n1613_43370# a_n1641_46494# 0.152421f
C4660 a_12861_44030# a_2324_44458# 0.95556f
C4661 a_13059_46348# a_13759_46122# 0.249771f
C4662 a_n1853_46287# a_n1991_46122# 0.737461f
C4663 a_19692_46634# a_6945_45028# 0.669658f
C4664 a_n1741_47186# VDD 0.912651f
C4665 a_4190_30871# a_7174_31319# 0.153555f
C4666 a_3065_45002# a_3080_42308# 0.171466f
C4667 a_22223_46124# a_20205_31679# 0.160234f
C4668 a_11415_45002# a_11823_42460# 0.349238f
C4669 a_13507_46334# a_11827_44484# 0.384415f
C4670 a_10193_42453# a_13575_42558# 0.175489f
C4671 a_1115_44172# a_1241_43940# 0.143754f
C4672 a_9290_44172# a_1307_43914# 0.122831f
C4673 a_12861_44030# a_19862_44208# 0.721035f
C4674 a_10586_45546# VDD 0.582083f
C4675 a_n1151_42308# a_12549_44172# 0.466584f
C4676 a_6151_47436# a_n1613_43370# 0.548675f
C4677 a_n97_42460# a_2982_43646# 0.180648f
C4678 a_2479_44172# a_2905_42968# 0.163227f
C4679 a_2063_45854# a_167_45260# 0.359284f
C4680 a_18597_46090# a_19123_46287# 0.188676f
C4681 C8_N_btm VREF 3.6701f
C4682 C9_N_btm VIN_N 1.82823f
C4683 C6_N_btm VCM 0.877241f
C4684 C7_N_btm VREF_GND 1.61142f
C4685 VDD EN_OFFSET_CAL 0.489629f
C4686 a_20301_43646# a_20556_43646# 0.114664f
C4687 a_5649_42852# a_5379_42460# 0.35554f
C4688 a_13720_44458# a_13857_44734# 0.126609f
C4689 a_n1613_43370# a_5111_44636# 0.601769f
C4690 a_768_44030# a_413_45260# 0.182253f
C4691 a_n743_46660# VDD 1.75634f
C4692 a_22612_30879# EN_OFFSET_CAL 0.118817f
C4693 a_17701_42308# VDD 0.243354f
C4694 a_13259_45724# a_11823_42460# 0.626941f
C4695 a_4185_45028# a_n913_45002# 0.855072f
C4696 a_4646_46812# a_6298_44484# 1.65052f
C4697 a_16327_47482# a_20512_43084# 0.118893f
C4698 a_11189_46129# VDD 0.944289f
C4699 a_1239_39043# comp_n 0.38743f
C4700 a_5937_45572# a_6109_44484# 0.163331f
C4701 a_2711_45572# a_14180_45002# 0.147337f
C4702 a_8016_46348# a_5891_43370# 0.183035f
C4703 a_n2661_46634# a_n2312_38680# 0.106815f
C4704 a_11530_34132# a_18194_35068# 0.4004f
C4705 VDAC_N RST_Z 0.154233f
C4706 a_8912_37509# VDD 18.3523f
C4707 a_15681_43442# a_15781_43660# 0.167615f
C4708 a_18834_46812# a_15227_44166# 0.231715f
C4709 a_15279_43071# a_5342_30871# 0.214197f
C4710 a_3537_45260# a_3905_42865# 0.258917f
C4711 a_9290_44172# a_13635_43156# 0.394766f
C4712 a_11750_44172# VDD 0.131662f
C4713 a_4791_45118# a_5111_44636# 1.11355f
C4714 a_21177_47436# VDD 0.179587f
C4715 COMP_P a_n1329_42308# 0.232443f
C4716 a_4361_42308# VDD 0.42717f
C4717 a_20841_46902# VDD 0.20446f
C4718 a_19511_42282# a_7174_31319# 0.240861f
C4719 a_1467_44172# a_1427_43646# 0.104539f
C4720 a_6761_42308# VDD 0.259312f
C4721 a_5742_30871# C6_P_btm 0.170624f
C4722 a_584_46384# a_3626_43646# 0.195961f
C4723 a_12549_44172# a_15493_43940# 0.932577f
C4724 a_13661_43548# a_18451_43940# 0.129334f
C4725 a_21496_47436# a_20916_46384# 0.113102f
C4726 a_3726_37500# a_4338_37500# 0.212154f
C4727 a_n4209_38502# VDD 0.811731f
C4728 a_16327_47482# a_18249_42858# 0.315855f
C4729 a_2382_45260# a_3232_43370# 0.239776f
C4730 a_9049_44484# a_8701_44490# 0.100038f
C4731 a_7499_43078# a_5883_43914# 0.100372f
C4732 a_4574_45260# a_4558_45348# 0.19344f
C4733 a_n1613_43370# a_n1423_46090# 0.15966f
C4734 a_11599_46634# a_13925_46122# 0.549622f
C4735 a_6151_47436# a_6945_45028# 0.335681f
C4736 a_n913_45002# a_11967_42832# 0.156551f
C4737 a_11599_46634# a_15599_45572# 0.26676f
C4738 a_n2157_46122# a_n1991_46122# 0.614266f
C4739 a_19692_46634# a_21137_46414# 0.242332f
C4740 a_n1920_47178# VDD 0.229556f
C4741 a_n2833_47464# CLK_DATA 0.331592f
C4742 a_14815_43914# a_14673_44172# 0.173231f
C4743 a_3877_44458# a_3065_45002# 0.287919f
C4744 a_5891_43370# a_8791_43396# 0.194389f
C4745 a_768_44030# a_644_44056# 0.177755f
C4746 a_5815_47464# a_n1613_43370# 0.360237f
C4747 a_18780_47178# a_18597_46090# 0.175179f
C4748 a_18479_47436# a_19386_47436# 0.219411f
C4749 a_7754_40130# a_7754_39964# 0.301877f
C4750 a_13661_43548# a_9145_43396# 0.135139f
C4751 a_n2293_46098# a_3905_42865# 0.237656f
C4752 a_2711_45572# a_18494_42460# 0.1183f
C4753 a_20447_31679# VDD 0.665681f
C4754 C7_N_btm VREF 1.818f
C4755 C8_N_btm VIN_N 0.907642f
C4756 VDD DATA[5] 0.504354f
C4757 C5_N_btm VCM 0.719982f
C4758 C6_N_btm VREF_GND 0.836236f
C4759 a_5205_44484# a_4223_44672# 0.235572f
C4760 a_3232_43370# a_5343_44458# 0.654021f
C4761 a_5891_43370# VDD 2.12137f
C4762 a_n1925_46634# a_8034_45724# 0.206805f
C4763 a_14537_43396# a_14955_43940# 0.104291f
C4764 a_18533_43940# VDD 0.182147f
C4765 a_10809_44734# a_22959_46124# 0.172346f
C4766 a_8953_45546# a_8049_45260# 0.156816f
C4767 a_22612_30879# a_20447_31679# 0.107874f
C4768 a_n1021_46688# VDD 0.226043f
C4769 a_n1630_35242# a_5742_30871# 1.85829f
C4770 a_4921_42308# a_5932_42308# 0.194195f
C4771 a_17595_43084# VDD 0.168112f
C4772 a_3218_45724# a_3175_45822# 0.132424f
C4773 a_4791_45118# a_3905_42865# 0.208831f
C4774 a_5937_45572# a_3357_43084# 0.257963f
C4775 a_n2293_46098# a_5147_45002# 0.211057f
C4776 a_9290_44172# VDD 2.74561f
C4777 a_n2956_38216# a_n2946_37984# 0.150404f
C4778 a_n443_46116# a_5129_47502# 0.10632f
C4779 a_7499_43078# a_3537_45260# 0.586701f
C4780 a_1823_45246# a_n2661_43922# 0.441151f
C4781 a_n2472_46634# a_n2293_46634# 0.163804f
C4782 a_5807_45002# a_2107_46812# 1.5594f
C4783 a_11530_34132# EN_VIN_BSTR_N 1.02927f
C4784 VDAC_N VDD 4.62327f
C4785 a_n3420_37440# VIN_P 0.143165f
C4786 a_n97_42460# a_7227_42852# 0.117893f
C4787 a_n237_47217# a_1848_45724# 0.232571f
C4788 a_5534_30871# a_5342_30871# 11.128201f
C4789 a_3537_45260# a_3600_43914# 0.157156f
C4790 a_10807_43548# VDD 0.68049f
C4791 a_n2472_46090# a_n2956_38680# 0.157373f
C4792 a_18479_47436# a_3357_43084# 0.292061f
C4793 a_4791_45118# a_5147_45002# 0.10845f
C4794 a_19787_47423# START 0.220891f
C4795 a_20990_47178# VDD 0.210484f
C4796 a_n2661_43922# a_n3674_39768# 0.152656f
C4797 a_18989_43940# a_18451_43940# 0.114286f
C4798 a_13467_32519# VDD 0.353373f
C4799 a_20273_46660# VDD 0.247553f
C4800 a_n1151_42308# a_n1557_42282# 0.214486f
C4801 a_n755_45592# a_n913_45002# 0.347782f
C4802 a_n971_45724# a_7577_46660# 0.523694f
C4803 a_13507_46334# a_20916_46384# 0.123008f
C4804 a_n4209_39304# VREF 0.195875f
C4805 a_2112_39137# VDD 0.284849f
C4806 a_3537_45260# a_4558_45348# 0.236111f
C4807 a_n881_46662# a_n1853_46287# 0.229188f
C4808 a_11599_46634# a_13759_46122# 0.262969f
C4809 a_n1059_45260# a_11967_42832# 0.627158f
C4810 a_22315_44484# VDD 0.213791f
C4811 a_n1613_43370# a_7499_43078# 0.324998f
C4812 a_n2157_46122# a_n1853_46287# 0.617317f
C4813 a_19692_46634# a_20708_46348# 0.318388f
C4814 a_n2293_46634# a_n443_42852# 2.09483f
C4815 a_n2109_47186# VDD 2.71791f
C4816 a_n357_42282# a_21356_42826# 0.156735f
C4817 a_12861_44030# a_15493_43396# 0.254093f
C4818 a_n1151_42308# a_11309_47204# 0.546434f
C4819 a_4915_47217# a_n881_46662# 1.23372f
C4820 a_18479_47436# a_18597_46090# 0.473843f
C4821 a_3754_39964# VDAC_Pi 0.296508f
C4822 a_2479_44172# a_1847_42826# 0.141223f
C4823 a_2437_43646# a_3357_43084# 0.424652f
C4824 a_22223_45572# a_19479_31679# 0.155323f
C4825 a_2711_45572# a_18184_42460# 0.367034f
C4826 a_3357_43084# SINGLE_ENDED 0.131897f
C4827 a_22959_45572# VDD 0.304443f
C4828 a_12465_44636# a_13059_46348# 0.163448f
C4829 a_10227_46804# a_20107_46660# 0.312495f
C4830 C6_N_btm VREF 1.41944f
C4831 C7_N_btm VIN_N 1.52449f
C4832 VDD DATA[4] 0.326957f
C4833 C4_N_btm VCM 0.716447f
C4834 C5_N_btm VREF_GND 0.676559f
C4835 a_4190_30871# a_743_42282# 0.18536f
C4836 a_18494_42460# a_20512_43084# 0.115057f
C4837 a_19319_43548# VDD 0.561461f
C4838 a_12465_44636# a_13556_45296# 0.248126f
C4839 a_2324_44458# a_526_44458# 0.279023f
C4840 a_5937_45572# a_8049_45260# 0.103218f
C4841 a_n1925_46634# VDD 0.783093f
C4842 a_2889_44172# a_2998_44172# 0.179664f
C4843 a_16795_42852# VDD 0.179044f
C4844 a_3218_45724# a_2711_45572# 0.1731f
C4845 a_4646_46812# a_5343_44458# 0.24395f
C4846 a_6755_46942# a_11691_44458# 0.192426f
C4847 a_10355_46116# VDD 0.222751f
C4848 a_n2810_45572# a_n2302_37984# 0.130495f
C4849 a_n2956_38216# a_n3420_37984# 0.208204f
C4850 a_n443_46116# a_4915_47217# 0.395101f
C4851 a_4791_45118# a_5129_47502# 0.240381f
C4852 a_4958_30871# VCM 0.642743f
C4853 a_7174_31319# RST_Z 0.216004f
C4854 a_1823_45246# a_n2661_42834# 0.174801f
C4855 a_n2472_46634# a_n2442_46660# 0.155358f
C4856 a_6886_37412# VDD 0.235486f
C4857 a_n97_42460# a_5755_42852# 0.149651f
C4858 a_n2661_46098# a_1176_45822# 0.144277f
C4859 a_2107_46812# a_3483_46348# 0.100707f
C4860 a_3232_43370# a_1414_42308# 0.248035f
C4861 a_10949_43914# VDD 0.797824f
C4862 a_5937_45572# a_8953_45546# 0.3871f
C4863 a_20894_47436# VDD 0.188358f
C4864 a_n2661_42834# a_n3674_39768# 0.150968f
C4865 a_9290_44172# a_10907_45822# 0.262972f
C4866 a_768_44030# a_742_44458# 0.216263f
C4867 a_20411_46873# VDD 0.348821f
C4868 a_19647_42308# a_13258_32519# 0.153411f
C4869 a_22775_42308# a_22465_38105# 0.330766f
C4870 a_3483_46348# a_n2661_44458# 1.44355f
C4871 a_12549_44172# a_11341_43940# 0.406618f
C4872 a_n755_45592# a_n1059_45260# 0.53237f
C4873 a_n357_42282# a_n913_45002# 0.309845f
C4874 a_n443_46116# a_1568_43370# 0.584982f
C4875 a_n1151_42308# a_4955_46873# 0.261025f
C4876 a_n356_44636# a_6123_31319# 0.169259f
C4877 a_3537_45260# a_4574_45260# 0.234297f
C4878 a_16327_47482# a_18083_42858# 0.591108f
C4879 a_11599_46634# a_13351_46090# 0.105205f
C4880 a_4646_46812# a_3090_45724# 0.199722f
C4881 a_n1613_43370# a_n1853_46287# 0.354256f
C4882 a_13507_46334# a_18907_42674# 0.202065f
C4883 a_18597_46090# a_19511_42282# 0.156698f
C4884 a_3422_30871# VDD 1.12305f
C4885 a_15227_44166# a_6945_45028# 0.548194f
C4886 a_n2288_47178# VDD 0.29372f
C4887 a_3090_45724# a_18479_45785# 0.259218f
C4888 a_3877_44458# a_2382_45260# 0.395451f
C4889 a_11415_45002# a_11652_45724# 0.128811f
C4890 a_11453_44696# a_17719_45144# 0.105851f
C4891 a_8953_45546# a_n443_42852# 0.134632f
C4892 a_2324_44458# a_8953_45002# 1.65784f
C4893 a_3090_45724# a_10057_43914# 0.230475f
C4894 a_n443_46116# a_n881_46662# 0.114922f
C4895 a_4915_47217# a_n1613_43370# 0.195064f
C4896 a_19963_31679# VDD 0.605279f
C4897 a_12861_44030# a_18280_46660# 0.140921f
C4898 a_n2661_46634# a_6755_46942# 1.40968f
C4899 C5_N_btm VREF 0.987144f
C4900 C6_N_btm VIN_N 0.391905f
C4901 VDD DATA[3] 0.309692f
C4902 C3_N_btm VCM 0.716273f
C4903 C4_N_btm VREF_GND 0.671882f
C4904 a_5111_44636# a_5518_44484# 0.124556f
C4905 a_7640_43914# VDD 0.196713f
C4906 a_768_44030# a_13259_45724# 0.315247f
C4907 a_13076_44458# a_13213_44734# 0.126609f
C4908 a_11823_42460# a_14205_43396# 0.176571f
C4909 a_4791_45118# a_n2661_43370# 0.408007f
C4910 a_n2312_38680# VDD 0.540248f
C4911 a_4921_42308# a_5755_42308# 0.175841f
C4912 a_2675_43914# a_2998_44172# 0.173844f
C4913 a_16414_43172# VDD 0.201389f
C4914 a_768_44030# a_n2661_43922# 1.9176f
C4915 a_12549_44172# a_n2293_43922# 0.194293f
C4916 a_9823_46155# VDD 0.102474f
C4917 a_4791_45118# a_4915_47217# 0.226891f
C4918 a_2063_45854# a_9863_47436# 0.12173f
C4919 a_7174_31319# VDD 0.669838f
C4920 a_12741_44636# a_14673_44172# 0.178572f
C4921 VDAC_N C10_N_btm 0.24639p
C4922 a_5700_37509# VDD 1.0734f
C4923 a_n237_47217# a_n755_45592# 0.286948f
C4924 a_10729_43914# VDD 0.681371f
C4925 a_n2840_46090# a_n2956_39304# 0.158668f
C4926 a_8199_44636# a_8953_45546# 0.71291f
C4927 a_10227_46804# a_3357_43084# 0.305304f
C4928 a_19787_47423# VDD 0.256911f
C4929 a_21487_43396# VDD 0.222231f
C4930 a_n1613_43370# a_5883_43914# 0.352323f
C4931 a_20107_46660# VDD 0.442554f
C4932 a_5934_30871# C5_N_btm 0.139996f
C4933 a_5932_42308# VDD 0.534416f
C4934 a_12549_44172# a_21115_43940# 0.211261f
C4935 a_n357_42282# a_n1059_45260# 7.3759f
C4936 a_12741_44636# a_12607_44458# 0.134974f
C4937 a_1609_45822# a_2437_43646# 0.189329f
C4938 a_16327_47482# a_n743_46660# 0.53683f
C4939 a_n971_45724# a_7411_46660# 0.567031f
C4940 a_n1613_43370# a_n881_46662# 1.06426f
C4941 a_10227_46804# a_5342_30871# 0.163388f
C4942 a_3357_43084# a_1307_43914# 0.197864f
C4943 a_1423_45028# VDD 4.06861f
C4944 a_n881_46662# a_n2293_46098# 0.291354f
C4945 a_n1613_43370# a_n2157_46122# 0.296124f
C4946 a_3877_44458# a_3090_45724# 0.23348f
C4947 a_4915_47217# a_6945_45028# 0.207881f
C4948 a_n743_46660# a_n356_45724# 0.223429f
C4949 a_12861_44030# a_15903_45785# 0.156145f
C4950 a_13059_46348# a_10903_43370# 0.11738f
C4951 a_n2497_47436# VDD 1.33346f
C4952 a_3090_45724# a_18175_45572# 0.130163f
C4953 a_n2293_46634# a_1307_43914# 0.184387f
C4954 a_13575_42558# a_14113_42308# 0.11418f
C4955 a_10193_42453# a_11551_42558# 0.228057f
C4956 a_2324_44458# a_8191_45002# 0.120399f
C4957 a_4791_45118# a_n881_46662# 0.429542f
C4958 a_n443_46116# a_n1613_43370# 0.410263f
C4959 a_12861_44030# a_11453_44696# 0.173308f
C4960 a_15493_43396# a_15743_43084# 0.517624f
C4961 a_2437_43646# a_22223_45572# 0.165664f
C4962 a_22591_45572# VDD 0.314172f
C4963 a_584_46384# a_1138_42852# 0.491749f
C4964 a_n443_46116# a_n2293_46098# 0.251135f
C4965 C4_N_btm VREF 0.98728f
C4966 C5_N_btm VIN_N 0.502041f
C4967 VDD DATA[2] 0.3216f
C4968 C2_N_btm VCM 0.716172f
C4969 C3_N_btm VREF_GND 0.67174f
C4970 a_5111_44636# a_5343_44458# 0.477401f
C4971 a_6109_44484# VDD 0.243629f
C4972 a_12549_44172# a_13259_45724# 0.110646f
C4973 a_n1151_42308# a_10193_42453# 0.238612f
C4974 a_11823_42460# a_14358_43442# 0.122636f
C4975 a_6945_45028# a_10809_44734# 0.953135f
C4976 a_21076_30879# a_20692_30879# 0.117886f
C4977 a_n2104_46634# VDD 0.286113f
C4978 a_15567_42826# VDD 0.163583f
C4979 a_768_44030# a_n2661_42834# 4.99505f
C4980 a_9569_46155# VDD 0.19288f
C4981 a_n2956_38216# a_n3565_38216# 0.307285f
C4982 a_4791_45118# a_n443_46116# 0.115639f
C4983 a_n3565_39304# a_n4209_38502# 5.79402f
C4984 a_20712_42282# VDD 0.282526f
C4985 a_7227_45028# a_6709_45028# 0.115677f
C4986 a_n2956_39768# a_n2442_46660# 6.5214f
C4987 a_10227_46804# a_6755_46942# 0.778648f
C4988 VDAC_N C9_N_btm 0.123386p
C4989 a_5088_37509# VDD 1.15925f
C4990 a_n1151_42308# a_n784_42308# 0.154055f
C4991 a_3065_45002# a_n2661_43370# 0.356646f
C4992 a_4185_45028# a_20974_43370# 0.184625f
C4993 a_n881_46662# a_6945_45028# 0.239384f
C4994 a_n746_45260# a_n755_45592# 0.172774f
C4995 a_14543_43071# a_5534_30871# 0.196814f
C4996 a_2382_45260# a_3905_42865# 0.291572f
C4997 a_10405_44172# VDD 0.408512f
C4998 a_4791_45118# a_3537_45260# 0.33264f
C4999 a_8016_46348# a_9625_46129# 0.128435f
C5000 a_8199_44636# a_5937_45572# 0.573373f
C5001 a_19386_47436# VDD 0.121241f
C5002 a_n1736_42282# a_n4318_37592# 0.153911f
C5003 a_20556_43646# VDD 0.34939f
C5004 a_19551_46910# VDD 0.226848f
C5005 a_n913_45002# a_1755_42282# 0.169955f
C5006 a_6171_42473# VDD 0.184622f
C5007 a_12549_44172# a_20935_43940# 0.110704f
C5008 a_n357_42282# a_n2017_45002# 0.580077f
C5009 a_n2293_45546# a_n967_45348# 0.119714f
C5010 a_n1151_42308# a_4646_46812# 0.330834f
C5011 a_12465_44636# a_13661_43548# 0.106973f
C5012 comp_n VDD 0.504719f
C5013 a_3429_45260# a_3537_45260# 0.138977f
C5014 a_11599_46634# a_12005_46116# 0.27095f
C5015 a_10467_46802# a_6755_46942# 0.256039f
C5016 a_4883_46098# a_4704_46090# 0.1774f
C5017 a_10193_42453# a_15493_43940# 0.597095f
C5018 a_20980_44850# VDD 0.132317f
C5019 a_13661_43548# a_2711_45572# 0.552383f
C5020 a_15227_44166# a_20708_46348# 0.106656f
C5021 a_n2833_47464# VDD 0.461379f
C5022 a_9313_44734# a_11967_42832# 0.216837f
C5023 a_4791_45118# a_8701_44490# 0.138973f
C5024 a_4185_45028# a_2711_45572# 0.102913f
C5025 a_13507_46334# a_18494_42460# 0.234442f
C5026 a_8034_45724# a_8049_45260# 0.141057f
C5027 a_11415_45002# a_11322_45546# 0.527707f
C5028 a_3483_46348# a_4099_45572# 0.15767f
C5029 a_6969_46634# VDD 0.154507f
C5030 a_13575_42558# a_13657_42558# 0.171361f
C5031 a_16922_45042# a_20749_43396# 0.106779f
C5032 a_10193_42453# a_5742_30871# 0.303452f
C5033 a_10903_43370# a_9482_43914# 1.20611f
C5034 a_n1151_42308# a_9804_47204# 0.108722f
C5035 a_4791_45118# a_n1613_43370# 0.223884f
C5036 a_18143_47464# a_18479_47436# 0.238309f
C5037 a_584_46384# a_768_44030# 0.105366f
C5038 a_2113_38308# VDAC_Pi 0.170908f
C5039 a_1209_43370# a_1049_43396# 0.194938f
C5040 a_n97_42460# a_n1557_42282# 0.149645f
C5041 a_13259_45724# a_13076_44458# 0.188498f
C5042 a_13059_46348# a_13483_43940# 0.124566f
C5043 a_17715_44484# a_17517_44484# 0.163303f
C5044 a_526_44458# a_3363_44484# 0.119556f
C5045 a_2437_43646# SINGLE_ENDED 0.117817f
C5046 a_3357_43084# VDD 1.66202f
C5047 a_4791_45118# a_n2293_46098# 0.411939f
C5048 C3_N_btm VREF 0.984942f
C5049 VDD DATA[1] 0.321585f
C5050 C4_N_btm VIN_N 0.50261f
C5051 C1_N_btm VCM 0.716121f
C5052 C2_N_btm VREF_GND 0.671742f
C5053 a_21259_43561# a_4190_30871# 0.198353f
C5054 a_3537_45260# a_8103_44636# 0.140404f
C5055 a_12891_46348# a_13259_45724# 1.04614f
C5056 a_17339_46660# a_18285_46348# 0.184197f
C5057 a_4361_42308# a_3823_42558# 0.114877f
C5058 a_11823_42460# a_14579_43548# 0.106967f
C5059 a_6945_45028# a_22223_46124# 0.17119f
C5060 a_765_45546# a_n443_42852# 0.232932f
C5061 a_n2293_46634# VDD 1.52629f
C5062 a_n784_42308# a_5742_30871# 0.550812f
C5063 a_n1761_44111# a_n1644_44306# 0.170098f
C5064 a_5342_30871# VDD 0.496295f
C5065 a_n443_46116# a_895_43940# 0.163929f
C5066 a_16375_45002# a_10193_42453# 0.125364f
C5067 a_9625_46129# VDD 0.996485f
C5068 a_4700_47436# a_n443_46116# 0.255594f
C5069 a_20107_42308# VDD 0.284252f
C5070 a_10227_46804# a_10249_46116# 0.137273f
C5071 VDAC_N C8_N_btm 61.723f
C5072 a_4338_37500# VDD 0.525635f
C5073 a_3726_37500# RST_Z 1.60318f
C5074 EN_VIN_BSTR_P a_n83_35174# 0.652984f
C5075 a_16237_45028# VDD 0.248452f
C5076 a_n971_45724# a_n755_45592# 0.347347f
C5077 a_2382_45260# a_3600_43914# 0.158274f
C5078 a_9672_43914# VDD 0.150499f
C5079 a_14035_46660# a_14180_46482# 0.157972f
C5080 a_18479_47436# START 0.313639f
C5081 a_18597_46090# VDD 0.930122f
C5082 a_n3674_38216# a_n4318_37592# 2.7294f
C5083 a_19279_43940# a_21398_44850# 0.183186f
C5084 a_743_42282# VDD 0.597869f
C5085 a_4646_46812# a_n2293_42834# 0.152973f
C5086 a_19123_46287# VDD 0.336379f
C5087 a_5755_42308# VDD 0.229304f
C5088 a_n755_45592# a_n2293_45010# 0.159033f
C5089 a_15143_45578# a_15037_45618# 0.13675f
C5090 a_2277_45546# VDD 0.209584f
C5091 a_12465_44636# a_5807_45002# 0.59474f
C5092 a_8530_39574# CAL_N 0.644218f
C5093 a_1736_39043# VDD 2.8939f
C5094 a_3065_45002# a_3537_45260# 0.162384f
C5095 a_10227_46804# a_5534_30871# 0.304847f
C5096 a_626_44172# VDD 0.621601f
C5097 a_10623_46897# a_10554_47026# 0.209641f
C5098 a_10428_46928# a_6755_46942# 0.155315f
C5099 a_10467_46802# a_10249_46116# 0.12624f
C5100 a_11599_46634# a_10903_43370# 0.439916f
C5101 a_n2661_46634# a_765_45546# 1.82448f
C5102 a_4791_45118# a_6945_45028# 0.493927f
C5103 a_526_44458# a_9803_43646# 0.170855f
C5104 a_14035_46660# a_13925_46122# 0.207108f
C5105 a_n2472_46090# a_n2293_46098# 0.176709f
C5106 w_11334_34010# VDD 1.90683f
C5107 a_13291_42460# a_14635_42282# 0.111986f
C5108 a_n2293_42282# a_n1630_35242# 0.18361f
C5109 a_5649_42852# a_4958_30871# 0.293366f
C5110 a_n913_45002# a_3539_42460# 0.359316f
C5111 a_13507_46334# a_18184_42460# 0.505552f
C5112 a_6755_46942# VDD 1.05713f
C5113 a_526_44458# a_n913_45002# 0.250864f
C5114 a_5937_45572# a_1307_43914# 0.101589f
C5115 a_8049_45260# VDD 1.89366f
C5116 a_n1151_42308# a_8128_46384# 0.328697f
C5117 a_11599_46634# a_4883_46098# 0.261488f
C5118 a_13717_47436# SMPL_ON_N 0.132417f
C5119 a_10227_46804# a_18479_47436# 1.40697f
C5120 a_19692_46634# a_15493_43940# 0.16692f
C5121 a_19479_31679# VDD 0.579914f
C5122 a_2437_43646# START 0.12936f
C5123 a_13507_46334# a_13059_46348# 0.192049f
C5124 a_n971_45724# a_3483_46348# 0.211534f
C5125 C2_N_btm VREF 0.987884f
C5126 VDD DATA[0] 1.05526f
C5127 C3_N_btm VIN_N 0.455045f
C5128 C0_N_btm VCM 0.717064f
C5129 C1_N_btm VREF_GND 0.673422f
C5130 a_2063_45854# a_11322_45546# 0.105268f
C5131 a_n743_46660# a_5066_45546# 0.124676f
C5132 a_14543_43071# a_13291_42460# 0.107887f
C5133 a_3232_43370# a_11341_43940# 0.112367f
C5134 a_11823_42460# a_13667_43396# 0.107673f
C5135 a_15037_43940# VDD 0.190221f
C5136 a_3090_45724# a_7499_43078# 0.23734f
C5137 a_n2442_46660# VDD 0.693209f
C5138 a_5379_42460# a_5932_42308# 0.761308f
C5139 a_11967_42832# a_15682_43940# 1.63211f
C5140 a_15279_43071# VDD 0.189193f
C5141 a_n3674_37592# a_n3420_37984# 0.172946f
C5142 a_11415_45002# a_6171_45002# 1.05801f
C5143 a_16327_47482# a_3422_30871# 0.220296f
C5144 a_n443_46116# a_2479_44172# 0.732848f
C5145 a_n755_45592# a_2711_45572# 0.168218f
C5146 a_6755_46942# a_11827_44484# 0.529579f
C5147 a_8953_45546# VDD 1.32809f
C5148 a_n2956_38216# a_n4209_38216# 0.232905f
C5149 a_4700_47436# a_4791_45118# 0.31818f
C5150 a_13258_32519# VDD 3.19231f
C5151 a_11415_45002# a_14673_44172# 0.229077f
C5152 a_10227_46804# a_10554_47026# 0.166977f
C5153 VDAC_N C7_N_btm 30.844f
C5154 a_3726_37500# VDD 0.341303f
C5155 a_n923_35174# a_n83_35174# 0.480251f
C5156 a_20193_45348# VDD 0.793111f
C5157 a_n971_45724# a_n357_42282# 0.271282f
C5158 a_584_46384# a_n2661_45546# 0.100439f
C5159 a_3090_45724# a_15227_44166# 0.428743f
C5160 a_n746_45260# a_310_45028# 0.378188f
C5161 a_9028_43914# VDD 0.17194f
C5162 a_10227_46804# a_2437_43646# 0.150025f
C5163 a_18780_47178# VDD 0.245515f
C5164 a_17701_42308# a_17531_42308# 0.109201f
C5165 a_11967_42832# a_20512_43084# 0.106819f
C5166 a_n1059_45260# a_15743_43084# 0.101833f
C5167 a_20301_43646# VDD 0.296691f
C5168 a_3090_45724# a_4558_45348# 0.147318f
C5169 a_18285_46348# VDD 0.259614f
C5170 a_6123_31319# C4_N_btm 0.132906f
C5171 a_20692_30879# a_413_45260# 0.111034f
C5172 a_1609_45822# VDD 0.270106f
C5173 a_20894_47436# a_20843_47204# 0.134298f
C5174 a_1239_39043# VDD 0.507578f
C5175 a_2437_43646# a_1307_43914# 0.160142f
C5176 a_n357_42282# a_9313_44734# 5.02008f
C5177 a_10428_46928# a_10249_46116# 0.704177f
C5178 a_n237_47217# a_n1925_42282# 0.109762f
C5179 a_10227_46804# a_8199_44636# 0.460391f
C5180 a_12465_44636# a_3483_46348# 0.210833f
C5181 a_4185_45028# a_5649_42852# 8.049951f
C5182 a_13507_46334# a_17303_42282# 1.68549f
C5183 a_14035_46660# a_13759_46122# 0.162408f
C5184 w_1575_34946# VDD 1.58877f
C5185 a_n2312_38680# a_n3565_39304# 0.418567f
C5186 a_n913_45002# a_3626_43646# 0.104422f
C5187 a_3232_43370# a_n97_42460# 0.113391f
C5188 a_3483_46348# a_2711_45572# 0.167588f
C5189 a_10249_46116# VDD 1.03004f
C5190 a_13717_47436# a_22731_47423# 0.109987f
C5191 a_10227_46804# a_18143_47464# 0.112443f
C5192 a_2063_45854# a_11309_47204# 0.141276f
C5193 a_n97_42460# a_4905_42826# 0.147727f
C5194 a_13259_45724# a_12607_44458# 0.132105f
C5195 a_22223_45572# VDD 0.287831f
C5196 a_n2109_47186# a_5164_46348# 0.603312f
C5197 a_584_46384# a_805_46414# 0.135394f
C5198 C1_N_btm VREF 0.98698f
C5199 VDD CLK_DATA 0.422202f
C5200 C2_N_btm VIN_N 0.502408f
C5201 C0_dummy_N_btm VCM 0.311452f
C5202 C0_N_btm VREF_GND 0.350401f
C5203 a_5111_44636# a_4223_44672# 0.418299f
C5204 a_17339_46660# a_765_45546# 0.244447f
C5205 a_n2312_39304# a_n3565_39590# 0.491833f
C5206 a_13565_43940# VDD 0.175245f
C5207 a_20820_30879# a_20692_30879# 8.973741f
C5208 a_8199_44636# a_8034_45724# 0.127067f
C5209 a_n2472_46634# VDD 0.287589f
C5210 a_5379_42460# a_6171_42473# 0.110293f
C5211 a_n913_45002# a_8037_42858# 0.316376f
C5212 a_5534_30871# VDD 0.513761f
C5213 a_3090_45724# a_n2661_43370# 0.101361f
C5214 a_n443_46116# a_2127_44172# 0.196411f
C5215 a_n2810_45572# a_n3565_38216# 0.104999f
C5216 a_5937_45572# VDD 2.20055f
C5217 a_19647_42308# VDD 0.227331f
C5218 a_n2840_46634# a_n2661_46634# 0.180867f
C5219 a_10227_46804# a_10623_46897# 0.180903f
C5220 VDAC_N C6_N_btm 15.440799f
C5221 a_n1532_35090# a_n83_35174# 0.558402f
C5222 a_n923_35174# EN_VIN_BSTR_P 1.02927f
C5223 a_n1151_42308# a_n961_42308# 0.109068f
C5224 a_5111_44636# a_n2293_42834# 0.110286f
C5225 a_11691_44458# VDD 3.25709f
C5226 a_10193_42453# a_n97_42460# 0.304653f
C5227 a_8333_44056# VDD 0.124235f
C5228 a_8016_46348# a_8199_44636# 0.33718f
C5229 a_18479_47436# VDD 1.47669f
C5230 a_n4318_38216# a_n4318_37592# 0.139499f
C5231 a_4190_30871# VDD 1.36846f
C5232 a_17829_46910# VDD 0.37446f
C5233 a_742_44458# a_2905_42968# 0.15065f
C5234 a_11341_43940# a_14021_43940# 3.06514f
C5235 a_n2956_38216# a_n2956_37592# 0.103811f
C5236 a_n863_45724# a_n913_45002# 0.565852f
C5237 a_n443_42852# VDD 3.69394f
C5238 a_4883_46098# a_5807_45002# 1.76125f
C5239 a_n97_42460# a_16137_43396# 0.134668f
C5240 a_n2293_43922# a_n784_42308# 1.67292f
C5241 a_10227_46804# a_13460_43230# 0.243111f
C5242 a_2382_45260# a_3537_45260# 0.250657f
C5243 a_3483_46348# a_15682_43940# 0.261013f
C5244 a_375_42282# VDD 0.591443f
C5245 a_10428_46928# a_10554_47026# 0.181217f
C5246 a_10467_46802# a_10623_46897# 0.107482f
C5247 a_12861_44030# a_12594_46348# 0.43362f
C5248 a_n237_47217# a_526_44458# 0.198088f
C5249 a_7715_46873# a_7832_46660# 0.157972f
C5250 a_11827_44484# a_11691_44458# 0.881979f
C5251 a_3232_43370# a_n2661_43922# 0.197944f
C5252 a_n4318_39304# a_n3420_39616# 0.256393f
C5253 a_12465_44636# a_13249_42308# 0.541909f
C5254 a_6655_43762# VDD 0.132357f
C5255 a_10554_47026# VDD 0.205847f
C5256 a_5891_43370# a_6293_42852# 0.107308f
C5257 a_10193_42453# a_10533_42308# 0.101629f
C5258 a_14635_42282# VDD 0.369964f
C5259 a_3090_45724# a_5883_43914# 0.132458f
C5260 a_16375_45002# a_16147_45260# 1.01554f
C5261 a_12861_44030# a_12465_44636# 0.242761f
C5262 a_11599_46634# a_13507_46334# 0.259318f
C5263 a_n97_42460# a_3080_42308# 0.353977f
C5264 a_14021_43940# a_10341_43396# 1.5617f
C5265 a_11967_42832# a_17333_42852# 0.14149f
C5266 a_2437_43646# VDD 1.17411f
C5267 a_n881_46662# a_3090_45724# 0.107805f
C5268 a_584_46384# a_472_46348# 0.31609f
C5269 C0_N_btm VREF 0.443884f
C5270 VDD SINGLE_ENDED 0.210835f
C5271 C1_N_btm VIN_N 0.39234f
C5272 C0_dummy_P_btm VCM 0.311452f
C5273 a_3537_45260# a_5343_44458# 0.378482f
C5274 a_12861_44030# a_2711_45572# 0.104124f
C5275 a_n1925_46634# a_5066_45546# 0.195997f
C5276 a_8975_43940# a_n2661_43922# 0.11532f
C5277 a_n2661_46634# VDD 2.23057f
C5278 a_2479_44172# a_895_43940# 0.318312f
C5279 a_n2472_43914# a_n3674_39768# 0.162742f
C5280 a_1414_42308# a_2998_44172# 0.447595f
C5281 a_14543_43071# VDD 0.18866f
C5282 a_13259_45724# a_10193_42453# 0.284945f
C5283 a_8199_44636# VDD 1.43837f
C5284 a_n1741_47186# a_11599_46634# 0.164599f
C5285 a_1343_38525# a_2112_39137# 0.22564f
C5286 a_19511_42282# VDD 0.244902f
C5287 a_11823_42460# a_n913_45002# 0.281323f
C5288 a_n2840_46634# a_n2956_39768# 0.156182f
C5289 a_n1613_43370# a_3524_46660# 0.28004f
C5290 a_10227_46804# a_10467_46802# 0.678578f
C5291 VDAC_N C5_N_btm 7.72452f
C5292 a_n1532_35090# EN_VIN_BSTR_P 0.340449f
C5293 a_n1151_42308# a_n1329_42308# 0.167748f
C5294 a_12549_44172# a_2324_44458# 0.506903f
C5295 a_n971_45724# a_n1099_45572# 0.508925f
C5296 a_13635_43156# a_13460_43230# 0.234322f
C5297 a_n97_42460# a_15764_42576# 0.174403f
C5298 a_8016_46348# a_8349_46414# 0.232167f
C5299 a_16327_47482# a_3357_43084# 0.114502f
C5300 a_3483_46348# a_10903_43370# 0.404121f
C5301 a_18143_47464# VDD 0.388551f
C5302 a_n2104_42282# a_n3674_38216# 0.155459f
C5303 a_21259_43561# VDD 0.192954f
C5304 a_3090_45724# a_3537_45260# 0.198803f
C5305 a_765_45546# VDD 2.19953f
C5306 a_21613_42308# a_22775_42308# 0.225363f
C5307 en_comp a_n1630_35242# 2.31448f
C5308 a_1467_44172# a_1756_43548# 0.100052f
C5309 a_4921_42308# VDD 0.214995f
C5310 a_1606_42308# VCM 0.152876f
C5311 a_12549_44172# a_19862_44208# 0.262561f
C5312 a_n2956_38216# a_n2810_45028# 5.73989f
C5313 a_n863_45724# a_n1059_45260# 0.162875f
C5314 a_509_45822# VDD 0.190119f
C5315 a_11599_46634# a_n743_46660# 0.248412f
C5316 a_9313_45822# a_2107_46812# 0.298046f
C5317 a_19787_47423# a_19594_46812# 0.108653f
C5318 a_8530_39574# a_8912_37509# 0.426772f
C5319 a_10227_46804# a_13635_43156# 0.320228f
C5320 a_2680_45002# a_3065_45002# 0.13328f
C5321 a_3483_46348# a_14955_43940# 0.242667f
C5322 a_16751_45260# VDD 0.121848f
C5323 a_10428_46928# a_10623_46897# 0.21686f
C5324 a_13507_46334# a_4185_45028# 0.479559f
C5325 a_4883_46098# a_3483_46348# 0.813604f
C5326 a_15743_43084# a_19339_43156# 0.128224f
C5327 a_3232_43370# a_n2661_42834# 0.127534f
C5328 a_n913_45002# a_2982_43646# 0.498826f
C5329 a_n699_43396# a_2998_44172# 0.127437f
C5330 a_5534_30871# a_n3420_39072# 0.339008f
C5331 a_2063_45854# a_8975_43940# 0.149528f
C5332 a_20202_43084# a_10193_42453# 0.296862f
C5333 a_10623_46897# VDD 0.189083f
C5334 a_13291_42460# VDD 0.546706f
C5335 a_10903_43370# a_11963_45334# 0.209081f
C5336 a_2324_44458# a_5205_44484# 0.523531f
C5337 a_9290_44172# a_9482_43914# 0.135239f
C5338 a_16327_47482# a_18597_46090# 1.28053f
C5339 a_17591_47464# a_10227_46804# 0.292864f
C5340 a_11967_42832# a_18083_42858# 0.472348f
C5341 a_7499_43078# a_n2293_42834# 0.352878f
C5342 a_21513_45002# VDD 0.416919f
C5343 a_584_46384# a_376_46348# 0.232754f
C5344 a_n237_47217# a_167_45260# 0.280171f
C5345 C0_P_btm VCM 0.717283f
C5346 C0_N_btm VIN_N 0.529671f
C5347 VDD START 0.114358f
C5348 a_n443_42852# a_n2661_42282# 0.133617f
C5349 a_15227_44166# a_12741_44636# 0.250453f
C5350 a_3090_45724# a_n2293_46098# 0.642755f
C5351 a_2063_45854# a_10193_42453# 0.114552f
C5352 a_11823_42460# a_9145_43396# 0.146085f
C5353 a_18184_42460# a_3422_30871# 0.649102f
C5354 a_4190_30871# a_n3420_39072# 0.10848f
C5355 a_8016_46348# a_8034_45724# 0.254614f
C5356 a_n2956_39768# VDD 0.697168f
C5357 a_n755_45592# a_6123_31319# 0.199766f
C5358 a_2127_44172# a_895_43940# 0.132679f
C5359 a_1414_42308# a_2889_44172# 0.128883f
C5360 a_13460_43230# VDD 0.276534f
C5361 a_n443_46116# a_1414_42308# 0.18376f
C5362 a_n2810_45572# a_n4209_38216# 0.195791f
C5363 a_8349_46414# VDD 0.209819f
C5364 a_n1151_42308# a_4915_47217# 0.1374f
C5365 a_n971_45724# a_n1435_47204# 2.23698f
C5366 a_n4064_39072# a_n2302_39072# 0.250408f
C5367 a_n356_44636# a_5342_30871# 0.133551f
C5368 a_11823_42460# a_n1059_45260# 0.100641f
C5369 a_4791_45118# a_3090_45724# 0.206257f
C5370 a_n1613_43370# a_3699_46634# 0.344308f
C5371 VDAC_N C4_N_btm 3.92765f
C5372 a_n1532_35090# a_n923_35174# 0.400297f
C5373 a_n1386_35608# EN_VIN_BSTR_P 0.573134f
C5374 a_5691_45260# a_5837_45028# 0.171361f
C5375 a_22959_45036# VDD 0.30999f
C5376 a_11813_46116# a_12156_46660# 0.157972f
C5377 a_16327_47482# a_8049_45260# 0.605463f
C5378 a_12545_42858# a_5534_30871# 0.17182f
C5379 a_n357_42282# a_8685_43396# 0.319118f
C5380 a_15227_44166# a_16375_45002# 0.117865f
C5381 a_584_46384# a_3232_43370# 0.277433f
C5382 a_10227_46804# VDD 2.77567f
C5383 a_n4318_38216# a_n3674_38216# 2.91597f
C5384 a_4190_30871# C10_N_btm 0.446355f
C5385 a_12594_46348# a_13527_45546# 0.100424f
C5386 a_6755_46942# a_14537_43396# 0.120241f
C5387 a_10903_43370# a_13249_42308# 0.211356f
C5388 a_17339_46660# VDD 0.555596f
C5389 a_9313_44734# a_15743_43084# 1.48048f
C5390 a_742_44458# a_1847_42826# 0.372436f
C5391 a_n3674_39768# a_n4318_39304# 2.75695f
C5392 a_5742_30871# EN_VIN_BSTR_N 0.643089f
C5393 a_10193_42453# a_15861_45028# 0.432483f
C5394 a_n863_45724# a_n2017_45002# 0.111825f
C5395 a_13507_46334# a_5807_45002# 1.64614f
C5396 a_7754_38470# a_8912_37509# 0.575911f
C5397 a_n2302_39072# VDD 0.355374f
C5398 a_n4064_39616# VREF_GND 0.241027f
C5399 a_2382_45260# a_3065_45002# 0.632538f
C5400 a_10227_46804# a_12895_43230# 0.152365f
C5401 a_3483_46348# a_13483_43940# 0.194464f
C5402 a_1307_43914# VDD 3.92807f
C5403 a_10428_46928# a_10467_46802# 0.820079f
C5404 a_n971_45724# a_526_44458# 0.21769f
C5405 a_12861_44030# a_10903_43370# 0.378457f
C5406 a_n1151_42308# a_10809_44734# 0.334692f
C5407 a_626_44172# a_n356_44636# 0.249281f
C5408 a_18579_44172# VDD 0.38178f
C5409 a_n2438_43548# a_n755_45592# 0.213107f
C5410 a_15227_44166# a_18985_46122# 0.287996f
C5411 a_4190_30871# a_19332_42282# 0.154377f
C5412 a_5111_44636# a_n97_42460# 0.211832f
C5413 a_9396_43370# VDD 0.288403f
C5414 a_16327_47482# a_20193_45348# 0.359904f
C5415 a_4791_45118# a_4743_44484# 0.165321f
C5416 a_10467_46802# VDD 0.401016f
C5417 a_13003_42852# VDD 0.132655f
C5418 a_8034_45724# VDD 0.812726f
C5419 a_n1151_42308# a_n881_46662# 1.41446f
C5420 a_2063_45854# a_9804_47204# 0.249806f
C5421 a_8696_44636# a_3232_43370# 0.169534f
C5422 a_n746_45260# a_167_45260# 0.234425f
C5423 C0_P_btm VREF_GND 0.350485f
C5424 C1_P_btm VCM 0.716121f
C5425 VDD RST_Z 4.72146f
C5426 C0_dummy_N_btm VIN_N 0.544204f
C5427 a_3080_42308# a_n2293_42282# 0.122474f
C5428 a_19692_46634# a_20202_43084# 0.172738f
C5429 a_n2661_46098# a_n2956_38680# 0.123968f
C5430 a_n2840_46634# VDD 0.306342f
C5431 COMP_P a_5742_30871# 0.1094f
C5432 a_2127_44172# a_2479_44172# 0.168988f
C5433 a_453_43940# a_895_43940# 0.420851f
C5434 a_1414_42308# a_2675_43914# 0.305556f
C5435 a_n2840_43914# a_n4318_39768# 0.170372f
C5436 a_13635_43156# VDD 0.463701f
C5437 a_3483_46348# CLK 0.408122f
C5438 a_8016_46348# VDD 1.42798f
C5439 a_3815_47204# a_4007_47204# 0.224415f
C5440 a_11682_45822# VDD 0.316586f
C5441 a_n1613_43370# a_2959_46660# 0.187029f
C5442 a_10227_46804# a_10150_46912# 0.236747f
C5443 a_5807_45002# a_n743_46660# 0.669712f
C5444 VDAC_N C3_N_btm 1.98783f
C5445 a_n1386_35608# a_n923_35174# 0.201937f
C5446 a_21513_45002# a_21359_45002# 0.289039f
C5447 a_413_45260# a_n2661_43370# 1.31746f
C5448 a_22223_45036# VDD 0.300162f
C5449 a_n746_45260# a_n863_45724# 0.664707f
C5450 a_5343_44458# a_6298_44484# 0.128602f
C5451 a_4223_44672# a_5883_43914# 0.967973f
C5452 a_3357_43084# a_3499_42826# 0.134316f
C5453 a_9290_44172# a_10835_43094# 0.172486f
C5454 a_413_45260# a_2998_44172# 0.161528f
C5455 a_7920_46348# a_8016_46348# 0.318386f
C5456 a_17591_47464# VDD 0.421992f
C5457 a_3090_45724# a_3065_45002# 0.475346f
C5458 a_526_44458# a_2711_45572# 0.392618f
C5459 a_19332_42282# a_19511_42282# 0.174683f
C5460 a_9028_43914# a_9165_43940# 0.126609f
C5461 a_3905_42558# VDD 0.176395f
C5462 a_10193_42453# a_8696_44636# 0.225102f
C5463 a_3754_38470# VDAC_P 0.323951f
C5464 a_7754_38470# VDAC_N 0.110573f
C5465 a_8530_39574# a_6886_37412# 0.616015f
C5466 a_n4064_39072# VDD 1.74897f
C5467 a_10227_46804# a_13113_42826# 0.159547f
C5468 a_16019_45002# VDD 0.174085f
C5469 a_10150_46912# a_10467_46802# 0.102355f
C5470 a_11827_44484# a_22223_45036# 0.179208f
C5471 a_13249_42308# a_13483_43940# 0.193724f
C5472 a_15227_44166# a_18819_46122# 0.288885f
C5473 a_8791_43396# VDD 0.191045f
C5474 a_16327_47482# a_11691_44458# 0.536141f
C5475 a_10428_46928# VDD 0.278873f
C5476 a_18494_42460# a_743_42282# 0.476713f
C5477 a_2324_44458# a_6171_45002# 2.73828f
C5478 a_10809_44734# a_413_45260# 0.333257f
C5479 a_n1151_42308# a_n1613_43370# 1.19311f
C5480 a_16327_47482# a_18479_47436# 0.723416f
C5481 a_16327_47482# a_4190_30871# 0.335014f
C5482 a_n237_47217# a_1823_45246# 0.370766f
C5483 C1_P_btm VREF_GND 0.673422f
C5484 C2_P_btm VCM 0.716172f
C5485 C0_P_btm VREF 0.443926f
C5486 a_3422_30871# a_4958_30871# 0.101017f
C5487 a_3537_45260# a_4223_44672# 0.1907f
C5488 a_22612_30879# VDD 3.2377f
C5489 a_1414_42308# a_895_43940# 0.208524f
C5490 a_12895_43230# VDD 0.212352f
C5491 a_18189_46348# a_16147_45260# 0.129202f
C5492 a_7920_46348# VDD 0.100184f
C5493 a_3785_47178# a_4007_47204# 0.106797f
C5494 a_n1151_42308# a_4791_45118# 1.16458f
C5495 a_2063_45854# a_6151_47436# 0.448977f
C5496 a_1736_39587# a_2112_39137# 0.269796f
C5497 a_20512_43084# a_15743_43084# 0.761578f
C5498 a_13661_43548# a_19319_43548# 0.189089f
C5499 a_n1613_43370# a_3177_46902# 0.209276f
C5500 a_10227_46804# a_9863_46634# 0.278164f
C5501 VDAC_N C2_N_btm 1.03255f
C5502 a_n2302_37690# VDD 0.350133f
C5503 a_3537_45260# a_n2293_42834# 0.195818f
C5504 a_4927_45028# a_5093_45028# 0.143754f
C5505 a_11827_44484# VDD 0.615802f
C5506 a_n971_45724# a_n863_45724# 0.199707f
C5507 a_3090_45724# a_15368_46634# 0.440843f
C5508 a_12379_42858# a_5534_30871# 0.128429f
C5509 a_12545_42858# a_13460_43230# 0.118423f
C5510 a_n97_42460# a_14113_42308# 0.356407f
C5511 a_7499_43078# a_n97_42460# 0.212833f
C5512 a_413_45260# a_2889_44172# 0.127135f
C5513 a_n443_46116# a_413_45260# 0.369976f
C5514 a_4646_46812# a_7227_45028# 0.305597f
C5515 a_20820_30879# a_10809_44734# 0.234047f
C5516 a_16588_47582# VDD 0.282243f
C5517 a_19279_43940# a_18579_44172# 0.372064f
C5518 a_n1059_45260# a_17499_43370# 0.385066f
C5519 a_2324_44458# a_8746_45002# 0.34917f
C5520 a_4958_30871# a_7174_31319# 0.107892f
C5521 a_21335_42336# a_21613_42308# 0.110671f
C5522 a_n2293_46098# a_4223_44672# 0.422068f
C5523 a_n2109_47186# a_5257_43370# 0.153164f
C5524 a_n443_46116# a_2609_46660# 0.349838f
C5525 a_7754_38470# a_6886_37412# 0.180842f
C5526 a_3754_38470# a_8912_37509# 1.88278f
C5527 a_n2946_39072# VDD 0.383374f
C5528 a_8530_39574# a_5700_37509# 0.947638f
C5529 a_n3420_39616# VREF_GND 0.117023f
C5530 a_18494_42460# a_13258_32519# 0.298557f
C5531 a_n443_42852# a_n356_44636# 0.262144f
C5532 a_15595_45028# VDD 0.156299f
C5533 a_10150_46912# a_10428_46928# 0.118759f
C5534 a_n2293_46634# a_13059_46348# 0.207934f
C5535 a_18494_42460# a_20193_45348# 0.116597f
C5536 a_n4318_40392# a_n4318_39768# 2.73673f
C5537 a_8147_43396# VDD 0.393534f
C5538 a_4791_45118# a_4223_44672# 0.399086f
C5539 a_n1613_43370# a_n2293_42834# 0.123758f
C5540 a_10150_46912# VDD 0.284144f
C5541 a_7499_43078# a_10533_42308# 0.225871f
C5542 a_18184_42460# a_743_42282# 0.126294f
C5543 a_2324_44458# a_3232_43370# 0.410727f
C5544 a_526_44458# a_n2661_45010# 0.703081f
C5545 a_12861_44030# a_12429_44172# 0.108591f
C5546 a_12861_44030# a_13507_46334# 0.315418f
C5547 a_22465_38105# a_22609_38406# 0.20695f
C5548 a_15493_43396# a_16409_43396# 0.566182f
C5549 a_4185_45028# a_3422_30871# 0.176529f
C5550 a_11599_46634# a_20107_46660# 0.266678f
C5551 C2_P_btm VREF_GND 0.671742f
C5552 C3_P_btm VCM 0.716273f
C5553 C1_P_btm VREF 0.98698f
C5554 C0_dummy_P_btm VIN_P 0.544204f
C5555 a_8953_45546# a_5066_45546# 0.191859f
C5556 a_21588_30879# VDD 1.78413f
C5557 a_742_44458# a_1756_43548# 0.152145f
C5558 a_1414_42308# a_2479_44172# 0.110442f
C5559 a_13113_42826# VDD 0.217254f
C5560 a_3785_47178# a_3815_47204# 0.270823f
C5561 a_2905_45572# a_n443_46116# 0.14923f
C5562 a_n1605_47204# a_n1435_47204# 0.110832f
C5563 a_1343_38525# a_1736_39043# 0.310247f
C5564 a_n3420_39072# a_n4064_39072# 4.93427f
C5565 a_18214_42558# VDD 0.295211f
C5566 a_15861_45028# a_16147_45260# 0.146279f
C5567 a_10907_45822# VDD 0.352181f
C5568 a_21588_30879# a_22612_30879# 7.53611f
C5569 a_n1613_43370# a_2609_46660# 0.631348f
C5570 a_5807_45002# a_n1925_46634# 0.933976f
C5571 VDAC_N C1_N_btm 0.55675f
C5572 a_n4064_37440# VDD 1.65981f
C5573 a_21359_45002# VDD 0.319372f
C5574 a_6755_46942# a_13059_46348# 0.239671f
C5575 a_3090_45724# a_14976_45028# 0.730613f
C5576 a_n746_45260# a_n2293_45546# 0.404324f
C5577 a_n971_45724# a_n1079_45724# 0.150623f
C5578 VCM VSS 40.3061f
C5579 VREF_GND VSS 17.4801f
C5580 VREF VSS 8.26148f
C5581 VIN_N VSS 13.1286f
C5582 VIN_P VSS 13.1075f
C5583 CLK VSS 1.55797f
C5584 EN_OFFSET_CAL VSS 0.505642f
C5585 DATA[5] VSS 0.561058f
C5586 DATA[4] VSS 0.755679f
C5587 DATA[3] VSS 1.01838f
C5588 DATA[2] VSS 0.536983f
C5589 DATA[1] VSS 0.550109f
C5590 DATA[0] VSS 0.616231f
C5591 CLK_DATA VSS 0.488979f
C5592 SINGLE_ENDED VSS 0.60168f
C5593 START VSS 0.991673f
C5594 RST_Z VSS 11.389f
C5595 VDD VSS 0.586439p
C5596 C10_N_btm VSS 0.264623p 
C5597 C9_N_btm VSS 0.114604p 
C5598 C8_N_btm VSS 60.275196f 
C5599 C7_N_btm VSS 32.1635f 
C5600 C6_N_btm VSS 17.8701f 
C5601 C5_N_btm VSS 10.4595f 
C5602 C4_N_btm VSS 7.67475f 
C5603 C3_N_btm VSS 5.70165f 
C5604 C2_N_btm VSS 4.38917f 
C5605 C1_N_btm VSS 3.94093f 
C5606 C0_N_btm VSS 5.62287f 
C5607 C0_dummy_N_btm VSS 4.25425f 
C5608 C0_dummy_P_btm VSS 4.26067f 
C5609 C0_P_btm VSS 5.63256f 
C5610 C1_P_btm VSS 3.96779f 
C5611 C2_P_btm VSS 4.40877f 
C5612 C3_P_btm VSS 5.70398f 
C5613 C4_P_btm VSS 7.68867f 
C5614 C5_P_btm VSS 10.4672f 
C5615 C6_P_btm VSS 17.865099f 
C5616 C7_P_btm VSS 32.1589f 
C5617 C8_P_btm VSS 60.269897f 
C5618 C9_P_btm VSS 0.114595p 
C5619 C10_P_btm VSS 0.264633p 
C5620 a_21589_35634# VSS 0.729455f 
C5621 a_19864_35138# VSS 1.75392f 
C5622 a_19120_35138# VSS 1.69667f 
C5623 a_18194_35068# VSS 2.11801f 
C5624 EN_VIN_BSTR_N VSS 9.03857f 
C5625 a_11530_34132# VSS 13.9862f 
C5626 a_n83_35174# VSS 1.72857f 
C5627 EN_VIN_BSTR_P VSS 9.263339f 
C5628 a_n923_35174# VSS 14.088f 
C5629 a_n1532_35090# VSS 2.16074f 
C5630 a_n1386_35608# VSS 1.75773f 
C5631 a_n1838_35608# VSS 0.737725f 
C5632 a_22609_37990# VSS 0.473213f 
C5633 a_22609_38406# VSS 0.588255f 
C5634 CAL_P VSS 11.418599f 
C5635 a_22469_39537# VSS 2.5954f 
C5636 a_22821_38993# VSS 0.55301f 
C5637 a_22545_38993# VSS 0.35571f 
C5638 a_22521_39511# VSS 1.85851f 
C5639 a_22459_39145# VSS 2.29285f 
C5640 a_22521_40055# VSS 1.21928f 
C5641 a_22469_40625# VSS 1.56643f 
C5642 a_22521_40599# VSS 1.85568f 
C5643 CAL_N VSS 8.69238f 
C5644 a_11206_38545# VSS 0.713084f 
C5645 VDAC_P VSS 79.0997f 
C5646 a_8912_37509# VSS 3.72815f 
C5647 VDAC_N VSS 79.6318f 
C5648 a_6886_37412# VSS 3.84457f 
C5649 a_5700_37509# VSS 2.08109f 
C5650 a_5088_37509# VSS 2.72043f 
C5651 a_4338_37500# VSS 2.61369f 
C5652 a_3726_37500# VSS 4.48332f 
C5653 a_n2302_37690# VSS 0.514508f 
C5654 a_n4064_37440# VSS 1.7233f 
C5655 a_n2946_37690# VSS 0.517242f 
C5656 a_n3420_37440# VSS 5.23286f 
C5657 a_n3690_37440# VSS 0.548488f 
C5658 a_n3565_37414# VSS 3.15906f 
C5659 a_n4334_37440# VSS 0.561497f 
C5660 a_n4209_37414# VSS 3.16282f 
C5661 a_8530_39574# VSS 2.76228f 
C5662 a_7754_38470# VSS 3.24598f 
C5663 a_3754_38470# VSS 4.77654f 
C5664 VDAC_Ni VSS 2.86404f 
C5665 a_7754_38636# VSS 0.353706f 
C5666 a_3754_38802# VSS 0.390074f 
C5667 a_7754_38968# VSS 0.330037f 
C5668 a_3754_39134# VSS 0.401983f 
C5669 a_7754_39300# VSS 0.330682f 
C5670 a_3754_39466# VSS 0.401172f 
C5671 a_7754_39632# VSS 0.340942f 
C5672 VDAC_Pi VSS 3.50355f 
C5673 a_7754_39964# VSS 2.62481f 
C5674 a_7754_40130# VSS 2.84104f 
C5675 a_3754_39964# VSS 0.671366f 
C5676 a_2113_38308# VSS 2.64372f 
C5677 a_n2302_37984# VSS 0.483504f 
C5678 a_n4064_37984# VSS 1.65074f 
C5679 a_n2946_37984# VSS 0.485942f 
C5680 a_n3420_37984# VSS 1.75918f 
C5681 a_n3690_38304# VSS 0.517812f 
C5682 a_n3565_38216# VSS 1.48743f 
C5683 a_n4334_38304# VSS 0.529531f 
C5684 a_n4209_38216# VSS 3.03366f 
C5685 a_2684_37794# VSS 0.414596f 
C5686 a_1177_38525# VSS 0.641945f 
C5687 a_n2302_38778# VSS 0.483515f 
C5688 a_n4064_38528# VSS 1.69554f 
C5689 a_n2946_38778# VSS 0.485895f 
C5690 a_n3420_38528# VSS 2.03238f 
C5691 a_n3690_38528# VSS 0.516979f 
C5692 a_n3565_38502# VSS 1.55586f 
C5693 a_n4334_38528# VSS 0.529888f 
C5694 a_n4209_38502# VSS 3.0175f 
C5695 a_2112_39137# VSS 0.414248f 
C5696 comp_n VSS 0.568772f 
C5697 a_1736_39043# VSS 0.897653f 
C5698 a_1239_39043# VSS 0.614001f 
C5699 a_n2302_39072# VSS 0.483504f 
C5700 a_n4064_39072# VSS 1.71745f 
C5701 a_n2946_39072# VSS 0.486447f 
C5702 a_n3420_39072# VSS 2.21624f 
C5703 a_n3690_39392# VSS 0.517965f 
C5704 a_n3565_39304# VSS 1.4403f 
C5705 a_n4334_39392# VSS 0.529516f 
C5706 a_n4209_39304# VSS 3.21429f 
C5707 a_1343_38525# VSS 3.5734f 
C5708 a_1736_39587# VSS 1.10676f 
C5709 a_1239_39587# VSS 0.634559f 
C5710 a_n2302_39866# VSS 0.483537f 
C5711 a_n4064_39616# VSS 2.17764f 
C5712 a_n2946_39866# VSS 0.527929f 
C5713 a_n3420_39616# VSS 2.11206f 
C5714 a_n3690_39616# VSS 0.574329f 
C5715 a_n3565_39590# VSS 2.04547f 
C5716 a_n4334_39616# VSS 0.529903f 
C5717 a_n4209_39590# VSS 3.92629f 
C5718 a_n2302_40160# VSS 0.522244f 
C5719 a_n4064_40160# VSS 3.2951f 
C5720 a_n4334_40480# VSS 0.578721f 
C5721 a_n4315_30879# VSS 4.84874f 
C5722 a_22465_38105# VSS 1.91115f 
C5723 a_22775_42308# VSS 0.602961f 
C5724 a_21613_42308# VSS 0.725408f 
C5725 a_21887_42336# VSS 0.234022f 
C5726 a_21335_42336# VSS 0.259392f 
C5727 a_7174_31319# VSS 5.51134f 
C5728 a_20712_42282# VSS 0.349662f 
C5729 a_20107_42308# VSS 0.344464f 
C5730 a_13258_32519# VSS 6.359931f 
C5731 a_19647_42308# VSS 0.313304f 
C5732 a_19511_42282# VSS 0.751141f 
C5733 a_19332_42282# VSS 0.31505f 
C5734 a_18907_42674# VSS 0.209311f 
C5735 a_18727_42674# VSS 0.233526f 
C5736 a_18057_42282# VSS 0.370712f 
C5737 a_17531_42308# VSS 0.253358f 
C5738 a_17303_42282# VSS 1.19698f 
C5739 a_4958_30871# VSS 5.01268f 
C5740 a_17124_42282# VSS 0.332693f 
C5741 a_15890_42674# VSS 0.180637f 
C5742 a_15959_42545# VSS 0.263128f 
C5743 a_15803_42450# VSS 0.566963f 
C5744 a_15764_42576# VSS 0.298494f 
C5745 a_15486_42560# VSS 0.263746f 
C5746 a_15051_42282# VSS 0.790649f 
C5747 a_14113_42308# VSS 1.42448f 
C5748 a_14456_42282# VSS 0.33927f 
C5749 a_13575_42558# VSS 0.370369f 
C5750 a_13070_42354# VSS 0.222095f 
C5751 a_12563_42308# VSS 0.330976f 
C5752 a_11551_42558# VSS 0.372919f 
C5753 a_5742_30871# VSS 8.193179f 
C5754 a_11323_42473# VSS 0.253445f 
C5755 a_10723_42308# VSS 0.342975f 
C5756 a_10533_42308# VSS 0.310658f 
C5757 a_9803_42558# VSS 0.370474f 
C5758 a_9223_42460# VSS 0.236204f 
C5759 a_8791_42308# VSS 0.301f 
C5760 a_8685_42308# VSS 0.163732f 
C5761 a_8325_42308# VSS 0.316205f 
C5762 a_8515_42308# VSS 0.250762f 
C5763 a_5934_30871# VSS 5.17381f 
C5764 a_7963_42308# VSS 0.256292f 
C5765 a_6123_31319# VSS 5.0238f 
C5766 a_7227_42308# VSS 0.359705f 
C5767 a_6761_42308# VSS 0.447596f 
C5768 a_5932_42308# VSS 5.11915f 
C5769 a_6171_42473# VSS 0.257988f 
C5770 a_5755_42308# VSS 0.314735f 
C5771 a_4921_42308# VSS 0.511258f 
C5772 a_5379_42460# VSS 0.564806f 
C5773 a_5267_42460# VSS 0.204309f 
C5774 a_3823_42558# VSS 0.381485f 
C5775 a_3318_42354# VSS 0.238394f 
C5776 a_2903_42308# VSS 0.340659f 
C5777 a_2713_42308# VSS 0.31991f 
C5778 a_2351_42308# VSS 0.210162f 
C5779 a_2123_42473# VSS 0.21778f 
C5780 a_1755_42282# VSS 3.17706f 
C5781 a_1606_42308# VSS 5.25438f 
C5782 a_961_42354# VSS 0.215753f 
C5783 a_1184_42692# VSS 0.222827f 
C5784 a_1576_42282# VSS 0.327109f 
C5785 a_1067_42314# VSS 0.32917f 
C5786 a_n1630_35242# VSS 10.134f 
C5787 a_564_42282# VSS 0.36802f 
C5788 a_n3674_37592# VSS 3.04613f 
C5789 a_n784_42308# VSS 6.50095f 
C5790 a_196_42282# VSS 0.343186f 
C5791 a_n473_42460# VSS 0.366068f 
C5792 a_n961_42308# VSS 0.328065f 
C5793 a_n1329_42308# VSS 0.30898f 
C5794 COMP_P VSS 11.0245f 
C5795 a_n4318_37592# VSS 1.00428f 
C5796 a_n1736_42282# VSS 0.320711f 
C5797 a_n3674_38216# VSS 1.68571f 
C5798 a_n2104_42282# VSS 0.346472f 
C5799 a_n4318_38216# VSS 0.964502f 
C5800 a_n2472_42282# VSS 0.335792f 
C5801 a_n3674_38680# VSS 0.881032f 
C5802 a_n2840_42282# VSS 0.343361f 
C5803 a_14097_32519# VSS 1.90783f 
C5804 a_22400_42852# VSS 2.02868f 
C5805 a_20256_43172# VSS 0.192089f 
C5806 a_14635_42282# VSS 0.336817f 
C5807 a_13291_42460# VSS 0.197331f 
C5808 a_n2293_42282# VSS 2.62914f 
C5809 a_22959_42860# VSS 0.34332f 
C5810 a_22223_42860# VSS 0.328988f 
C5811 a_22165_42308# VSS 0.354098f 
C5812 a_21671_42860# VSS 0.316857f 
C5813 a_21195_42852# VSS 0.277519f 
C5814 a_21356_42826# VSS 0.304166f 
C5815 a_20922_43172# VSS 0.266814f 
C5816 a_19987_42826# VSS 0.378798f 
C5817 a_19164_43230# VSS 0.264863f 
C5818 a_19339_43156# VSS 0.471496f 
C5819 a_18599_43230# VSS 0.266382f 
C5820 a_18817_42826# VSS 0.182139f 
C5821 a_18249_42858# VSS 0.302863f 
C5822 a_17333_42852# VSS 0.29982f 
C5823 a_18083_42858# VSS 0.578693f 
C5824 a_17701_42308# VSS 0.179963f 
C5825 a_17595_43084# VSS 0.205109f 
C5826 a_16795_42852# VSS 0.362281f 
C5827 a_16414_43172# VSS 0.270304f 
C5828 a_15567_42826# VSS 0.316627f 
C5829 a_5342_30871# VSS 4.18054f 
C5830 a_15279_43071# VSS 0.248252f 
C5831 a_5534_30871# VSS 4.58413f 
C5832 a_14543_43071# VSS 0.246071f 
C5833 a_13460_43230# VSS 0.259861f 
C5834 a_13635_43156# VSS 0.7696f 
C5835 a_12895_43230# VSS 0.250159f 
C5836 a_13113_42826# VSS 0.174096f 
C5837 a_12545_42858# VSS 0.287468f 
C5838 a_12089_42308# VSS 0.283874f 
C5839 a_12379_42858# VSS 0.549229f 
C5840 a_10341_42308# VSS 0.317389f 
C5841 a_10922_42852# VSS 0.176112f 
C5842 a_10991_42826# VSS 0.261283f 
C5843 a_10796_42968# VSS 0.29877f 
C5844 a_10835_43094# VSS 0.59174f 
C5845 a_10518_42984# VSS 0.260322f 
C5846 a_10083_42826# VSS 0.762957f 
C5847 a_8952_43230# VSS 0.261046f 
C5848 a_9127_43156# VSS 0.77314f 
C5849 a_8387_43230# VSS 0.255573f 
C5850 a_8605_42826# VSS 0.181157f 
C5851 a_8037_42858# VSS 0.293593f 
C5852 a_7765_42852# VSS 0.252651f 
C5853 a_7871_42858# VSS 0.503534f 
C5854 a_7227_42852# VSS 0.36607f 
C5855 a_5755_42852# VSS 0.383967f 
C5856 a_5111_42852# VSS 0.354197f 
C5857 a_4520_42826# VSS 0.334784f 
C5858 a_3935_42891# VSS 0.26911f 
C5859 a_3681_42891# VSS 0.301094f 
C5860 a_2905_42968# VSS 0.305424f 
C5861 a_2075_43172# VSS 0.537699f 
C5862 a_1847_42826# VSS 0.670072f 
C5863 a_791_42968# VSS 0.335942f 
C5864 a_685_42968# VSS 0.220885f 
C5865 a_n4318_38680# VSS 1.39087f 
C5866 a_n3674_39304# VSS 1.06639f 
C5867 a_n13_43084# VSS 0.368998f 
C5868 a_n1076_43230# VSS 0.263204f 
C5869 a_n901_43156# VSS 0.76245f 
C5870 a_n1641_43230# VSS 0.256397f 
C5871 a_n1423_42826# VSS 0.1805f 
C5872 a_n1991_42858# VSS 0.295941f 
C5873 a_n1853_43023# VSS 1.30078f 
C5874 a_n2157_42858# VSS 0.556569f 
C5875 a_n2472_42826# VSS 0.301801f 
C5876 a_n2840_42826# VSS 0.327636f 
C5877 a_20749_43396# VSS 0.253248f 
C5878 a_17364_32525# VSS 1.89349f 
C5879 a_22959_43396# VSS 0.345439f 
C5880 a_14209_32519# VSS 2.01016f 
C5881 a_22591_43396# VSS 0.335697f 
C5882 a_13887_32519# VSS 1.94312f 
C5883 a_22223_43396# VSS 0.333609f 
C5884 a_5649_42852# VSS 1.95364f 
C5885 a_13678_32519# VSS 2.06126f 
C5886 a_21855_43396# VSS 0.334538f 
C5887 a_4361_42308# VSS 1.30251f 
C5888 a_13467_32519# VSS 2.22551f 
C5889 a_19095_43396# VSS 0.132304f 
C5890 a_21487_43396# VSS 0.293844f 
C5891 a_743_42282# VSS 1.36822f 
C5892 a_4190_30871# VSS 7.37741f 
C5893 a_21259_43561# VSS 0.217667f 
C5894 a_16823_43084# VSS 1.23251f 
C5895 a_19700_43370# VSS 0.335707f 
C5896 a_19268_43646# VSS 0.242693f 
C5897 a_15743_43084# VSS 1.49489f 
C5898 a_18783_43370# VSS 0.360096f 
C5899 a_18525_43370# VSS 0.361236f 
C5900 a_18429_43548# VSS 0.222219f 
C5901 a_17324_43396# VSS 0.258017f 
C5902 a_17499_43370# VSS 0.762886f 
C5903 a_16759_43396# VSS 0.252915f 
C5904 a_16977_43638# VSS 0.178776f 
C5905 a_16409_43396# VSS 0.290743f 
C5906 a_16547_43609# VSS 0.561468f 
C5907 a_16243_43396# VSS 0.562369f 
C5908 a_16137_43396# VSS 0.635905f 
C5909 a_15781_43660# VSS 0.234761f 
C5910 a_15681_43442# VSS 0.20154f 
C5911 a_12281_43396# VSS 0.691406f 
C5912 a_10341_43396# VSS 0.796012f 
C5913 a_14955_43396# VSS 0.266041f 
C5914 a_15095_43370# VSS 0.436411f 
C5915 a_14205_43396# VSS 0.2933f 
C5916 a_14358_43442# VSS 0.198188f 
C5917 a_14579_43548# VSS 0.293668f 
C5918 a_13667_43396# VSS 0.265557f 
C5919 a_10695_43548# VSS 0.279385f 
C5920 a_9803_43646# VSS 0.371929f 
C5921 a_9145_43396# VSS 0.437647f 
C5922 a_8685_43396# VSS 1.0146f 
C5923 a_3457_43396# VSS 0.379621f 
C5924 a_2813_43396# VSS 0.412407f 
C5925 a_9396_43370# VSS 0.338475f 
C5926 a_8791_43396# VSS 0.235222f 
C5927 a_8147_43396# VSS 0.256103f 
C5928 a_7112_43396# VSS 0.256956f 
C5929 a_7287_43370# VSS 0.754599f 
C5930 a_6547_43396# VSS 0.253718f 
C5931 a_6765_43638# VSS 0.174622f 
C5932 a_6197_43396# VSS 0.290517f 
C5933 a_6293_42852# VSS 0.473619f 
C5934 a_6031_43396# VSS 0.541083f 
C5935 a_648_43396# VSS 0.231254f 
C5936 a_3539_42460# VSS 0.337918f 
C5937 a_3626_43646# VSS 1.9807f 
C5938 a_2982_43646# VSS 3.25953f 
C5939 a_n1557_42282# VSS 0.870257f 
C5940 a_4905_42826# VSS 0.781685f 
C5941 a_3080_42308# VSS 5.07176f 
C5942 a_4699_43561# VSS 0.267684f 
C5943 a_4235_43370# VSS 0.33553f 
C5944 a_4093_43548# VSS 0.320586f 
C5945 a_1756_43548# VSS 0.322408f 
C5946 a_1568_43370# VSS 0.63594f 
C5947 a_1049_43396# VSS 0.216408f 
C5948 a_1209_43370# VSS 0.281234f 
C5949 a_458_43396# VSS 0.252302f 
C5950 a_104_43370# VSS 0.297328f 
C5951 a_n97_42460# VSS 6.9914f 
C5952 a_n447_43370# VSS 0.269574f 
C5953 a_n1352_43396# VSS 0.260107f 
C5954 a_n1177_43370# VSS 0.478516f 
C5955 a_n1917_43396# VSS 0.258245f 
C5956 a_n1699_43638# VSS 0.175452f 
C5957 a_n2267_43396# VSS 0.297246f 
C5958 a_n2129_43609# VSS 1.07965f 
C5959 a_n2433_43396# VSS 0.56533f 
C5960 a_n4318_39304# VSS 0.959585f 
C5961 a_n2840_43370# VSS 0.316787f 
C5962 a_17538_32519# VSS 1.8877f 
C5963 a_20974_43370# VSS 0.458091f 
C5964 a_14401_32519# VSS 2.32323f 
C5965 a_21381_43940# VSS 0.358332f 
C5966 a_19319_43548# VSS 0.229395f 
C5967 a_14021_43940# VSS 0.387813f 
C5968 a_11173_44260# VSS 0.219946f 
C5969 a_10555_44260# VSS 0.346315f 
C5970 a_22959_43948# VSS 0.341565f 
C5971 a_15493_43940# VSS 0.460801f 
C5972 a_22223_43948# VSS 0.31992f 
C5973 a_11341_43940# VSS 0.365183f 
C5974 a_21115_43940# VSS 0.204633f 
C5975 a_20935_43940# VSS 0.222887f 
C5976 a_20623_43914# VSS 0.371294f 
C5977 a_20365_43914# VSS 0.359455f 
C5978 a_20269_44172# VSS 0.225063f 
C5979 a_19862_44208# VSS 0.562087f 
C5980 a_19478_44306# VSS 0.278384f 
C5981 a_15493_43396# VSS 0.277875f 
C5982 a_19328_44172# VSS 0.2031f 
C5983 a_18451_43940# VSS 0.377396f 
C5984 a_18326_43940# VSS 0.276559f 
C5985 a_18079_43940# VSS 0.21121f 
C5986 a_17973_43940# VSS 0.359917f 
C5987 a_17737_43940# VSS 0.386318f 
C5988 a_15682_43940# VSS 1.9643f 
C5989 a_14955_43940# VSS 0.365393f 
C5990 a_13483_43940# VSS 0.376442f 
C5991 a_12429_44172# VSS 0.389129f 
C5992 a_11750_44172# VSS 0.221782f 
C5993 a_10807_43548# VSS 0.451031f 
C5994 a_10949_43914# VSS 0.257331f 
C5995 a_10729_43914# VSS 0.34307f 
C5996 a_10405_44172# VSS 0.142993f 
C5997 a_9672_43914# VSS 0.323006f 
C5998 a_9028_43914# VSS 0.398016f 
C5999 a_8333_44056# VSS 0.331632f 
C6000 a_n2661_42282# VSS 1.51789f 
C6001 a_3499_42826# VSS 0.380221f 
C6002 a_n3674_39768# VSS 0.890487f 
C6003 a_n4318_39768# VSS 1.09976f 
C6004 a_7845_44172# VSS 0.239173f 
C6005 a_7542_44172# VSS 0.283767f 
C6006 a_7281_43914# VSS 0.271121f 
C6007 a_6453_43914# VSS 0.26639f 
C6008 a_5663_43940# VSS 0.488325f 
C6009 a_5495_43940# VSS 0.212229f 
C6010 a_5013_44260# VSS 0.279924f 
C6011 a_5244_44056# VSS 0.216368f 
C6012 a_3905_42865# VSS 0.9893f 
C6013 a_3600_43914# VSS 0.422049f 
C6014 a_2998_44172# VSS 0.503048f 
C6015 a_2889_44172# VSS 0.217034f 
C6016 a_2675_43914# VSS 0.2974f 
C6017 a_895_43940# VSS 0.237723f 
C6018 a_2479_44172# VSS 0.817462f 
C6019 a_2127_44172# VSS 0.517911f 
C6020 a_453_43940# VSS 0.285192f 
C6021 a_1414_42308# VSS 1.07452f 
C6022 a_1467_44172# VSS 0.187431f 
C6023 a_1115_44172# VSS 0.52592f 
C6024 a_644_44056# VSS 0.227493f 
C6025 a_175_44278# VSS 0.226801f 
C6026 a_n984_44318# VSS 0.27358f 
C6027 a_n809_44244# VSS 0.785904f 
C6028 a_n1549_44318# VSS 0.264547f 
C6029 a_n1331_43914# VSS 0.185087f 
C6030 a_n1899_43946# VSS 0.299008f 
C6031 a_n1761_44111# VSS 0.392075f 
C6032 a_n2065_43946# VSS 0.658803f 
C6033 a_n2472_43914# VSS 0.3103f 
C6034 a_n2840_43914# VSS 0.345355f 
C6035 a_19237_31679# VSS 1.48755f 
C6036 a_22959_44484# VSS 0.343897f 
C6037 a_17730_32519# VSS 2.45301f 
C6038 a_22591_44484# VSS 0.315361f 
C6039 a_22485_44484# VSS 0.590119f 
C6040 a_20512_43084# VSS 0.561552f 
C6041 a_22315_44484# VSS 0.238239f 
C6042 a_3422_30871# VSS 9.01786f 
C6043 a_18579_44172# VSS 0.812679f 
C6044 a_19279_43940# VSS 1.69633f 
C6045 a_20766_44850# VSS 0.177656f 
C6046 a_20835_44721# VSS 0.260406f 
C6047 a_20679_44626# VSS 0.58931f 
C6048 a_20640_44752# VSS 0.296084f 
C6049 a_20362_44736# VSS 0.255907f 
C6050 a_20159_44458# VSS 0.483669f 
C6051 a_19615_44636# VSS 0.238459f 
C6052 a_11967_42832# VSS 6.11191f 
C6053 a_17517_44484# VSS 0.244051f 
C6054 a_14673_44172# VSS 0.290001f 
C6055 a_11541_44484# VSS 0.139071f 
C6056 a_15433_44458# VSS 0.301508f 
C6057 a_14815_43914# VSS 0.445698f 
C6058 a_n2293_43922# VSS 3.31971f 
C6059 a_n2661_43922# VSS 1.51991f 
C6060 a_n2661_42834# VSS 1.20196f 
C6061 a_9159_44484# VSS 0.158168f 
C6062 a_10617_44484# VSS 0.119149f 
C6063 a_5708_44484# VSS 0.231649f 
C6064 a_3363_44484# VSS 0.27629f 
C6065 a_556_44484# VSS 0.201935f 
C6066 a_9313_44734# VSS 1.31461f 
C6067 a_5891_43370# VSS 2.82295f 
C6068 a_8375_44464# VSS 0.211867f 
C6069 a_7640_43914# VSS 0.542377f 
C6070 a_6109_44484# VSS 0.648821f 
C6071 a_n23_44458# VSS 0.278255f 
C6072 a_n356_44636# VSS 2.91333f 
C6073 a_18989_43940# VSS 0.423174f 
C6074 a_18374_44850# VSS 0.179731f 
C6075 a_18443_44721# VSS 0.253971f 
C6076 a_18287_44626# VSS 0.507939f 
C6077 a_18248_44752# VSS 0.294917f 
C6078 a_17970_44736# VSS 0.26161f 
C6079 a_17767_44458# VSS 0.474097f 
C6080 a_16979_44734# VSS 0.363013f 
C6081 a_14539_43914# VSS 1.18088f 
C6082 a_16112_44458# VSS 0.326339f 
C6083 a_15004_44636# VSS 0.254778f 
C6084 a_13720_44458# VSS 0.403209f 
C6085 a_13076_44458# VSS 0.38829f 
C6086 a_12883_44458# VSS 0.287544f 
C6087 a_12607_44458# VSS 0.499331f 
C6088 a_8975_43940# VSS 0.652857f 
C6089 a_10057_43914# VSS 0.654189f 
C6090 a_10440_44484# VSS 0.210149f 
C6091 a_10334_44484# VSS 0.210217f 
C6092 a_10157_44484# VSS 0.208916f 
C6093 a_9838_44484# VSS 0.276258f 
C6094 a_5883_43914# VSS 0.792825f 
C6095 a_8701_44490# VSS 0.358059f 
C6096 a_8103_44636# VSS 0.340824f 
C6097 a_6298_44484# VSS 1.93814f 
C6098 a_5518_44484# VSS 0.242995f 
C6099 a_5343_44458# VSS 1.28071f 
C6100 a_4743_44484# VSS 0.327178f 
C6101 a_n699_43396# VSS 1.82142f 
C6102 a_4223_44672# VSS 0.659279f 
C6103 a_2779_44458# VSS 0.532137f 
C6104 a_949_44458# VSS 1.97734f 
C6105 a_742_44458# VSS 1.02263f 
C6106 a_n452_44636# VSS 0.254732f 
C6107 a_n1352_44484# VSS 0.269853f 
C6108 a_n1177_44458# VSS 0.493891f 
C6109 a_n1917_44484# VSS 0.280038f 
C6110 a_n1699_44726# VSS 0.197478f 
C6111 a_n2267_44484# VSS 0.308908f 
C6112 a_n2129_44697# VSS 0.307327f 
C6113 a_n2433_44484# VSS 0.679598f 
C6114 a_n2661_44458# VSS 0.487677f 
C6115 a_n4318_40392# VSS 0.995833f 
C6116 a_n2840_44458# VSS 0.316322f 
C6117 a_19721_31679# VSS 1.61485f 
C6118 a_18114_32519# VSS 3.10957f 
C6119 a_20193_45348# VSS 1.70015f 
C6120 a_11691_44458# VSS 1.78467f 
C6121 a_19113_45348# VSS 0.367248f 
C6122 a_22959_45036# VSS 0.345334f 
C6123 a_22223_45036# VSS 0.354178f 
C6124 a_11827_44484# VSS 1.28091f 
C6125 a_21359_45002# VSS 0.397791f 
C6126 a_21101_45002# VSS 0.35202f 
C6127 a_21005_45260# VSS 0.212992f 
C6128 a_20567_45036# VSS 0.31908f 
C6129 a_18494_42460# VSS 1.15626f 
C6130 a_18184_42460# VSS 0.838573f 
C6131 a_19778_44110# VSS 0.599421f 
C6132 a_18911_45144# VSS 0.307008f 
C6133 a_18587_45118# VSS 0.214925f 
C6134 a_18315_45260# VSS 0.334834f 
C6135 a_17719_45144# VSS 0.331229f 
C6136 a_17613_45144# VSS 0.244364f 
C6137 a_17023_45118# VSS 0.20885f 
C6138 a_16922_45042# VSS 0.818675f 
C6139 a_n2661_43370# VSS 0.820606f 
C6140 a_8560_45348# VSS 0.185033f 
C6141 a_n2293_42834# VSS 1.1151f 
C6142 a_2304_45348# VSS 0.182367f 
C6143 a_1423_45028# VSS 0.980773f 
C6144 a_626_44172# VSS 0.67926f 
C6145 a_375_42282# VSS 0.447027f 
C6146 a_16751_45260# VSS 0.316547f 
C6147 a_1307_43914# VSS 2.30311f 
C6148 a_16019_45002# VSS 0.25377f 
C6149 a_15595_45028# VSS 0.214111f 
C6150 a_15415_45028# VSS 0.221991f 
C6151 a_14797_45144# VSS 0.249222f 
C6152 a_14537_43396# VSS 1.73146f 
C6153 a_14180_45002# VSS 0.327485f 
C6154 a_13777_45326# VSS 0.272936f 
C6155 a_13556_45296# VSS 1.01916f 
C6156 a_9482_43914# VSS 3.42654f 
C6157 a_13348_45260# VSS 0.243533f 
C6158 a_13159_45002# VSS 0.265737f 
C6159 a_13017_45260# VSS 0.362048f 
C6160 a_11963_45334# VSS 0.226884f 
C6161 a_11787_45002# VSS 0.212512f 
C6162 a_10951_45334# VSS 0.228638f 
C6163 a_10775_45002# VSS 0.204487f 
C6164 a_8953_45002# VSS 1.94941f 
C6165 a_8191_45002# VSS 0.325964f 
C6166 a_7705_45326# VSS 0.273009f 
C6167 a_6709_45028# VSS 0.354418f 
C6168 a_7229_43940# VSS 0.786182f 
C6169 a_7276_45260# VSS 0.251523f 
C6170 a_5205_44484# VSS 0.546179f 
C6171 a_6431_45366# VSS 0.233718f 
C6172 a_6171_45002# VSS 0.700605f 
C6173 a_3232_43370# VSS 2.99721f 
C6174 a_5691_45260# VSS 0.370273f 
C6175 a_4927_45028# VSS 0.520892f 
C6176 a_5111_44636# VSS 3.44603f 
C6177 a_5147_45002# VSS 0.803306f 
C6178 a_4558_45348# VSS 0.446148f 
C6179 a_4574_45260# VSS 0.208274f 
C6180 a_3537_45260# VSS 2.45782f 
C6181 a_3429_45260# VSS 0.274034f 
C6182 a_3065_45002# VSS 0.864786f 
C6183 a_2680_45002# VSS 0.321351f 
C6184 a_2382_45260# VSS 1.03422f 
C6185 a_2274_45254# VSS 0.187307f 
C6186 a_1667_45002# VSS 0.345429f 
C6187 a_327_44734# VSS 0.419171f 
C6188 a_413_45260# VSS 4.87522f 
C6189 a_n37_45144# VSS 0.321746f 
C6190 a_n143_45144# VSS 0.209896f 
C6191 a_n467_45028# VSS 0.311181f 
C6192 a_n967_45348# VSS 0.453992f 
C6193 en_comp VSS 7.869411f 
C6194 a_n2956_37592# VSS 2.90302f 
C6195 a_n2810_45028# VSS 1.52635f 
C6196 a_n745_45366# VSS 0.257282f 
C6197 a_n913_45002# VSS 5.04726f 
C6198 a_n1059_45260# VSS 2.30619f 
C6199 a_n2017_45002# VSS 1.09013f 
C6200 a_n2109_45247# VSS 0.252392f 
C6201 a_n2293_45010# VSS 0.614925f 
C6202 a_n2472_45002# VSS 0.298945f 
C6203 a_n2661_45010# VSS 0.839496f 
C6204 a_n2840_45002# VSS 0.340687f 
C6205 a_20447_31679# VSS 1.48786f 
C6206 a_22959_45572# VSS 0.34535f 
C6207 a_19963_31679# VSS 1.43433f 
C6208 a_22591_45572# VSS 0.363695f 
C6209 a_3357_43084# VSS 2.42707f 
C6210 a_19479_31679# VSS 1.66892f 
C6211 a_22223_45572# VSS 0.334964f 
C6212 a_2437_43646# VSS 6.25635f 
C6213 a_21513_45002# VSS 0.669089f 
C6214 a_21188_45572# VSS 0.284872f 
C6215 a_21363_45546# VSS 0.515994f 
C6216 a_20623_45572# VSS 0.256236f 
C6217 a_20841_45814# VSS 0.180037f 
C6218 a_20273_45572# VSS 0.288513f 
C6219 a_20107_45572# VSS 0.541125f 
C6220 a_17668_45572# VSS 0.217142f 
C6221 a_19256_45572# VSS 0.257674f 
C6222 a_19431_45546# VSS 0.487121f 
C6223 a_18691_45572# VSS 0.255356f 
C6224 a_18909_45814# VSS 0.178658f 
C6225 a_18341_45572# VSS 0.291608f 
C6226 a_18479_45785# VSS 1.15946f 
C6227 a_18175_45572# VSS 0.516981f 
C6228 a_16147_45260# VSS 0.506229f 
C6229 a_17478_45572# VSS 0.232341f 
C6230 a_15861_45028# VSS 0.449058f 
C6231 a_8696_44636# VSS 0.917254f 
C6232 a_16680_45572# VSS 0.258674f 
C6233 a_16855_45546# VSS 0.471485f 
C6234 a_16115_45572# VSS 0.253972f 
C6235 a_16333_45814# VSS 0.178165f 
C6236 a_15765_45572# VSS 0.291326f 
C6237 a_15903_45785# VSS 0.4164f 
C6238 a_15599_45572# VSS 0.50233f 
C6239 a_15037_45618# VSS 0.209713f 
C6240 a_11136_45572# VSS 0.17156f 
C6241 a_9159_45572# VSS 0.151638f 
C6242 a_8192_45572# VSS 0.17002f 
C6243 a_10907_45822# VSS 0.547001f 
C6244 a_15143_45578# VSS 0.315994f 
C6245 a_14495_45572# VSS 0.325874f 
C6246 a_13249_42308# VSS 1.08648f 
C6247 a_13904_45546# VSS 0.327907f 
C6248 a_13527_45546# VSS 0.245514f 
C6249 a_13163_45724# VSS 0.180841f 
C6250 a_12791_45546# VSS 0.237787f 
C6251 a_11823_42460# VSS 2.45644f 
C6252 a_12427_45724# VSS 0.190531f 
C6253 a_11962_45724# VSS 0.218739f 
C6254 a_11652_45724# VSS 0.258015f 
C6255 a_11525_45546# VSS 0.346102f 
C6256 a_11322_45546# VSS 0.62914f 
C6257 a_10490_45724# VSS 0.972668f 
C6258 a_8746_45002# VSS 0.547616f 
C6259 a_10193_42453# VSS 3.59848f 
C6260 a_10180_45724# VSS 0.281135f 
C6261 a_10053_45546# VSS 0.373668f 
C6262 a_9049_44484# VSS 0.249658f 
C6263 a_7499_43078# VSS 3.22587f 
C6264 a_8568_45546# VSS 0.317032f 
C6265 a_8162_45546# VSS 0.376225f 
C6266 a_4880_45572# VSS 0.182839f 
C6267 a_3775_45552# VSS 0.209244f 
C6268 a_7227_45028# VSS 0.439395f 
C6269 a_6598_45938# VSS 0.185967f 
C6270 a_6667_45809# VSS 0.264656f 
C6271 a_6511_45714# VSS 0.647716f 
C6272 a_6472_45840# VSS 0.310105f 
C6273 a_6194_45824# VSS 0.2717f 
C6274 a_5907_45546# VSS 0.592148f 
C6275 a_5263_45724# VSS 0.250928f 
C6276 a_4099_45572# VSS 0.33915f 
C6277 a_2711_45572# VSS 1.77517f 
C6278 a_2277_45546# VSS 0.303704f 
C6279 a_1609_45822# VSS 0.5528f 
C6280 a_n443_42852# VSS 4.64762f 
C6281 a_n23_45546# VSS 0.281189f 
C6282 a_n356_45724# VSS 0.32306f 
C6283 a_3503_45724# VSS 0.322319f 
C6284 a_3316_45546# VSS 0.336134f 
C6285 a_3218_45724# VSS 0.379893f 
C6286 a_2957_45546# VSS 0.276358f 
C6287 a_1848_45724# VSS 0.245258f 
C6288 a_997_45618# VSS 0.248122f 
C6289 a_n755_45592# VSS 5.8889f 
C6290 a_n357_42282# VSS 2.46134f 
C6291 a_310_45028# VSS 0.207165f 
C6292 a_n1099_45572# VSS 0.339525f 
C6293 a_380_45546# VSS 0.337145f 
C6294 a_n452_45724# VSS 0.253614f 
C6295 a_n863_45724# VSS 3.49288f 
C6296 a_n1079_45724# VSS 0.289271f 
C6297 a_n2293_45546# VSS 0.879703f 
C6298 a_n2956_38216# VSS 1.49846f 
C6299 a_n2472_45546# VSS 0.340801f 
C6300 a_n2661_45546# VSS 1.58481f 
C6301 a_n2810_45572# VSS 1.43198f 
C6302 a_n2840_45546# VSS 0.344757f 
C6303 a_20692_30879# VSS 1.59585f 
C6304 a_20205_31679# VSS 1.45349f 
C6305 a_16375_45002# VSS 1.44161f 
C6306 a_13259_45724# VSS 4.49011f 
C6307 a_12638_46436# VSS 0.162178f 
C6308 a_12379_46436# VSS 0.275423f 
C6309 a_10586_45546# VSS 0.542658f 
C6310 a_8049_45260# VSS 0.741927f 
C6311 a_8034_45724# VSS 0.299594f 
C6312 a_5066_45546# VSS 0.436834f 
C6313 a_n1925_42282# VSS 1.34109f 
C6314 a_526_44458# VSS 6.44493f 
C6315 a_n2956_38680# VSS 1.34225f 
C6316 a_n2956_39304# VSS 1.60721f 
C6317 a_22959_46124# VSS 0.345245f 
C6318 a_10809_44734# VSS 1.05002f 
C6319 a_22223_46124# VSS 0.354467f 
C6320 a_6945_45028# VSS 0.978274f 
C6321 a_21137_46414# VSS 0.340736f 
C6322 a_20708_46348# VSS 0.268156f 
C6323 a_19900_46494# VSS 0.26164f 
C6324 a_20075_46420# VSS 0.475201f 
C6325 a_19335_46494# VSS 0.260378f 
C6326 a_19553_46090# VSS 0.179968f 
C6327 a_18985_46122# VSS 0.297132f 
C6328 a_18819_46122# VSS 0.545109f 
C6329 a_17957_46116# VSS 0.309446f 
C6330 a_18189_46348# VSS 0.296366f 
C6331 a_17715_44484# VSS 0.55862f 
C6332 a_17583_46090# VSS 0.307562f 
C6333 a_15682_46116# VSS 1.96743f 
C6334 a_2324_44458# VSS 6.12227f 
C6335 a_14840_46494# VSS 0.263367f 
C6336 a_15015_46420# VSS 0.472948f 
C6337 a_14275_46494# VSS 0.258968f 
C6338 a_14493_46090# VSS 0.176122f 
C6339 a_13925_46122# VSS 0.294602f 
C6340 a_13759_46122# VSS 0.518292f 
C6341 a_13351_46090# VSS 0.304427f 
C6342 a_12594_46348# VSS 0.284494f 
C6343 a_12005_46116# VSS 0.381711f 
C6344 a_10903_43370# VSS 2.66576f 
C6345 a_11387_46155# VSS 0.260117f 
C6346 a_11133_46155# VSS 0.299642f 
C6347 a_11189_46129# VSS 0.32558f 
C6348 a_9290_44172# VSS 4.78398f 
C6349 a_10355_46116# VSS 0.290668f 
C6350 a_9823_46155# VSS 0.261206f 
C6351 a_9569_46155# VSS 0.304755f 
C6352 a_9625_46129# VSS 0.369694f 
C6353 a_8953_45546# VSS 1.00397f 
C6354 a_5937_45572# VSS 1.8333f 
C6355 a_8199_44636# VSS 2.29742f 
C6356 a_8349_46414# VSS 0.273442f 
C6357 a_8016_46348# VSS 0.539696f 
C6358 a_7920_46348# VSS 0.269852f 
C6359 a_6419_46155# VSS 0.273686f 
C6360 a_6165_46155# VSS 0.303989f 
C6361 a_5497_46414# VSS 0.304684f 
C6362 a_5204_45822# VSS 0.338817f 
C6363 a_5164_46348# VSS 0.419282f 
C6364 a_5068_46348# VSS 0.25855f 
C6365 a_4704_46090# VSS 0.296767f 
C6366 a_4419_46090# VSS 0.357571f 
C6367 a_4185_45028# VSS 2.50501f 
C6368 a_3699_46348# VSS 0.226584f 
C6369 a_3483_46348# VSS 4.80498f 
C6370 a_3147_46376# VSS 0.52775f 
C6371 a_2804_46116# VSS 0.222855f 
C6372 a_2698_46116# VSS 0.215567f 
C6373 a_2521_46116# VSS 0.220999f 
C6374 a_167_45260# VSS 1.32487f 
C6375 a_2202_46116# VSS 0.273578f 
C6376 a_1823_45246# VSS 2.36307f 
C6377 a_1138_42852# VSS 0.456566f 
C6378 a_1176_45822# VSS 0.278365f 
C6379 a_1208_46090# VSS 0.348206f 
C6380 a_805_46414# VSS 0.27506f 
C6381 a_472_46348# VSS 0.32751f 
C6382 a_376_46348# VSS 0.285607f 
C6383 a_n1076_46494# VSS 0.262147f 
C6384 a_n901_46420# VSS 0.762523f 
C6385 a_n1641_46494# VSS 0.256945f 
C6386 a_n1423_46090# VSS 0.176189f 
C6387 a_n1991_46122# VSS 0.305274f 
C6388 a_n1853_46287# VSS 0.341802f 
C6389 a_n2157_46122# VSS 0.525314f 
C6390 a_n2293_46098# VSS 0.690447f 
C6391 a_n2472_46090# VSS 0.290925f 
C6392 a_n2840_46090# VSS 0.340313f 
C6393 a_21076_30879# VSS 2.00065f 
C6394 a_22959_46660# VSS 0.338967f 
C6395 a_12741_44636# VSS 0.979225f 
C6396 a_20820_30879# VSS 1.64286f 
C6397 a_22591_46660# VSS 0.292786f 
C6398 a_11415_45002# VSS 1.63684f 
C6399 a_20202_43084# VSS 1.05073f 
C6400 a_22365_46825# VSS 0.208388f 
C6401 a_18280_46660# VSS 0.29316f 
C6402 a_17639_46660# VSS 0.308795f 
C6403 a_22000_46634# VSS 0.295895f 
C6404 a_21188_46660# VSS 0.261124f 
C6405 a_21363_46634# VSS 0.488515f 
C6406 a_20623_46660# VSS 0.258464f 
C6407 a_20841_46902# VSS 0.180869f 
C6408 a_20273_46660# VSS 0.309206f 
C6409 a_20411_46873# VSS 0.393328f 
C6410 a_20107_46660# VSS 0.575208f 
C6411 a_19123_46287# VSS 0.477642f 
C6412 a_18285_46348# VSS 0.577053f 
C6413 a_765_45546# VSS 0.902406f 
C6414 a_17339_46660# VSS 0.927636f 
C6415 a_16721_46634# VSS 0.305539f 
C6416 a_16388_46812# VSS 1.42609f 
C6417 a_13059_46348# VSS 2.36107f 
C6418 a_14513_46634# VSS 0.29862f 
C6419 a_14180_46812# VSS 0.368158f 
C6420 a_14035_46660# VSS 0.322858f 
C6421 a_13885_46660# VSS 0.297377f 
C6422 a_19692_46634# VSS 1.97188f 
C6423 a_19466_46812# VSS 0.675335f 
C6424 a_19333_46634# VSS 0.289568f 
C6425 a_15227_44166# VSS 2.80559f 
C6426 a_18834_46812# VSS 0.198054f 
C6427 a_17609_46634# VSS 0.205547f 
C6428 a_16292_46812# VSS 0.271203f 
C6429 a_15559_46634# VSS 0.394779f 
C6430 a_15368_46634# VSS 0.278142f 
C6431 a_14976_45028# VSS 0.479565f 
C6432 a_3090_45724# VSS 2.6372f 
C6433 a_15009_46634# VSS 0.270859f 
C6434 a_14084_46812# VSS 0.251005f 
C6435 a_13607_46688# VSS 0.218935f 
C6436 a_12816_46660# VSS 0.260317f 
C6437 a_12991_46634# VSS 0.475827f 
C6438 a_12251_46660# VSS 0.270927f 
C6439 a_12469_46902# VSS 0.193369f 
C6440 a_11901_46660# VSS 0.303844f 
C6441 a_11813_46116# VSS 0.563718f 
C6442 a_11735_46660# VSS 0.520568f 
C6443 a_8270_45546# VSS 0.779033f 
C6444 a_6969_46634# VSS 0.289597f 
C6445 a_6755_46942# VSS 3.33348f 
C6446 a_10249_46116# VSS 0.414443f 
C6447 a_10554_47026# VSS 0.191251f 
C6448 a_10623_46897# VSS 0.283572f 
C6449 a_10467_46802# VSS 0.523954f 
C6450 a_10428_46928# VSS 0.314538f 
C6451 a_10150_46912# VSS 0.276624f 
C6452 a_9863_46634# VSS 0.607398f 
C6453 a_8492_46660# VSS 0.283316f 
C6454 a_8667_46634# VSS 0.596387f 
C6455 a_7927_46660# VSS 0.269867f 
C6456 a_8145_46902# VSS 0.179735f 
C6457 a_7577_46660# VSS 0.314978f 
C6458 a_7715_46873# VSS 0.546182f 
C6459 a_7411_46660# VSS 0.532412f 
C6460 a_5257_43370# VSS 1.42323f 
C6461 a_6540_46812# VSS 0.248814f 
C6462 a_5732_46660# VSS 0.260482f 
C6463 a_5907_46634# VSS 0.473347f 
C6464 a_5167_46660# VSS 0.263586f 
C6465 a_5385_46902# VSS 0.17737f 
C6466 a_4817_46660# VSS 0.296797f 
C6467 a_4955_46873# VSS 0.365781f 
C6468 a_4651_46660# VSS 0.548065f 
C6469 a_4646_46812# VSS 2.12519f 
C6470 a_3877_44458# VSS 2.8543f 
C6471 a_3524_46660# VSS 0.267612f 
C6472 a_3699_46634# VSS 0.499647f 
C6473 a_2959_46660# VSS 0.261026f 
C6474 a_3177_46902# VSS 0.184239f 
C6475 a_2609_46660# VSS 0.302878f 
C6476 a_2443_46660# VSS 0.657702f 
C6477 a_n2661_46098# VSS 2.05975f 
C6478 a_1799_45572# VSS 0.30194f 
C6479 a_1983_46706# VSS 0.205951f 
C6480 a_2107_46812# VSS 1.13475f 
C6481 a_948_46660# VSS 0.263413f 
C6482 a_1123_46634# VSS 0.776627f 
C6483 a_383_46660# VSS 0.269735f 
C6484 a_601_46902# VSS 0.192316f 
C6485 a_33_46660# VSS 0.309712f 
C6486 a_171_46873# VSS 0.579977f 
C6487 a_n133_46660# VSS 0.576523f 
C6488 a_n2438_43548# VSS 2.99787f 
C6489 a_n743_46660# VSS 3.29885f 
C6490 a_n1021_46688# VSS 0.271211f 
C6491 a_n1925_46634# VSS 1.33202f 
C6492 a_n2312_38680# VSS 2.0221f 
C6493 a_n2104_46634# VSS 0.340006f 
C6494 a_n2293_46634# VSS 1.52366f 
C6495 a_n2442_46660# VSS 1.32617f 
C6496 a_n2472_46634# VSS 0.323981f 
C6497 a_n2661_46634# VSS 0.742038f 
C6498 a_n2956_39768# VSS 1.30197f 
C6499 a_n2840_46634# VSS 0.328049f 
C6500 a_22612_30879# VSS 3.18235f 
C6501 a_21588_30879# VSS 2.65298f 
C6502 a_20916_46384# VSS 0.827544f 
C6503 a_20843_47204# VSS 0.121976f 
C6504 a_19594_46812# VSS 0.277274f 
C6505 a_19321_45002# VSS 1.15234f 
C6506 a_13747_46662# VSS 2.11905f 
C6507 a_13661_43548# VSS 2.82749f 
C6508 a_5807_45002# VSS 2.5828f 
C6509 a_768_44030# VSS 3.03052f 
C6510 a_12549_44172# VSS 2.68201f 
C6511 a_12891_46348# VSS 1.22195f 
C6512 a_11309_47204# VSS 0.423399f 
C6513 a_9804_47204# VSS 0.528639f 
C6514 a_8128_46384# VSS 0.573494f 
C6515 a_n881_46662# VSS 4.56296f 
C6516 a_n1613_43370# VSS 4.90074f 
C6517 a_2747_46873# VSS 0.287894f 
C6518 a_n2312_39304# VSS 1.49307f 
C6519 a_n2312_40392# VSS 2.25565f 
C6520 a_22959_47212# VSS 0.322938f 
C6521 a_11453_44696# VSS 0.689179f 
C6522 SMPL_ON_N VSS 2.60102f 
C6523 a_22731_47423# VSS 0.227778f 
C6524 a_22223_47212# VSS 0.332189f 
C6525 a_12465_44636# VSS 5.61685f 
C6526 a_21811_47423# VSS 0.23358f 
C6527 a_4883_46098# VSS 1.54736f 
C6528 a_21496_47436# VSS 0.249536f 
C6529 a_13507_46334# VSS 4.83849f 
C6530 a_21177_47436# VSS 0.223524f 
C6531 a_20990_47178# VSS 0.224581f 
C6532 a_20894_47436# VSS 0.233111f 
C6533 a_19787_47423# VSS 0.258015f 
C6534 a_19386_47436# VSS 0.209882f 
C6535 a_18597_46090# VSS 2.82344f 
C6536 a_18780_47178# VSS 0.319719f 
C6537 a_18479_47436# VSS 1.19826f 
C6538 a_18143_47464# VSS 0.579061f 
C6539 a_10227_46804# VSS 8.12328f 
C6540 a_17591_47464# VSS 0.576556f 
C6541 a_16588_47582# VSS 0.263715f 
C6542 a_16763_47508# VSS 0.587861f 
C6543 a_16023_47582# VSS 0.264352f 
C6544 a_16327_47482# VSS 5.17799f 
C6545 a_16241_47178# VSS 0.18232f 
C6546 a_15673_47210# VSS 0.315684f 
C6547 a_15811_47375# VSS 0.349499f 
C6548 a_15507_47210# VSS 0.556554f 
C6549 a_11599_46634# VSS 2.84967f 
C6550 a_14955_47212# VSS 0.358339f 
C6551 a_14311_47204# VSS 0.248858f 
C6552 a_13487_47204# VSS 0.643275f 
C6553 a_12861_44030# VSS 3.64545f 
C6554 a_13717_47436# VSS 1.02478f 
C6555 a_n1435_47204# VSS 9.72476f 
C6556 a_13381_47204# VSS 0.225132f 
C6557 a_11459_47204# VSS 0.553679f 
C6558 a_9313_45822# VSS 1.04727f 
C6559 a_11031_47542# VSS 0.247302f 
C6560 a_9863_47436# VSS 0.265619f 
C6561 a_9067_47204# VSS 0.606182f 
C6562 a_6575_47204# VSS 0.798434f 
C6563 a_7903_47542# VSS 0.258657f 
C6564 a_7227_47204# VSS 0.610401f 
C6565 a_6851_47204# VSS 0.346433f 
C6566 a_6491_46660# VSS 0.343406f 
C6567 a_6545_47178# VSS 0.597936f 
C6568 a_6151_47436# VSS 2.12954f 
C6569 a_5815_47464# VSS 0.594449f 
C6570 a_5129_47502# VSS 0.361487f 
C6571 a_4915_47217# VSS 2.79467f 
C6572 a_n443_46116# VSS 4.167f 
C6573 a_4791_45118# VSS 2.65418f 
C6574 a_4700_47436# VSS 0.271201f 
C6575 a_4007_47204# VSS 0.628996f 
C6576 a_3815_47204# VSS 0.440491f 
C6577 a_3785_47178# VSS 0.541893f 
C6578 a_3381_47502# VSS 0.320926f 
C6579 a_n1151_42308# VSS 3.78206f 
C6580 a_3160_47472# VSS 0.607125f 
C6581 a_2905_45572# VSS 0.47073f 
C6582 a_2952_47436# VSS 0.275026f 
C6583 a_2553_47502# VSS 0.294118f 
C6584 a_2063_45854# VSS 1.92678f 
C6585 a_584_46384# VSS 2.10508f 
C6586 a_2124_47436# VSS 0.276508f 
C6587 a_1431_47204# VSS 0.595895f 
C6588 a_1239_47204# VSS 0.33333f 
C6589 a_1209_47178# VSS 0.474725f 
C6590 a_327_47204# VSS 0.581187f 
C6591 a_n785_47204# VSS 0.361759f 
C6592 a_n23_47502# VSS 0.278861f 
C6593 a_n237_47217# VSS 3.05697f 
C6594 a_n746_45260# VSS 0.993718f 
C6595 a_n971_45724# VSS 4.81311f 
C6596 a_n452_47436# VSS 0.28781f 
C6597 a_n815_47178# VSS 0.513835f 
C6598 a_n1605_47204# VSS 0.250546f 
C6599 SMPL_ON_P VSS 4.94844f 
C6600 a_n1741_47186# VSS 1.81488f 
C6601 a_n1920_47178# VSS 0.310881f 
C6602 a_n2109_47186# VSS 0.936844f 
C6603 a_n2288_47178# VSS 0.346995f 
C6604 a_n2497_47436# VSS 2.31207f 
C6605 a_n2833_47464# VSS 0.602779f 
C6606 w_11334_34010# VSS 51.3801f 
C6607 w_1575_34946# VSS 51.6622f 
.ends
