magic
tech sky130A
magscale 1 2
timestamp 1717107273
<< nwell >>
rect 9837 1950 10810 2516
rect 9729 862 10833 1428
<< locali >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2830 10170 2870
rect 3700 2810 10170 2830
rect 3700 2770 3800 2810
rect 3700 -1770 3710 2770
rect 3780 -1770 3800 2770
rect 10330 -830 10360 -770
rect 3700 -1830 3800 -1770
rect 3700 -1840 10140 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1890 10140 -1840
rect 3700 -1900 10140 -1890
<< viali >>
rect 3830 2830 10100 2870
rect 3710 -1770 3780 2770
rect 10130 -540 10170 2740
rect 10428 2514 10494 2562
rect 10579 2512 10645 2562
rect 10748 2512 10815 2566
rect 10348 2410 10398 2470
rect 10668 2350 10718 2410
rect 10348 2077 10398 2127
rect 10430 1904 10491 1953
rect 10579 1904 10646 1954
rect 10748 1900 10815 1954
rect 10587 1789 10648 1838
rect 10348 1520 10408 1580
rect 10697 1570 10731 1604
rect 10428 1426 10494 1474
rect 10575 1424 10638 1490
rect 10688 1430 10748 1490
rect 10864 1430 10924 1500
rect 10428 961 10493 1009
rect 10702 977 10767 1025
rect 10346 816 10411 864
rect 10622 816 10687 864
rect 10270 -830 10330 -770
rect 3820 -1890 10100 -1840
<< metal1 >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2830 10170 2870
rect 3700 2810 10170 2830
rect 10282 2810 11720 2900
rect 3700 2770 3800 2810
rect 3700 -1770 3710 2770
rect 3780 1840 3800 2770
rect 10130 2752 10170 2810
rect 6880 2740 6890 2750
rect 3900 2690 6890 2740
rect 6950 2740 6960 2750
rect 10124 2740 10176 2752
rect 6950 2690 10020 2740
rect 10124 1840 10130 2740
rect 3780 1500 10130 1840
rect 3780 -600 3800 1500
rect 6880 610 6890 620
rect 3890 560 6890 610
rect 6950 610 6960 620
rect 6950 560 10010 610
rect 6880 410 6890 420
rect 3890 360 6890 410
rect 6950 410 6960 420
rect 6950 360 10010 410
rect 9730 70 9740 130
rect 9800 70 9810 130
rect 9750 -460 9790 70
rect 10124 -70 10130 1500
rect 10170 2280 10176 2740
rect 10738 2572 10748 2580
rect 10578 2568 10588 2570
rect 10416 2562 10506 2568
rect 10416 2514 10428 2562
rect 10494 2514 10506 2562
rect 10416 2508 10506 2514
rect 10567 2562 10588 2568
rect 10567 2512 10579 2562
rect 10567 2510 10588 2512
rect 10648 2510 10658 2570
rect 10736 2510 10748 2572
rect 10818 2510 10828 2580
rect 11020 2520 11030 2580
rect 11090 2520 11100 2580
rect 10342 2470 10404 2482
rect 10318 2410 10328 2470
rect 10398 2410 10404 2470
rect 10342 2398 10404 2410
rect 10446 2392 10478 2508
rect 10567 2506 10657 2510
rect 10736 2506 10827 2510
rect 10662 2410 10724 2422
rect 10662 2400 10668 2410
rect 10718 2400 10724 2410
rect 10648 2392 10658 2400
rect 10446 2347 10658 2392
rect 10648 2340 10658 2347
rect 10718 2340 10728 2400
rect 10662 2338 10724 2340
rect 10170 2190 10338 2280
rect 10170 1190 10176 2190
rect 10338 2133 10348 2137
rect 10336 2077 10348 2133
rect 10408 2077 10418 2137
rect 10336 2071 10410 2077
rect 11050 1960 11080 2520
rect 11120 2430 11130 2490
rect 11190 2430 11200 2490
rect 10418 1953 10503 1959
rect 10418 1904 10430 1953
rect 10491 1904 10503 1953
rect 10418 1898 10503 1904
rect 10567 1900 10578 1960
rect 10638 1954 10658 1960
rect 10646 1904 10658 1954
rect 10638 1900 10658 1904
rect 10567 1898 10658 1900
rect 10458 1830 10488 1898
rect 10736 1894 10748 1960
rect 10738 1890 10748 1894
rect 10818 1890 10828 1960
rect 11020 1900 11030 1960
rect 11090 1900 11100 1960
rect 10578 1844 10588 1850
rect 10575 1838 10588 1844
rect 10648 1844 10658 1850
rect 10575 1830 10587 1838
rect 10458 1800 10587 1830
rect 10575 1789 10587 1800
rect 10648 1789 10660 1844
rect 10940 1790 10950 1850
rect 11010 1790 11020 1850
rect 10575 1783 10660 1789
rect 10818 1650 10828 1720
rect 10898 1650 10908 1720
rect 10665 1604 10747 1611
rect 10665 1600 10697 1604
rect 10731 1600 10747 1604
rect 10665 1590 10688 1600
rect 10336 1580 10420 1586
rect 10336 1520 10348 1580
rect 10408 1520 10420 1580
rect 10336 1514 10420 1520
rect 10468 1560 10688 1590
rect 10468 1480 10498 1560
rect 10678 1540 10688 1560
rect 10748 1540 10758 1600
rect 10569 1500 10644 1502
rect 10858 1500 10930 1512
rect 10558 1490 10648 1500
rect 10416 1474 10506 1480
rect 10416 1426 10428 1474
rect 10494 1426 10506 1474
rect 10416 1420 10506 1426
rect 10558 1424 10575 1490
rect 10638 1424 10648 1490
rect 10676 1490 10760 1496
rect 10858 1490 10864 1500
rect 10676 1430 10688 1490
rect 10748 1430 10760 1490
rect 10856 1430 10864 1490
rect 10924 1430 10930 1500
rect 10676 1424 10760 1430
rect 10558 1406 10648 1424
rect 10558 1340 10568 1406
rect 10631 1340 10648 1406
rect 10708 1290 10738 1424
rect 10858 1418 10930 1430
rect 10878 1417 10928 1418
rect 10878 1300 10918 1417
rect 10608 1230 10618 1290
rect 10678 1240 10738 1290
rect 10850 1240 10860 1300
rect 10920 1240 10930 1300
rect 10678 1230 10688 1240
rect 10170 1100 10328 1190
rect 10170 150 10176 1100
rect 10690 1030 10779 1031
rect 10418 1015 10428 1020
rect 10416 960 10428 1015
rect 10488 1015 10498 1020
rect 10488 1009 10505 1015
rect 10493 961 10505 1009
rect 10688 970 10698 1030
rect 10768 971 10779 1030
rect 10768 970 10778 971
rect 10488 960 10505 961
rect 10416 955 10505 960
rect 10334 864 10423 870
rect 10334 860 10346 864
rect 10328 816 10346 860
rect 10411 816 10423 864
rect 10328 810 10423 816
rect 10608 810 10618 870
rect 10678 864 10699 870
rect 10687 816 10699 864
rect 10678 810 10699 816
rect 10328 740 10418 810
rect 10328 680 10338 740
rect 10398 690 10418 740
rect 10398 680 10408 690
rect 10788 630 10808 649
rect 10748 560 10758 630
rect 10828 560 10838 630
rect 10590 380 10600 440
rect 10660 380 10670 440
rect 10390 180 10400 250
rect 10470 180 10480 250
rect 10610 190 10640 380
rect 10170 60 10280 150
rect 10348 132 10408 142
rect 10456 132 10516 142
rect 10690 80 10800 110
rect 10348 62 10364 72
rect 10456 62 10516 72
rect 10170 -70 10176 60
rect 10290 -40 10300 20
rect 10360 -40 10370 20
rect 10110 -130 10120 -70
rect 10180 -130 10190 -70
rect 9730 -520 9740 -460
rect 9800 -520 9810 -460
rect 10124 -540 10130 -130
rect 10170 -270 10176 -130
rect 10310 -220 10360 -40
rect 10500 -170 10560 20
rect 10770 -70 10800 80
rect 10840 70 10850 130
rect 10910 70 10920 130
rect 10750 -130 10760 -70
rect 10820 -130 10830 -70
rect 10490 -230 10500 -170
rect 10560 -230 10570 -170
rect 10170 -360 10280 -270
rect 10348 -280 10408 -270
rect 10456 -280 10516 -270
rect 10770 -300 10800 -130
rect 10680 -330 10800 -300
rect 10348 -350 10364 -340
rect 10456 -350 10516 -340
rect 10170 -440 10176 -360
rect 10170 -540 10180 -440
rect 10390 -460 10400 -390
rect 10470 -460 10480 -390
rect 10124 -600 10180 -540
rect 10610 -580 10640 -410
rect 3780 -940 10180 -600
rect 10580 -640 10590 -580
rect 10650 -640 10660 -580
rect 10260 -670 10350 -660
rect 10260 -730 10280 -670
rect 10340 -730 10350 -670
rect 10750 -730 10760 -670
rect 10820 -730 10830 -670
rect 10260 -764 10350 -730
rect 10258 -770 10350 -764
rect 10258 -830 10270 -770
rect 10330 -830 10350 -770
rect 10600 -830 10610 -770
rect 10670 -830 10680 -770
rect 10258 -836 10350 -830
rect 10260 -840 10350 -836
rect 10410 -930 10420 -870
rect 10480 -930 10490 -870
rect 10620 -930 10650 -830
rect 3780 -1770 3800 -940
rect 10359 -986 10419 -976
rect 10467 -986 10527 -976
rect 10760 -1000 10800 -730
rect 10680 -1030 10800 -1000
rect 10359 -1056 10375 -1046
rect 10467 -1056 10527 -1046
rect 10510 -1180 10570 -1090
rect 10500 -1240 10510 -1180
rect 10570 -1240 10580 -1180
rect 10510 -1340 10570 -1240
rect 10359 -1386 10419 -1376
rect 10467 -1386 10527 -1376
rect 10760 -1400 10800 -1030
rect 10860 -990 10890 70
rect 10960 -160 10990 1790
rect 11050 870 11080 1900
rect 11030 810 11040 870
rect 11100 810 11110 870
rect 11040 520 11100 530
rect 11040 450 11100 460
rect 11050 250 11080 450
rect 11030 190 11040 250
rect 11100 190 11110 250
rect 10920 -220 10930 -160
rect 10990 -220 11000 -160
rect 10920 -340 10930 -280
rect 10990 -340 11000 -280
rect 10860 -1050 10870 -990
rect 10930 -1050 10940 -990
rect 10970 -1380 11000 -340
rect 11050 -400 11080 190
rect 11030 -460 11040 -400
rect 11100 -460 11110 -400
rect 11140 -580 11170 2430
rect 11210 2340 11220 2400
rect 11280 2340 11290 2400
rect 11220 430 11250 2340
rect 11290 2087 11300 2147
rect 11360 2087 11370 2147
rect 11310 740 11340 2087
rect 11650 1720 11720 2810
rect 11640 1650 11650 1720
rect 11720 1650 11730 1720
rect 11470 1540 11480 1600
rect 11540 1540 11550 1600
rect 11380 1370 11440 1380
rect 11380 1300 11440 1310
rect 11290 680 11300 740
rect 11360 680 11370 740
rect 11200 370 11210 430
rect 11270 370 11280 430
rect 11100 -640 11110 -580
rect 11170 -640 11180 -580
rect 11030 -910 11040 -850
rect 11100 -910 11110 -850
rect 10680 -1430 10800 -1400
rect 10940 -1440 10950 -1380
rect 11010 -1440 11020 -1380
rect 10359 -1456 10375 -1446
rect 10467 -1456 10527 -1446
rect 11050 -1490 11080 -910
rect 10400 -1560 10410 -1500
rect 10470 -1560 10480 -1500
rect 10620 -1630 10650 -1500
rect 11030 -1550 11040 -1490
rect 11100 -1550 11110 -1490
rect 11140 -1630 11170 -640
rect 11220 -760 11250 370
rect 11200 -820 11210 -760
rect 11270 -820 11280 -760
rect 11310 -1190 11340 680
rect 11400 40 11430 1300
rect 11490 520 11520 1540
rect 11560 1490 11620 1500
rect 11560 1420 11620 1430
rect 11460 460 11470 520
rect 11530 460 11540 520
rect 11570 140 11600 1420
rect 11650 630 11720 1650
rect 11640 560 11650 630
rect 11720 560 11730 630
rect 11550 130 11600 140
rect 11520 70 11530 130
rect 11590 70 11600 130
rect 11380 30 11440 40
rect 11380 -40 11440 -30
rect 11570 -860 11600 70
rect 11650 -670 11720 560
rect 11710 -730 11720 -670
rect 11650 -780 11720 -730
rect 11530 -920 11540 -860
rect 11600 -920 11610 -860
rect 11290 -1250 11300 -1190
rect 11360 -1250 11370 -1190
rect 10590 -1690 10600 -1630
rect 10660 -1690 10670 -1630
rect 11090 -1690 11100 -1630
rect 11160 -1690 11170 -1630
rect 3700 -1830 3800 -1770
rect 3890 -1780 6890 -1720
rect 6950 -1780 10030 -1720
rect 3700 -1840 10140 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1890 10140 -1840
rect 3700 -1900 10140 -1890
<< via1 >>
rect 6890 2690 6950 2750
rect 6890 560 6950 620
rect 6890 360 6950 420
rect 9740 70 9800 130
rect 10588 2562 10648 2570
rect 10588 2512 10645 2562
rect 10645 2512 10648 2562
rect 10588 2510 10648 2512
rect 10748 2566 10818 2580
rect 10748 2512 10815 2566
rect 10815 2512 10818 2566
rect 10748 2510 10818 2512
rect 11030 2520 11090 2580
rect 10328 2410 10348 2470
rect 10348 2410 10388 2470
rect 10658 2350 10668 2400
rect 10668 2350 10718 2400
rect 10658 2340 10718 2350
rect 10348 2127 10408 2137
rect 10348 2077 10398 2127
rect 10398 2077 10408 2127
rect 11130 2430 11190 2490
rect 10578 1954 10638 1960
rect 10578 1904 10579 1954
rect 10579 1904 10638 1954
rect 10578 1900 10638 1904
rect 10748 1954 10818 1960
rect 10748 1900 10815 1954
rect 10815 1900 10818 1954
rect 10748 1890 10818 1900
rect 11030 1900 11090 1960
rect 10588 1838 10648 1850
rect 10588 1790 10648 1838
rect 10950 1790 11010 1850
rect 10828 1650 10898 1720
rect 10348 1520 10408 1580
rect 10688 1570 10697 1600
rect 10697 1570 10731 1600
rect 10731 1570 10748 1600
rect 10688 1540 10748 1570
rect 10568 1340 10631 1406
rect 10618 1230 10678 1290
rect 10860 1240 10920 1300
rect 10428 1009 10488 1020
rect 10428 961 10488 1009
rect 10698 1025 10768 1030
rect 10698 977 10702 1025
rect 10702 977 10767 1025
rect 10767 977 10768 1025
rect 10698 970 10768 977
rect 10428 960 10488 961
rect 10618 864 10678 870
rect 10618 816 10622 864
rect 10622 816 10678 864
rect 10618 810 10678 816
rect 10338 680 10398 740
rect 10758 560 10828 630
rect 10600 380 10660 440
rect 10400 180 10470 250
rect 10348 72 10408 132
rect 10456 72 10516 132
rect 10300 -40 10360 20
rect 10120 -130 10130 -70
rect 10130 -130 10170 -70
rect 10170 -130 10180 -70
rect 9740 -520 9800 -460
rect 10850 70 10910 130
rect 10760 -130 10820 -70
rect 10500 -230 10560 -170
rect 10348 -340 10408 -280
rect 10456 -340 10516 -280
rect 10400 -460 10470 -390
rect 10590 -640 10650 -580
rect 10280 -730 10340 -670
rect 10760 -730 10820 -670
rect 10610 -830 10670 -770
rect 10420 -930 10480 -870
rect 10359 -1046 10419 -986
rect 10467 -1046 10527 -986
rect 10510 -1240 10570 -1180
rect 10359 -1446 10419 -1386
rect 10467 -1446 10527 -1386
rect 11040 810 11100 870
rect 11040 460 11100 520
rect 11040 190 11100 250
rect 10930 -220 10990 -160
rect 10930 -340 10990 -280
rect 10870 -1050 10930 -990
rect 11040 -460 11100 -400
rect 11220 2340 11280 2400
rect 11300 2087 11360 2147
rect 11650 1650 11720 1720
rect 11480 1540 11540 1600
rect 11380 1310 11440 1370
rect 11300 680 11360 740
rect 11210 370 11270 430
rect 11110 -640 11170 -580
rect 11040 -910 11100 -850
rect 10950 -1440 11010 -1380
rect 10410 -1560 10470 -1500
rect 11040 -1550 11100 -1490
rect 11210 -820 11270 -760
rect 11560 1430 11620 1490
rect 11470 460 11530 520
rect 11650 560 11720 630
rect 11530 70 11590 130
rect 11380 -30 11440 30
rect 11650 -730 11710 -670
rect 11540 -920 11600 -860
rect 11300 -1250 11360 -1190
rect 10600 -1690 10660 -1630
rect 11100 -1690 11160 -1630
rect 6890 -1780 6950 -1720
<< metal2 >>
rect 6890 2750 6950 2760
rect 6890 620 6950 2690
rect 10608 2625 11770 2655
rect 10608 2580 10638 2625
rect 10748 2580 10818 2590
rect 10588 2570 10648 2580
rect 10588 2500 10648 2510
rect 11030 2580 11090 2590
rect 10818 2530 11030 2560
rect 11090 2530 11770 2560
rect 11030 2510 11090 2520
rect 10748 2500 10818 2510
rect 11130 2490 11190 2500
rect 10328 2470 10388 2480
rect 10388 2440 11130 2470
rect 11130 2420 11190 2430
rect 10328 2400 10388 2410
rect 10658 2400 10718 2410
rect 11220 2400 11280 2410
rect 10718 2360 11220 2390
rect 10658 2330 10718 2340
rect 11220 2330 11280 2340
rect 11300 2147 11360 2157
rect 10348 2137 10408 2147
rect 10408 2087 11300 2117
rect 11300 2077 11360 2087
rect 10348 2067 10408 2077
rect 10598 2010 11770 2040
rect 10598 1970 10628 2010
rect 10578 1960 10638 1970
rect 10578 1890 10638 1900
rect 10748 1960 10818 1970
rect 11030 1960 11090 1970
rect 10818 1900 11030 1930
rect 11030 1890 11090 1900
rect 10748 1880 10818 1890
rect 10588 1850 10648 1860
rect 10950 1850 11010 1860
rect 10648 1810 10950 1840
rect 10588 1780 10648 1790
rect 10950 1780 11010 1790
rect 10828 1720 10898 1730
rect 11650 1720 11720 1730
rect 10898 1650 11650 1720
rect 10828 1640 10898 1650
rect 11650 1640 11720 1650
rect 10688 1600 10748 1610
rect 10348 1580 10408 1590
rect 11480 1600 11540 1610
rect 10748 1550 11480 1580
rect 10688 1530 10748 1540
rect 11480 1530 11540 1540
rect 10348 1510 10408 1520
rect 10358 1480 10388 1510
rect 11560 1490 11620 1500
rect 10358 1450 11560 1480
rect 11560 1420 11620 1430
rect 10568 1406 10631 1416
rect 10631 1370 10648 1380
rect 11380 1370 11440 1380
rect 10631 1340 11380 1370
rect 10568 1330 10631 1340
rect 10860 1300 10920 1310
rect 11380 1300 11440 1310
rect 10618 1290 10678 1300
rect 10860 1230 10920 1240
rect 10618 1220 10678 1230
rect 10428 1020 10488 1030
rect 10628 1020 10658 1220
rect 10488 980 10658 1020
rect 10698 1030 10768 1040
rect 10878 1020 10918 1230
rect 10768 980 10918 1020
rect 10698 960 10768 970
rect 10428 950 10488 960
rect 10618 870 10678 880
rect 11040 870 11100 880
rect 10678 820 11040 850
rect 10618 800 10678 810
rect 11040 800 11100 810
rect 10338 740 10398 750
rect 11300 740 11360 750
rect 10398 680 11300 720
rect 10338 670 10398 680
rect 11300 670 11360 680
rect 3610 560 6890 600
rect 10758 630 10828 640
rect 11650 630 11720 640
rect 6950 560 7610 600
rect 6890 550 6950 560
rect 6890 420 6950 430
rect 6890 -290 6950 360
rect 7570 120 7610 560
rect 10828 560 11650 630
rect 10758 550 10828 560
rect 11650 550 11720 560
rect 11040 520 11100 530
rect 11470 520 11530 530
rect 11100 470 11470 500
rect 11040 450 11100 460
rect 11470 450 11530 460
rect 10600 440 10660 450
rect 11210 430 11270 440
rect 10660 390 11210 420
rect 10600 370 10660 380
rect 11210 360 11270 370
rect 10400 250 10470 260
rect 11040 250 11100 260
rect 10470 200 11040 240
rect 11040 180 11100 190
rect 10400 170 10470 180
rect 9740 130 9800 140
rect 7570 80 9740 120
rect 10348 132 10408 142
rect 9800 80 10348 120
rect 9740 60 9800 70
rect 10348 62 10408 72
rect 10456 132 10516 142
rect 10850 130 10910 140
rect 10516 80 10850 120
rect 10456 62 10516 72
rect 10850 60 10910 70
rect 11530 130 11590 140
rect 11530 60 11590 70
rect 11380 30 11440 40
rect 10300 20 10360 30
rect 10360 -20 11380 10
rect 11440 -20 11770 10
rect 11380 -40 11440 -30
rect 10300 -50 10360 -40
rect 10120 -70 10180 -60
rect 10760 -70 10820 -60
rect 10180 -120 10760 -80
rect 10120 -140 10180 -130
rect 10760 -140 10820 -130
rect 10930 -160 10990 -150
rect 10500 -170 10560 -160
rect 10560 -210 10930 -180
rect 10930 -230 10990 -220
rect 10500 -240 10560 -230
rect 10348 -280 10408 -270
rect 3610 -330 10348 -290
rect 6890 -1720 6950 -330
rect 9600 -1400 9640 -330
rect 10348 -350 10408 -340
rect 10456 -280 10516 -270
rect 10930 -280 10990 -270
rect 10516 -330 10930 -300
rect 10456 -350 10516 -340
rect 10930 -350 10990 -340
rect 10400 -390 10470 -380
rect 9740 -460 9800 -450
rect 11040 -400 11100 -390
rect 10470 -450 11040 -410
rect 10400 -470 10470 -460
rect 11040 -470 11100 -460
rect 9740 -530 9800 -520
rect 9750 -1000 9790 -530
rect 10590 -580 10650 -570
rect 11110 -580 11170 -570
rect 10650 -630 11110 -600
rect 10590 -650 10650 -640
rect 11110 -650 11170 -640
rect 10280 -670 10340 -660
rect 10760 -670 10820 -660
rect 10340 -720 10760 -680
rect 10280 -740 10340 -730
rect 11650 -670 11710 -660
rect 10820 -720 11650 -680
rect 10760 -740 10820 -730
rect 11650 -740 11710 -730
rect 11210 -760 11270 -750
rect 10610 -770 10670 -760
rect 10670 -810 11210 -780
rect 11210 -830 11270 -820
rect 10610 -840 10670 -830
rect 11040 -850 11100 -840
rect 10420 -870 10480 -860
rect 10480 -900 11040 -870
rect 11540 -860 11600 -850
rect 11100 -900 11540 -870
rect 11040 -920 11100 -910
rect 11540 -930 11600 -920
rect 10420 -940 10480 -930
rect 10359 -986 10419 -976
rect 9750 -1040 10359 -1000
rect 10359 -1056 10419 -1046
rect 10467 -986 10527 -976
rect 10870 -990 10930 -980
rect 10527 -1030 10870 -1000
rect 10467 -1056 10527 -1046
rect 10870 -1060 10930 -1050
rect 10510 -1180 10570 -1170
rect 11300 -1190 11360 -1180
rect 10570 -1230 11300 -1200
rect 10510 -1250 10570 -1240
rect 11300 -1260 11360 -1250
rect 10359 -1386 10419 -1376
rect 9600 -1440 10359 -1400
rect 10359 -1456 10419 -1446
rect 10467 -1386 10527 -1376
rect 10950 -1380 11010 -1370
rect 10527 -1430 10950 -1390
rect 10467 -1456 10527 -1446
rect 10950 -1450 11010 -1440
rect 11040 -1490 11100 -1480
rect 10410 -1500 10470 -1490
rect 10470 -1550 11040 -1530
rect 10470 -1560 11100 -1550
rect 10410 -1570 10470 -1560
rect 10600 -1630 10660 -1620
rect 11100 -1630 11160 -1620
rect 10660 -1670 11100 -1640
rect 10600 -1700 10660 -1690
rect 11100 -1700 11160 -1690
rect 6890 -1790 6950 -1780
use sky130_fd_pr__pfet_01v8_lvt_B59788  sky130_fd_pr__pfet_01v8_lvt_B59788_0
timestamp 1717106919
transform 1 0 6954 0 1 -681
box -3254 -1219 3254 1219
use sky130_fd_pr__pfet_01v8_M4CK9Z  sky130_fd_pr__pfet_01v8_M4CK9Z_0
timestamp 1717106919
transform 1 0 10481 0 -1 -313
box -359 -261 359 261
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 10834 0 1 1689
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1710522493
transform 1 0 10834 0 -1 2777
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1710522493
transform 1 0 10834 0 1 601
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10834 0 -1 2777
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1710522493
transform -1 0 10834 0 1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10558 0 -1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1710522493
transform -1 0 10558 0 -1 2777
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1710522493
transform -1 0 10558 0 1 1689
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1710522493
transform 1 0 10282 0 1 601
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1710522493
transform 1 0 10558 0 1 601
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform -1 0 10926 0 -1 1689
box -38 -48 406 592
use sky130_fd_pr__pfet_01v8_lvt_B59788  XM24
timestamp 1717106919
transform 1 0 6954 0 1 1651
box -3254 -1219 3254 1219
use sky130_fd_pr__nfet_01v8_75Z3GH  XM27
timestamp 1717106919
transform 1 0 10541 0 1 -1416
box -311 -252 311 252
use sky130_fd_pr__pfet_01v8_M4CK9Z  XM29
timestamp 1717106919
transform 1 0 10481 0 1 103
box -359 -261 359 261
use sky130_fd_pr__nfet_01v8_75Z3GH  XM37
timestamp 1717106919
transform 1 0 10541 0 -1 -1018
box -311 -252 311 252
<< labels >>
rlabel metal2 3610 -330 3650 -290 1 CAL_P
port 3 n
rlabel metal2 3610 560 3650 600 1 CAL_N
port 4 n
rlabel metal1 9980 2820 10140 2880 1 VDD
port 0 n
flabel metal1 11050 305 11080 335 0 FreeSans 80 0 0 0 LOAD_CAL_Z
flabel metal1 10960 300 10990 330 0 FreeSans 80 0 0 0 EN_COMP_Z
flabel metal1 11140 310 11170 340 0 FreeSans 80 0 0 0 CAL_RESULTi
flabel metal1 11220 480 11250 510 0 FreeSans 80 0 0 0 CAL_RESULT_Z
flabel metal1 11310 460 11340 490 0 FreeSans 80 0 0 0 EN_COMPi
rlabel metal2 11740 2530 11770 2560 1 CAL_CYCLE
port 7 n
rlabel metal2 11740 2625 11770 2655 1 CAL_RESULT
port 1 n
rlabel metal2 11735 2010 11765 2040 1 EN_COMP
port 2 n
rlabel metal2 11735 -20 11765 10 1 EN
port 5 n
rlabel metal1 10348 2820 10508 2880 1 VSS
port 6 n
<< end >>
