magic
tech sky130A
magscale 1 2
timestamp 1717106919
<< error_p >>
rect -77 281 -19 287
rect 115 281 173 287
rect -77 247 -65 281
rect 115 247 127 281
rect -77 241 -19 247
rect 115 241 173 247
rect -173 -247 -115 -241
rect 19 -247 77 -241
rect -173 -281 -161 -247
rect 19 -281 31 -247
rect -173 -287 -115 -281
rect 19 -287 77 -281
<< nwell >>
rect -359 -419 359 419
<< pmoshvt >>
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
<< pdiff >>
rect -221 188 -159 200
rect -221 -188 -209 188
rect -175 -188 -159 188
rect -221 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 221 200
rect 159 -188 175 188
rect 209 -188 221 188
rect 159 -200 221 -188
<< pdiffc >>
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
<< nsubdiff >>
rect -323 349 -227 383
rect 227 349 323 383
rect -323 287 -289 349
rect 289 287 323 349
rect -323 -349 -289 -287
rect 289 -349 323 -287
rect -323 -383 -227 -349
rect 227 -383 323 -349
<< nsubdiffcont >>
rect -227 349 227 383
rect -323 -287 -289 287
rect 289 -287 323 287
rect -227 -383 227 -349
<< poly >>
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
<< polycont >>
rect -65 247 -31 281
rect 127 247 161 281
rect -161 -281 -127 -247
rect 31 -281 65 -247
<< locali >>
rect -323 349 -227 383
rect 227 349 323 383
rect -323 287 -289 349
rect 289 287 323 349
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect -323 -349 -289 -287
rect 289 -349 323 -287
rect -323 -383 -227 -349
rect 227 -383 323 -349
<< viali >>
rect -65 247 -31 281
rect 127 247 161 281
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect -161 -281 -127 -247
rect 31 -281 65 -247
<< metal1 >>
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
<< properties >>
string FIXED_BBOX -306 -366 306 366
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 2 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
