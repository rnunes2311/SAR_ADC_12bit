magic
tech sky130A
magscale 1 2
timestamp 1711821647
<< error_p >>
rect 74 1542 132 1548
rect 74 1508 86 1542
rect 74 1502 132 1508
rect 74 1139 132 1145
rect 74 1105 86 1139
rect 74 1099 132 1105
rect 76 706 134 712
rect 76 672 88 706
rect 76 666 134 672
rect -764 316 -706 322
rect -554 316 -496 322
rect -344 316 -286 322
rect -134 316 -76 322
rect 76 316 134 322
rect -764 282 -752 316
rect -554 282 -542 316
rect -344 282 -332 316
rect -134 282 -122 316
rect 76 282 88 316
rect -764 276 -706 282
rect -554 276 -496 282
rect -344 276 -286 282
rect -134 276 -76 282
rect 76 276 134 282
<< pwell >>
rect 70 1492 136 1558
rect -768 266 -702 332
rect -348 266 -282 332
rect 72 266 138 332
<< nmos >>
rect 88 1270 118 1470
rect 88 867 118 1067
rect 90 434 120 634
rect -750 44 -720 244
rect -540 44 -510 244
rect -330 44 -300 244
rect -120 44 -90 244
rect 90 44 120 244
<< ndiff >>
rect 26 1458 88 1470
rect 26 1282 38 1458
rect 72 1282 88 1458
rect 26 1270 88 1282
rect 118 1458 180 1470
rect 118 1282 134 1458
rect 168 1282 180 1458
rect 118 1270 180 1282
rect 26 1055 88 1067
rect 26 879 38 1055
rect 72 879 88 1055
rect 26 867 88 879
rect 118 1055 180 1067
rect 118 879 134 1055
rect 168 879 180 1055
rect 118 867 180 879
rect 28 622 90 634
rect 28 446 40 622
rect 74 446 90 622
rect 28 434 90 446
rect 120 622 182 634
rect 120 446 136 622
rect 170 446 182 622
rect 120 434 182 446
rect -812 232 -750 244
rect -812 56 -800 232
rect -766 56 -750 232
rect -812 44 -750 56
rect -720 232 -658 244
rect -720 56 -704 232
rect -670 56 -658 232
rect -720 44 -658 56
rect -602 232 -540 244
rect -602 56 -590 232
rect -556 56 -540 232
rect -602 44 -540 56
rect -510 232 -448 244
rect -510 56 -494 232
rect -460 56 -448 232
rect -510 44 -448 56
rect -392 232 -330 244
rect -392 56 -380 232
rect -346 56 -330 232
rect -392 44 -330 56
rect -300 232 -238 244
rect -300 56 -284 232
rect -250 56 -238 232
rect -300 44 -238 56
rect -182 232 -120 244
rect -182 56 -170 232
rect -136 56 -120 232
rect -182 44 -120 56
rect -90 232 -28 244
rect -90 56 -74 232
rect -40 56 -28 232
rect -90 44 -28 56
rect 28 232 90 244
rect 28 56 40 232
rect 74 56 90 232
rect 28 44 90 56
rect 120 232 182 244
rect 120 56 136 232
rect 170 56 182 232
rect 120 44 182 56
<< ndiffc >>
rect 38 1282 72 1458
rect 134 1282 168 1458
rect 38 879 72 1055
rect 134 879 168 1055
rect 40 446 74 622
rect 136 446 170 622
rect -800 56 -766 232
rect -704 56 -670 232
rect -590 56 -556 232
rect -494 56 -460 232
rect -380 56 -346 232
rect -284 56 -250 232
rect -170 56 -136 232
rect -74 56 -40 232
rect 40 56 74 232
rect 136 56 170 232
<< poly >>
rect 70 1542 136 1558
rect 70 1508 86 1542
rect 120 1508 136 1542
rect 70 1492 136 1508
rect 88 1470 118 1492
rect 88 1244 118 1270
rect 70 1139 136 1155
rect 70 1105 86 1139
rect 120 1105 136 1139
rect 70 1089 136 1105
rect 88 1067 118 1089
rect 88 841 118 867
rect 72 706 138 722
rect 72 672 88 706
rect 122 672 138 706
rect 72 656 138 672
rect 90 634 120 656
rect 90 408 120 434
rect -768 316 -702 332
rect -768 282 -752 316
rect -718 282 -702 316
rect -768 266 -702 282
rect -558 316 -492 332
rect -558 282 -542 316
rect -508 282 -492 316
rect -558 266 -492 282
rect -348 316 -282 332
rect -348 282 -332 316
rect -298 282 -282 316
rect -348 266 -282 282
rect -138 316 -72 332
rect -138 282 -122 316
rect -88 282 -72 316
rect -138 266 -72 282
rect 72 316 138 332
rect 72 282 88 316
rect 122 282 138 316
rect 72 266 138 282
rect -750 244 -720 266
rect -540 244 -510 266
rect -330 244 -300 266
rect -120 244 -90 266
rect 90 244 120 266
rect -750 18 -720 44
rect -540 18 -510 44
rect -330 18 -300 44
rect -120 18 -90 44
rect 90 18 120 44
<< polycont >>
rect 86 1508 120 1542
rect 86 1105 120 1139
rect 88 672 122 706
rect -752 282 -718 316
rect -542 282 -508 316
rect -332 282 -298 316
rect -122 282 -88 316
rect 88 282 122 316
<< locali >>
rect 70 1508 86 1542
rect 120 1508 136 1542
rect 38 1458 72 1474
rect 38 1266 72 1282
rect 134 1458 168 1474
rect 134 1266 168 1282
rect 70 1105 86 1139
rect 120 1105 136 1139
rect 38 1055 72 1071
rect 38 863 72 879
rect 134 1055 168 1071
rect 134 863 168 879
rect 72 672 88 706
rect 122 672 138 706
rect 40 622 74 638
rect 40 430 74 446
rect 136 622 170 638
rect 136 430 170 446
rect -768 282 -752 316
rect -718 282 -702 316
rect -558 282 -542 316
rect -508 282 -492 316
rect -348 282 -332 316
rect -298 282 -282 316
rect -138 282 -122 316
rect -88 282 -72 316
rect 72 282 88 316
rect 122 282 138 316
rect -800 232 -766 248
rect -800 40 -766 56
rect -704 232 -670 248
rect -704 40 -670 56
rect -590 232 -556 248
rect -590 40 -556 56
rect -494 232 -460 248
rect -494 40 -460 56
rect -380 232 -346 248
rect -380 40 -346 56
rect -284 232 -250 248
rect -284 40 -250 56
rect -170 232 -136 248
rect -170 40 -136 56
rect -74 232 -40 248
rect -74 40 -40 56
rect 40 232 74 248
rect 40 40 74 56
rect 136 232 170 248
rect 136 40 170 56
<< viali >>
rect 86 1508 120 1542
rect 38 1282 72 1458
rect 134 1282 168 1458
rect 86 1105 120 1139
rect 38 879 72 1055
rect 134 879 168 1055
rect 88 672 122 706
rect 40 446 74 622
rect 136 446 170 622
rect -752 282 -718 316
rect -542 282 -508 316
rect -332 282 -298 316
rect -122 282 -88 316
rect 88 282 122 316
rect -800 56 -766 232
rect -704 56 -670 232
rect -590 56 -556 232
rect -494 56 -460 232
rect -380 56 -346 232
rect -284 56 -250 232
rect -170 56 -136 232
rect -74 56 -40 232
rect 40 56 74 232
rect 136 56 170 232
<< metal1 >>
rect 74 1542 132 1548
rect 74 1508 86 1542
rect 120 1508 132 1542
rect 74 1502 132 1508
rect 32 1458 78 1470
rect 32 1282 38 1458
rect 72 1282 78 1458
rect 32 1270 78 1282
rect 128 1458 174 1470
rect 128 1282 134 1458
rect 168 1282 174 1458
rect 128 1270 174 1282
rect 74 1139 132 1145
rect 74 1105 86 1139
rect 120 1105 132 1139
rect 74 1099 132 1105
rect 32 1055 78 1067
rect 32 879 38 1055
rect 72 879 78 1055
rect 32 867 78 879
rect 128 1055 174 1067
rect 128 879 134 1055
rect 168 879 174 1055
rect 128 867 174 879
rect 76 706 134 712
rect 76 672 88 706
rect 122 672 134 706
rect 76 666 134 672
rect 34 622 80 634
rect 34 446 40 622
rect 74 446 80 622
rect 34 434 80 446
rect 130 622 176 634
rect 130 446 136 622
rect 170 446 176 622
rect 130 434 176 446
rect -764 316 -706 322
rect -764 282 -752 316
rect -718 282 -706 316
rect -764 276 -706 282
rect -554 316 -496 322
rect -554 282 -542 316
rect -508 282 -496 316
rect -554 276 -496 282
rect -344 316 -286 322
rect -344 282 -332 316
rect -298 282 -286 316
rect -344 276 -286 282
rect -134 316 -76 322
rect -134 282 -122 316
rect -88 282 -76 316
rect -134 276 -76 282
rect 76 316 134 322
rect 76 282 88 316
rect 122 282 134 316
rect 76 276 134 282
rect -806 232 -760 244
rect -806 56 -800 232
rect -766 56 -760 232
rect -806 44 -760 56
rect -710 232 -664 244
rect -710 56 -704 232
rect -670 56 -664 232
rect -710 44 -664 56
rect -596 232 -550 244
rect -596 56 -590 232
rect -556 56 -550 232
rect -596 44 -550 56
rect -500 232 -454 244
rect -500 56 -494 232
rect -460 56 -454 232
rect -500 44 -454 56
rect -386 232 -340 244
rect -386 56 -380 232
rect -346 56 -340 232
rect -386 44 -340 56
rect -290 232 -244 244
rect -290 56 -284 232
rect -250 56 -244 232
rect -290 44 -244 56
rect -176 232 -130 244
rect -176 56 -170 232
rect -136 56 -130 232
rect -176 44 -130 56
rect -80 232 -34 244
rect -80 56 -74 232
rect -40 56 -34 232
rect -80 44 -34 56
rect 34 232 80 244
rect 34 56 40 232
rect 74 56 80 232
rect 34 44 80 56
rect 130 232 176 244
rect 130 56 136 232
rect 170 56 176 232
rect 130 44 176 56
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
