magic
tech sky130A
magscale 1 2
timestamp 1713891259
<< viali >>
rect -220 940 -170 990
rect -770 854 -720 904
rect -650 860 -600 910
rect -40 854 10 904
rect 130 864 180 914
rect 240 674 290 724
rect 240 420 290 470
rect -770 240 -720 290
rect -660 240 -610 290
rect -40 240 10 290
rect 130 230 180 280
rect -220 160 -170 210
<< metal1 >>
rect -232 990 -158 996
rect -232 934 -220 990
rect -160 979 -150 990
rect -160 949 168 979
rect -230 930 -220 934
rect -160 930 -150 949
rect 138 920 168 949
rect -662 910 -588 916
rect 118 914 192 920
rect -782 904 -708 910
rect -790 844 -780 904
rect -720 848 -708 904
rect -662 860 -650 910
rect -600 860 -588 910
rect -662 854 -588 860
rect -60 854 -50 914
rect 10 910 20 914
rect 10 854 22 910
rect 118 864 130 914
rect 180 864 192 914
rect 118 858 192 864
rect -720 844 -710 848
rect -635 810 -605 854
rect -52 848 22 854
rect -660 750 -650 810
rect -590 750 -580 810
rect -635 714 -605 750
rect 228 724 302 730
rect 228 714 240 724
rect -635 684 240 714
rect 228 674 240 684
rect 290 674 302 724
rect 228 668 302 674
rect 228 470 302 476
rect 228 460 240 470
rect -650 430 240 460
rect -790 240 -780 300
rect -720 296 -710 300
rect -650 296 -620 430
rect 228 420 240 430
rect 290 420 302 470
rect 228 414 302 420
rect -720 240 -708 296
rect -782 234 -708 240
rect -672 290 -598 296
rect -52 290 22 296
rect -672 240 -660 290
rect -610 240 -598 290
rect -672 234 -598 240
rect -650 200 -620 234
rect -60 230 -50 290
rect 10 234 22 290
rect 118 280 192 286
rect 10 230 20 234
rect 118 230 130 280
rect 180 230 192 280
rect 118 224 192 230
rect -230 216 -220 220
rect -670 140 -660 200
rect -600 140 -590 200
rect -232 160 -220 216
rect -160 195 -150 220
rect 138 195 168 224
rect -160 165 168 195
rect -160 160 -150 165
rect -232 154 -158 160
<< via1 >>
rect -220 940 -170 990
rect -170 940 -160 990
rect -220 930 -160 940
rect -780 854 -770 904
rect -770 854 -720 904
rect -780 844 -720 854
rect -50 904 10 914
rect -50 854 -40 904
rect -40 854 10 904
rect -650 750 -590 810
rect -780 290 -720 300
rect -780 240 -770 290
rect -770 240 -720 290
rect -50 240 -40 290
rect -40 240 10 290
rect -50 230 10 240
rect -660 140 -600 200
rect -220 210 -160 220
rect -220 160 -170 210
rect -170 160 -160 210
<< metal2 >>
rect -890 1028 -5 1058
rect -220 990 -160 1000
rect -890 914 -745 934
rect -220 920 -160 930
rect -35 924 -5 1028
rect -890 904 -720 914
rect -780 834 -720 844
rect -650 810 -590 820
rect -890 750 -650 780
rect -650 740 -590 750
rect -645 627 -615 660
rect -210 627 -180 920
rect -50 914 10 924
rect -50 844 10 854
rect -890 597 -180 627
rect -890 435 -615 465
rect -890 310 -745 340
rect -780 300 -720 310
rect -645 300 -615 435
rect -645 290 10 300
rect -645 270 -50 290
rect -780 230 -720 240
rect -220 220 -160 230
rect -50 220 10 230
rect -660 200 -600 210
rect -890 170 -660 200
rect -220 150 -160 160
rect -660 130 -600 140
rect -205 100 -175 150
rect -890 70 -175 100
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -792 0 -1 1116
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_1
timestamp 1710522493
transform 1 0 -792 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -56 0 -1 1116
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_1
timestamp 1710522493
transform 1 0 -56 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -148 0 -1 1116
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1710522493
transform 1 0 -148 0 1 28
box -38 -48 130 592
<< end >>
