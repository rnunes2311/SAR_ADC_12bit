magic
tech sky130A
magscale 1 2
timestamp 1714249130
<< metal1 >>
rect -445 28135 -415 31492
rect -385 28225 -355 31492
rect -325 28315 -295 31492
rect -265 28405 -235 31492
rect -205 28495 -175 31492
rect -145 28585 -115 31492
rect -85 28675 -55 31492
rect -25 28855 5 31492
rect 35 28945 65 31492
rect 95 29035 125 31492
rect 155 29125 185 31492
rect 215 29215 245 31492
rect 275 29305 305 31492
rect 335 29395 365 31492
rect 395 29485 425 31492
rect 455 29575 485 31492
rect 515 29665 545 31492
rect 575 29755 605 31492
rect 635 29845 665 31492
rect 695 29935 725 31492
rect 755 30025 785 31492
rect 815 30140 845 31492
rect 905 31410 935 31492
rect 880 31350 890 31410
rect 950 31350 960 31410
rect 995 30795 1025 31492
rect 995 30765 3025 30795
rect 815 30130 875 30140
rect 815 30060 875 30070
rect 2345 30040 2405 30050
rect 755 29995 2345 30025
rect 2345 29970 2405 29980
rect 3350 29935 3360 29950
rect 695 29905 3360 29935
rect 3350 29890 3360 29905
rect 3420 29890 3430 29950
rect 3870 29845 3880 29860
rect 635 29815 3880 29845
rect 3870 29800 3880 29815
rect 3940 29800 3950 29860
rect 4120 29755 4130 29770
rect 575 29725 4130 29755
rect 4120 29710 4130 29725
rect 4190 29710 4200 29770
rect 4360 29665 4370 29680
rect 515 29635 4370 29665
rect 4360 29620 4370 29635
rect 4430 29620 4440 29680
rect 4610 29575 4620 29590
rect 455 29545 4620 29575
rect 4610 29530 4620 29545
rect 4680 29530 4690 29590
rect 4850 29485 4860 29500
rect 395 29455 4860 29485
rect 4850 29440 4860 29455
rect 4920 29440 4930 29500
rect 5090 29395 5100 29410
rect 335 29365 5100 29395
rect 5090 29350 5100 29365
rect 5160 29350 5170 29410
rect 5340 29305 5350 29320
rect 275 29275 5350 29305
rect 5340 29260 5350 29275
rect 5410 29260 5420 29320
rect 5570 29215 5580 29230
rect 215 29185 5580 29215
rect 5570 29170 5580 29185
rect 5640 29170 5650 29230
rect 8090 29170 8100 29230
rect 8160 29215 8170 29230
rect 8160 29185 15040 29215
rect 8160 29170 8170 29185
rect 6120 29125 6130 29140
rect 155 29095 6130 29125
rect 6120 29080 6130 29095
rect 6190 29080 6200 29140
rect 8860 29080 8870 29140
rect 8930 29125 8940 29140
rect 8930 29095 15040 29125
rect 8930 29080 8940 29095
rect 6890 29035 6900 29050
rect 95 29005 6900 29035
rect 6890 28990 6900 29005
rect 6960 28990 6970 29050
rect 9630 28990 9640 29050
rect 9700 29035 9710 29050
rect 9700 29005 15040 29035
rect 9700 28990 9710 29005
rect 7280 28945 7290 28960
rect 35 28915 7290 28945
rect 7280 28900 7290 28915
rect 7350 28900 7360 28960
rect 10010 28900 10020 28960
rect 10080 28945 10090 28960
rect 10080 28915 15040 28945
rect 10080 28900 10090 28915
rect 7450 28855 7460 28870
rect -25 28825 7460 28855
rect 7450 28810 7460 28825
rect 7520 28810 7530 28870
rect 10200 28810 10210 28870
rect 10270 28855 10280 28870
rect 10270 28825 15040 28855
rect 10270 28810 10280 28825
rect 5940 28720 5950 28780
rect 6010 28765 6020 28780
rect 7670 28765 7680 28780
rect 6010 28735 7680 28765
rect 6010 28720 6020 28735
rect 7670 28720 7680 28735
rect 7740 28720 7750 28780
rect 11690 28720 11700 28780
rect 11760 28765 11770 28780
rect 11760 28735 15040 28765
rect 11760 28720 11770 28735
rect 10410 28675 10420 28690
rect -85 28645 10420 28675
rect 10410 28630 10420 28645
rect 10480 28630 10490 28690
rect 11850 28630 11860 28690
rect 11920 28675 11930 28690
rect 11920 28645 15040 28675
rect 11920 28630 11930 28645
rect 10600 28585 10610 28600
rect -145 28555 10610 28585
rect 10600 28540 10610 28555
rect 10670 28540 10680 28600
rect 12010 28540 12020 28600
rect 12080 28585 12090 28600
rect 12080 28555 15040 28585
rect 12080 28540 12090 28555
rect 10720 28495 10730 28510
rect -205 28465 10730 28495
rect 10720 28450 10730 28465
rect 10790 28450 10800 28510
rect 12170 28450 12180 28510
rect 12240 28495 12250 28510
rect 12240 28465 15040 28495
rect 12240 28450 12250 28465
rect 10930 28405 10940 28420
rect -265 28375 10940 28405
rect 10930 28360 10940 28375
rect 11000 28360 11010 28420
rect 11770 28360 11780 28420
rect 11840 28405 11850 28420
rect 11840 28375 15040 28405
rect 11840 28360 11850 28375
rect 11140 28315 11150 28330
rect -325 28285 11150 28315
rect 11140 28270 11150 28285
rect 11210 28270 11220 28330
rect 11930 28270 11940 28330
rect 12000 28315 12010 28330
rect 12000 28285 15040 28315
rect 12000 28270 12010 28285
rect 11350 28225 11360 28240
rect -385 28195 11360 28225
rect 11350 28180 11360 28195
rect 11420 28180 11430 28240
rect 12090 28180 12100 28240
rect 12160 28225 12170 28240
rect 12160 28195 15040 28225
rect 12160 28180 12170 28195
rect 11560 28135 11570 28150
rect -445 28105 11570 28135
rect 11560 28090 11570 28105
rect 11630 28090 11640 28150
rect 12250 28090 12260 28150
rect 12320 28135 12330 28150
rect 12320 28105 15040 28135
rect 12320 28090 12330 28105
rect 13730 25945 13740 25960
rect 13630 25915 13740 25945
rect 13730 25900 13740 25915
rect 13800 25900 13810 25960
rect 13820 25855 13830 25870
rect 13625 25825 13830 25855
rect 13820 25810 13830 25825
rect 13890 25810 13900 25870
rect 13910 25765 13920 25780
rect 13625 25735 13920 25765
rect 13910 25720 13920 25735
rect 13980 25720 13990 25780
rect 14000 25675 14010 25690
rect 13630 25645 14010 25675
rect 14000 25630 14010 25645
rect 14070 25630 14080 25690
rect 14090 25585 14100 25600
rect 13605 25555 14100 25585
rect 14090 25540 14100 25555
rect 14160 25540 14170 25600
rect 14180 25495 14190 25510
rect 13615 25465 14190 25495
rect 14180 25450 14190 25465
rect 14250 25450 14260 25510
rect 14270 25405 14280 25420
rect 13615 25375 14280 25405
rect 14270 25360 14280 25375
rect 14340 25360 14350 25420
rect 14720 25315 14730 25330
rect 13625 25285 14730 25315
rect 14720 25270 14730 25285
rect 14790 25270 14800 25330
rect 14360 25225 14370 25240
rect 13615 25195 14370 25225
rect 14360 25180 14370 25195
rect 14430 25180 14440 25240
rect 14630 25135 14640 25150
rect 13625 25105 14640 25135
rect 14630 25090 14640 25105
rect 14700 25090 14710 25150
rect 14540 25045 14550 25060
rect 13615 25015 14550 25045
rect 14540 25000 14550 25015
rect 14610 25000 14620 25060
rect 14450 24955 14460 24970
rect 13625 24925 14460 24955
rect 14450 24910 14460 24925
rect 14520 24910 14530 24970
rect 14718 13160 14802 13166
rect 14718 13150 14730 13160
rect 13656 13110 14730 13150
rect 14718 13100 14730 13110
rect 14790 13100 14802 13160
rect 14718 13094 14802 13100
rect 14628 12790 14712 12796
rect 14628 12780 14640 12790
rect 13678 12740 14640 12780
rect 14628 12730 14640 12740
rect 14700 12730 14712 12790
rect 14628 12724 14712 12730
rect 14538 12420 14622 12426
rect 14538 12410 14550 12420
rect 13688 12370 14550 12410
rect 14538 12360 14550 12370
rect 14610 12360 14622 12420
rect 14538 12354 14622 12360
rect 14448 12050 14532 12056
rect 14448 12040 14460 12050
rect 13666 12000 14460 12040
rect 14448 11990 14460 12000
rect 14520 11990 14532 12050
rect 14448 11984 14532 11990
rect 14358 11680 14442 11686
rect 14358 11670 14370 11680
rect 13682 11630 14370 11670
rect 14358 11620 14370 11630
rect 14430 11620 14442 11680
rect 14358 11614 14442 11620
rect 14268 11310 14352 11316
rect 14268 11300 14280 11310
rect 13650 11260 14280 11300
rect 14268 11250 14280 11260
rect 14340 11250 14352 11310
rect 14268 11244 14352 11250
rect 14178 10570 14262 10576
rect 14178 10560 14190 10570
rect 13672 10520 14190 10560
rect 14178 10510 14190 10520
rect 14250 10510 14262 10570
rect 14178 10504 14262 10510
rect 14088 10200 14172 10206
rect 14088 10190 14100 10200
rect 13654 10150 14100 10190
rect 14088 10140 14100 10150
rect 14160 10140 14172 10200
rect 14088 10134 14172 10140
rect 13998 9460 14082 9466
rect 13998 9450 14010 9460
rect 13684 9410 14010 9450
rect 13998 9400 14010 9410
rect 14070 9400 14082 9460
rect 13998 9394 14082 9400
rect 13908 8350 13992 8356
rect 13908 8340 13920 8350
rect 13654 8300 13920 8340
rect 13908 8290 13920 8300
rect 13980 8290 13992 8350
rect 13908 8284 13992 8290
rect 13818 6500 13902 6506
rect 13818 6490 13830 6500
rect 13680 6450 13830 6490
rect 13818 6440 13830 6450
rect 13890 6440 13902 6500
rect 13818 6434 13902 6440
rect 13728 4280 13812 4286
rect 13728 4220 13740 4280
rect 13800 4220 13812 4280
rect 13728 4214 13812 4220
<< via1 >>
rect 890 31350 950 31410
rect 815 30070 875 30130
rect 2345 29980 2405 30040
rect 3360 29890 3420 29950
rect 3880 29800 3940 29860
rect 4130 29710 4190 29770
rect 4370 29620 4430 29680
rect 4620 29530 4680 29590
rect 4860 29440 4920 29500
rect 5100 29350 5160 29410
rect 5350 29260 5410 29320
rect 5580 29170 5640 29230
rect 8100 29170 8160 29230
rect 6130 29080 6190 29140
rect 8870 29080 8930 29140
rect 6900 28990 6960 29050
rect 9640 28990 9700 29050
rect 7290 28900 7350 28960
rect 10020 28900 10080 28960
rect 7460 28810 7520 28870
rect 10210 28810 10270 28870
rect 5950 28720 6010 28780
rect 7680 28720 7740 28780
rect 11700 28720 11760 28780
rect 10420 28630 10480 28690
rect 11860 28630 11920 28690
rect 10610 28540 10670 28600
rect 12020 28540 12080 28600
rect 10730 28450 10790 28510
rect 12180 28450 12240 28510
rect 10940 28360 11000 28420
rect 11780 28360 11840 28420
rect 11150 28270 11210 28330
rect 11940 28270 12000 28330
rect 11360 28180 11420 28240
rect 12100 28180 12160 28240
rect 11570 28090 11630 28150
rect 12260 28090 12320 28150
rect 13740 25900 13800 25960
rect 13830 25810 13890 25870
rect 13920 25720 13980 25780
rect 14010 25630 14070 25690
rect 14100 25540 14160 25600
rect 14190 25450 14250 25510
rect 14280 25360 14340 25420
rect 14730 25270 14790 25330
rect 14370 25180 14430 25240
rect 14640 25090 14700 25150
rect 14550 25000 14610 25060
rect 14460 24910 14520 24970
rect 14730 13100 14790 13160
rect 14640 12730 14700 12790
rect 14550 12360 14610 12420
rect 14460 11990 14520 12050
rect 14370 11620 14430 11680
rect 14280 11250 14340 11310
rect 14190 10510 14250 10570
rect 14100 10140 14160 10200
rect 14010 9400 14070 9460
rect 13920 8290 13980 8350
rect 13830 6440 13890 6500
rect 13740 4220 13800 4280
<< metal2 >>
rect -380 31720 -320 31730
rect -320 31660 2810 31670
rect -380 31620 2810 31660
rect -320 31610 2810 31620
rect -380 31550 -320 31560
rect 890 31410 950 31420
rect 950 31400 965 31410
rect 950 31360 2710 31400
rect 950 31350 965 31360
rect 890 31340 950 31350
rect -510 31230 -450 31240
rect -450 31180 4080 31220
rect -510 31160 -450 31170
rect 5950 31170 6010 31180
rect 5950 31100 6010 31110
rect -120 30590 -50 30600
rect -60 30556 -50 30590
rect -60 30530 2941 30556
rect -120 30500 2941 30530
rect -60 30440 2941 30500
rect -120 30410 2941 30440
rect -60 30380 2941 30410
rect -60 30350 -50 30380
rect -120 30340 -50 30350
rect 5950 30170 6010 30180
rect 805 30120 815 30130
rect 300 30080 815 30120
rect 300 28000 340 30080
rect 805 30070 815 30080
rect 875 30070 885 30130
rect 5950 30100 6010 30110
rect 2345 30040 2405 30050
rect 2345 29970 2405 29980
rect 2345 28050 2385 29970
rect 3360 29950 3420 29960
rect 3360 29880 3420 29890
rect 3370 28040 3410 29880
rect 3880 29860 3940 29870
rect 3880 29790 3940 29800
rect 3890 28060 3930 29790
rect 4130 29770 4190 29780
rect 4130 29700 4190 29710
rect 4140 28040 4180 29700
rect 4370 29680 4430 29690
rect 4370 29610 4430 29620
rect 4380 28040 4420 29610
rect 4620 29590 4680 29600
rect 4620 29520 4680 29530
rect 4630 28040 4670 29520
rect 4860 29500 4920 29510
rect 4860 29430 4920 29440
rect 4870 28040 4910 29430
rect 5100 29410 5160 29420
rect 5100 29340 5160 29350
rect 5110 28060 5150 29340
rect 5350 29320 5410 29330
rect 5350 29250 5410 29260
rect 5360 28080 5400 29250
rect 5580 29230 5640 29240
rect 5580 29160 5640 29170
rect 5590 28060 5630 29160
rect 5960 28790 6000 30100
rect 8100 29230 8160 29240
rect 8100 29160 8160 29170
rect 6130 29140 6190 29150
rect 6130 29070 6190 29080
rect 5950 28780 6010 28790
rect 5950 28710 6010 28720
rect 6140 28050 6180 29070
rect 6900 29050 6960 29060
rect 6900 28980 6960 28990
rect 6910 28040 6950 28980
rect 7290 28960 7350 28970
rect 7290 28890 7350 28900
rect 7300 28050 7340 28890
rect 7460 28870 7520 28880
rect 7460 28800 7520 28810
rect 7470 28020 7510 28800
rect 7680 28780 7740 28790
rect 7680 28710 7740 28720
rect 7690 28050 7730 28710
rect 8110 28080 8150 29160
rect 8870 29140 8930 29150
rect 8870 29070 8930 29080
rect 8880 28090 8920 29070
rect 9640 29050 9700 29060
rect 9640 28980 9700 28990
rect 9650 28080 9690 28980
rect 10020 28960 10080 28970
rect 10020 28890 10080 28900
rect 10030 28080 10070 28890
rect 10210 28870 10270 28880
rect 10210 28800 10270 28810
rect 10220 28080 10260 28800
rect 11700 28780 11760 28790
rect 11700 28710 11760 28720
rect 10420 28690 10480 28700
rect 10420 28620 10480 28630
rect 10430 28060 10470 28620
rect 10610 28600 10670 28610
rect 10610 28530 10670 28540
rect 10620 28060 10660 28530
rect 10730 28510 10790 28520
rect 10730 28440 10790 28450
rect 10740 28060 10780 28440
rect 10940 28420 11000 28430
rect 10940 28350 11000 28360
rect 10950 28040 10990 28350
rect 11150 28330 11210 28340
rect 11150 28260 11210 28270
rect 11160 28060 11200 28260
rect 11360 28240 11420 28250
rect 11360 28170 11420 28180
rect 11370 28050 11410 28170
rect 11570 28150 11630 28160
rect 11570 28080 11630 28090
rect 11710 28080 11750 28710
rect 11860 28690 11920 28700
rect 11860 28620 11920 28630
rect 11780 28420 11840 28430
rect 11780 28350 11840 28360
rect 11790 28080 11830 28350
rect 11870 28080 11910 28620
rect 12020 28600 12080 28610
rect 12020 28530 12080 28540
rect 11940 28330 12000 28340
rect 11940 28260 12000 28270
rect 11950 28080 11990 28260
rect 12030 28080 12070 28530
rect 12180 28510 12240 28520
rect 12180 28440 12240 28450
rect 12100 28240 12160 28250
rect 12100 28170 12160 28180
rect 12110 28080 12150 28170
rect 12190 28080 12230 28440
rect 12260 28150 12320 28160
rect 12260 28080 12320 28090
rect 10 27740 70 27750
rect 70 27695 90 27735
rect 10 27670 70 27680
rect -120 27440 -60 27450
rect -60 27395 90 27435
rect -120 27370 -60 27380
rect -250 27130 -190 27140
rect -190 27085 90 27125
rect -250 27060 -190 27070
rect -380 26720 -320 26730
rect -320 26675 90 26715
rect -380 26650 -320 26660
rect -510 26590 -450 26600
rect -450 26545 90 26585
rect -510 26520 -450 26530
rect 13740 25960 13800 25970
rect 13740 25890 13800 25900
rect 13750 4290 13790 25890
rect 13830 25870 13890 25880
rect 13830 25800 13890 25810
rect 13840 6510 13880 25800
rect 13920 25780 13980 25790
rect 13920 25710 13980 25720
rect 13930 8360 13970 25710
rect 14010 25690 14070 25700
rect 14010 25620 14070 25630
rect 14020 9470 14060 25620
rect 14100 25600 14160 25610
rect 14100 25530 14160 25540
rect 14110 10210 14150 25530
rect 14190 25510 14250 25520
rect 14190 25440 14250 25450
rect 14200 10580 14240 25440
rect 14280 25420 14340 25430
rect 14280 25350 14340 25360
rect 14290 11320 14330 25350
rect 14730 25330 14790 25340
rect 14730 25260 14790 25270
rect 14370 25240 14430 25250
rect 14370 25170 14430 25180
rect 14380 11690 14420 25170
rect 14640 25150 14700 25160
rect 14640 25080 14700 25090
rect 14550 25060 14610 25070
rect 14550 24990 14610 25000
rect 14460 24970 14520 24980
rect 14460 24900 14520 24910
rect 14470 12060 14510 24900
rect 14560 12430 14600 24990
rect 14650 12800 14690 25080
rect 14740 13170 14780 25260
rect 14730 13160 14790 13170
rect 14730 13090 14790 13100
rect 14640 12790 14700 12800
rect 14640 12720 14700 12730
rect 14550 12420 14610 12430
rect 14550 12350 14610 12360
rect 14460 12050 14520 12060
rect 14460 11980 14520 11990
rect 14370 11680 14430 11690
rect 14370 11610 14430 11620
rect 14280 11310 14340 11320
rect 14280 11240 14340 11250
rect 14190 10570 14250 10580
rect 14190 10500 14250 10510
rect 14100 10200 14160 10210
rect 14100 10130 14160 10140
rect 14010 9460 14070 9470
rect 14010 9390 14070 9400
rect 13920 8350 13980 8360
rect 13920 8280 13980 8290
rect 13830 6500 13890 6510
rect 13830 6430 13890 6440
rect 13740 4280 13800 4290
rect 13740 4210 13800 4220
<< via2 >>
rect -380 31660 -320 31720
rect -380 31560 -320 31620
rect -510 31170 -450 31230
rect 5950 31110 6010 31170
rect -120 30530 -60 30590
rect -120 30440 -60 30500
rect -120 30350 -60 30410
rect 5950 30110 6010 30170
rect 10 27680 70 27740
rect -120 27380 -60 27440
rect -250 27070 -190 27130
rect -380 26660 -320 26720
rect -510 26530 -450 26590
<< metal3 >>
rect -510 31235 -450 31800
rect -380 31725 -320 31800
rect -390 31720 -310 31725
rect -390 31660 -380 31720
rect -320 31660 -310 31720
rect -390 31620 -310 31660
rect -390 31560 -380 31620
rect -320 31560 -310 31620
rect -390 31555 -310 31560
rect -520 31230 -440 31235
rect -520 31170 -510 31230
rect -450 31170 -440 31230
rect -520 31165 -440 31170
rect -510 26595 -450 31165
rect -380 26725 -320 31555
rect -250 27135 -190 31800
rect -120 30595 -60 31800
rect -130 30590 -50 30595
rect -130 30530 -120 30590
rect -60 30530 -50 30590
rect -130 30500 -50 30530
rect -130 30440 -120 30500
rect -60 30440 -50 30500
rect -130 30410 -50 30440
rect -130 30350 -120 30410
rect -60 30350 -50 30410
rect -130 30345 -50 30350
rect -120 27445 -60 30345
rect 10 27745 70 31800
rect 5940 31170 6020 31180
rect 5940 31110 5950 31170
rect 6010 31110 6020 31170
rect 5940 31100 6020 31110
rect 5950 30180 6010 31100
rect 5940 30170 6020 30180
rect 5940 30110 5950 30170
rect 6010 30110 6020 30170
rect 5940 30100 6020 30110
rect 0 27740 80 27745
rect 0 27680 10 27740
rect 70 27680 80 27740
rect 0 27675 80 27680
rect -130 27440 -50 27445
rect -130 27380 -120 27440
rect -60 27380 -50 27440
rect -130 27375 -50 27380
rect -260 27130 -180 27135
rect -260 27070 -250 27130
rect -190 27070 -180 27130
rect -260 27065 -180 27070
rect -390 26720 -310 26725
rect -390 26660 -380 26720
rect -320 26660 -310 26720
rect -390 26655 -310 26660
rect -520 26590 -440 26595
rect -520 26530 -510 26590
rect -450 26530 -440 26590
rect -520 26525 -440 26530
use bootstrap  bootstrap_0 ~/Desktop/SAR_ADC_12bit/layout/../bootstrap/layout
timestamp 1711831820
transform -1 0 22799 0 -1 31768
box 9245 72 20179 2258
use CDAC_mim_12bit  CDAC_mim_12bit_1 ~/Desktop/SAR_ADC_12bit/layout/../CDAC
timestamp 1712086820
transform 1 0 400 0 1 370
box -400 -370 13390 24200
use switches  switches_0 ~/Desktop/SAR_ADC_12bit/layout/../switches/layout
timestamp 1711974700
transform 1 0 220 0 1 24045
box -200 855 13477 4090
<< end >>
