magic
tech sky130A
timestamp 1711975147
<< error_p >>
rect -67 86 -38 89
rect 143 86 172 89
rect -67 69 -61 86
rect 143 69 149 86
rect -67 66 -38 69
rect 143 66 172 69
rect -172 -69 -143 -66
rect 38 -69 67 -66
rect -172 -86 -166 -69
rect 38 -86 44 -69
rect -172 -89 -143 -86
rect 38 -89 67 -86
<< pwell >>
rect -265 -155 265 155
<< nmoslvt >>
rect -165 -50 -150 50
rect -60 -50 -45 50
rect 45 -50 60 50
rect 150 -50 165 50
<< ndiff >>
rect -196 44 -165 50
rect -196 -44 -190 44
rect -173 -44 -165 44
rect -196 -50 -165 -44
rect -150 44 -119 50
rect -150 -44 -142 44
rect -125 -44 -119 44
rect -150 -50 -119 -44
rect -91 44 -60 50
rect -91 -44 -85 44
rect -68 -44 -60 44
rect -91 -50 -60 -44
rect -45 44 -14 50
rect -45 -44 -37 44
rect -20 -44 -14 44
rect -45 -50 -14 -44
rect 14 44 45 50
rect 14 -44 20 44
rect 37 -44 45 44
rect 14 -50 45 -44
rect 60 44 91 50
rect 60 -44 68 44
rect 85 -44 91 44
rect 60 -50 91 -44
rect 119 44 150 50
rect 119 -44 125 44
rect 142 -44 150 44
rect 119 -50 150 -44
rect 165 44 196 50
rect 165 -44 173 44
rect 190 -44 196 44
rect 165 -50 196 -44
<< ndiffc >>
rect -190 -44 -173 44
rect -142 -44 -125 44
rect -85 -44 -68 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 68 -44 85 44
rect 125 -44 142 44
rect 173 -44 190 44
<< psubdiff >>
rect -247 120 -199 137
rect 199 120 247 137
rect -247 89 -230 120
rect 230 89 247 120
rect -247 -120 -230 -89
rect 230 -120 247 -89
rect -247 -137 -199 -120
rect 199 -137 247 -120
<< psubdiffcont >>
rect -199 120 199 137
rect -247 -89 -230 89
rect 230 -89 247 89
rect -199 -137 199 -120
<< poly >>
rect -69 86 -36 94
rect -69 69 -61 86
rect -44 69 -36 86
rect -165 50 -150 63
rect -69 61 -36 69
rect 141 86 174 94
rect 141 69 149 86
rect 166 69 174 86
rect -60 50 -45 61
rect 45 50 60 63
rect 141 61 174 69
rect 150 50 165 61
rect -165 -61 -150 -50
rect -174 -69 -141 -61
rect -60 -63 -45 -50
rect 45 -61 60 -50
rect -174 -86 -166 -69
rect -149 -86 -141 -69
rect -174 -94 -141 -86
rect 36 -69 69 -61
rect 150 -63 165 -50
rect 36 -86 44 -69
rect 61 -86 69 -69
rect 36 -94 69 -86
<< polycont >>
rect -61 69 -44 86
rect 149 69 166 86
rect -166 -86 -149 -69
rect 44 -86 61 -69
<< locali >>
rect -247 120 -199 137
rect 199 120 247 137
rect -247 89 -230 120
rect 230 89 247 120
rect -69 69 -61 86
rect -44 69 -36 86
rect 141 69 149 86
rect 166 69 174 86
rect -190 44 -173 52
rect -190 -52 -173 -44
rect -142 44 -125 52
rect -142 -52 -125 -44
rect -85 44 -68 52
rect -85 -52 -68 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 68 44 85 52
rect 68 -52 85 -44
rect 125 44 142 52
rect 125 -52 142 -44
rect 173 44 190 52
rect 173 -52 190 -44
rect -174 -86 -166 -69
rect -149 -86 -141 -69
rect 36 -86 44 -69
rect 61 -86 69 -69
rect -247 -120 -230 -89
rect 230 -120 247 -89
rect -247 -137 -199 -120
rect 199 -137 247 -120
<< viali >>
rect -61 69 -44 86
rect 149 69 166 86
rect -190 -44 -173 44
rect -142 -44 -125 44
rect -85 -44 -68 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 68 -44 85 44
rect 125 -44 142 44
rect 173 -44 190 44
rect -166 -86 -149 -69
rect 44 -86 61 -69
<< metal1 >>
rect -67 86 -38 89
rect -67 69 -61 86
rect -44 69 -38 86
rect -67 66 -38 69
rect 143 86 172 89
rect 143 69 149 86
rect 166 69 172 86
rect 143 66 172 69
rect -193 44 -170 50
rect -193 -44 -190 44
rect -173 -44 -170 44
rect -193 -50 -170 -44
rect -145 44 -122 50
rect -145 -44 -142 44
rect -125 -44 -122 44
rect -145 -50 -122 -44
rect -88 44 -65 50
rect -88 -44 -85 44
rect -68 -44 -65 44
rect -88 -50 -65 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 65 44 88 50
rect 65 -44 68 44
rect 85 -44 88 44
rect 65 -50 88 -44
rect 122 44 145 50
rect 122 -44 125 44
rect 142 -44 145 44
rect 122 -50 145 -44
rect 170 44 193 50
rect 170 -44 173 44
rect 190 -44 193 44
rect 170 -50 193 -44
rect -172 -69 -143 -66
rect -172 -86 -166 -69
rect -149 -86 -143 -69
rect -172 -89 -143 -86
rect 38 -69 67 -66
rect 38 -86 44 -69
rect 61 -86 67 -69
rect 38 -89 67 -86
<< properties >>
string FIXED_BBOX -238 -128 238 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
