magic
tech sky130A
magscale 1 2
timestamp 1715383943
<< pwell >>
rect -400 23970 -220 24000
rect -115 23970 70 24000
rect -400 23940 70 23970
rect 12740 23940 13140 24000
rect -400 -330 13140 23940
<< psubdiff >>
rect -304 23840 -280 23880
rect 13000 23840 13024 23880
rect -370 23740 -330 23770
rect -370 -100 -330 -70
rect -304 -210 -280 -170
rect 13000 -210 13024 -170
<< psubdiffcont >>
rect -280 23840 13000 23880
rect -370 -70 -330 23740
rect -280 -210 13000 -170
<< locali >>
rect -215 24130 -155 24170
rect -205 23880 -165 24130
rect 12980 24075 13040 24115
rect 12995 23880 13035 24075
rect -370 23740 -330 23880
rect -296 23840 -280 23880
rect 13000 23840 13035 23880
rect -370 -140 -330 -70
rect -296 -210 -280 -170
rect 13000 -210 13016 -170
<< viali >>
rect -255 24130 -215 24170
rect -155 24130 -115 24170
rect 12940 24075 12980 24115
rect 13040 24075 13080 24115
rect -270 23840 12910 23880
rect -370 -50 -330 23740
rect -220 -210 12960 -170
<< metal1 >>
rect -275 24120 -265 24180
rect -205 23886 -165 24180
rect -105 24120 -95 24180
rect 12920 24065 12930 24125
rect 12990 24025 13030 24125
rect 13090 24065 13100 24125
rect -282 23880 12922 23886
rect 12995 23880 13035 24025
rect -370 23793 -330 23880
rect -300 23840 -270 23880
rect 12910 23840 13035 23880
rect -282 23834 12922 23840
rect -376 23783 -330 23793
rect -376 23740 -324 23783
rect -376 -50 -370 23740
rect -330 -50 -324 23740
rect 30 23510 70 23540
rect 430 23510 470 23540
rect 830 23510 870 23540
rect 1230 23510 1270 23540
rect 1630 23510 1670 23540
rect 2030 23510 2070 23540
rect 2430 23510 2470 23540
rect 3230 23510 3270 23540
rect 3630 23510 3670 23540
rect 4030 23510 4070 23540
rect 4430 23510 4470 23540
rect 4830 23510 4870 23540
rect 5230 23510 5270 23540
rect 5630 23510 5670 23540
rect 6030 23510 6070 23540
rect 6430 23510 6470 23540
rect 6830 23510 6870 23540
rect 7230 23510 7270 23540
rect 7630 23510 7670 23540
rect 8030 23510 8070 23540
rect 8430 23510 8470 23540
rect 8830 23510 8870 23540
rect 9230 23510 9270 23540
rect 9630 23510 9670 23540
rect 10030 23510 10070 23540
rect 10430 23510 10470 23540
rect 10830 23510 10870 23540
rect 11230 23510 11270 23540
rect 11630 23510 11670 23540
rect 12030 23510 12070 23540
rect 12430 23510 12470 23540
rect 30 23470 12960 23510
rect 30 23140 70 23470
rect 430 23140 470 23470
rect 830 23140 870 23470
rect 1230 23140 1270 23470
rect 1630 23140 1670 23470
rect 2030 23140 2070 23470
rect 2430 23140 2470 23470
rect 2830 23140 2870 23470
rect 3230 23140 3270 23470
rect 3630 23140 3670 23470
rect 4030 23140 4070 23470
rect 4430 23140 4470 23470
rect 4830 23140 4870 23470
rect 5230 23140 5270 23470
rect 5630 23140 5670 23470
rect 6030 23140 6070 23470
rect 6430 23140 6470 23470
rect 6830 23140 6870 23470
rect 7230 23140 7270 23470
rect 7630 23140 7670 23470
rect 8030 23140 8070 23470
rect 8430 23140 8470 23470
rect 8830 23140 8870 23470
rect 9230 23140 9270 23470
rect 9630 23140 9670 23470
rect 10030 23140 10070 23470
rect 10430 23140 10470 23470
rect 10830 23140 10870 23470
rect 11230 23140 11270 23470
rect 11630 23140 11670 23470
rect 12030 23140 12070 23470
rect 12430 23140 12470 23470
rect 30 23100 12960 23140
rect 30 22770 70 23100
rect 430 22770 470 23100
rect 830 22770 870 23100
rect 1230 22770 1270 23100
rect 1630 22770 1670 23100
rect 2030 22770 2070 23100
rect 2430 22770 2470 23100
rect 2830 22770 2870 23100
rect 3230 22770 3270 23100
rect 3630 22770 3670 23100
rect 4030 22770 4070 23100
rect 4430 22770 4470 23100
rect 4830 22770 4870 23100
rect 5230 22770 5270 23100
rect 5630 22770 5670 23100
rect 6030 22770 6070 23100
rect 6430 22770 6470 23100
rect 6830 22770 6870 23100
rect 7230 22770 7270 23100
rect 7630 22770 7670 23100
rect 8030 22770 8070 23100
rect 8430 22770 8470 23100
rect 8830 22770 8870 23100
rect 9230 22770 9270 23100
rect 9630 22770 9670 23100
rect 10030 22770 10070 23100
rect 10430 22770 10470 23100
rect 10830 22770 10870 23100
rect 11230 22770 11270 23100
rect 11630 22770 11670 23100
rect 12030 22770 12070 23100
rect 12430 22770 12470 23100
rect 30 22730 12960 22770
rect 30 22400 70 22730
rect 430 22400 470 22730
rect 830 22400 870 22730
rect 1230 22400 1270 22730
rect 1630 22400 1670 22730
rect 2030 22400 2070 22730
rect 2430 22400 2470 22730
rect 2830 22400 2870 22730
rect 3230 22400 3270 22730
rect 3630 22400 3670 22730
rect 4030 22400 4070 22730
rect 4430 22400 4470 22730
rect 4830 22400 4870 22730
rect 5230 22400 5270 22730
rect 5630 22400 5670 22730
rect 6030 22400 6070 22730
rect 6430 22400 6470 22730
rect 6830 22400 6870 22730
rect 7230 22400 7270 22730
rect 7630 22400 7670 22730
rect 8030 22400 8070 22730
rect 8430 22400 8470 22730
rect 8830 22400 8870 22730
rect 9230 22400 9270 22730
rect 9630 22400 9670 22730
rect 10030 22400 10070 22730
rect 10430 22400 10470 22730
rect 10830 22400 10870 22730
rect 11230 22400 11270 22730
rect 11630 22400 11670 22730
rect 12030 22400 12070 22730
rect 12430 22400 12470 22730
rect 30 22360 12960 22400
rect 30 22030 70 22360
rect 430 22030 470 22360
rect 830 22030 870 22360
rect 1230 22030 1270 22360
rect 1630 22030 1670 22360
rect 2030 22030 2070 22360
rect 2430 22030 2470 22360
rect 2830 22030 2870 22360
rect 3230 22030 3270 22360
rect 3630 22030 3670 22360
rect 4030 22030 4070 22360
rect 4430 22030 4470 22360
rect 4830 22030 4870 22360
rect 5230 22030 5270 22360
rect 5630 22030 5670 22360
rect 6030 22030 6070 22360
rect 6430 22030 6470 22360
rect 6830 22030 6870 22360
rect 7230 22030 7270 22360
rect 7630 22030 7670 22360
rect 8030 22030 8070 22360
rect 8430 22030 8470 22360
rect 8830 22030 8870 22360
rect 9230 22030 9270 22360
rect 9630 22030 9670 22360
rect 10030 22030 10070 22360
rect 10430 22030 10470 22360
rect 10830 22030 10870 22360
rect 11230 22030 11270 22360
rect 11630 22030 11670 22360
rect 12030 22030 12070 22360
rect 12430 22030 12470 22360
rect 30 21990 12960 22030
rect 30 21660 70 21990
rect 430 21660 470 21990
rect 830 21660 870 21990
rect 1230 21660 1270 21990
rect 1630 21660 1670 21990
rect 2030 21660 2070 21990
rect 2430 21660 2470 21990
rect 2830 21660 2870 21990
rect 3230 21660 3270 21990
rect 3630 21660 3670 21990
rect 4030 21660 4070 21990
rect 4430 21660 4470 21990
rect 4830 21660 4870 21990
rect 5230 21660 5270 21990
rect 5630 21660 5670 21990
rect 6030 21660 6070 21990
rect 6430 21660 6470 21990
rect 6830 21660 6870 21990
rect 7230 21660 7270 21990
rect 7630 21660 7670 21990
rect 8030 21660 8070 21990
rect 8430 21660 8470 21990
rect 8830 21660 8870 21990
rect 9230 21660 9270 21990
rect 9630 21660 9670 21990
rect 10030 21660 10070 21990
rect 10430 21660 10470 21990
rect 10830 21660 10870 21990
rect 11230 21660 11270 21990
rect 11630 21660 11670 21990
rect 12030 21660 12070 21990
rect 12430 21660 12470 21990
rect 30 21620 12960 21660
rect 30 21290 70 21620
rect 430 21290 470 21620
rect 830 21290 870 21620
rect 1230 21290 1270 21620
rect 1630 21290 1670 21620
rect 2030 21290 2070 21620
rect 2430 21290 2470 21620
rect 2830 21290 2870 21620
rect 3230 21290 3270 21620
rect 3630 21290 3670 21620
rect 4030 21290 4070 21620
rect 4430 21290 4470 21620
rect 4830 21290 4870 21620
rect 5230 21290 5270 21620
rect 5630 21290 5670 21620
rect 6030 21290 6070 21620
rect 6430 21290 6470 21620
rect 6830 21290 6870 21620
rect 7230 21290 7270 21620
rect 7630 21290 7670 21620
rect 8030 21290 8070 21620
rect 8430 21290 8470 21620
rect 8830 21290 8870 21620
rect 9230 21290 9270 21620
rect 9630 21290 9670 21620
rect 10030 21290 10070 21620
rect 10430 21290 10470 21620
rect 10830 21290 10870 21620
rect 11230 21290 11270 21620
rect 11630 21290 11670 21620
rect 12030 21290 12070 21620
rect 12430 21290 12470 21620
rect 30 21250 12960 21290
rect 30 20920 70 21250
rect 430 20920 470 21250
rect 830 20920 870 21250
rect 1230 20920 1270 21250
rect 1630 20920 1670 21250
rect 2030 20920 2070 21250
rect 2430 20920 2470 21250
rect 2830 20920 2870 21250
rect 3230 20920 3270 21250
rect 3630 20920 3670 21250
rect 4030 20920 4070 21250
rect 4430 20920 4470 21250
rect 4830 20920 4870 21250
rect 5230 20920 5270 21250
rect 5630 20920 5670 21250
rect 6030 20920 6070 21250
rect 6430 20920 6470 21250
rect 6830 20920 6870 21250
rect 7230 20920 7270 21250
rect 7630 20920 7670 21250
rect 8030 20920 8070 21250
rect 8430 20920 8470 21250
rect 8830 20920 8870 21250
rect 9230 20920 9270 21250
rect 9630 20920 9670 21250
rect 10030 20920 10070 21250
rect 10430 20920 10470 21250
rect 10830 20920 10870 21250
rect 11230 20920 11270 21250
rect 11630 20920 11670 21250
rect 12030 20920 12070 21250
rect 12430 20920 12470 21250
rect 30 20880 12960 20920
rect 30 20550 70 20880
rect 430 20550 470 20880
rect 830 20550 870 20880
rect 1230 20550 1270 20880
rect 1630 20550 1670 20880
rect 2030 20550 2070 20880
rect 2430 20550 2470 20880
rect 2830 20550 2870 20880
rect 3230 20550 3270 20880
rect 3630 20550 3670 20880
rect 4030 20550 4070 20880
rect 4430 20550 4470 20880
rect 4830 20550 4870 20880
rect 5230 20550 5270 20880
rect 5630 20550 5670 20880
rect 6030 20550 6070 20880
rect 6430 20550 6470 20880
rect 6830 20550 6870 20880
rect 7230 20550 7270 20880
rect 7630 20550 7670 20880
rect 8030 20550 8070 20880
rect 8430 20550 8470 20880
rect 8830 20550 8870 20880
rect 9230 20550 9270 20880
rect 9630 20550 9670 20880
rect 10030 20550 10070 20880
rect 10430 20550 10470 20880
rect 10830 20550 10870 20880
rect 11230 20550 11270 20880
rect 11630 20550 11670 20880
rect 12030 20550 12070 20880
rect 12430 20550 12470 20880
rect 30 20510 12960 20550
rect 30 20180 70 20510
rect 430 20180 470 20510
rect 830 20180 870 20510
rect 1230 20180 1270 20510
rect 1630 20180 1670 20510
rect 2030 20180 2070 20510
rect 2430 20180 2470 20510
rect 2830 20180 2870 20510
rect 3230 20180 3270 20510
rect 3630 20180 3670 20510
rect 4030 20180 4070 20510
rect 4430 20180 4470 20510
rect 4830 20180 4870 20510
rect 5230 20180 5270 20510
rect 5630 20180 5670 20510
rect 6030 20180 6070 20510
rect 6430 20180 6470 20510
rect 6830 20180 6870 20510
rect 7230 20180 7270 20510
rect 7630 20180 7670 20510
rect 8030 20180 8070 20510
rect 8430 20180 8470 20510
rect 8830 20180 8870 20510
rect 9230 20180 9270 20510
rect 9630 20180 9670 20510
rect 10030 20180 10070 20510
rect 10430 20180 10470 20510
rect 10830 20180 10870 20510
rect 11230 20180 11270 20510
rect 11630 20180 11670 20510
rect 12030 20180 12070 20510
rect 12430 20180 12470 20510
rect 30 20140 12960 20180
rect 30 19810 70 20140
rect 430 19810 470 20140
rect 830 19810 870 20140
rect 1230 19810 1270 20140
rect 1630 19810 1670 20140
rect 2030 19810 2070 20140
rect 2430 19810 2470 20140
rect 2830 19810 2870 20140
rect 3230 19810 3270 20140
rect 3630 19810 3670 20140
rect 4030 19810 4070 20140
rect 4430 19810 4470 20140
rect 4830 19810 4870 20140
rect 5230 19810 5270 20140
rect 5630 19810 5670 20140
rect 6030 19810 6070 20140
rect 6430 19810 6470 20140
rect 6830 19810 6870 20140
rect 7230 19810 7270 20140
rect 7630 19810 7670 20140
rect 8030 19810 8070 20140
rect 8430 19810 8470 20140
rect 8830 19810 8870 20140
rect 9230 19810 9270 20140
rect 9630 19810 9670 20140
rect 10030 19810 10070 20140
rect 10430 19810 10470 20140
rect 10830 19810 10870 20140
rect 11230 19810 11270 20140
rect 11630 19810 11670 20140
rect 12030 19810 12070 20140
rect 12430 19810 12470 20140
rect 30 19770 12960 19810
rect 30 19440 70 19770
rect 430 19440 470 19770
rect 830 19440 870 19770
rect 1230 19440 1270 19770
rect 1630 19440 1670 19770
rect 2030 19440 2070 19770
rect 2430 19440 2470 19770
rect 2830 19440 2870 19770
rect 3230 19740 3270 19770
rect 3630 19740 3670 19770
rect 4030 19740 4070 19770
rect 4430 19740 4470 19770
rect 4830 19740 4870 19770
rect 5230 19740 5270 19770
rect 5630 19740 5670 19770
rect 6030 19740 6070 19770
rect 6430 19740 6470 19770
rect 6830 19740 6870 19770
rect 7230 19740 7270 19770
rect 7630 19740 7670 19770
rect 8030 19740 8070 19770
rect 8430 19740 8470 19770
rect 8830 19740 8870 19770
rect 9230 19740 9270 19770
rect 9630 19740 9670 19770
rect 10030 19740 10070 19770
rect 10430 19740 10470 19770
rect 10830 19740 10870 19770
rect 11230 19740 11270 19770
rect 11630 19740 11670 19770
rect 12030 19740 12070 19770
rect 12430 19740 12470 19770
rect 30 19400 3140 19440
rect 30 19070 70 19400
rect 430 19070 470 19400
rect 830 19070 870 19400
rect 1230 19070 1270 19400
rect 1630 19070 1670 19400
rect 2030 19070 2070 19400
rect 2430 19070 2470 19400
rect 2830 19070 2870 19400
rect 3230 19070 3270 19470
rect 3630 19440 3670 19470
rect 4030 19440 4070 19470
rect 4430 19440 4470 19470
rect 4830 19440 4870 19470
rect 5230 19440 5270 19470
rect 5630 19440 5670 19470
rect 6030 19440 6070 19470
rect 6430 19440 6470 19470
rect 6830 19440 6870 19470
rect 7230 19440 7270 19470
rect 7630 19440 7670 19470
rect 8030 19440 8070 19470
rect 8430 19440 8470 19470
rect 8830 19440 8870 19470
rect 9230 19440 9270 19470
rect 9630 19440 9670 19470
rect 10030 19440 10070 19470
rect 10430 19440 10470 19470
rect 10830 19440 10870 19470
rect 11230 19440 11270 19470
rect 11630 19440 11670 19470
rect 12030 19440 12070 19470
rect 12430 19440 12470 19470
rect 3480 19400 12500 19440
rect 12690 19400 12960 19440
rect 3630 19070 3670 19400
rect 4030 19070 4070 19400
rect 4430 19070 4470 19400
rect 4830 19070 4870 19400
rect 5230 19070 5270 19400
rect 5630 19070 5670 19400
rect 6030 19070 6070 19400
rect 6430 19070 6470 19400
rect 6830 19070 6870 19400
rect 7230 19070 7270 19400
rect 7630 19070 7670 19400
rect 8030 19070 8070 19400
rect 8430 19070 8470 19400
rect 8830 19070 8870 19400
rect 9230 19070 9270 19400
rect 9630 19070 9670 19400
rect 10030 19070 10070 19400
rect 10430 19070 10470 19400
rect 10830 19070 10870 19400
rect 11230 19070 11270 19400
rect 11630 19070 11670 19400
rect 12030 19070 12070 19400
rect 12430 19070 12470 19400
rect 30 19030 3140 19070
rect 3230 19030 12960 19070
rect 30 18700 70 19030
rect 430 18700 470 19030
rect 830 18700 870 19030
rect 1230 18700 1270 19030
rect 1630 18700 1670 19030
rect 2030 18700 2070 19030
rect 2430 18700 2470 19030
rect 2830 18700 2870 19030
rect 3230 18700 3270 19030
rect 3630 18700 3670 19030
rect 4030 18700 4070 19030
rect 4430 18700 4470 19030
rect 4830 18700 4870 19030
rect 5230 18700 5270 19030
rect 5630 18700 5670 19030
rect 6030 18700 6070 19030
rect 6430 18700 6470 19030
rect 6830 18700 6870 19030
rect 7230 18700 7270 19030
rect 7630 18700 7670 19030
rect 8030 18700 8070 19030
rect 8430 18700 8470 19030
rect 8830 18700 8870 19030
rect 9230 18700 9270 19030
rect 9630 18700 9670 19030
rect 10030 18700 10070 19030
rect 10430 18700 10470 19030
rect 10830 18700 10870 19030
rect 11230 18700 11270 19030
rect 11630 18700 11670 19030
rect 12030 18700 12070 19030
rect 12430 18700 12470 19030
rect 30 18660 3140 18700
rect 3230 18660 12960 18700
rect 30 18330 70 18660
rect 430 18330 470 18660
rect 830 18330 870 18660
rect 1230 18330 1270 18660
rect 1630 18330 1670 18660
rect 2030 18330 2070 18660
rect 2430 18330 2470 18660
rect 2830 18330 2870 18660
rect 3230 18330 3270 18660
rect 3630 18330 3670 18660
rect 4030 18330 4070 18660
rect 4430 18330 4470 18660
rect 4830 18330 4870 18660
rect 5230 18330 5270 18660
rect 5630 18330 5670 18660
rect 6030 18330 6070 18660
rect 6430 18330 6470 18660
rect 6830 18330 6870 18660
rect 7230 18330 7270 18660
rect 7630 18330 7670 18660
rect 8030 18330 8070 18660
rect 8430 18330 8470 18660
rect 8830 18330 8870 18660
rect 9230 18330 9270 18660
rect 9630 18330 9670 18660
rect 10030 18330 10070 18660
rect 10430 18330 10470 18660
rect 10830 18330 10870 18660
rect 11230 18330 11270 18660
rect 11630 18330 11670 18660
rect 12030 18330 12070 18660
rect 12430 18330 12470 18660
rect 30 18290 3140 18330
rect 3230 18290 12960 18330
rect 30 17960 70 18290
rect 430 17960 470 18290
rect 830 17960 870 18290
rect 1230 17960 1270 18290
rect 1630 17960 1670 18290
rect 2030 17960 2070 18290
rect 2430 17960 2470 18290
rect 2830 17960 2870 18290
rect 3230 17960 3270 18290
rect 3630 17960 3670 18290
rect 4030 17960 4070 18290
rect 4430 17960 4470 18290
rect 4830 17960 4870 18290
rect 5230 17960 5270 18290
rect 5630 17960 5670 18290
rect 6030 17960 6070 18290
rect 6430 17960 6470 18290
rect 6830 17960 6870 18290
rect 7230 17960 7270 18290
rect 7630 17960 7670 18290
rect 8030 17960 8070 18290
rect 8430 17960 8470 18290
rect 8830 17960 8870 18290
rect 9230 17960 9270 18290
rect 9630 17960 9670 18290
rect 10030 17960 10070 18290
rect 10430 17960 10470 18290
rect 10830 17960 10870 18290
rect 11230 17960 11270 18290
rect 11630 17960 11670 18290
rect 12030 17960 12070 18290
rect 12430 17960 12470 18290
rect 30 17920 3140 17960
rect 3230 17920 12960 17960
rect 30 17590 70 17920
rect 430 17590 470 17920
rect 830 17590 870 17920
rect 1230 17590 1270 17920
rect 1630 17590 1670 17920
rect 2030 17590 2070 17920
rect 2430 17590 2470 17920
rect 2830 17590 2870 17920
rect 3230 17590 3270 17920
rect 3630 17590 3670 17920
rect 4030 17590 4070 17920
rect 4430 17590 4470 17920
rect 4830 17590 4870 17920
rect 5230 17590 5270 17920
rect 5630 17590 5670 17920
rect 6030 17590 6070 17920
rect 6430 17590 6470 17920
rect 6830 17590 6870 17920
rect 7230 17590 7270 17920
rect 7630 17590 7670 17920
rect 8030 17590 8070 17920
rect 8430 17590 8470 17920
rect 8830 17590 8870 17920
rect 9230 17590 9270 17920
rect 9630 17590 9670 17920
rect 10030 17590 10070 17920
rect 10430 17590 10470 17920
rect 10830 17590 10870 17920
rect 11230 17590 11270 17920
rect 11630 17590 11670 17920
rect 12030 17590 12070 17920
rect 12430 17590 12470 17920
rect 30 17550 3140 17590
rect 3230 17550 12960 17590
rect 30 17220 70 17550
rect 430 17220 470 17550
rect 830 17220 870 17550
rect 1230 17220 1270 17550
rect 1630 17220 1670 17550
rect 2030 17220 2070 17550
rect 2430 17220 2470 17550
rect 2830 17220 2870 17550
rect 3230 17220 3270 17550
rect 3630 17220 3670 17550
rect 4030 17220 4070 17550
rect 4430 17220 4470 17550
rect 4830 17220 4870 17550
rect 5230 17220 5270 17550
rect 5630 17220 5670 17550
rect 6030 17520 6070 17550
rect 6430 17520 6470 17550
rect 6830 17520 6870 17550
rect 7230 17520 7270 17550
rect 7630 17520 7670 17550
rect 8030 17520 8070 17550
rect 8430 17520 8470 17550
rect 8830 17520 8870 17550
rect 9230 17520 9270 17550
rect 9630 17520 9670 17550
rect 10030 17520 10070 17550
rect 10430 17520 10470 17550
rect 10830 17520 10870 17550
rect 11230 17520 11270 17550
rect 11630 17520 11670 17550
rect 12030 17520 12070 17550
rect 12430 17520 12470 17550
rect 6430 17220 6470 17250
rect 6830 17220 6870 17250
rect 7230 17220 7270 17250
rect 8030 17220 8070 17250
rect 8430 17220 8470 17250
rect 8830 17220 8870 17250
rect 9230 17220 9270 17250
rect 9630 17220 9670 17250
rect 10030 17220 10070 17250
rect 10430 17220 10470 17250
rect 10830 17220 10870 17250
rect 11230 17220 11270 17250
rect 11630 17220 11670 17250
rect 12030 17220 12070 17250
rect 12430 17220 12470 17250
rect 30 17180 3140 17220
rect 3230 17180 5940 17220
rect 6030 17180 12960 17220
rect 30 16850 70 17180
rect 430 16850 470 17180
rect 830 16850 870 17180
rect 1230 16850 1270 17180
rect 1630 16850 1670 17180
rect 2030 16850 2070 17180
rect 2430 16850 2470 17180
rect 2830 16850 2870 17180
rect 3230 16850 3270 17180
rect 3630 16850 3670 17180
rect 4030 16850 4070 17180
rect 4430 16850 4470 17180
rect 4830 16850 4870 17180
rect 5230 16850 5270 17180
rect 5630 16850 5670 17180
rect 6030 16850 6070 17180
rect 6430 16850 6470 17180
rect 6830 16850 6870 17180
rect 7230 16850 7270 17180
rect 7630 16850 7670 17180
rect 8030 16850 8070 17180
rect 8430 16850 8470 17180
rect 8830 16850 8870 17180
rect 9230 16850 9270 17180
rect 9630 16850 9670 17180
rect 10030 16850 10070 17180
rect 10430 16850 10470 17180
rect 10830 16850 10870 17180
rect 11230 16850 11270 17180
rect 11630 16850 11670 17180
rect 12030 16850 12070 17180
rect 12430 16850 12470 17180
rect 30 16810 3140 16850
rect 3230 16810 5940 16850
rect 6030 16810 12960 16850
rect 30 16480 70 16810
rect 430 16480 470 16810
rect 830 16480 870 16810
rect 1230 16480 1270 16810
rect 1630 16480 1670 16810
rect 2030 16480 2070 16810
rect 2430 16480 2470 16810
rect 2830 16480 2870 16810
rect 3230 16480 3270 16810
rect 3630 16480 3670 16810
rect 4030 16480 4070 16810
rect 4430 16480 4470 16810
rect 4830 16480 4870 16810
rect 5230 16480 5270 16810
rect 5630 16480 5670 16810
rect 6030 16480 6070 16810
rect 6430 16480 6470 16810
rect 6830 16480 6870 16810
rect 7230 16480 7270 16810
rect 7630 16480 7670 16810
rect 8030 16480 8070 16810
rect 8430 16480 8470 16810
rect 8830 16480 8870 16810
rect 9230 16480 9270 16810
rect 9630 16480 9670 16810
rect 10030 16480 10070 16810
rect 10430 16480 10470 16810
rect 10830 16480 10870 16810
rect 11230 16480 11270 16810
rect 11630 16480 11670 16810
rect 12030 16480 12070 16810
rect 12430 16480 12470 16810
rect 30 16440 3140 16480
rect 3230 16440 5940 16480
rect 6030 16440 12960 16480
rect 30 16110 70 16440
rect 430 16110 470 16440
rect 830 16110 870 16440
rect 1230 16110 1270 16440
rect 1630 16110 1670 16440
rect 2030 16110 2070 16440
rect 2430 16110 2470 16440
rect 2830 16110 2870 16440
rect 3230 16110 3270 16440
rect 3630 16110 3670 16440
rect 4030 16110 4070 16440
rect 4430 16110 4470 16440
rect 4830 16110 4870 16440
rect 5230 16110 5270 16440
rect 5630 16110 5670 16440
rect 6030 16110 6070 16440
rect 6430 16110 6470 16440
rect 6830 16110 6870 16440
rect 7230 16110 7270 16440
rect 7630 16110 7670 16440
rect 8030 16110 8070 16440
rect 8430 16110 8470 16440
rect 8830 16110 8870 16440
rect 9230 16110 9270 16440
rect 9630 16110 9670 16440
rect 10030 16110 10070 16440
rect 10430 16110 10470 16440
rect 10830 16110 10870 16440
rect 11230 16110 11270 16440
rect 11630 16110 11670 16440
rect 12030 16110 12070 16440
rect 12430 16110 12470 16440
rect 30 16070 3140 16110
rect 3230 16070 5940 16110
rect 6030 16070 12960 16110
rect 30 15740 70 16070
rect 430 15740 470 16070
rect 830 15740 870 16070
rect 1230 15740 1270 16070
rect 1630 15740 1670 16070
rect 2030 15740 2070 16070
rect 2430 15740 2470 16070
rect 2830 15740 2870 16070
rect 3230 15740 3270 16070
rect 3630 15740 3670 16070
rect 4030 15740 4070 16070
rect 4430 15740 4470 16070
rect 4830 15740 4870 16070
rect 5230 15740 5270 16070
rect 5630 15740 5670 16070
rect 6030 15740 6070 16070
rect 6430 15740 6470 16070
rect 6830 15740 6870 16070
rect 7230 15740 7270 16070
rect 7630 15740 7670 16070
rect 8030 15740 8070 16070
rect 8430 15740 8470 16070
rect 8830 15740 8870 16070
rect 9230 15740 9270 16070
rect 9630 15740 9670 16070
rect 10030 15740 10070 16070
rect 10430 15740 10470 16070
rect 10830 15740 10870 16070
rect 11230 15740 11270 16070
rect 11630 15740 11670 16070
rect 12030 15740 12070 16070
rect 12430 15740 12470 16070
rect 30 15700 3140 15740
rect 3230 15700 5940 15740
rect 6030 15700 12960 15740
rect 30 15370 70 15700
rect 430 15370 470 15700
rect 830 15370 870 15700
rect 1230 15370 1270 15700
rect 1630 15370 1670 15700
rect 2030 15370 2070 15700
rect 2430 15370 2470 15700
rect 2830 15370 2870 15700
rect 3230 15370 3270 15700
rect 3630 15370 3670 15700
rect 4030 15370 4070 15700
rect 4430 15370 4470 15700
rect 4830 15370 4870 15700
rect 5230 15370 5270 15700
rect 5630 15370 5670 15700
rect 6030 15370 6070 15700
rect 6430 15370 6470 15700
rect 6830 15370 6870 15700
rect 7230 15370 7270 15700
rect 7630 15370 7670 15700
rect 8030 15670 8070 15700
rect 8430 15670 8470 15700
rect 8830 15670 8870 15700
rect 9230 15670 9270 15700
rect 9630 15670 9670 15700
rect 10030 15670 10070 15700
rect 10430 15670 10470 15700
rect 10830 15670 10870 15700
rect 11230 15670 11270 15700
rect 11630 15670 11670 15700
rect 12030 15670 12070 15700
rect 12430 15670 12470 15700
rect 30 15330 3140 15370
rect 3230 15330 5940 15370
rect 6030 15330 7850 15370
rect 8030 15330 12960 15370
rect 30 15000 70 15330
rect 430 15000 470 15330
rect 830 15000 870 15330
rect 1230 15000 1270 15330
rect 1630 15000 1670 15330
rect 2030 15000 2070 15330
rect 2430 15000 2470 15330
rect 2830 15000 2870 15330
rect 3230 15000 3270 15330
rect 3630 15000 3670 15330
rect 4030 15000 4070 15330
rect 4430 15000 4470 15330
rect 4830 15000 4870 15330
rect 5230 15000 5270 15330
rect 5630 15000 5670 15330
rect 6030 15000 6070 15330
rect 6430 15000 6470 15330
rect 6830 15000 6870 15330
rect 7230 15000 7270 15330
rect 7630 15000 7670 15330
rect 8030 15000 8070 15330
rect 8430 15000 8470 15330
rect 8830 15000 8870 15300
rect 9230 15000 9270 15330
rect 9630 15000 9670 15330
rect 10030 15000 10070 15330
rect 10430 15000 10470 15330
rect 10830 15000 10870 15330
rect 11230 15000 11270 15330
rect 11630 15000 11670 15330
rect 12030 15000 12070 15330
rect 12430 15000 12470 15330
rect 30 14960 2930 15000
rect 3230 14960 5940 15000
rect 6030 14960 7810 15000
rect 8030 14960 12960 15000
rect 30 14630 70 14960
rect 430 14630 470 14960
rect 830 14630 870 14960
rect 1230 14630 1270 14960
rect 1630 14630 1670 14960
rect 2030 14630 2070 14960
rect 2430 14630 2470 14960
rect 3230 14630 3270 14960
rect 3630 14630 3670 14960
rect 4030 14630 4070 14960
rect 4430 14630 4470 14960
rect 4830 14630 4870 14960
rect 5230 14630 5270 14960
rect 5630 14630 5670 14960
rect 6030 14630 6070 14960
rect 6430 14630 6470 14960
rect 6830 14630 6870 14960
rect 7230 14630 7270 14960
rect 8030 14630 8070 14960
rect 8430 14630 8470 14960
rect 8830 14630 8870 14960
rect 9230 14630 9270 14960
rect 9630 14630 9670 14960
rect 10030 14630 10070 14960
rect 10430 14630 10470 14960
rect 10830 14630 10870 14960
rect 11230 14630 11270 14960
rect 11630 14630 11670 14960
rect 12030 14630 12070 14960
rect 12430 14630 12470 14960
rect 30 14590 2740 14630
rect 30 14260 70 14590
rect 430 14260 470 14590
rect 830 14260 870 14590
rect 1230 14260 1270 14590
rect 1630 14260 1670 14590
rect 2030 14260 2070 14590
rect 2430 14260 2470 14590
rect 30 14220 2740 14260
rect 30 13890 70 14220
rect 430 13890 470 14220
rect 830 13890 870 14220
rect 1230 13890 1270 14220
rect 1630 13890 1670 14220
rect 2030 13890 2070 14220
rect 2430 13890 2470 14220
rect 30 13850 2740 13890
rect 30 13520 70 13850
rect 430 13520 470 13850
rect 830 13520 870 13850
rect 1230 13520 1270 13850
rect 1630 13520 1670 13850
rect 2030 13520 2070 13850
rect 2430 13520 2470 13850
rect 30 13480 2740 13520
rect 30 13150 70 13480
rect 430 13150 470 13480
rect 830 13150 870 13480
rect 1230 13150 1270 13480
rect 1630 13150 1670 13480
rect 2030 13150 2070 13480
rect 2430 13150 2470 13480
rect 30 13110 2740 13150
rect 30 12780 70 13110
rect 430 12780 470 13110
rect 830 12780 870 13110
rect 1230 12780 1270 13110
rect 1630 12780 1670 13110
rect 2030 12780 2070 13110
rect 2430 12780 2470 13110
rect 30 12740 2740 12780
rect 30 12410 70 12740
rect 430 12410 470 12740
rect 830 12410 870 12740
rect 1230 12410 1270 12740
rect 1630 12410 1670 12740
rect 2030 12410 2070 12740
rect 2430 12410 2470 12740
rect 30 12370 2740 12410
rect 30 12040 70 12370
rect 430 12040 470 12370
rect 830 12040 870 12370
rect 1230 12040 1270 12370
rect 1630 12040 1670 12370
rect 2030 12040 2070 12370
rect 2430 12040 2470 12370
rect 2830 12040 2870 14600
rect 3080 14590 5940 14630
rect 6030 14590 7540 14630
rect 3230 14260 3270 14590
rect 3630 14260 3670 14590
rect 4030 14260 4070 14590
rect 4430 14260 4470 14590
rect 4830 14260 4870 14590
rect 5230 14260 5270 14590
rect 5630 14260 5670 14590
rect 6030 14260 6070 14590
rect 6430 14260 6470 14590
rect 6830 14260 6870 14590
rect 7230 14260 7270 14590
rect 3090 14220 5940 14260
rect 6030 14220 7540 14260
rect 3230 13890 3270 14220
rect 3630 13890 3670 14220
rect 4030 13890 4070 14220
rect 4430 13890 4470 14220
rect 4830 13890 4870 14220
rect 5230 13890 5270 14220
rect 5630 13890 5670 14220
rect 6030 13890 6070 14220
rect 6430 13890 6470 14220
rect 6830 13890 6870 14220
rect 7230 13890 7270 14220
rect 3080 13850 5940 13890
rect 6030 13850 7540 13890
rect 3230 13520 3270 13850
rect 3630 13520 3670 13850
rect 4030 13520 4070 13850
rect 4430 13520 4470 13850
rect 4830 13520 4870 13850
rect 5230 13520 5270 13850
rect 5630 13520 5670 13850
rect 6030 13520 6070 13850
rect 6430 13520 6470 13850
rect 6830 13520 6870 13850
rect 7230 13520 7270 13850
rect 3100 13480 5940 13520
rect 6030 13480 7540 13520
rect 3230 13150 3270 13480
rect 3630 13150 3670 13480
rect 4030 13150 4070 13480
rect 4430 13150 4470 13480
rect 4830 13150 4870 13480
rect 5230 13150 5270 13480
rect 5630 13150 5670 13480
rect 6030 13150 6070 13480
rect 6430 13150 6470 13480
rect 6830 13150 6870 13480
rect 7230 13150 7270 13480
rect 3120 13110 5940 13150
rect 6030 13110 7540 13150
rect 3230 12780 3270 13110
rect 3630 12780 3670 13110
rect 4030 12780 4070 13110
rect 4430 12780 4470 13110
rect 4830 12780 4870 13110
rect 5230 12780 5270 13110
rect 5630 12780 5670 13110
rect 6030 12780 6070 13110
rect 6430 12780 6470 13110
rect 6830 12780 6870 13110
rect 7230 12780 7270 13110
rect 3120 12740 5940 12780
rect 6030 12740 7540 12780
rect 3230 12410 3270 12740
rect 3630 12410 3670 12740
rect 4030 12410 4070 12740
rect 4430 12410 4470 12740
rect 4830 12410 4870 12740
rect 5230 12410 5270 12740
rect 5630 12460 5670 12740
rect 6030 12410 6070 12740
rect 6430 12410 6470 12740
rect 6830 12410 6870 12740
rect 7230 12410 7270 12740
rect 3110 12370 5940 12410
rect 6030 12370 7540 12410
rect 3230 12040 3270 12370
rect 3630 12040 3670 12370
rect 4030 12040 4070 12370
rect 4430 12040 4470 12370
rect 4830 12040 4870 12370
rect 5230 12040 5270 12370
rect 6030 12040 6070 12370
rect 6430 12040 6470 12370
rect 6830 12040 6870 12370
rect 7230 12040 7270 12370
rect 30 12000 2740 12040
rect 2830 12000 5440 12040
rect 5870 12000 7540 12040
rect 30 11670 70 12000
rect 430 11670 470 12000
rect 830 11670 870 12000
rect 1230 11670 1270 12000
rect 1630 11670 1670 12000
rect 2030 11670 2070 12000
rect 2430 11670 2470 12000
rect 2830 11670 2870 12000
rect 3230 11670 3270 12000
rect 3630 11670 3670 12000
rect 4030 11670 4070 12000
rect 4430 11670 4470 12000
rect 4830 11670 4870 12000
rect 5230 11670 5270 12000
rect 5630 11670 5670 12000
rect 6030 11670 6070 12000
rect 6430 11670 6470 12000
rect 6830 11670 6870 12000
rect 7230 11670 7270 12000
rect 30 11630 2740 11670
rect 2830 11630 5430 11670
rect 5820 11630 7540 11670
rect 30 11300 70 11630
rect 430 11300 470 11630
rect 830 11300 870 11630
rect 1230 11300 1270 11630
rect 1630 11300 1670 11630
rect 2030 11300 2070 11630
rect 2430 11300 2470 11630
rect 30 11260 2740 11300
rect 30 10930 70 11260
rect 430 10930 470 11260
rect 830 10930 870 11260
rect 1230 10930 1270 11260
rect 1630 10930 1670 11260
rect 2030 10930 2070 11260
rect 2430 10930 2470 11260
rect 30 10890 2740 10930
rect 30 10560 70 10890
rect 430 10560 470 10890
rect 830 10560 870 10890
rect 1230 10560 1270 10890
rect 1630 10560 1670 10890
rect 2030 10560 2070 10890
rect 2430 10560 2470 10890
rect 30 10520 2740 10560
rect 30 10190 70 10520
rect 430 10190 470 10520
rect 830 10190 870 10520
rect 1230 10190 1270 10520
rect 1630 10190 1670 10520
rect 2030 10190 2070 10520
rect 2430 10190 2470 10520
rect 30 10150 2740 10190
rect 30 9820 70 10150
rect 430 9820 470 10150
rect 830 9820 870 10150
rect 1230 9820 1270 10150
rect 1630 9820 1670 10150
rect 2030 9820 2070 10150
rect 2430 9820 2470 10150
rect 30 9780 2740 9820
rect 30 9450 70 9780
rect 430 9450 470 9780
rect 830 9450 870 9780
rect 1230 9450 1270 9780
rect 1630 9450 1670 9780
rect 2030 9450 2070 9780
rect 2430 9450 2470 9780
rect 30 9410 2740 9450
rect 30 8710 70 9410
rect 430 9080 470 9410
rect 830 9080 870 9410
rect 1230 9080 1270 9410
rect 1630 9080 1670 9410
rect 2030 9080 2070 9410
rect 2430 9080 2470 9410
rect 310 9040 2540 9080
rect 2830 9060 2870 11630
rect 3230 11300 3270 11630
rect 3630 11300 3670 11630
rect 4030 11300 4070 11630
rect 4430 11300 4470 11630
rect 4830 11300 4870 11630
rect 5230 11300 5270 11630
rect 6030 11300 6070 11630
rect 6430 11300 6470 11630
rect 6830 11300 6870 11630
rect 7230 11300 7270 11630
rect 3090 11260 5940 11300
rect 6030 11260 7540 11300
rect 3230 10930 3270 11260
rect 3630 10930 3670 11260
rect 4030 10930 4070 11260
rect 4430 10930 4470 11260
rect 4830 10930 4870 11260
rect 5230 10930 5270 11260
rect 5630 10930 5670 11260
rect 6030 10930 6070 11260
rect 6430 10930 6470 11260
rect 6830 10930 6870 11260
rect 7230 10930 7270 11260
rect 3090 10890 5940 10930
rect 6030 10890 7540 10930
rect 3230 10560 3270 10890
rect 3630 10560 3670 10890
rect 4030 10560 4070 10890
rect 4430 10560 4470 10890
rect 4830 10560 4870 10890
rect 5230 10560 5270 10890
rect 5630 10560 5670 10890
rect 6030 10560 6070 10890
rect 6430 10560 6470 10890
rect 6830 10560 6870 10890
rect 7230 10560 7270 10890
rect 3100 10520 5940 10560
rect 6030 10520 7540 10560
rect 3230 10190 3270 10520
rect 3630 10190 3670 10520
rect 4030 10190 4070 10520
rect 4430 10190 4470 10520
rect 4830 10190 4870 10520
rect 5230 10190 5270 10520
rect 5630 10190 5670 10520
rect 6030 10190 6070 10520
rect 6430 10190 6470 10520
rect 6830 10190 6870 10520
rect 7230 10190 7270 10520
rect 3100 10150 5940 10190
rect 6030 10150 7540 10190
rect 3230 9820 3270 10150
rect 3630 9820 3670 10150
rect 4030 9820 4070 10150
rect 4430 9820 4470 10150
rect 4830 9820 4870 10150
rect 5230 9820 5270 10150
rect 5630 9820 5670 10150
rect 6030 9820 6070 10150
rect 6430 9820 6470 10150
rect 6830 9820 6870 10150
rect 7230 9820 7270 10150
rect 3110 9780 5940 9820
rect 6030 9780 7540 9820
rect 3230 9450 3270 9780
rect 3630 9450 3670 9780
rect 4030 9450 4070 9780
rect 4430 9450 4470 9780
rect 4830 9450 4870 9780
rect 5230 9450 5270 9780
rect 5630 9450 5670 9780
rect 6030 9450 6070 9780
rect 6430 9450 6470 9780
rect 6830 9450 6870 9780
rect 7230 9450 7270 9780
rect 3100 9410 5940 9450
rect 6030 9410 7540 9450
rect 3230 9080 3270 9410
rect 3630 9080 3670 9410
rect 4030 9080 4070 9410
rect 4430 9080 4470 9410
rect 4830 9080 4870 9410
rect 5230 9080 5270 9410
rect 5630 9080 5670 9410
rect 3110 9040 5940 9080
rect 430 8710 470 9040
rect 830 8710 870 9040
rect 1230 8710 1270 9040
rect 1630 8710 1670 9040
rect 2030 8710 2070 9040
rect 2430 8710 2470 9040
rect 2830 8710 2870 8720
rect 3230 8710 3270 9040
rect 3630 8710 3670 9040
rect 4030 8710 4070 9040
rect 4430 8710 4470 9040
rect 4830 8710 4870 9040
rect 5230 8710 5270 9040
rect 5630 8710 5670 9040
rect 6030 8710 6070 9410
rect 6430 9080 6470 9410
rect 6830 9080 6870 9410
rect 7230 9080 7270 9410
rect 6170 9040 7410 9080
rect 7630 9040 7670 14600
rect 7840 14590 12960 14630
rect 8030 14260 8070 14590
rect 7840 14220 8120 14260
rect 8030 13890 8070 14220
rect 7840 13850 8120 13890
rect 8030 13520 8070 13850
rect 7840 13480 8120 13520
rect 8030 13150 8070 13480
rect 7840 13110 8120 13150
rect 8030 12780 8070 13110
rect 7840 12740 8120 12780
rect 8030 12410 8070 12740
rect 7840 12370 8120 12410
rect 8030 12040 8070 12370
rect 7840 12000 8120 12040
rect 8030 11670 8070 12000
rect 7840 11630 8120 11670
rect 8030 11300 8070 11630
rect 7840 11260 8120 11300
rect 8030 10930 8070 11260
rect 7840 10890 8120 10930
rect 8030 10560 8070 10890
rect 7840 10520 8120 10560
rect 8030 10190 8070 10520
rect 7840 10150 8120 10190
rect 8030 9820 8070 10150
rect 7840 9780 8120 9820
rect 8030 9450 8070 9780
rect 7840 9410 8120 9450
rect 8030 9080 8070 9410
rect 8430 9080 8470 14590
rect 8830 12350 8870 14590
rect 9460 14220 9740 14260
rect 9860 14220 10140 14260
rect 10260 14220 10540 14260
rect 10660 14220 10940 14260
rect 11060 14220 11340 14260
rect 11460 14220 11740 14260
rect 11860 14220 12140 14260
rect 12260 14220 12540 14260
rect 12690 14220 12960 14260
rect 9230 13870 9270 14210
rect 9630 13890 9670 14220
rect 10030 13890 10070 14220
rect 10430 13890 10470 14220
rect 10830 13890 10870 14220
rect 11230 13890 11270 14220
rect 11630 13890 11670 14220
rect 12030 13890 12070 14220
rect 12430 13890 12470 14220
rect 9460 13850 9740 13890
rect 9900 13850 12960 13890
rect 9230 13500 9270 13840
rect 9630 13520 9670 13850
rect 10030 13520 10070 13850
rect 10430 13840 10470 13850
rect 10830 13840 10870 13850
rect 11230 13840 11270 13850
rect 11630 13840 11670 13850
rect 12030 13840 12070 13850
rect 12430 13840 12470 13850
rect 9460 13480 9740 13520
rect 9880 13480 10080 13520
rect 9230 13130 9270 13470
rect 9630 13150 9670 13480
rect 10030 13150 10070 13480
rect 9460 13110 9740 13150
rect 9890 13110 10090 13150
rect 9230 12760 9270 13100
rect 9630 12780 9670 13110
rect 10030 12780 10070 13110
rect 9460 12740 9740 12780
rect 9890 12740 10090 12780
rect 9230 12390 9270 12730
rect 9630 12410 9670 12740
rect 10430 12410 10470 13550
rect 10720 13480 10850 13520
rect 11120 13480 12650 13520
rect 12690 13480 12960 13520
rect 10830 13150 10870 13480
rect 10720 13110 10870 13150
rect 10830 12780 10870 13110
rect 10720 12740 10870 12780
rect 10830 12410 10870 12740
rect 9460 12370 9740 12410
rect 9230 12040 9270 12360
rect 9630 12040 9670 12370
rect 9120 12000 9300 12040
rect 9460 12000 9740 12040
rect 8830 11680 8870 12000
rect 9230 11670 9270 11990
rect 9630 11670 9670 12000
rect 9130 11630 9310 11670
rect 9460 11630 9740 11670
rect 8830 9080 8870 11290
rect 9230 11280 9270 11620
rect 9630 11300 9670 11630
rect 10030 11300 10070 12380
rect 10310 12370 10470 12410
rect 10720 12370 10870 12410
rect 10430 12040 10470 12370
rect 10830 12040 10870 12370
rect 10310 12000 10470 12040
rect 10710 12000 10870 12040
rect 10430 11670 10470 12000
rect 10830 11670 10870 12000
rect 10310 11630 10470 11670
rect 10730 11630 10870 11670
rect 10430 11300 10470 11630
rect 10830 11300 10870 11630
rect 9460 11260 9740 11300
rect 10310 11260 10470 11300
rect 10720 11260 10870 11300
rect 9230 10910 9270 11250
rect 9630 10930 9670 11260
rect 10030 10930 10070 10940
rect 9460 10890 9740 10930
rect 9900 10890 10080 10930
rect 9230 10540 9270 10880
rect 9630 10560 9670 10890
rect 10030 10560 10070 10890
rect 9490 10520 10100 10560
rect 9230 10170 9270 10510
rect 9630 10190 9670 10520
rect 10030 10190 10070 10520
rect 9520 10150 10090 10190
rect 10430 10160 10470 11260
rect 10830 10930 10870 11260
rect 10730 10890 10870 10930
rect 10830 10560 10870 10890
rect 11230 10560 11270 13150
rect 11510 13110 12960 13150
rect 11630 10900 11670 12760
rect 11890 12740 13390 12780
rect 12340 12370 13390 12410
rect 12740 12000 13390 12040
rect 12030 11740 12070 11930
rect 12740 11630 13390 11670
rect 12030 11370 12070 11560
rect 12340 11260 13390 11300
rect 12340 10890 13390 10930
rect 12030 10630 12070 10820
rect 12430 10630 12470 10820
rect 10700 10520 10870 10560
rect 11500 10520 12090 10560
rect 12340 10520 12440 10560
rect 12690 10520 12960 10560
rect 10830 10190 10870 10520
rect 10710 10150 13390 10190
rect 9230 9800 9270 10140
rect 9630 9890 9670 10150
rect 10030 9880 10070 10150
rect 9510 9780 12670 9820
rect 12740 9780 13390 9820
rect 9230 9430 9270 9770
rect 9630 9450 9670 9770
rect 10030 9450 10070 9770
rect 10430 9450 10470 9770
rect 10830 9450 10870 9770
rect 11230 9450 11270 9770
rect 11630 9450 11670 9770
rect 12030 9450 12070 9770
rect 12430 9450 12470 9770
rect 9450 9410 12960 9450
rect 7840 9040 8120 9080
rect 8300 9040 12610 9080
rect 12740 9040 13390 9080
rect 6430 8710 6470 9040
rect 6830 8710 6870 9040
rect 7230 8710 7270 9040
rect 7630 8710 7670 8720
rect 30 8670 3140 8710
rect 3230 8670 5940 8710
rect 6030 8670 7860 8710
rect 30 8340 70 8670
rect 430 8340 470 8670
rect 830 8340 870 8670
rect 1230 8340 1270 8670
rect 1630 8340 1670 8670
rect 2030 8340 2070 8670
rect 2430 8340 2470 8670
rect 2830 8340 2870 8670
rect 3230 8340 3270 8670
rect 3630 8340 3670 8670
rect 4030 8340 4070 8670
rect 4430 8340 4470 8670
rect 4830 8340 4870 8670
rect 5230 8340 5270 8670
rect 5630 8340 5670 8670
rect 6030 8340 6070 8670
rect 6430 8340 6470 8670
rect 6830 8340 6870 8670
rect 7230 8340 7270 8670
rect 7630 8340 7670 8670
rect 30 8300 3140 8340
rect 3230 8300 5940 8340
rect 6030 8300 7830 8340
rect 8030 8300 8070 9040
rect 8430 8710 8470 9040
rect 8830 8710 8870 9040
rect 9230 8710 9270 9040
rect 9630 8710 9670 9040
rect 10030 8710 10070 9040
rect 10430 8710 10470 9040
rect 10830 8710 10870 9040
rect 11230 8710 11270 9040
rect 11630 8710 11670 9040
rect 12030 8710 12070 9040
rect 12430 8710 12470 9040
rect 8300 8670 12610 8710
rect 12690 8670 12960 8710
rect 8430 8340 8470 8670
rect 8830 8340 8870 8670
rect 9230 8340 9270 8670
rect 9630 8340 9670 8670
rect 10030 8340 10070 8670
rect 10430 8340 10470 8670
rect 10830 8340 10870 8670
rect 11230 8340 11270 8670
rect 11630 8340 11670 8670
rect 12030 8340 12070 8670
rect 12430 8340 12470 8670
rect 8300 8300 12610 8340
rect 12690 8300 12960 8340
rect 30 7970 70 8300
rect 430 7970 470 8300
rect 830 7970 870 8300
rect 1230 7970 1270 8300
rect 1630 7970 1670 8300
rect 2030 7970 2070 8300
rect 2430 7970 2470 8300
rect 2830 7970 2870 8300
rect 3230 7970 3270 8300
rect 3630 7970 3670 8300
rect 4030 7970 4070 8300
rect 4430 7970 4470 8300
rect 4830 7970 4870 8300
rect 5230 7970 5270 8300
rect 5630 7970 5670 8300
rect 30 7930 3140 7970
rect 3230 7930 5940 7970
rect 30 7600 70 7930
rect 430 7600 470 7930
rect 830 7600 870 7930
rect 1230 7600 1270 7930
rect 1630 7600 1670 7930
rect 2030 7600 2070 7930
rect 2430 7600 2470 7930
rect 2830 7600 2870 7930
rect 3230 7600 3270 7930
rect 3630 7600 3670 7930
rect 4030 7600 4070 7930
rect 4430 7600 4470 7930
rect 4830 7600 4870 7930
rect 5230 7600 5270 7930
rect 5630 7600 5670 7930
rect 30 7560 3140 7600
rect 3230 7560 5940 7600
rect 30 7230 70 7560
rect 430 7230 470 7560
rect 830 7230 870 7560
rect 1230 7230 1270 7560
rect 1630 7230 1670 7560
rect 2030 7230 2070 7560
rect 2430 7230 2470 7560
rect 2830 7230 2870 7560
rect 3230 7230 3270 7560
rect 3630 7230 3670 7560
rect 4030 7230 4070 7560
rect 4430 7230 4470 7560
rect 4830 7230 4870 7560
rect 5230 7230 5270 7560
rect 5630 7230 5670 7560
rect 6030 7230 6070 8300
rect 6430 7970 6470 8300
rect 6830 7970 6870 8300
rect 7230 7970 7270 8300
rect 7630 7970 7670 8300
rect 9230 8230 9270 8300
rect 9630 8230 9670 8300
rect 10030 8230 10070 8300
rect 10430 8230 10470 8300
rect 10830 8230 10870 8300
rect 11230 8230 11270 8300
rect 11630 8230 11670 8300
rect 12030 8230 12070 8300
rect 12430 8230 12470 8300
rect 8030 7970 8070 8000
rect 8430 7970 8470 8000
rect 8830 7970 8870 8000
rect 9230 7970 9270 8000
rect 9630 7970 9670 8000
rect 10030 7970 10070 8000
rect 10430 7970 10470 8000
rect 10830 7970 10870 8000
rect 11230 7970 11270 8000
rect 11630 7970 11670 8000
rect 12030 7970 12070 8000
rect 6330 7930 12470 7970
rect 12740 7930 13390 7970
rect 6430 7600 6470 7930
rect 6830 7600 6870 7930
rect 7230 7600 7270 7930
rect 7630 7600 7670 7930
rect 8030 7600 8070 7930
rect 8430 7600 8470 7930
rect 8830 7600 8870 7930
rect 9230 7600 9270 7930
rect 9630 7600 9670 7930
rect 10030 7600 10070 7930
rect 10430 7600 10470 7930
rect 10830 7600 10870 7930
rect 11230 7600 11270 7930
rect 11630 7600 11670 7930
rect 12030 7600 12070 7930
rect 12430 7630 12470 7930
rect 6280 7560 12490 7600
rect 12690 7560 12960 7600
rect 6430 7230 6470 7560
rect 6830 7230 6870 7560
rect 7230 7230 7270 7560
rect 7630 7230 7670 7560
rect 8030 7230 8070 7560
rect 8430 7230 8470 7560
rect 8830 7230 8870 7560
rect 9230 7230 9270 7560
rect 9630 7230 9670 7560
rect 10030 7230 10070 7560
rect 10430 7230 10470 7560
rect 10830 7230 10870 7560
rect 11230 7230 11270 7560
rect 11630 7230 11670 7560
rect 12030 7230 12070 7560
rect 12430 7230 12470 7560
rect 30 7190 3140 7230
rect 3230 7190 5940 7230
rect 6030 7190 12960 7230
rect 30 6860 70 7190
rect 430 6860 470 7190
rect 830 6860 870 7190
rect 1230 6860 1270 7190
rect 1630 6860 1670 7190
rect 2030 6860 2070 7190
rect 2430 6860 2470 7190
rect 2830 6860 2870 7190
rect 3230 6860 3270 7190
rect 3630 6860 3670 7190
rect 4030 6860 4070 7190
rect 4430 6860 4470 7190
rect 4830 6860 4870 7190
rect 5230 6860 5270 7190
rect 5630 6860 5670 7190
rect 6030 6860 6070 7190
rect 6430 6860 6470 7190
rect 6830 6860 6870 7190
rect 7230 6860 7270 7190
rect 7630 6860 7670 7190
rect 8030 6860 8070 7190
rect 8430 6860 8470 7190
rect 8830 6860 8870 7190
rect 9230 6860 9270 7190
rect 9630 6860 9670 7190
rect 10030 6860 10070 7190
rect 10430 6860 10470 7190
rect 10830 6860 10870 7190
rect 11230 6860 11270 7190
rect 11630 6860 11670 7190
rect 12030 6860 12070 7190
rect 12430 6860 12470 7190
rect 30 6820 3140 6860
rect 3230 6820 5940 6860
rect 6030 6820 12960 6860
rect 30 6490 70 6820
rect 430 6490 470 6820
rect 830 6490 870 6820
rect 1230 6490 1270 6820
rect 1630 6490 1670 6820
rect 2030 6490 2070 6820
rect 2430 6490 2470 6820
rect 2830 6490 2870 6820
rect 3230 6490 3270 6820
rect 3630 6490 3670 6820
rect 4030 6490 4070 6820
rect 4430 6490 4470 6820
rect 4830 6490 4870 6820
rect 5230 6490 5270 6820
rect 5630 6490 5670 6820
rect 6030 6490 6070 6820
rect 6430 6490 6470 6820
rect 6830 6490 6870 6820
rect 7230 6490 7270 6820
rect 7630 6490 7670 6820
rect 8030 6490 8070 6820
rect 8430 6490 8470 6820
rect 8830 6490 8870 6820
rect 9230 6490 9270 6820
rect 9630 6490 9670 6820
rect 10030 6490 10070 6820
rect 10430 6490 10470 6820
rect 10830 6490 10870 6820
rect 11230 6490 11270 6820
rect 11630 6490 11670 6820
rect 12030 6490 12070 6820
rect 12430 6490 12470 6820
rect 30 6450 3140 6490
rect 3230 6450 5780 6490
rect 6030 6450 12960 6490
rect 30 6120 70 6450
rect 430 6120 470 6450
rect 830 6120 870 6450
rect 1230 6120 1270 6450
rect 1630 6120 1670 6450
rect 2030 6120 2070 6450
rect 2430 6120 2470 6450
rect 2830 6120 2870 6450
rect 30 6080 3140 6120
rect 30 5750 70 6080
rect 430 5750 470 6080
rect 830 5750 870 6080
rect 1230 5750 1270 6080
rect 1630 5750 1670 6080
rect 2030 5750 2070 6080
rect 2430 5750 2470 6080
rect 2830 5750 2870 6080
rect 30 5710 3140 5750
rect 30 5380 70 5710
rect 430 5380 470 5710
rect 830 5380 870 5710
rect 1230 5380 1270 5710
rect 1630 5380 1670 5710
rect 2030 5380 2070 5710
rect 2430 5380 2470 5710
rect 2830 5380 2870 5710
rect 3230 5380 3270 6450
rect 3630 6120 3670 6450
rect 4030 6120 4070 6450
rect 4430 6120 4470 6450
rect 4830 6120 4870 6450
rect 5230 6120 5270 6450
rect 5630 6120 5670 6450
rect 6030 6410 6070 6450
rect 6430 6410 6470 6450
rect 6830 6410 6870 6450
rect 7230 6410 7270 6450
rect 7630 6410 7670 6450
rect 8030 6410 8070 6450
rect 8430 6410 8470 6450
rect 8830 6410 8870 6450
rect 9230 6410 9270 6450
rect 9630 6410 9670 6450
rect 10030 6410 10070 6450
rect 10430 6410 10470 6450
rect 10830 6410 10870 6450
rect 11230 6410 11270 6450
rect 11630 6410 11670 6450
rect 12030 6410 12070 6450
rect 3500 6100 12450 6120
rect 3500 6080 12470 6100
rect 12740 6080 13390 6120
rect 3630 5750 3670 6080
rect 4030 5750 4070 6080
rect 4430 5750 4470 6080
rect 4830 5750 4870 6080
rect 5230 5750 5270 6080
rect 5630 5750 5670 6080
rect 6030 5750 6070 6080
rect 6430 5750 6470 6080
rect 6830 5750 6870 6080
rect 7230 5750 7270 6080
rect 7630 5750 7670 6080
rect 8030 5750 8070 6080
rect 8430 5750 8470 6080
rect 8830 5750 8870 6080
rect 9230 5750 9270 6080
rect 9630 5750 9670 6080
rect 10030 5750 10070 6080
rect 10430 5750 10470 6080
rect 10830 5750 10870 6080
rect 11230 5750 11270 6080
rect 11630 5750 11670 6080
rect 12030 5750 12070 6080
rect 12430 5750 12470 6080
rect 3500 5710 12470 5750
rect 12690 5710 12960 5750
rect 3630 5380 3670 5710
rect 4030 5380 4070 5710
rect 4430 5380 4470 5710
rect 4830 5380 4870 5710
rect 5230 5380 5270 5710
rect 5630 5380 5670 5710
rect 6030 5380 6070 5710
rect 6430 5380 6470 5710
rect 6830 5380 6870 5710
rect 7230 5380 7270 5710
rect 7630 5380 7670 5710
rect 8030 5380 8070 5710
rect 8430 5380 8470 5710
rect 8830 5380 8870 5710
rect 9230 5380 9270 5710
rect 9630 5380 9670 5710
rect 10030 5380 10070 5710
rect 10430 5380 10470 5710
rect 10830 5380 10870 5710
rect 11230 5380 11270 5710
rect 11630 5380 11670 5710
rect 12030 5380 12070 5710
rect 12430 5380 12470 5710
rect 30 5340 3140 5380
rect 3230 5340 12960 5380
rect 30 5010 70 5340
rect 430 5010 470 5340
rect 830 5010 870 5340
rect 1230 5010 1270 5340
rect 1630 5010 1670 5340
rect 2030 5010 2070 5340
rect 2430 5010 2470 5340
rect 2830 5010 2870 5340
rect 3230 5010 3270 5340
rect 3630 5010 3670 5340
rect 4030 5010 4070 5340
rect 4430 5010 4470 5340
rect 4830 5010 4870 5340
rect 5230 5010 5270 5340
rect 5630 5010 5670 5340
rect 6030 5010 6070 5340
rect 6430 5010 6470 5340
rect 6830 5010 6870 5340
rect 7230 5010 7270 5340
rect 7630 5010 7670 5340
rect 8030 5010 8070 5340
rect 8430 5010 8470 5340
rect 8830 5010 8870 5340
rect 9230 5010 9270 5340
rect 9630 5010 9670 5340
rect 10030 5010 10070 5340
rect 10430 5010 10470 5340
rect 10830 5010 10870 5340
rect 11230 5010 11270 5340
rect 11630 5010 11670 5340
rect 12030 5010 12070 5340
rect 12430 5010 12470 5340
rect 30 4970 3140 5010
rect 3230 4970 12960 5010
rect 30 4640 70 4970
rect 430 4640 470 4970
rect 830 4640 870 4970
rect 1230 4640 1270 4970
rect 1630 4640 1670 4970
rect 2030 4640 2070 4970
rect 2430 4640 2470 4970
rect 2830 4640 2870 4970
rect 3230 4640 3270 4970
rect 3630 4640 3670 4970
rect 4030 4640 4070 4970
rect 4430 4640 4470 4970
rect 4830 4640 4870 4970
rect 5230 4640 5270 4970
rect 5630 4640 5670 4970
rect 6030 4640 6070 4970
rect 6430 4640 6470 4970
rect 6830 4640 6870 4970
rect 7230 4640 7270 4970
rect 7630 4640 7670 4970
rect 8030 4640 8070 4970
rect 8430 4640 8470 4970
rect 8830 4640 8870 4970
rect 9230 4640 9270 4970
rect 9630 4640 9670 4970
rect 10030 4640 10070 4970
rect 10430 4640 10470 4970
rect 10830 4640 10870 4970
rect 11230 4640 11270 4970
rect 11630 4640 11670 4970
rect 12030 4640 12070 4970
rect 12430 4640 12470 4970
rect 30 4600 3140 4640
rect 3230 4600 12960 4640
rect 30 3900 70 4600
rect 430 4270 470 4600
rect 830 4270 870 4600
rect 1230 4270 1270 4600
rect 1630 4270 1670 4600
rect 2030 4270 2070 4600
rect 2430 4270 2470 4600
rect 2830 4270 2870 4600
rect 3230 4270 3270 4600
rect 3630 4270 3670 4600
rect 4030 4270 4070 4600
rect 4430 4270 4470 4600
rect 4830 4270 4870 4600
rect 5230 4270 5270 4600
rect 5630 4270 5670 4600
rect 6030 4270 6070 4600
rect 6430 4270 6470 4600
rect 6830 4270 6870 4600
rect 7230 4270 7270 4600
rect 7630 4270 7670 4600
rect 8030 4270 8070 4600
rect 8430 4270 8470 4600
rect 8830 4270 8870 4600
rect 9230 4270 9270 4600
rect 9630 4270 9670 4600
rect 10030 4270 10070 4600
rect 10430 4270 10470 4600
rect 10830 4270 10870 4600
rect 11230 4270 11270 4600
rect 11630 4270 11670 4600
rect 12030 4270 12070 4600
rect 12430 4270 12470 4600
rect 100 4230 2960 4270
rect 3230 4230 12960 4270
rect 430 3900 470 4230
rect 830 3900 870 4230
rect 1230 3900 1270 4230
rect 1630 3900 1670 4230
rect 2030 3900 2070 4230
rect 2430 3900 2470 4230
rect 2830 3900 2870 4230
rect 3230 4200 3270 4230
rect 3630 4200 3670 4230
rect 4030 4200 4070 4230
rect 4430 4200 4470 4230
rect 4830 4200 4870 4230
rect 5230 4200 5270 4230
rect 5630 4200 5670 4230
rect 6030 4210 6070 4230
rect 6430 4210 6470 4230
rect 6830 4210 6870 4230
rect 7230 4210 7270 4230
rect 7630 4210 7670 4230
rect 8030 4210 8070 4230
rect 8430 4210 8470 4230
rect 8830 4210 8870 4230
rect 9230 4210 9270 4230
rect 9630 4210 9670 4230
rect 10030 4210 10070 4230
rect 10430 4210 10470 4230
rect 10830 4210 10870 4230
rect 11230 4210 11270 4230
rect 11630 4210 11670 4230
rect 12030 4210 12070 4230
rect 12430 4210 12470 4230
rect 30 3860 13390 3900
rect 30 3530 70 3860
rect 430 3530 470 3860
rect 830 3530 870 3860
rect 1230 3530 1270 3860
rect 1630 3530 1670 3860
rect 2030 3530 2070 3860
rect 2430 3530 2470 3860
rect 2830 3530 2870 3860
rect 3230 3530 3270 3860
rect 3630 3530 3670 3860
rect 4030 3530 4070 3860
rect 4430 3530 4470 3860
rect 4830 3530 4870 3860
rect 5230 3530 5270 3860
rect 5630 3530 5670 3860
rect 6030 3530 6070 3860
rect 6430 3530 6470 3860
rect 6830 3530 6870 3860
rect 7230 3530 7270 3860
rect 7630 3530 7670 3860
rect 8030 3530 8070 3860
rect 8430 3530 8470 3860
rect 8830 3530 8870 3860
rect 9230 3530 9270 3860
rect 9630 3530 9670 3860
rect 10030 3530 10070 3860
rect 10430 3530 10470 3860
rect 10830 3530 10870 3860
rect 11230 3530 11270 3860
rect 11630 3530 11670 3860
rect 12030 3530 12070 3860
rect 12430 3530 12470 3860
rect 30 3490 12960 3530
rect 30 3160 70 3490
rect 430 3160 470 3490
rect 830 3160 870 3490
rect 1230 3160 1270 3490
rect 1630 3160 1670 3490
rect 2030 3160 2070 3490
rect 2430 3160 2470 3490
rect 2830 3160 2870 3490
rect 3230 3160 3270 3490
rect 3630 3160 3670 3490
rect 4030 3160 4070 3490
rect 4430 3160 4470 3490
rect 4830 3160 4870 3490
rect 5230 3160 5270 3490
rect 5630 3160 5670 3490
rect 6030 3160 6070 3490
rect 6430 3160 6470 3490
rect 6830 3160 6870 3490
rect 7230 3160 7270 3490
rect 7630 3160 7670 3490
rect 8030 3160 8070 3490
rect 8430 3160 8470 3490
rect 8830 3160 8870 3490
rect 9230 3160 9270 3490
rect 9630 3160 9670 3490
rect 10030 3160 10070 3490
rect 10430 3160 10470 3490
rect 10830 3160 10870 3490
rect 11230 3160 11270 3490
rect 11630 3160 11670 3490
rect 12030 3160 12070 3490
rect 12430 3160 12470 3490
rect 30 3120 12960 3160
rect 30 2790 70 3120
rect 430 2790 470 3120
rect 830 2790 870 3120
rect 1230 2790 1270 3120
rect 1630 2790 1670 3120
rect 2030 2790 2070 3120
rect 2430 2790 2470 3120
rect 2830 2790 2870 3120
rect 3230 2790 3270 3120
rect 3630 2790 3670 3120
rect 4030 2790 4070 3120
rect 4430 2790 4470 3120
rect 4830 2790 4870 3120
rect 5230 2790 5270 3120
rect 5630 2790 5670 3120
rect 6030 2790 6070 3120
rect 6430 2790 6470 3120
rect 6830 2790 6870 3120
rect 7230 2790 7270 3120
rect 7630 2790 7670 3120
rect 8030 2790 8070 3120
rect 8430 2790 8470 3120
rect 8830 2790 8870 3120
rect 9230 2790 9270 3120
rect 9630 2790 9670 3120
rect 10030 2790 10070 3120
rect 10430 2790 10470 3120
rect 10830 2790 10870 3120
rect 11230 2790 11270 3120
rect 11630 2790 11670 3120
rect 12030 2790 12070 3120
rect 12430 2790 12470 3120
rect 30 2750 12960 2790
rect 30 2420 70 2750
rect 430 2420 470 2750
rect 830 2420 870 2750
rect 1230 2420 1270 2750
rect 1630 2420 1670 2750
rect 2030 2420 2070 2750
rect 2430 2420 2470 2750
rect 2830 2420 2870 2750
rect 3230 2420 3270 2750
rect 3630 2420 3670 2750
rect 4030 2420 4070 2750
rect 4430 2420 4470 2750
rect 4830 2420 4870 2750
rect 5230 2420 5270 2750
rect 5630 2420 5670 2750
rect 6030 2420 6070 2750
rect 6430 2420 6470 2750
rect 6830 2420 6870 2750
rect 7230 2420 7270 2750
rect 7630 2420 7670 2750
rect 8030 2420 8070 2750
rect 8430 2420 8470 2750
rect 8830 2420 8870 2750
rect 9230 2420 9270 2750
rect 9630 2420 9670 2750
rect 10030 2420 10070 2750
rect 10430 2420 10470 2750
rect 10830 2420 10870 2750
rect 11230 2420 11270 2750
rect 11630 2420 11670 2750
rect 12030 2420 12070 2750
rect 12430 2420 12470 2750
rect 30 2380 12960 2420
rect 30 2050 70 2380
rect 430 2050 470 2380
rect 830 2050 870 2380
rect 1230 2050 1270 2380
rect 1630 2050 1670 2380
rect 2030 2050 2070 2380
rect 2430 2050 2470 2380
rect 2830 2050 2870 2380
rect 3230 2050 3270 2380
rect 3630 2050 3670 2380
rect 4030 2050 4070 2380
rect 4430 2050 4470 2380
rect 4830 2050 4870 2380
rect 5230 2050 5270 2380
rect 5630 2050 5670 2380
rect 6030 2050 6070 2380
rect 6430 2050 6470 2380
rect 6830 2050 6870 2380
rect 7230 2050 7270 2380
rect 7630 2050 7670 2380
rect 8030 2050 8070 2380
rect 8430 2050 8470 2380
rect 8830 2050 8870 2380
rect 9230 2050 9270 2380
rect 9630 2050 9670 2380
rect 10030 2050 10070 2380
rect 10430 2050 10470 2380
rect 10830 2050 10870 2380
rect 11230 2050 11270 2380
rect 11630 2050 11670 2380
rect 12030 2050 12070 2380
rect 12430 2050 12470 2380
rect 30 2010 12960 2050
rect 30 1680 70 2010
rect 430 1680 470 2010
rect 830 1680 870 2010
rect 1230 1680 1270 2010
rect 1630 1680 1670 2010
rect 2030 1680 2070 2010
rect 2430 1680 2470 2010
rect 2830 1680 2870 2010
rect 3230 1680 3270 2010
rect 3630 1680 3670 2010
rect 4030 1680 4070 2010
rect 4430 1680 4470 2010
rect 4830 1680 4870 2010
rect 5230 1680 5270 2010
rect 5630 1680 5670 2010
rect 6030 1680 6070 2010
rect 6430 1680 6470 2010
rect 6830 1680 6870 2010
rect 7230 1680 7270 2010
rect 7630 1680 7670 2010
rect 8030 1680 8070 2010
rect 8430 1680 8470 2010
rect 8830 1680 8870 2010
rect 9230 1680 9270 2010
rect 9630 1680 9670 2010
rect 10030 1680 10070 2010
rect 10430 1680 10470 2010
rect 10830 1680 10870 2010
rect 11230 1680 11270 2010
rect 11630 1680 11670 2010
rect 12030 1680 12070 2010
rect 12430 1680 12470 2010
rect 30 1640 12960 1680
rect 30 1310 70 1640
rect 430 1310 470 1640
rect 830 1310 870 1640
rect 1230 1310 1270 1640
rect 1630 1310 1670 1640
rect 2030 1310 2070 1640
rect 2430 1310 2470 1640
rect 2830 1310 2870 1640
rect 3230 1310 3270 1640
rect 3630 1310 3670 1640
rect 4030 1310 4070 1640
rect 4430 1310 4470 1640
rect 4830 1310 4870 1640
rect 5230 1310 5270 1640
rect 5630 1310 5670 1640
rect 6030 1310 6070 1640
rect 6430 1310 6470 1640
rect 6830 1310 6870 1640
rect 7230 1310 7270 1640
rect 7630 1310 7670 1640
rect 8030 1310 8070 1640
rect 8430 1310 8470 1640
rect 8830 1310 8870 1640
rect 9230 1310 9270 1640
rect 9630 1310 9670 1640
rect 10030 1310 10070 1640
rect 10430 1310 10470 1640
rect 10830 1310 10870 1640
rect 11230 1310 11270 1640
rect 11630 1310 11670 1640
rect 12030 1310 12070 1640
rect 12430 1310 12470 1640
rect 30 1270 12960 1310
rect 30 940 70 1270
rect 430 940 470 1270
rect 830 940 870 1270
rect 1230 940 1270 1270
rect 1630 940 1670 1270
rect 2030 940 2070 1270
rect 2430 940 2470 1270
rect 2830 940 2870 1270
rect 3230 940 3270 1270
rect 3630 940 3670 1270
rect 4030 940 4070 1270
rect 4430 940 4470 1270
rect 4830 940 4870 1270
rect 5230 940 5270 1270
rect 5630 940 5670 1270
rect 6030 940 6070 1270
rect 6430 940 6470 1270
rect 6830 940 6870 1270
rect 7230 940 7270 1270
rect 7630 940 7670 1270
rect 8030 940 8070 1270
rect 8430 940 8470 1270
rect 8830 940 8870 1270
rect 9230 940 9270 1270
rect 9630 940 9670 1270
rect 10030 940 10070 1270
rect 10430 940 10470 1270
rect 10830 940 10870 1270
rect 11230 940 11270 1270
rect 11630 940 11670 1270
rect 12030 940 12070 1270
rect 12430 940 12470 1270
rect 30 900 12960 940
rect 30 570 70 900
rect 430 570 470 900
rect 830 570 870 900
rect 1230 570 1270 900
rect 1630 570 1670 900
rect 2030 570 2070 900
rect 2430 570 2470 900
rect 2830 570 2870 900
rect 3230 570 3270 900
rect 3630 570 3670 900
rect 4030 570 4070 900
rect 4430 570 4470 900
rect 4830 570 4870 900
rect 5230 570 5270 900
rect 5630 570 5670 900
rect 6030 570 6070 900
rect 6430 570 6470 900
rect 6830 570 6870 900
rect 7230 570 7270 900
rect 7630 570 7670 900
rect 8030 570 8070 900
rect 8430 570 8470 900
rect 8830 570 8870 900
rect 9230 570 9270 900
rect 9630 570 9670 900
rect 10030 570 10070 900
rect 10430 570 10470 900
rect 10830 570 10870 900
rect 11230 570 11270 900
rect 11630 570 11670 900
rect 12030 570 12070 900
rect 12430 570 12470 900
rect 30 530 12960 570
rect 30 130 70 530
rect 430 200 470 530
rect 830 200 870 530
rect 1230 200 1270 530
rect 1630 200 1670 530
rect 2030 200 2070 530
rect 2430 200 2470 530
rect 2830 200 2870 530
rect 3230 200 3270 530
rect 3630 200 3670 530
rect 4030 200 4070 530
rect 4430 200 4470 530
rect 4830 200 4870 530
rect 5230 200 5270 530
rect 5630 200 5670 530
rect 6030 200 6070 530
rect 6430 200 6470 530
rect 6830 200 6870 530
rect 7230 200 7270 530
rect 7630 200 7670 530
rect 8030 200 8070 530
rect 8430 200 8470 530
rect 8830 200 8870 530
rect 9230 200 9270 530
rect 9630 200 9670 530
rect 10030 200 10070 530
rect 10430 200 10470 530
rect 10830 200 10870 530
rect 11230 200 11270 530
rect 11630 200 11670 530
rect 12030 200 12070 530
rect 12430 200 12470 530
rect 310 160 12590 200
rect 12700 160 12970 200
rect 430 130 470 160
rect 830 130 870 160
rect 1230 130 1270 160
rect 1630 130 1670 160
rect 2030 130 2070 160
rect 2430 130 2470 160
rect 2830 130 2870 160
rect -376 -103 -324 -50
rect -370 -116 -324 -103
rect -370 -140 -330 -116
rect -232 -170 12972 -164
rect -300 -210 -220 -170
rect 12960 -210 13020 -170
rect -232 -216 12972 -210
<< via1 >>
rect -265 24170 -205 24180
rect -265 24130 -255 24170
rect -255 24130 -215 24170
rect -215 24130 -205 24170
rect -265 24120 -205 24130
rect -165 24170 -105 24180
rect -165 24130 -155 24170
rect -155 24130 -115 24170
rect -115 24130 -105 24170
rect -165 24120 -105 24130
rect 12930 24115 12990 24125
rect 12930 24075 12940 24115
rect 12940 24075 12980 24115
rect 12980 24075 12990 24115
rect 12930 24065 12990 24075
rect 13030 24115 13090 24125
rect 13030 24075 13040 24115
rect 13040 24075 13080 24115
rect 13080 24075 13090 24115
rect 13030 24065 13090 24075
<< metal2 >>
rect -275 24180 -95 24190
rect -275 24120 -265 24180
rect -205 24120 -165 24180
rect -105 24120 -95 24180
rect -275 24110 -95 24120
rect 12915 24125 13105 24135
rect 12990 24065 13030 24125
rect 12915 24055 13105 24065
<< via2 >>
rect -265 24120 -205 24180
rect -165 24120 -105 24180
rect 12915 24065 12930 24125
rect 12930 24065 12975 24125
rect 13045 24065 13090 24125
rect 13090 24065 13105 24125
<< metal3 >>
rect -275 24180 -95 24185
rect -275 24120 -265 24180
rect -205 24120 -165 24180
rect -105 24120 -95 24180
rect -275 24115 -95 24120
rect -215 23980 -155 24115
rect 12895 24055 12905 24135
rect 12985 24055 13035 24135
rect 13115 24055 13125 24135
rect 12985 23980 13045 24055
rect 170 23875 180 23945
rect 250 23875 260 23945
rect 570 23875 580 23945
rect 650 23875 660 23945
rect 970 23875 980 23945
rect 1050 23875 1060 23945
rect 1370 23875 1380 23945
rect 1450 23875 1460 23945
rect 1770 23875 1780 23945
rect 1850 23875 1860 23945
rect 2170 23875 2180 23945
rect 2250 23875 2260 23945
rect 2570 23875 2580 23945
rect 2650 23875 2660 23945
rect 2970 23875 2980 23945
rect 3050 23875 3060 23945
rect 3370 23875 3380 23945
rect 3450 23875 3460 23945
rect 3770 23875 3780 23945
rect 3850 23875 3860 23945
rect 4170 23875 4180 23945
rect 4250 23875 4260 23945
rect 4570 23875 4580 23945
rect 4650 23875 4660 23945
rect 4970 23875 4980 23945
rect 5050 23875 5060 23945
rect 5370 23875 5380 23945
rect 5450 23875 5460 23945
rect 5770 23875 5780 23945
rect 5850 23875 5860 23945
rect 6170 23875 6180 23945
rect 6250 23875 6260 23945
rect 6570 23875 6580 23945
rect 6650 23875 6660 23945
rect 6970 23875 6980 23945
rect 7050 23875 7060 23945
rect 7370 23875 7380 23945
rect 7450 23875 7460 23945
rect 7770 23875 7780 23945
rect 7850 23875 7860 23945
rect 8170 23875 8180 23945
rect 8250 23875 8260 23945
rect 8570 23875 8580 23945
rect 8650 23875 8660 23945
rect 8970 23875 8980 23945
rect 9050 23875 9060 23945
rect 9370 23875 9380 23945
rect 9450 23875 9460 23945
rect 9770 23875 9780 23945
rect 9850 23875 9860 23945
rect 10170 23875 10180 23945
rect 10250 23875 10260 23945
rect 10570 23875 10580 23945
rect 10650 23875 10660 23945
rect 10970 23875 10980 23945
rect 11050 23875 11060 23945
rect 11370 23875 11380 23945
rect 11450 23875 11460 23945
rect 11770 23875 11780 23945
rect 11850 23875 11860 23945
rect 12170 23875 12180 23945
rect 12250 23875 12260 23945
rect 12570 23875 12580 23945
rect 12650 23875 12660 23945
<< via3 >>
rect 12905 24125 12985 24135
rect 12905 24065 12915 24125
rect 12915 24065 12975 24125
rect 12975 24065 12985 24125
rect 12905 24055 12985 24065
rect 13035 24125 13115 24135
rect 13035 24065 13045 24125
rect 13045 24065 13105 24125
rect 13105 24065 13115 24125
rect 13035 24055 13115 24065
rect 180 23875 250 23945
rect 580 23875 650 23945
rect 980 23875 1050 23945
rect 1380 23875 1450 23945
rect 1780 23875 1850 23945
rect 2180 23875 2250 23945
rect 2580 23875 2650 23945
rect 2980 23875 3050 23945
rect 3380 23875 3450 23945
rect 3780 23875 3850 23945
rect 4180 23875 4250 23945
rect 4580 23875 4650 23945
rect 4980 23875 5050 23945
rect 5380 23875 5450 23945
rect 5780 23875 5850 23945
rect 6180 23875 6250 23945
rect 6580 23875 6650 23945
rect 6980 23875 7050 23945
rect 7380 23875 7450 23945
rect 7780 23875 7850 23945
rect 8180 23875 8250 23945
rect 8580 23875 8650 23945
rect 8980 23875 9050 23945
rect 9380 23875 9450 23945
rect 9780 23875 9850 23945
rect 10180 23875 10250 23945
rect 10580 23875 10650 23945
rect 10980 23875 11050 23945
rect 11380 23875 11450 23945
rect 11780 23875 11850 23945
rect 12180 23875 12250 23945
rect 12580 23875 12650 23945
<< metal4 >>
rect 180 24075 12650 24145
rect 180 23946 250 24075
rect 580 23946 650 24075
rect 980 23946 1050 24075
rect 1380 23946 1450 24075
rect 1780 23946 1850 24075
rect 2180 23946 2250 24075
rect 2580 23946 2650 24075
rect 2980 23946 3050 24075
rect 3380 23946 3450 24075
rect 3780 23946 3850 24075
rect 4180 23946 4250 24075
rect 4580 23946 4650 24075
rect 4980 23946 5050 24075
rect 5380 23946 5450 24075
rect 5780 23946 5850 24075
rect 6180 23946 6250 24075
rect 6580 23946 6650 24075
rect 6980 23946 7050 24075
rect 7380 23946 7450 24075
rect 7780 23946 7850 24075
rect 8180 23946 8250 24075
rect 8580 23946 8650 24075
rect 8980 23946 9050 24075
rect 9380 23946 9450 24075
rect 9780 23946 9850 24075
rect 10180 23946 10250 24075
rect 10580 23946 10650 24075
rect 10980 23946 11050 24075
rect 11380 23946 11450 24075
rect 11780 23946 11850 24075
rect 12180 23946 12250 24075
rect 12580 23946 12650 24075
rect 12895 24135 13125 24145
rect 12895 24055 12905 24135
rect 12985 24055 13035 24135
rect 13115 24055 13125 24135
rect 12895 24045 13125 24055
rect 179 23945 251 23946
rect 179 23875 180 23945
rect 250 23875 251 23945
rect 179 23874 251 23875
rect 579 23945 651 23946
rect 579 23875 580 23945
rect 650 23875 651 23945
rect 579 23874 651 23875
rect 979 23945 1051 23946
rect 979 23875 980 23945
rect 1050 23875 1051 23945
rect 979 23874 1051 23875
rect 1379 23945 1451 23946
rect 1379 23875 1380 23945
rect 1450 23875 1451 23945
rect 1379 23874 1451 23875
rect 1779 23945 1851 23946
rect 1779 23875 1780 23945
rect 1850 23875 1851 23945
rect 1779 23874 1851 23875
rect 2179 23945 2251 23946
rect 2179 23875 2180 23945
rect 2250 23875 2251 23945
rect 2179 23874 2251 23875
rect 2579 23945 2651 23946
rect 2579 23875 2580 23945
rect 2650 23875 2651 23945
rect 2579 23874 2651 23875
rect 2979 23945 3051 23946
rect 2979 23875 2980 23945
rect 3050 23875 3051 23945
rect 2979 23874 3051 23875
rect 3379 23945 3451 23946
rect 3379 23875 3380 23945
rect 3450 23875 3451 23945
rect 3379 23874 3451 23875
rect 3779 23945 3851 23946
rect 3779 23875 3780 23945
rect 3850 23875 3851 23945
rect 3779 23874 3851 23875
rect 4179 23945 4251 23946
rect 4179 23875 4180 23945
rect 4250 23875 4251 23945
rect 4179 23874 4251 23875
rect 4579 23945 4651 23946
rect 4579 23875 4580 23945
rect 4650 23875 4651 23945
rect 4579 23874 4651 23875
rect 4979 23945 5051 23946
rect 4979 23875 4980 23945
rect 5050 23875 5051 23945
rect 4979 23874 5051 23875
rect 5379 23945 5451 23946
rect 5379 23875 5380 23945
rect 5450 23875 5451 23945
rect 5379 23874 5451 23875
rect 5779 23945 5851 23946
rect 5779 23875 5780 23945
rect 5850 23875 5851 23945
rect 5779 23874 5851 23875
rect 6179 23945 6251 23946
rect 6179 23875 6180 23945
rect 6250 23875 6251 23945
rect 6179 23874 6251 23875
rect 6579 23945 6651 23946
rect 6579 23875 6580 23945
rect 6650 23875 6651 23945
rect 6579 23874 6651 23875
rect 6979 23945 7051 23946
rect 6979 23875 6980 23945
rect 7050 23875 7051 23945
rect 6979 23874 7051 23875
rect 7379 23945 7451 23946
rect 7379 23875 7380 23945
rect 7450 23875 7451 23945
rect 7379 23874 7451 23875
rect 7779 23945 7851 23946
rect 7779 23875 7780 23945
rect 7850 23875 7851 23945
rect 7779 23874 7851 23875
rect 8179 23945 8251 23946
rect 8179 23875 8180 23945
rect 8250 23875 8251 23945
rect 8179 23874 8251 23875
rect 8579 23945 8651 23946
rect 8579 23875 8580 23945
rect 8650 23875 8651 23945
rect 8579 23874 8651 23875
rect 8979 23945 9051 23946
rect 8979 23875 8980 23945
rect 9050 23875 9051 23945
rect 8979 23874 9051 23875
rect 9379 23945 9451 23946
rect 9379 23875 9380 23945
rect 9450 23875 9451 23945
rect 9379 23874 9451 23875
rect 9779 23945 9851 23946
rect 9779 23875 9780 23945
rect 9850 23875 9851 23945
rect 9779 23874 9851 23875
rect 10179 23945 10251 23946
rect 10179 23875 10180 23945
rect 10250 23875 10251 23945
rect 10179 23874 10251 23875
rect 10579 23945 10651 23946
rect 10579 23875 10580 23945
rect 10650 23875 10651 23945
rect 10579 23874 10651 23875
rect 10979 23945 11051 23946
rect 10979 23875 10980 23945
rect 11050 23875 11051 23945
rect 10979 23874 11051 23875
rect 11379 23945 11451 23946
rect 11379 23875 11380 23945
rect 11450 23875 11451 23945
rect 11379 23874 11451 23875
rect 11779 23945 11851 23946
rect 11779 23875 11780 23945
rect 11850 23875 11851 23945
rect 11779 23874 11851 23875
rect 12179 23945 12251 23946
rect 12179 23875 12180 23945
rect 12250 23875 12251 23945
rect 12179 23874 12251 23875
rect 12579 23945 12651 23946
rect 12579 23875 12580 23945
rect 12650 23875 12651 23945
rect 12579 23874 12651 23875
use unit_cap  unit_cap_0
array 0 31 400 0 63 370
timestamp 1715382157
transform 1 0 -1225 0 1 -1450
box 1255 1440 1625 1810
use unit_cap  unit_cap_1
array 0 0 340 0 65 370
timestamp 1715382157
transform 1 0 -1625 0 1 -1820
box 1255 1440 1625 1810
use unit_cap  unit_cap_2
array 0 31 400 0 0 370
timestamp 1715382157
transform 1 0 -1225 0 1 -1820
box 1255 1440 1625 1810
use unit_cap  unit_cap_4
array 0 0 340 0 65 370
timestamp 1715382157
transform 1 0 11575 0 1 -1820
box 1255 1440 1625 1810
use unit_cap  unit_cap_5
array 0 31 400 0 0 370
timestamp 1715382157
transform 1 0 -1225 0 1 22230
box 1255 1440 1625 1810
<< labels >>
rlabel metal1 13360 3870 13380 3890 1 C10
port 12 n
rlabel metal1 13360 6090 13380 6110 1 C9
port 11 n
rlabel metal1 13360 7940 13380 7960 1 C8
port 10 n
rlabel metal1 13360 9050 13380 9070 1 C7
port 9 n
rlabel metal1 13360 9790 13380 9810 1 C6
port 8 n
rlabel metal1 13360 10160 13380 10180 1 C5
port 7 n
rlabel metal1 13360 10900 13380 10920 1 C4
port 6 n
rlabel metal1 13360 12750 13380 12770 1 C3
port 5 n
rlabel metal1 13360 11270 13380 11290 1 C2
port 4 n
rlabel metal1 13360 12380 13380 12400 1 C1
port 3 n
rlabel metal1 13360 12010 13380 12030 1 C0
port 2 n
rlabel metal1 13360 11640 13380 11660 1 C0_dummy
port 1 n
rlabel metal4 12975 24065 13035 24125 1 VSS
port 14 n
rlabel metal4 12390 24090 12495 24135 1 Ctop
port 15 n
<< end >>
