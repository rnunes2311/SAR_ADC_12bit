magic
tech sky130A
magscale 1 2
timestamp 1717107273
<< viali >>
rect -1400 870 -1350 920
rect -1290 860 -1240 910
rect 606 901 657 961
rect 770 860 820 910
rect -860 770 -810 820
rect 1150 790 1200 840
rect -1410 290 -1360 340
rect -860 330 -810 380
rect -220 324 -170 374
rect -1290 234 -1240 284
rect -760 234 -710 284
rect -650 234 -600 284
rect -40 234 10 284
rect 130 234 180 284
rect 504 234 554 284
rect 770 234 820 284
rect 1150 244 1200 294
rect 606 181 656 231
<< metal1 >>
rect -1285 1010 1200 1040
rect -1412 920 -1338 926
rect -1430 860 -1420 920
rect -1350 870 -1338 920
rect -1285 916 -1255 1010
rect 600 961 663 973
rect -1360 864 -1338 870
rect -1302 910 -1228 916
rect -1360 860 -1350 864
rect -1302 860 -1290 910
rect -1240 860 -1228 910
rect 600 901 606 961
rect 657 960 663 961
rect 600 900 610 901
rect 670 900 680 960
rect 758 910 832 916
rect 600 889 663 900
rect -1302 854 -1228 860
rect 758 860 770 910
rect 820 860 832 910
rect 758 854 832 860
rect -872 820 -798 826
rect -872 780 -860 820
rect -880 770 -860 780
rect -810 780 -798 820
rect -810 770 -790 780
rect -880 750 -790 770
rect -880 690 -870 750
rect -810 690 -790 750
rect -880 680 -790 690
rect 775 680 805 854
rect 1170 850 1200 1010
rect 1140 846 1150 850
rect 1138 790 1150 846
rect 1210 790 1220 850
rect 1138 784 1212 790
rect -880 650 805 680
rect -1420 430 -1410 490
rect -1350 430 -1340 490
rect -855 464 805 494
rect -1400 346 -1370 430
rect -855 386 -825 464
rect -872 380 -798 386
rect -1422 340 -1348 346
rect -1422 290 -1410 340
rect -1360 290 -1348 340
rect -872 330 -860 380
rect -810 330 -798 380
rect -232 374 -158 380
rect -872 324 -798 330
rect -1422 284 -1348 290
rect -1302 284 -1228 290
rect -1302 234 -1290 284
rect -1240 234 -1228 284
rect -860 250 -830 324
rect -240 314 -230 374
rect -170 364 -158 374
rect 600 370 610 430
rect 670 370 680 430
rect -170 334 170 364
rect -170 318 -158 334
rect -170 314 -160 318
rect -1302 228 -1228 234
rect -1285 134 -1255 228
rect -890 190 -880 250
rect -820 190 -810 250
rect -780 234 -770 294
rect -710 290 -700 294
rect 140 290 170 334
rect -710 234 -698 290
rect -772 228 -698 234
rect -662 284 -588 290
rect -662 234 -650 284
rect -600 234 -588 284
rect -662 228 -588 234
rect -52 284 22 290
rect 118 284 192 290
rect -52 228 -40 284
rect -640 192 -610 228
rect -50 224 -40 228
rect 20 224 30 284
rect 118 234 130 284
rect 180 234 192 284
rect 492 284 566 290
rect 492 240 504 284
rect 118 228 192 234
rect 480 192 490 240
rect 554 234 566 284
rect 620 237 650 370
rect 775 290 805 464
rect 1138 294 1212 300
rect 758 284 832 290
rect -640 180 490 192
rect 550 228 566 234
rect 594 231 668 237
rect 550 180 560 228
rect 594 181 606 231
rect 656 181 668 231
rect 758 234 770 284
rect 820 234 832 284
rect 1138 238 1150 294
rect 1140 234 1150 238
rect 1210 234 1220 294
rect 758 228 832 234
rect -640 162 539 180
rect 594 175 668 181
rect 1170 134 1200 234
rect -1285 104 1200 134
<< via1 >>
rect -1420 870 -1400 920
rect -1400 870 -1360 920
rect -1420 860 -1360 870
rect 610 901 657 960
rect 657 901 670 960
rect 610 900 670 901
rect -870 690 -810 750
rect 1150 840 1210 850
rect 1150 790 1200 840
rect 1200 790 1210 840
rect -1410 430 -1350 490
rect -230 324 -220 374
rect -220 324 -170 374
rect 610 370 670 430
rect -230 314 -170 324
rect -880 190 -820 250
rect -770 284 -710 294
rect -770 234 -760 284
rect -760 234 -710 284
rect -40 234 10 284
rect 10 234 20 284
rect -40 224 20 234
rect 490 234 504 240
rect 504 234 550 240
rect 490 180 550 234
rect 1150 244 1200 294
rect 1200 244 1210 294
rect 1150 234 1210 244
<< metal2 >>
rect 620 1000 1290 1030
rect -1500 960 -1375 990
rect 620 970 650 1000
rect -1405 930 -1375 960
rect 610 960 670 970
rect -1420 920 -1360 930
rect 610 890 670 900
rect -1420 850 -1360 860
rect 1150 850 1210 860
rect 1210 800 1290 830
rect 1150 780 1210 790
rect -870 750 -810 760
rect -1500 720 -870 750
rect -870 680 -810 690
rect -1500 500 -1355 524
rect -1500 494 -1350 500
rect -1410 490 -1350 494
rect 625 484 1290 514
rect 625 440 655 484
rect -1410 420 -1350 430
rect 610 430 670 440
rect -230 374 -170 384
rect -1500 334 -740 364
rect -770 304 -740 334
rect 610 360 670 370
rect 1035 375 1290 405
rect 1035 319 1065 375
rect -230 304 -170 314
rect -770 294 -710 304
rect -880 250 -820 260
rect -1500 204 -880 234
rect -770 224 -710 234
rect -880 180 -820 190
rect -215 114 -185 304
rect -30 294 1065 319
rect -40 289 1065 294
rect 1150 294 1210 304
rect -40 284 20 289
rect -40 214 20 224
rect 490 240 550 250
rect 1210 254 1290 284
rect 1150 224 1210 234
rect 490 170 550 180
rect -1500 84 -185 114
rect 505 134 535 170
rect 505 104 1290 134
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -1436 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_1
timestamp 1710522493
transform 1 0 -792 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_2
timestamp 1710522493
transform 1 0 -1436 0 -1 1116
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 312 0 -1 1116
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -792 0 -1 1116
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 588 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_1
timestamp 1710522493
transform 1 0 -56 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_2
timestamp 1710522493
transform 1 0 588 0 -1 1116
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -148 0 1 28
box -38 -48 130 592
<< end >>
