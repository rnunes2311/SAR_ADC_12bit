magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< pwell >>
rect -201 -2382 201 2382
<< psubdiff >>
rect -165 2312 -69 2346
rect 69 2312 165 2346
rect -165 2250 -131 2312
rect 131 2250 165 2312
rect -165 -2312 -131 -2250
rect 131 -2312 165 -2250
rect -165 -2346 -69 -2312
rect 69 -2346 165 -2312
<< psubdiffcont >>
rect -69 2312 69 2346
rect -165 -2250 -131 2250
rect 131 -2250 165 2250
rect -69 -2346 69 -2312
<< xpolycontact >>
rect -35 1784 35 2216
rect -35 -2216 35 -1784
<< ppolyres >>
rect -35 -1784 35 1784
<< locali >>
rect -165 2312 -69 2346
rect 69 2312 165 2346
rect -165 2250 -131 2312
rect 131 2250 165 2312
rect -165 -2312 -131 -2250
rect 131 -2312 165 -2250
rect -165 -2346 -69 -2312
rect 69 -2346 165 -2312
<< viali >>
rect -19 1801 19 2198
rect -19 -2198 19 -1801
<< metal1 >>
rect -25 2198 25 2210
rect -25 1801 -19 2198
rect 19 1801 25 2198
rect -25 1789 25 1801
rect -25 -1801 25 -1789
rect -25 -2198 -19 -1801
rect 19 -2198 25 -1801
rect -25 -2210 25 -2198
<< properties >>
string FIXED_BBOX -148 -2329 148 2329
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 18.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 17.56k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
