magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< nwell >>
rect -641 -2855 641 2855
<< pmos >>
rect -445 1036 -345 2636
rect -287 1036 -187 2636
rect -129 1036 -29 2636
rect 29 1036 129 2636
rect 187 1036 287 2636
rect 345 1036 445 2636
rect -445 -800 -345 800
rect -287 -800 -187 800
rect -129 -800 -29 800
rect 29 -800 129 800
rect 187 -800 287 800
rect 345 -800 445 800
rect -445 -2636 -345 -1036
rect -287 -2636 -187 -1036
rect -129 -2636 -29 -1036
rect 29 -2636 129 -1036
rect 187 -2636 287 -1036
rect 345 -2636 445 -1036
<< pdiff >>
rect -503 2624 -445 2636
rect -503 1048 -491 2624
rect -457 1048 -445 2624
rect -503 1036 -445 1048
rect -345 2624 -287 2636
rect -345 1048 -333 2624
rect -299 1048 -287 2624
rect -345 1036 -287 1048
rect -187 2624 -129 2636
rect -187 1048 -175 2624
rect -141 1048 -129 2624
rect -187 1036 -129 1048
rect -29 2624 29 2636
rect -29 1048 -17 2624
rect 17 1048 29 2624
rect -29 1036 29 1048
rect 129 2624 187 2636
rect 129 1048 141 2624
rect 175 1048 187 2624
rect 129 1036 187 1048
rect 287 2624 345 2636
rect 287 1048 299 2624
rect 333 1048 345 2624
rect 287 1036 345 1048
rect 445 2624 503 2636
rect 445 1048 457 2624
rect 491 1048 503 2624
rect 445 1036 503 1048
rect -503 788 -445 800
rect -503 -788 -491 788
rect -457 -788 -445 788
rect -503 -800 -445 -788
rect -345 788 -287 800
rect -345 -788 -333 788
rect -299 -788 -287 788
rect -345 -800 -287 -788
rect -187 788 -129 800
rect -187 -788 -175 788
rect -141 -788 -129 788
rect -187 -800 -129 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 129 788 187 800
rect 129 -788 141 788
rect 175 -788 187 788
rect 129 -800 187 -788
rect 287 788 345 800
rect 287 -788 299 788
rect 333 -788 345 788
rect 287 -800 345 -788
rect 445 788 503 800
rect 445 -788 457 788
rect 491 -788 503 788
rect 445 -800 503 -788
rect -503 -1048 -445 -1036
rect -503 -2624 -491 -1048
rect -457 -2624 -445 -1048
rect -503 -2636 -445 -2624
rect -345 -1048 -287 -1036
rect -345 -2624 -333 -1048
rect -299 -2624 -287 -1048
rect -345 -2636 -287 -2624
rect -187 -1048 -129 -1036
rect -187 -2624 -175 -1048
rect -141 -2624 -129 -1048
rect -187 -2636 -129 -2624
rect -29 -1048 29 -1036
rect -29 -2624 -17 -1048
rect 17 -2624 29 -1048
rect -29 -2636 29 -2624
rect 129 -1048 187 -1036
rect 129 -2624 141 -1048
rect 175 -2624 187 -1048
rect 129 -2636 187 -2624
rect 287 -1048 345 -1036
rect 287 -2624 299 -1048
rect 333 -2624 345 -1048
rect 287 -2636 345 -2624
rect 445 -1048 503 -1036
rect 445 -2624 457 -1048
rect 491 -2624 503 -1048
rect 445 -2636 503 -2624
<< pdiffc >>
rect -491 1048 -457 2624
rect -333 1048 -299 2624
rect -175 1048 -141 2624
rect -17 1048 17 2624
rect 141 1048 175 2624
rect 299 1048 333 2624
rect 457 1048 491 2624
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect -491 -2624 -457 -1048
rect -333 -2624 -299 -1048
rect -175 -2624 -141 -1048
rect -17 -2624 17 -1048
rect 141 -2624 175 -1048
rect 299 -2624 333 -1048
rect 457 -2624 491 -1048
<< nsubdiff >>
rect -605 2785 -509 2819
rect 509 2785 605 2819
rect -605 2723 -571 2785
rect 571 2723 605 2785
rect -605 -2785 -571 -2723
rect 571 -2785 605 -2723
rect -605 -2819 -509 -2785
rect 509 -2819 605 -2785
<< nsubdiffcont >>
rect -509 2785 509 2819
rect -605 -2723 -571 2723
rect 571 -2723 605 2723
rect -509 -2819 509 -2785
<< poly >>
rect -445 2717 -345 2733
rect -445 2683 -429 2717
rect -361 2683 -345 2717
rect -445 2636 -345 2683
rect -287 2717 -187 2733
rect -287 2683 -271 2717
rect -203 2683 -187 2717
rect -287 2636 -187 2683
rect -129 2717 -29 2733
rect -129 2683 -113 2717
rect -45 2683 -29 2717
rect -129 2636 -29 2683
rect 29 2717 129 2733
rect 29 2683 45 2717
rect 113 2683 129 2717
rect 29 2636 129 2683
rect 187 2717 287 2733
rect 187 2683 203 2717
rect 271 2683 287 2717
rect 187 2636 287 2683
rect 345 2717 445 2733
rect 345 2683 361 2717
rect 429 2683 445 2717
rect 345 2636 445 2683
rect -445 989 -345 1036
rect -445 955 -429 989
rect -361 955 -345 989
rect -445 939 -345 955
rect -287 989 -187 1036
rect -287 955 -271 989
rect -203 955 -187 989
rect -287 939 -187 955
rect -129 989 -29 1036
rect -129 955 -113 989
rect -45 955 -29 989
rect -129 939 -29 955
rect 29 989 129 1036
rect 29 955 45 989
rect 113 955 129 989
rect 29 939 129 955
rect 187 989 287 1036
rect 187 955 203 989
rect 271 955 287 989
rect 187 939 287 955
rect 345 989 445 1036
rect 345 955 361 989
rect 429 955 445 989
rect 345 939 445 955
rect -445 881 -345 897
rect -445 847 -429 881
rect -361 847 -345 881
rect -445 800 -345 847
rect -287 881 -187 897
rect -287 847 -271 881
rect -203 847 -187 881
rect -287 800 -187 847
rect -129 881 -29 897
rect -129 847 -113 881
rect -45 847 -29 881
rect -129 800 -29 847
rect 29 881 129 897
rect 29 847 45 881
rect 113 847 129 881
rect 29 800 129 847
rect 187 881 287 897
rect 187 847 203 881
rect 271 847 287 881
rect 187 800 287 847
rect 345 881 445 897
rect 345 847 361 881
rect 429 847 445 881
rect 345 800 445 847
rect -445 -847 -345 -800
rect -445 -881 -429 -847
rect -361 -881 -345 -847
rect -445 -897 -345 -881
rect -287 -847 -187 -800
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -287 -897 -187 -881
rect -129 -847 -29 -800
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect -129 -897 -29 -881
rect 29 -847 129 -800
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 29 -897 129 -881
rect 187 -847 287 -800
rect 187 -881 203 -847
rect 271 -881 287 -847
rect 187 -897 287 -881
rect 345 -847 445 -800
rect 345 -881 361 -847
rect 429 -881 445 -847
rect 345 -897 445 -881
rect -445 -955 -345 -939
rect -445 -989 -429 -955
rect -361 -989 -345 -955
rect -445 -1036 -345 -989
rect -287 -955 -187 -939
rect -287 -989 -271 -955
rect -203 -989 -187 -955
rect -287 -1036 -187 -989
rect -129 -955 -29 -939
rect -129 -989 -113 -955
rect -45 -989 -29 -955
rect -129 -1036 -29 -989
rect 29 -955 129 -939
rect 29 -989 45 -955
rect 113 -989 129 -955
rect 29 -1036 129 -989
rect 187 -955 287 -939
rect 187 -989 203 -955
rect 271 -989 287 -955
rect 187 -1036 287 -989
rect 345 -955 445 -939
rect 345 -989 361 -955
rect 429 -989 445 -955
rect 345 -1036 445 -989
rect -445 -2683 -345 -2636
rect -445 -2717 -429 -2683
rect -361 -2717 -345 -2683
rect -445 -2733 -345 -2717
rect -287 -2683 -187 -2636
rect -287 -2717 -271 -2683
rect -203 -2717 -187 -2683
rect -287 -2733 -187 -2717
rect -129 -2683 -29 -2636
rect -129 -2717 -113 -2683
rect -45 -2717 -29 -2683
rect -129 -2733 -29 -2717
rect 29 -2683 129 -2636
rect 29 -2717 45 -2683
rect 113 -2717 129 -2683
rect 29 -2733 129 -2717
rect 187 -2683 287 -2636
rect 187 -2717 203 -2683
rect 271 -2717 287 -2683
rect 187 -2733 287 -2717
rect 345 -2683 445 -2636
rect 345 -2717 361 -2683
rect 429 -2717 445 -2683
rect 345 -2733 445 -2717
<< polycont >>
rect -429 2683 -361 2717
rect -271 2683 -203 2717
rect -113 2683 -45 2717
rect 45 2683 113 2717
rect 203 2683 271 2717
rect 361 2683 429 2717
rect -429 955 -361 989
rect -271 955 -203 989
rect -113 955 -45 989
rect 45 955 113 989
rect 203 955 271 989
rect 361 955 429 989
rect -429 847 -361 881
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect 361 847 429 881
rect -429 -881 -361 -847
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect 361 -881 429 -847
rect -429 -989 -361 -955
rect -271 -989 -203 -955
rect -113 -989 -45 -955
rect 45 -989 113 -955
rect 203 -989 271 -955
rect 361 -989 429 -955
rect -429 -2717 -361 -2683
rect -271 -2717 -203 -2683
rect -113 -2717 -45 -2683
rect 45 -2717 113 -2683
rect 203 -2717 271 -2683
rect 361 -2717 429 -2683
<< locali >>
rect -605 2785 -509 2819
rect 509 2785 605 2819
rect -605 2723 -571 2785
rect 571 2723 605 2785
rect -445 2683 -429 2717
rect -361 2683 -345 2717
rect -287 2683 -271 2717
rect -203 2683 -187 2717
rect -129 2683 -113 2717
rect -45 2683 -29 2717
rect 29 2683 45 2717
rect 113 2683 129 2717
rect 187 2683 203 2717
rect 271 2683 287 2717
rect 345 2683 361 2717
rect 429 2683 445 2717
rect -491 2624 -457 2640
rect -491 1032 -457 1048
rect -333 2624 -299 2640
rect -333 1032 -299 1048
rect -175 2624 -141 2640
rect -175 1032 -141 1048
rect -17 2624 17 2640
rect -17 1032 17 1048
rect 141 2624 175 2640
rect 141 1032 175 1048
rect 299 2624 333 2640
rect 299 1032 333 1048
rect 457 2624 491 2640
rect 457 1032 491 1048
rect -445 955 -429 989
rect -361 955 -345 989
rect -287 955 -271 989
rect -203 955 -187 989
rect -129 955 -113 989
rect -45 955 -29 989
rect 29 955 45 989
rect 113 955 129 989
rect 187 955 203 989
rect 271 955 287 989
rect 345 955 361 989
rect 429 955 445 989
rect -445 847 -429 881
rect -361 847 -345 881
rect -287 847 -271 881
rect -203 847 -187 881
rect -129 847 -113 881
rect -45 847 -29 881
rect 29 847 45 881
rect 113 847 129 881
rect 187 847 203 881
rect 271 847 287 881
rect 345 847 361 881
rect 429 847 445 881
rect -491 788 -457 804
rect -491 -804 -457 -788
rect -333 788 -299 804
rect -333 -804 -299 -788
rect -175 788 -141 804
rect -175 -804 -141 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 141 788 175 804
rect 141 -804 175 -788
rect 299 788 333 804
rect 299 -804 333 -788
rect 457 788 491 804
rect 457 -804 491 -788
rect -445 -881 -429 -847
rect -361 -881 -345 -847
rect -287 -881 -271 -847
rect -203 -881 -187 -847
rect -129 -881 -113 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 113 -881 129 -847
rect 187 -881 203 -847
rect 271 -881 287 -847
rect 345 -881 361 -847
rect 429 -881 445 -847
rect -445 -989 -429 -955
rect -361 -989 -345 -955
rect -287 -989 -271 -955
rect -203 -989 -187 -955
rect -129 -989 -113 -955
rect -45 -989 -29 -955
rect 29 -989 45 -955
rect 113 -989 129 -955
rect 187 -989 203 -955
rect 271 -989 287 -955
rect 345 -989 361 -955
rect 429 -989 445 -955
rect -491 -1048 -457 -1032
rect -491 -2640 -457 -2624
rect -333 -1048 -299 -1032
rect -333 -2640 -299 -2624
rect -175 -1048 -141 -1032
rect -175 -2640 -141 -2624
rect -17 -1048 17 -1032
rect -17 -2640 17 -2624
rect 141 -1048 175 -1032
rect 141 -2640 175 -2624
rect 299 -1048 333 -1032
rect 299 -2640 333 -2624
rect 457 -1048 491 -1032
rect 457 -2640 491 -2624
rect -445 -2717 -429 -2683
rect -361 -2717 -345 -2683
rect -287 -2717 -271 -2683
rect -203 -2717 -187 -2683
rect -129 -2717 -113 -2683
rect -45 -2717 -29 -2683
rect 29 -2717 45 -2683
rect 113 -2717 129 -2683
rect 187 -2717 203 -2683
rect 271 -2717 287 -2683
rect 345 -2717 361 -2683
rect 429 -2717 445 -2683
rect -605 -2785 -571 -2723
rect 571 -2785 605 -2723
rect -605 -2819 -509 -2785
rect 509 -2819 605 -2785
<< viali >>
rect -429 2683 -361 2717
rect -271 2683 -203 2717
rect -113 2683 -45 2717
rect 45 2683 113 2717
rect 203 2683 271 2717
rect 361 2683 429 2717
rect -491 1048 -457 2624
rect -333 1048 -299 2624
rect -175 1048 -141 2624
rect -17 1048 17 2624
rect 141 1048 175 2624
rect 299 1048 333 2624
rect 457 1048 491 2624
rect -429 955 -361 989
rect -271 955 -203 989
rect -113 955 -45 989
rect 45 955 113 989
rect 203 955 271 989
rect 361 955 429 989
rect -429 847 -361 881
rect -271 847 -203 881
rect -113 847 -45 881
rect 45 847 113 881
rect 203 847 271 881
rect 361 847 429 881
rect -491 -788 -457 788
rect -333 -788 -299 788
rect -175 -788 -141 788
rect -17 -788 17 788
rect 141 -788 175 788
rect 299 -788 333 788
rect 457 -788 491 788
rect -429 -881 -361 -847
rect -271 -881 -203 -847
rect -113 -881 -45 -847
rect 45 -881 113 -847
rect 203 -881 271 -847
rect 361 -881 429 -847
rect -429 -989 -361 -955
rect -271 -989 -203 -955
rect -113 -989 -45 -955
rect 45 -989 113 -955
rect 203 -989 271 -955
rect 361 -989 429 -955
rect -491 -2624 -457 -1048
rect -333 -2624 -299 -1048
rect -175 -2624 -141 -1048
rect -17 -2624 17 -1048
rect 141 -2624 175 -1048
rect 299 -2624 333 -1048
rect 457 -2624 491 -1048
rect -429 -2717 -361 -2683
rect -271 -2717 -203 -2683
rect -113 -2717 -45 -2683
rect 45 -2717 113 -2683
rect 203 -2717 271 -2683
rect 361 -2717 429 -2683
<< metal1 >>
rect -441 2717 -349 2723
rect -441 2683 -429 2717
rect -361 2683 -349 2717
rect -441 2677 -349 2683
rect -283 2717 -191 2723
rect -283 2683 -271 2717
rect -203 2683 -191 2717
rect -283 2677 -191 2683
rect -125 2717 -33 2723
rect -125 2683 -113 2717
rect -45 2683 -33 2717
rect -125 2677 -33 2683
rect 33 2717 125 2723
rect 33 2683 45 2717
rect 113 2683 125 2717
rect 33 2677 125 2683
rect 191 2717 283 2723
rect 191 2683 203 2717
rect 271 2683 283 2717
rect 191 2677 283 2683
rect 349 2717 441 2723
rect 349 2683 361 2717
rect 429 2683 441 2717
rect 349 2677 441 2683
rect -497 2624 -451 2636
rect -497 1048 -491 2624
rect -457 1048 -451 2624
rect -497 1036 -451 1048
rect -339 2624 -293 2636
rect -339 1048 -333 2624
rect -299 1048 -293 2624
rect -339 1036 -293 1048
rect -181 2624 -135 2636
rect -181 1048 -175 2624
rect -141 1048 -135 2624
rect -181 1036 -135 1048
rect -23 2624 23 2636
rect -23 1048 -17 2624
rect 17 1048 23 2624
rect -23 1036 23 1048
rect 135 2624 181 2636
rect 135 1048 141 2624
rect 175 1048 181 2624
rect 135 1036 181 1048
rect 293 2624 339 2636
rect 293 1048 299 2624
rect 333 1048 339 2624
rect 293 1036 339 1048
rect 451 2624 497 2636
rect 451 1048 457 2624
rect 491 1048 497 2624
rect 451 1036 497 1048
rect -441 989 -349 995
rect -441 955 -429 989
rect -361 955 -349 989
rect -441 949 -349 955
rect -283 989 -191 995
rect -283 955 -271 989
rect -203 955 -191 989
rect -283 949 -191 955
rect -125 989 -33 995
rect -125 955 -113 989
rect -45 955 -33 989
rect -125 949 -33 955
rect 33 989 125 995
rect 33 955 45 989
rect 113 955 125 989
rect 33 949 125 955
rect 191 989 283 995
rect 191 955 203 989
rect 271 955 283 989
rect 191 949 283 955
rect 349 989 441 995
rect 349 955 361 989
rect 429 955 441 989
rect 349 949 441 955
rect -441 881 -349 887
rect -441 847 -429 881
rect -361 847 -349 881
rect -441 841 -349 847
rect -283 881 -191 887
rect -283 847 -271 881
rect -203 847 -191 881
rect -283 841 -191 847
rect -125 881 -33 887
rect -125 847 -113 881
rect -45 847 -33 881
rect -125 841 -33 847
rect 33 881 125 887
rect 33 847 45 881
rect 113 847 125 881
rect 33 841 125 847
rect 191 881 283 887
rect 191 847 203 881
rect 271 847 283 881
rect 191 841 283 847
rect 349 881 441 887
rect 349 847 361 881
rect 429 847 441 881
rect 349 841 441 847
rect -497 788 -451 800
rect -497 -788 -491 788
rect -457 -788 -451 788
rect -497 -800 -451 -788
rect -339 788 -293 800
rect -339 -788 -333 788
rect -299 -788 -293 788
rect -339 -800 -293 -788
rect -181 788 -135 800
rect -181 -788 -175 788
rect -141 -788 -135 788
rect -181 -800 -135 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 135 788 181 800
rect 135 -788 141 788
rect 175 -788 181 788
rect 135 -800 181 -788
rect 293 788 339 800
rect 293 -788 299 788
rect 333 -788 339 788
rect 293 -800 339 -788
rect 451 788 497 800
rect 451 -788 457 788
rect 491 -788 497 788
rect 451 -800 497 -788
rect -441 -847 -349 -841
rect -441 -881 -429 -847
rect -361 -881 -349 -847
rect -441 -887 -349 -881
rect -283 -847 -191 -841
rect -283 -881 -271 -847
rect -203 -881 -191 -847
rect -283 -887 -191 -881
rect -125 -847 -33 -841
rect -125 -881 -113 -847
rect -45 -881 -33 -847
rect -125 -887 -33 -881
rect 33 -847 125 -841
rect 33 -881 45 -847
rect 113 -881 125 -847
rect 33 -887 125 -881
rect 191 -847 283 -841
rect 191 -881 203 -847
rect 271 -881 283 -847
rect 191 -887 283 -881
rect 349 -847 441 -841
rect 349 -881 361 -847
rect 429 -881 441 -847
rect 349 -887 441 -881
rect -441 -955 -349 -949
rect -441 -989 -429 -955
rect -361 -989 -349 -955
rect -441 -995 -349 -989
rect -283 -955 -191 -949
rect -283 -989 -271 -955
rect -203 -989 -191 -955
rect -283 -995 -191 -989
rect -125 -955 -33 -949
rect -125 -989 -113 -955
rect -45 -989 -33 -955
rect -125 -995 -33 -989
rect 33 -955 125 -949
rect 33 -989 45 -955
rect 113 -989 125 -955
rect 33 -995 125 -989
rect 191 -955 283 -949
rect 191 -989 203 -955
rect 271 -989 283 -955
rect 191 -995 283 -989
rect 349 -955 441 -949
rect 349 -989 361 -955
rect 429 -989 441 -955
rect 349 -995 441 -989
rect -497 -1048 -451 -1036
rect -497 -2624 -491 -1048
rect -457 -2624 -451 -1048
rect -497 -2636 -451 -2624
rect -339 -1048 -293 -1036
rect -339 -2624 -333 -1048
rect -299 -2624 -293 -1048
rect -339 -2636 -293 -2624
rect -181 -1048 -135 -1036
rect -181 -2624 -175 -1048
rect -141 -2624 -135 -1048
rect -181 -2636 -135 -2624
rect -23 -1048 23 -1036
rect -23 -2624 -17 -1048
rect 17 -2624 23 -1048
rect -23 -2636 23 -2624
rect 135 -1048 181 -1036
rect 135 -2624 141 -1048
rect 175 -2624 181 -1048
rect 135 -2636 181 -2624
rect 293 -1048 339 -1036
rect 293 -2624 299 -1048
rect 333 -2624 339 -1048
rect 293 -2636 339 -2624
rect 451 -1048 497 -1036
rect 451 -2624 457 -1048
rect 491 -2624 497 -1048
rect 451 -2636 497 -2624
rect -441 -2683 -349 -2677
rect -441 -2717 -429 -2683
rect -361 -2717 -349 -2683
rect -441 -2723 -349 -2717
rect -283 -2683 -191 -2677
rect -283 -2717 -271 -2683
rect -203 -2717 -191 -2683
rect -283 -2723 -191 -2717
rect -125 -2683 -33 -2677
rect -125 -2717 -113 -2683
rect -45 -2717 -33 -2683
rect -125 -2723 -33 -2717
rect 33 -2683 125 -2677
rect 33 -2717 45 -2683
rect 113 -2717 125 -2683
rect 33 -2723 125 -2717
rect 191 -2683 283 -2677
rect 191 -2717 203 -2683
rect 271 -2717 283 -2683
rect 191 -2723 283 -2717
rect 349 -2683 441 -2677
rect 349 -2717 361 -2683
rect 429 -2717 441 -2683
rect 349 -2723 441 -2717
<< properties >>
string FIXED_BBOX -588 -2802 588 2802
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.5 m 3 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
