magic
tech sky130A
magscale 1 2
timestamp 1711310191
<< metal3 >>
rect -986 1262 986 1290
rect -986 -1262 902 1262
rect 966 -1262 986 1262
rect -986 -1290 986 -1262
<< via3 >>
rect 902 -1262 966 1262
<< mimcap >>
rect -946 1210 654 1250
rect -946 -1210 -906 1210
rect 614 -1210 654 1210
rect -946 -1250 654 -1210
<< mimcapcontact >>
rect -906 -1210 614 1210
<< metal4 >>
rect 886 1262 982 1278
rect -907 1210 615 1211
rect -907 -1210 -906 1210
rect 614 -1210 615 1210
rect -907 -1211 615 -1210
rect 886 -1262 902 1262
rect 966 -1262 982 1262
rect 886 -1278 982 -1262
<< properties >>
string FIXED_BBOX -986 -1290 694 1290
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 8 l 12.5 val 207.79 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
