magic
tech sky130A
magscale 1 2
timestamp 1712048491
<< nwell >>
rect 1764 1494 3312 1620
rect 1790 1460 3312 1494
rect 1790 1450 3290 1460
<< nsubdiff >>
rect 1830 1520 1880 1580
rect 3170 1520 3230 1580
<< nsubdiffcont >>
rect 1880 1520 3170 1580
<< locali >>
rect 1840 1580 3210 1590
rect 1840 1520 1880 1580
rect 3170 1520 3210 1580
rect 1840 1460 3210 1520
rect 1865 1131 1884 1181
rect 2689 1131 2883 1181
rect 2372 810 2708 824
rect 2372 732 2390 810
rect 2700 732 2708 810
rect 2372 721 2708 732
rect 2635 -550 2647 -516
rect 2685 -550 2741 -516
rect 2152 -1606 3237 -1531
rect 2152 -1688 2196 -1606
rect 2780 -1610 2860 -1606
rect 3211 -1688 3237 -1606
rect 2152 -1715 3237 -1688
<< viali >>
rect 2940 1244 2993 1359
rect 1764 1131 1865 1181
rect 1930 1060 1970 1220
rect 2050 1131 2180 1171
rect 2280 1131 2320 1171
rect 2360 1131 2400 1171
rect 2480 1131 2610 1181
rect 2390 732 2700 810
rect 2647 -550 2685 -516
rect 2196 -1610 2780 -1606
rect 2860 -1610 3211 -1606
rect 2196 -1688 3211 -1610
<< metal1 >>
rect 1810 1570 3260 1620
rect 1810 1550 3250 1570
rect 1810 1540 2250 1550
rect 1810 1480 1860 1540
rect 1920 1480 2050 1540
rect 2110 1490 2250 1540
rect 2310 1490 2450 1550
rect 2510 1490 2680 1550
rect 2740 1490 3140 1550
rect 3200 1490 3250 1550
rect 3360 1540 3400 1580
rect 2110 1480 3250 1490
rect 1810 1440 3250 1480
rect 1810 1420 3260 1440
rect 3570 1400 3610 1432
rect 2920 1320 2930 1380
rect 2990 1359 3000 1380
rect 2920 1300 2940 1320
rect 2920 1240 2930 1300
rect 2993 1244 3000 1359
rect 3090 1260 3100 1320
rect 3160 1310 3170 1320
rect 3200 1310 3210 1320
rect 3160 1270 3210 1310
rect 3160 1260 3170 1270
rect 3200 1260 3210 1270
rect 3270 1310 3280 1320
rect 3504 1312 3610 1400
rect 3716 1312 3822 1432
rect 3900 1330 3910 1390
rect 3970 1330 3980 1390
rect 3270 1270 3380 1310
rect 3270 1260 3280 1270
rect 2990 1240 3000 1244
rect 3900 1240 3910 1300
rect 3970 1240 3980 1300
rect 2934 1232 2999 1240
rect 1924 1220 1976 1232
rect 1924 1210 1930 1220
rect 1970 1210 1976 1220
rect 1752 1181 1877 1187
rect 1752 1131 1764 1181
rect 1865 1131 1877 1181
rect 1910 1150 1920 1210
rect 1980 1150 1990 1210
rect 2040 1180 2190 1190
rect 2460 1181 2630 1200
rect 1752 1125 1877 1131
rect 1924 1120 1930 1150
rect 1970 1120 1976 1150
rect 2030 1120 2040 1180
rect 2100 1171 2130 1180
rect 2100 1120 2130 1131
rect 2190 1120 2200 1180
rect 2260 1121 2270 1181
rect 2330 1121 2360 1181
rect 2420 1121 2430 1181
rect 2460 1131 2480 1181
rect 2610 1170 2630 1181
rect 2840 1170 2850 1180
rect 2610 1140 2850 1170
rect 2610 1131 2630 1140
rect 2460 1120 2630 1131
rect 2840 1120 2850 1140
rect 2910 1120 2930 1180
rect 2990 1170 3000 1180
rect 2990 1140 3040 1170
rect 2990 1120 3000 1140
rect 1910 1060 1920 1120
rect 1980 1060 1990 1120
rect 2040 1110 2190 1120
rect 1924 1048 1976 1060
rect 2060 -1280 2150 920
rect 2351 810 2712 816
rect 2351 732 2390 810
rect 2700 800 2712 810
rect 2710 740 2720 800
rect 2700 732 2720 740
rect 2351 726 2720 732
rect 2351 100 2412 726
rect 2660 600 2720 726
rect 2750 680 2760 740
rect 2820 680 2860 740
rect 2920 680 3100 740
rect 2750 670 3100 680
rect 2660 530 2830 600
rect 3090 520 3100 580
rect 3160 520 3170 580
rect 2440 221 2487 479
rect 2595 465 2740 495
rect 2520 270 2530 330
rect 2590 270 2610 330
rect 2670 270 2680 330
rect 2440 174 2670 221
rect 2639 112 2670 174
rect 2351 -80 2500 100
rect 2595 83 2670 112
rect 2604 41 2670 83
rect 2200 -350 2210 -290
rect 2270 -350 2280 -290
rect 2200 -380 2280 -350
rect 2200 -440 2210 -380
rect 2270 -440 2280 -380
rect 2520 -390 2560 -150
rect 2710 -305 2740 465
rect 3090 430 3100 490
rect 3160 430 3170 490
rect 2770 170 2780 230
rect 2840 170 2850 230
rect 2970 170 2980 230
rect 3040 170 3050 230
rect 2770 80 2780 140
rect 2840 80 2850 140
rect 2970 80 2980 140
rect 3040 80 3050 140
rect 2880 -60 2890 0
rect 2950 -60 2960 0
rect 3070 -60 3080 0
rect 3140 -60 3150 0
rect 2880 -150 2890 -90
rect 2950 -150 2960 -90
rect 3070 -150 3080 -90
rect 3140 -150 3150 -90
rect 2830 -305 2840 -280
rect 2710 -335 2840 -305
rect 2830 -340 2840 -335
rect 2900 -340 2930 -280
rect 2990 -340 3000 -280
rect 2520 -430 3070 -390
rect 2230 -1170 2260 -440
rect 2620 -550 2630 -490
rect 2690 -550 2720 -490
rect 2780 -550 2790 -490
rect 2620 -560 2790 -550
rect 2860 -570 2870 -510
rect 2940 -570 2950 -510
rect 2860 -600 2950 -570
rect 2860 -660 2870 -600
rect 2940 -660 2950 -600
rect 3030 -570 3070 -430
rect 3030 -620 3260 -570
rect 2650 -730 2660 -670
rect 2720 -730 2730 -670
rect 2650 -820 2660 -760
rect 2720 -820 2730 -760
rect 2890 -880 2920 -660
rect 3180 -680 3190 -620
rect 3250 -680 3260 -620
rect 3180 -720 3260 -680
rect 3180 -780 3190 -720
rect 3250 -780 3260 -720
rect 2290 -1000 2300 -920
rect 2370 -1000 2390 -920
rect 2460 -1000 2470 -920
rect 2860 -950 2870 -880
rect 2940 -950 2950 -880
rect 3080 -940 3090 -880
rect 3150 -940 3160 -880
rect 2860 -980 2950 -950
rect 3090 -970 3160 -940
rect 2230 -1220 2370 -1170
rect 2400 -1250 2430 -1000
rect 2860 -1050 2870 -980
rect 2940 -1050 2950 -980
rect 3080 -1030 3090 -970
rect 3150 -1030 3160 -970
rect 2060 -1420 2280 -1280
rect 2360 -1320 2430 -1250
rect 2370 -1370 2430 -1320
rect 2470 -1160 2589 -1134
rect 2470 -1340 2610 -1160
rect 2470 -1388 2600 -1340
rect 2470 -1390 2616 -1388
rect 2060 -1527 2150 -1420
rect 2470 -1527 2550 -1390
rect 2780 -1527 2860 -1164
rect 2930 -1420 3020 -1160
rect 2930 -1527 3010 -1420
rect 2060 -1606 3237 -1527
rect 3388 -1590 3494 -1470
rect 3612 -1590 3718 -1470
rect 3842 -1590 3948 -1470
rect 2060 -1620 2196 -1606
rect 2780 -1610 2860 -1606
rect 2060 -1680 2180 -1620
rect 2060 -1688 2196 -1680
rect 3211 -1688 3237 -1606
rect 2060 -1740 3237 -1688
<< via1 >>
rect 1860 1480 1920 1540
rect 2050 1480 2110 1540
rect 2250 1490 2310 1550
rect 2450 1490 2510 1550
rect 2680 1490 2740 1550
rect 3140 1490 3200 1550
rect 2930 1359 2990 1380
rect 2930 1320 2940 1359
rect 2940 1320 2990 1359
rect 2930 1244 2940 1300
rect 2940 1244 2990 1300
rect 3100 1260 3160 1320
rect 3210 1260 3270 1320
rect 3910 1330 3970 1390
rect 2930 1240 2990 1244
rect 3910 1240 3970 1300
rect 1920 1150 1930 1210
rect 1930 1150 1970 1210
rect 1970 1150 1980 1210
rect 2040 1171 2100 1180
rect 2130 1171 2190 1180
rect 2040 1131 2050 1171
rect 2050 1131 2100 1171
rect 2130 1131 2180 1171
rect 2180 1131 2190 1171
rect 2040 1120 2100 1131
rect 2130 1120 2190 1131
rect 2270 1171 2330 1181
rect 2270 1131 2280 1171
rect 2280 1131 2320 1171
rect 2320 1131 2330 1171
rect 2270 1121 2330 1131
rect 2360 1171 2420 1181
rect 2360 1131 2400 1171
rect 2400 1131 2420 1171
rect 2360 1121 2420 1131
rect 2850 1120 2910 1180
rect 2930 1120 2990 1180
rect 1920 1060 1930 1120
rect 1930 1060 1970 1120
rect 1970 1060 1980 1120
rect 2400 740 2460 800
rect 2530 740 2590 800
rect 2650 740 2700 800
rect 2700 740 2710 800
rect 2760 680 2820 740
rect 2860 680 2920 740
rect 3100 520 3160 580
rect 2530 270 2590 330
rect 2610 270 2670 330
rect 2210 -350 2270 -290
rect 2210 -440 2270 -380
rect 3100 430 3160 490
rect 2780 170 2840 230
rect 2980 170 3040 230
rect 2780 80 2840 140
rect 2980 80 3040 140
rect 2890 -60 2950 0
rect 3080 -60 3140 0
rect 2890 -150 2950 -90
rect 3080 -150 3140 -90
rect 2840 -340 2900 -280
rect 2930 -340 2990 -280
rect 2630 -516 2690 -490
rect 2630 -550 2647 -516
rect 2647 -550 2685 -516
rect 2685 -550 2690 -516
rect 2720 -550 2780 -490
rect 2870 -570 2940 -510
rect 2870 -660 2940 -600
rect 2660 -730 2720 -670
rect 2660 -820 2720 -760
rect 3190 -680 3250 -620
rect 3190 -780 3250 -720
rect 2300 -1000 2370 -920
rect 2390 -1000 2460 -920
rect 2870 -950 2940 -880
rect 3090 -940 3150 -880
rect 2870 -1050 2940 -980
rect 3090 -1030 3150 -970
rect 2180 -1680 2196 -1620
rect 2196 -1680 2240 -1620
rect 2380 -1680 2440 -1620
rect 2600 -1680 2660 -1620
rect 2810 -1680 2870 -1620
rect 3050 -1680 3110 -1620
<< metal2 >>
rect 1810 1550 2846 1620
rect 1810 1540 2250 1550
rect 1810 1480 1860 1540
rect 1920 1480 2050 1540
rect 2110 1490 2250 1540
rect 2310 1490 2450 1550
rect 2510 1490 2680 1550
rect 2740 1490 2846 1550
rect 2110 1480 2846 1490
rect 1810 1420 2846 1480
rect 3056 1550 3260 1620
rect 3056 1490 3140 1550
rect 3200 1490 3260 1550
rect 3056 1420 3260 1490
rect 1930 1260 2280 1290
rect 1930 1220 1970 1260
rect 1920 1210 1980 1220
rect 2240 1191 2280 1260
rect 1920 1120 1980 1150
rect 1920 1050 1980 1060
rect 2040 1180 2190 1190
rect 2100 1120 2130 1180
rect 2040 1110 2190 1120
rect 2240 1181 2420 1191
rect 2240 1121 2270 1181
rect 2330 1121 2360 1181
rect 2240 1111 2420 1121
rect 2040 -940 2080 1110
rect 2240 710 2280 1111
rect 2630 810 2710 1420
rect 3910 1400 4020 1430
rect 3910 1390 3950 1400
rect 2930 1380 2990 1390
rect 2930 1300 2990 1320
rect 3100 1320 3160 1330
rect 3210 1320 3270 1330
rect 3160 1270 3210 1310
rect 3100 1250 3160 1260
rect 3210 1250 3270 1260
rect 3910 1300 4020 1330
rect 2930 1230 2990 1240
rect 2850 1180 2990 1190
rect 2910 1120 2930 1180
rect 2850 1110 2990 1120
rect 2400 800 2710 810
rect 2460 740 2530 800
rect 2590 740 2650 800
rect 2400 730 2710 740
rect 2760 740 2920 750
rect 2120 700 2280 710
rect 2120 680 2760 700
rect 2820 680 2860 740
rect 2120 670 2920 680
rect 2120 -510 2160 670
rect 2530 330 2670 340
rect 2220 270 2530 310
rect 2590 270 2610 330
rect 2950 310 2990 1110
rect 3220 730 3260 1250
rect 3910 1230 3950 1240
rect 3910 1190 4020 1230
rect 3110 690 3260 730
rect 3110 590 3150 690
rect 3100 580 3160 590
rect 3100 490 3160 520
rect 3100 420 3160 430
rect 2670 270 2990 310
rect 2220 -280 2260 270
rect 2530 260 2670 270
rect 2780 230 2840 240
rect 2980 230 3040 240
rect 2840 170 2980 210
rect 2780 140 3040 170
rect 2840 90 2980 140
rect 2780 70 2840 80
rect 2980 70 3040 80
rect 2890 0 2950 10
rect 3080 0 3140 10
rect 2950 -60 3080 -20
rect 2890 -90 3140 -60
rect 2950 -140 3080 -90
rect 2890 -160 2950 -150
rect 3080 -160 3140 -150
rect 2840 -280 2990 -270
rect 2210 -290 2270 -280
rect 2900 -340 2930 -280
rect 2840 -350 2990 -340
rect 2210 -380 2270 -350
rect 2210 -450 2270 -440
rect 2630 -490 2780 -480
rect 2120 -550 2630 -510
rect 2690 -550 2720 -490
rect 2880 -500 2930 -350
rect 2630 -560 2780 -550
rect 2870 -510 2940 -500
rect 2870 -600 2940 -570
rect 2660 -670 2720 -660
rect 2870 -670 2940 -660
rect 3190 -620 3250 -610
rect 3190 -720 3250 -680
rect 2660 -760 3190 -730
rect 2720 -770 3190 -760
rect 3920 -730 3960 1190
rect 3250 -770 3960 -730
rect 3190 -790 3250 -780
rect 2660 -830 2720 -820
rect 2870 -880 2940 -870
rect 2300 -920 2460 -910
rect 2040 -980 2300 -940
rect 2370 -1000 2390 -920
rect 2460 -950 2870 -930
rect 3090 -880 3150 -870
rect 2940 -940 3090 -930
rect 2940 -950 3150 -940
rect 2460 -970 3150 -950
rect 2460 -980 3090 -970
rect 2460 -1000 2870 -980
rect 2300 -1010 2460 -1000
rect 2940 -1000 3090 -980
rect 3090 -1040 3150 -1030
rect 2870 -1060 2940 -1050
rect 2120 -1620 3237 -1527
rect 2120 -1680 2180 -1620
rect 2240 -1680 2380 -1620
rect 2440 -1680 2600 -1620
rect 2660 -1680 2810 -1620
rect 2870 -1680 2910 -1620
rect 2970 -1680 3050 -1620
rect 3110 -1680 3237 -1620
rect 2120 -1740 3237 -1680
<< via2 >>
rect 3950 1390 4020 1400
rect 3950 1330 3970 1390
rect 3970 1330 4020 1390
rect 3950 1240 3970 1300
rect 3970 1240 4020 1300
rect 3950 1230 4020 1240
rect 2810 -1680 2870 -1620
rect 2910 -1680 2970 -1620
<< metal3 >>
rect 3940 1400 4030 1420
rect 3940 1330 3950 1400
rect 4020 1330 4030 1400
rect 3940 1300 4030 1330
rect 3940 1230 3950 1300
rect 4020 1230 4030 1300
rect 3940 1210 4030 1230
rect 2790 -1610 2990 -1600
rect 2790 -1690 2800 -1610
rect 2880 -1690 2900 -1610
rect 2980 -1690 2990 -1610
<< via3 >>
rect 3950 1330 4020 1400
rect 3950 1230 4020 1300
rect 2800 -1620 2880 -1610
rect 2800 -1680 2810 -1620
rect 2810 -1680 2870 -1620
rect 2870 -1680 2880 -1620
rect 2800 -1690 2880 -1680
rect 2900 -1620 2980 -1610
rect 2900 -1680 2910 -1620
rect 2910 -1680 2970 -1620
rect 2970 -1680 2980 -1620
rect 2900 -1690 2980 -1680
<< metal4 >>
rect 3940 1400 4030 1420
rect 3940 1360 3950 1400
rect 3720 1330 3950 1360
rect 4020 1330 4030 1400
rect 3720 1300 4030 1330
rect 3720 1260 3950 1300
rect 3940 1230 3950 1260
rect 4020 1230 4030 1300
rect 3940 1210 4030 1230
rect 2840 -1600 2940 -1330
rect 2790 -1610 2990 -1600
rect 2790 -1690 2800 -1610
rect 2880 -1690 2900 -1610
rect 2980 -1690 2990 -1610
rect 2790 -1700 2990 -1690
use sky130_fd_pr__pfet_01v8_LG57AL  sky130_fd_pr__pfet_01v8_LG57AL_0
timestamp 1711315072
transform -1 0 2546 0 1 431
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LG57AL  sky130_fd_pr__pfet_01v8_LG57AL_1
timestamp 1711315072
transform -1 0 2546 0 1 -31
box -211 -284 211 284
use sky130_fd_pr__res_high_po_0p35_GKNPGE  sky130_fd_pr__res_high_po_0p35_GKNPGE_0
timestamp 1711308867
transform 1 0 3942 0 1 -71
box -35 -1666 35 1666
use sky130_fd_sc_hd__inv_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 1802 0 1 916
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 2078 0 1 916
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  x3
timestamp 1710522493
transform 1 0 2538 0 1 916
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 2814 0 1 916
box -38 -48 498 592
use sky130_fd_pr__cap_mim_m3_1_U4WBBP  XC2
timestamp 1711312488
transform 0 1 3020 -1 0 56
box -1436 -840 1436 840
use sky130_fd_pr__nfet_01v8_6ENSLP  XM1
timestamp 1711313579
transform 1 0 2695 0 1 -988
box -263 -610 263 610
use sky130_fd_pr__pfet_01v8_XGJYDL  XM2
timestamp 1711314126
transform 1 0 2963 0 1 241
box -311 -619 311 619
use sky130_fd_pr__nfet_01v8_J4Y94J  XM4
timestamp 1711311798
transform 1 0 3063 0 1 -1019
box -211 -579 211 579
use sky130_fd_pr__nfet_01v8_8XY3SE  XM6
timestamp 1711315072
transform -1 0 2327 0 1 -1319
box -211 -279 211 279
use sky130_fd_pr__res_high_po_0p35_GKNPGE  XR1
timestamp 1711308867
transform 1 0 3382 0 1 -71
box -35 -1666 35 1666
use sky130_fd_pr__res_high_po_0p35_GKNPGE  XR2
timestamp 1711308867
transform 1 0 3494 0 1 -71
box -35 -1666 35 1666
use sky130_fd_pr__res_high_po_0p35_GKNPGE  XR3
timestamp 1711308867
transform 1 0 3606 0 1 -71
box -35 -1666 35 1666
use sky130_fd_pr__res_high_po_0p35_GKNPGE  XR4
timestamp 1711308867
transform 1 0 3718 0 1 -71
box -35 -1666 35 1666
use sky130_fd_pr__res_high_po_0p35_GKNPGE  XR5
timestamp 1711308867
transform 1 0 3830 0 1 -71
box -35 -1666 35 1666
<< labels >>
rlabel metal1 3360 1540 3400 1580 1 t_10ns
port 1 n
rlabel metal1 3410 -1550 3470 -1500 1 t_8p5ns
port 2 n
rlabel metal1 3520 1330 3580 1370 1 t_7ns
port 3 n
rlabel metal1 3630 -1550 3690 -1510 1 t_5p3ns
port 4 n
rlabel metal1 3740 1350 3800 1390 1 t_3p7ns
port 5 n
rlabel metal1 3850 -1550 3910 -1510 1 t_2p1ns
port 6 n
flabel metal2 2220 -1730 2420 -1530 0 FreeSans 1280 0 0 0 VSS
port 9 nsew
flabel metal1 1910 1420 2110 1620 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
rlabel metal1 1764 1131 1819 1181 1 IN
port 8 n
rlabel metal2 2930 1280 2990 1340 1 OUT
port 7 n
<< end >>
