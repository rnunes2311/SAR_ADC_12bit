magic
tech sky130A
magscale 1 2
timestamp 1713726127
<< metal1 >>
rect 3760 10430 3770 10530
rect 3940 10430 3950 10530
rect 4090 9890 4100 9990
rect 4270 9890 4280 9990
rect 3760 9340 3770 9440
rect 3940 9340 3950 9440
rect 4090 8800 4100 8900
rect 4270 8800 4280 8900
rect 3760 8250 3770 8350
rect 3940 8250 3950 8350
rect 4090 7710 4100 7810
rect 4270 7710 4280 7810
rect 3760 7170 3770 7270
rect 3940 7170 3950 7270
<< via1 >>
rect 3770 10430 3940 10530
rect 4100 9890 4270 9990
rect 3770 9340 3940 9440
rect 4100 8800 4270 8900
rect 3770 8250 3940 8350
rect 4100 7710 4270 7810
rect 3770 7170 3940 7270
<< metal2 >>
rect 3770 10530 3940 10540
rect 3770 9440 3940 10430
rect 3770 8350 3940 9340
rect 3770 7270 3940 8250
rect 4100 9990 4270 10000
rect 4100 8900 4270 9890
rect 4100 7810 4270 8800
rect 4100 7700 4270 7710
rect 3770 7160 3940 7170
use bbm_unit  bbm_unit_0
timestamp 1713724235
transform -1 0 4607 0 1 9363
box -890 -20 626 620
use bbm_unit_x2  bbm_unit_x2_2
array 0 0 1516 0 2 1088
timestamp 1713724073
transform 1 0 3431 0 1 7187
box -890 -20 626 1164
use bbm_unit_x2  bbm_unit_x2_3
array 0 0 1516 0 1 1088
timestamp 1713724073
transform -1 0 4607 0 1 7187
box -890 -20 626 1164
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5123 0 -1 10479
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 4019 0 -1 10479
box -38 -48 1142 592
<< end >>
