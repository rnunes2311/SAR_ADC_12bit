** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/top_level_differential_sim.sch

* Skywater 130 nm PDK models
.lib /opt/pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ff

* Models for diodes, resistors, capacitors
*.include /opt/pdk/share/pdk/sky130A/libs.tech/combined/continuous/models_diodes.spice

*.include /opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sky130_fd_pr__model__r+c.model.spice

* Models for standard digital cells
.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

* C extraction spice netlist for CDAC
.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/subcells/CDAC/CDAC_mim_12bit_flat.spice

* Spice netlist for state machine generated by openlane
.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/subcells/state_machine/state_machine_openlane_generated.spice

* C or RC extraction of the SAR ADC
*.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/SAR_ADC_12bit_flat.spice

**.subckt top_level_differential_sim
V1 VDD VSS {VDD}
.save i(v1)
V2 net1 VSS {VCM}
.save i(v2)
V3 net2 VSS {VREF}
.save i(v3)
V4 VSS GND 0
V7 START VSS pulse(0 1.8 20n 1n 1n 100n 1u)
V8 RST_Z VSS pwl(0 0 10n 0 10.1n 1.8)
V5 net4 VSS pwl(0 0.4000 1u 0.4000 1.001u 0.8000 2u 0.8000 2.001u 0.9599 3u 0.9599 3.001u 0.2401 4u 0.2401 4.001u 0.0186 5u 0.0186
+ 5.001u 1.1814 6u 1.1814)
x1 VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START EN_OFFSET_CAL CLK VREF_GND
+ SINGLE_ENDED SAR_ADC_12bit
R1 net1 VCM 500 m=1
V9 CLK VSS pulse(0 1.8 0 1n 1n 40n 50n)
V6 net5 VSS pwl(0 0.8000 1u 0.8000 1.001u 0.4000 2u 0.4000 2.001u 0.2401 3u 0.2401 3.001u 0.9599 4u 0.9599 4.001u 1.1814 5u 1.1814
+ 5.001u 0.0186 6u 0.0186)
V10 net3 VSS {VREF_GND}
.save i(v10)
R6 net2 VREF 500 m=1
R7 net3 VREF_GND 500 m=1
R8 net4 VIN_P 500 m=1
R9 net5 VIN_N 500 m=1
V11 EN_OFFSET_CAL VSS pwl(0 0 3u 0 3.001u 1.8)
V12 SINGLE_ENDED VSS 0
**** begin user architecture code


* Supply, common mode and reference voltage
.param VDD = 1.7
.param VREF = 1.2
.param VREF_GND = 0
.param VCM = 0.5

*.save all

* Control signals
.save start rst_z clk en_offset_cal

* Input signals
.save vin_p vin_n

* Reference, supply
.save vref vref_gnd vcm vdd

* Output signals
.save clk_data data[5] data[4] data[3] data[2] data[1] data[0]

* Internal signals
.save x1.vdac_p x1.vdac_n x1.vdac_pi x1.vdac_ni x1.smpl x1.en_comp x1.comp_p x1.comp_n x1.cal_p x1.cal_n
.save x1.en_vin_bstr_p x1.en_vin_bstr_n
.save x1.c10_p_btm x1.c9_p_btm x1.c8_p_btm x1.c7_p_btm x1.c6_p_btm x1.c5_p_btm x1.c4_p_btm x1.c3_p_btm x1.c2_p_btm x1.c1_p_btm x1.c0_p_btm x1.C0_dummy_p_btm
.save x1.c10_n_btm x1.c9_n_btm x1.c8_n_btm x1.c7_n_btm x1.c6_n_btm x1.c5_n_btm x1.c4_n_btm x1.c3_n_btm x1.c2_n_btm x1.c1_n_btm x1.c0_n_btm x1.C0_dummy_n_btm

.option GMIN=1e-12 reltol=1e-5
.control
		set temp = 0
		set tnom = 0
		set num_threads=8
		tran 10n 6u
		write top_level_differential_sim.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  ../schematic/SAR_ADC_12bit.sym # of pins=14
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/SAR_ADC_12bit.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/SAR_ADC_12bit.sch
.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START
+ EN_OFFSET_CAL CLK VREF_GND SINGLE_ENDED
*.ipin VIN_P
*.ipin VDD
*.ipin VREF
*.ipin VCM
*.ipin VSS
*.ipin VIN_N
*.ipin RST_Z
*.ipin START
*.opin CLK_DATA
*.opin DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]
*.ipin EN_OFFSET_CAL
*.ipin CLK
*.ipin VREF_GND
*.ipin SINGLE_ENDED
x1 C0_dummy_N_btm C0_N_btm C1_N_btm C2_N_btm C3_N_btm C4_N_btm C5_N_btm C6_N_btm C7_N_btm C8_N_btm C9_N_btm C10_N_btm VDAC_N VSS
+ CDAC_12bit
x2 C0_dummy_P_btm C0_P_btm C1_P_btm C2_P_btm C3_P_btm C4_P_btm C5_P_btm C6_P_btm C7_P_btm C8_P_btm C9_P_btm C10_P_btm VDAC_P VSS
+ CDAC_12bit
x3 VCM VREF_GND VREF VIN_P EN_VIN_BSTR_P EN_REF_Z_P[10] EN_REF_Z_P[9] EN_REF_Z_P[8] EN_REF_Z_P[7] EN_REF_Z_P[6] EN_REF_Z_P[5]
+ EN_REF_Z_P[4] EN_REF_Z_P[3] EN_REF_Z_P[2] EN_REF_Z_P[1] EN_REF_Z_P[0] EN_VSS_P[10] EN_VSS_P[9] EN_VSS_P[8] EN_VSS_P[7] EN_VSS_P[6] EN_VSS_P[5]
+ EN_VSS_P[4] EN_VSS_P[3] EN_VSS_P[2] EN_VSS_P[1] EN_VSS_P[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3]
+ EN_VCM[2] EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY C8_P_btm C7_P_btm C0_P_btm C6_P_btm C5_P_btm C0_dummy_P_btm C4_P_btm C3_P_btm VDAC_P
+ C10_P_btm C9_P_btm C2_P_btm C1_P_btm VDD VSS switches
x4 VCM VREF_GND VREF VIN_N EN_VIN_BSTR_N EN_REF_Z_N[10] EN_REF_Z_N[9] EN_REF_Z_N[8] EN_REF_Z_N[7] EN_REF_Z_N[6] EN_REF_Z_N[5]
+ EN_REF_Z_N[4] EN_REF_Z_N[3] EN_REF_Z_N[2] EN_REF_Z_N[1] EN_REF_Z_N[0] EN_VSS_N[10] EN_VSS_N[9] EN_VSS_N[8] EN_VSS_N[7] EN_VSS_N[6] EN_VSS_N[5]
+ EN_VSS_N[4] EN_VSS_N[3] EN_VSS_N[2] EN_VSS_N[1] EN_VSS_N[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3]
+ EN_VCM[2] EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY C8_N_btm C7_N_btm C0_N_btm C6_N_btm C5_N_btm C0_dummy_N_btm C4_N_btm C3_N_btm VDAC_N
+ C10_N_btm C9_N_btm C2_N_btm C1_N_btm VDD VSS switches
x5 VDAC_N VDAC_P VDD RST_Z VDAC_Pi VDAC_Ni VSS CAL_P CAL_N preamplifier
x6 VDD VDAC_Pi VDAC_Ni EN_COMP COMP_P COMP_N VSS latched_comparator
x7 VDD COMP_P EN_COMP CAL_P CAL_N EN_VOS_CAL VSS OFFSET_CAL_CYCLE offset_calibration
x8 VDD VSS RST_Z START COMP_P SMPL EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2]
+ EN_VCM[1] EN_VCM[0] EN_COMP SMPL_ON_P SMPL_ON_N EN_VCM_DUMMY EN_VCM_SW EN_OFFSET_CAL OFFSET_CAL_CYCLE EN_VOS_CAL CLK_DATA DATA[5] DATA[4]
+ DATA[3] DATA[2] DATA[1] DATA[0] EN_VSS_N[10] EN_VSS_N[9] EN_VSS_N[8] EN_VSS_N[7] EN_VSS_N[6] EN_VSS_N[5] EN_VSS_N[4] EN_VSS_N[3]
+ EN_VSS_N[2] EN_VSS_N[1] EN_VSS_N[0] EN_REF_Z_N[10] EN_REF_Z_N[9] EN_REF_Z_N[8] EN_REF_Z_N[7] EN_REF_Z_N[6] EN_REF_Z_N[5] EN_REF_Z_N[4]
+ EN_REF_Z_N[3] EN_REF_Z_N[2] EN_REF_Z_N[1] EN_REF_Z_N[0] EN_VSS_P_BBM[10] EN_VSS_P_BBM[9] EN_VSS_P_BBM[8] EN_VSS_P_BBM[7] EN_VSS_P_BBM[6]
+ EN_VSS_P_BBM[5] EN_VSS_P_BBM[4] EN_VSS_P_BBM[3] EN_VSS_P_BBM[2] EN_VSS_P_BBM[1] EN_VSS_P_BBM[0] EN_REF_Z_P_BBM[10] EN_REF_Z_P_BBM[9]
+ EN_REF_Z_P_BBM[8] EN_REF_Z_P_BBM[7] EN_REF_Z_P_BBM[6] EN_REF_Z_P_BBM[5] EN_REF_Z_P_BBM[4] EN_REF_Z_P_BBM[3] EN_REF_Z_P_BBM[2] EN_REF_Z_P_BBM[1]
+ EN_REF_Z_P_BBM[0] CLK EN_VCM_SW EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2] EN_VCM[1] EN_VCM[0]
+ SINGLE_ENDED state_machine
x11 VDD VSS VIN_P SMPL_ON_P SMPL EN_VIN_BSTR_P bootstrap
x12 VDD VSS VIN_N SMPL_ON_N SMPL EN_VIN_BSTR_N bootstrap
x9 EN_VSS_P_BBM[10] EN_VSS_P_BBM[9] EN_VSS_P_BBM[8] EN_VSS_P_BBM[7] EN_VSS_P_BBM[6] EN_VSS_P_BBM[5] EN_VSS_P_BBM[4]
+ EN_VSS_P_BBM[3] EN_VSS_P_BBM[2] EN_VSS_P_BBM[1] EN_VSS_P_BBM[0] VDD VSS EN_VSS_P[10] EN_VSS_P[9] EN_VSS_P[8] EN_VSS_P[7] EN_VSS_P[6] EN_VSS_P[5]
+ EN_VSS_P[4] EN_VSS_P[3] EN_VSS_P[2] EN_VSS_P[1] EN_VSS_P[0] EN_REF_Z_P[10] EN_REF_Z_P[9] EN_REF_Z_P[8] EN_REF_Z_P[7] EN_REF_Z_P[6]
+ EN_REF_Z_P[5] EN_REF_Z_P[4] EN_REF_Z_P[3] EN_REF_Z_P[2] EN_REF_Z_P[1] EN_REF_Z_P[0] EN_REF_Z_P_BBM[10] EN_REF_Z_P_BBM[9] EN_REF_Z_P_BBM[8]
+ EN_REF_Z_P_BBM[7] EN_REF_Z_P_BBM[6] EN_REF_Z_P_BBM[5] EN_REF_Z_P_BBM[4] EN_REF_Z_P_BBM[3] EN_REF_Z_P_BBM[2] EN_REF_Z_P_BBM[1] EN_REF_Z_P_BBM[0]
+ break_before_make
.ends


* expanding   symbol:  subcells/switches/switches.sym # of pins=25
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/switches/switches.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/switches/switches.sch
.subckt switches VCM VREF_GND VREF VIN EN_VIN EN_VREF_Z[10] EN_VREF_Z[9] EN_VREF_Z[8] EN_VREF_Z[7] EN_VREF_Z[6] EN_VREF_Z[5]
+ EN_VREF_Z[4] EN_VREF_Z[3] EN_VREF_Z[2] EN_VREF_Z[1] EN_VREF_Z[0] EN_VSS[10] EN_VSS[9] EN_VSS[8] EN_VSS[7] EN_VSS[6] EN_VSS[5] EN_VSS[4]
+ EN_VSS[3] EN_VSS[2] EN_VSS[1] EN_VSS[0] EN_VCM[10] EN_VCM[9] EN_VCM[8] EN_VCM[7] EN_VCM[6] EN_VCM[5] EN_VCM[4] EN_VCM[3] EN_VCM[2]
+ EN_VCM[1] EN_VCM[0] EN_VCM_SW EN_VCM_DUMMY Cbtm_8 Cbtm_7 Cbtm_0 Cbtm_6 Cbtm_5 Cbtm_0_dummy Cbtm_4 Cbtm_3 VDAC Cbtm_10 Cbtm_9 Cbtm_2 Cbtm_1
+ VDD VSS
*.ipin VCM
*.ipin VREF_GND
*.ipin VREF
*.ipin VIN
*.ipin VDD
*.opin Cbtm_0_dummy
*.opin Cbtm_0
*.opin Cbtm_1
*.opin Cbtm_2
*.opin Cbtm_3
*.opin Cbtm_4
*.opin Cbtm_5
*.opin Cbtm_6
*.opin Cbtm_7
*.opin Cbtm_8
*.opin Cbtm_9
*.opin Cbtm_10
*.opin VDAC
*.ipin EN_VIN
*.ipin
*+ EN_VREF_Z[10],EN_VREF_Z[9],EN_VREF_Z[8],EN_VREF_Z[7],EN_VREF_Z[6],EN_VREF_Z[5],EN_VREF_Z[4],EN_VREF_Z[3],EN_VREF_Z[2],EN_VREF_Z[1],EN_VREF_Z[0]
*.ipin EN_VSS[10],EN_VSS[9],EN_VSS[8],EN_VSS[7],EN_VSS[6],EN_VSS[5],EN_VSS[4],EN_VSS[3],EN_VSS[2],EN_VSS[1],EN_VSS[0]
*.ipin EN_VCM[10],EN_VCM[9],EN_VCM[8],EN_VCM[7],EN_VCM[6],EN_VCM[5],EN_VCM[4],EN_VCM[3],EN_VCM[2],EN_VCM[1],EN_VCM[0]
*.ipin EN_VCM_DUMMY
*.ipin EN_VCM_SW
*.ipin VSS
x1 VCM EN_VCM_SW VDAC VDD VSS switch_VCM
x2 VCM VREF_GND VIN VREF EN_VCM[10] EN_VREF_Z[10] Cbtm_10 VDD EN_VSS[10] EN_VIN VSS switch_C10
x3 VCM VREF_GND VIN VREF EN_VCM[9] EN_VREF_Z[9] Cbtm_9 VDD EN_VSS[9] EN_VIN VSS switch_C9
x4 VCM VREF_GND VIN VREF EN_VCM[8] EN_VREF_Z[8] Cbtm_8 VDD EN_VSS[8] EN_VIN VSS switch_C8
x5 VCM VREF_GND VIN VREF EN_VCM[7] EN_VREF_Z[7] Cbtm_7 VDD EN_VSS[7] EN_VIN VSS switch_C7
x6 VCM VREF_GND VIN VREF EN_VCM[6] EN_VREF_Z[6] Cbtm_6 VDD EN_VSS[6] EN_VIN VSS switch_C6
x7 VCM VREF_GND VIN VREF EN_VCM[5] EN_VREF_Z[5] Cbtm_5 VDD EN_VSS[5] EN_VIN VSS switch_C5
x8 VCM VREF_GND VIN VREF EN_VCM[4] EN_VREF_Z[4] Cbtm_4 VDD EN_VSS[4] EN_VIN VSS switch_C5
x9 VCM VREF_GND VIN VREF EN_VCM[3] EN_VREF_Z[3] Cbtm_3 VDD EN_VSS[3] EN_VIN VSS switch_C5
x10 VCM VREF_GND VIN VREF EN_VCM[2] EN_VREF_Z[2] Cbtm_2 VDD EN_VSS[2] EN_VIN VSS switch_C5
x11 VCM VREF_GND VIN VREF EN_VCM[1] EN_VREF_Z[1] Cbtm_1 VDD EN_VSS[1] EN_VIN VSS switch_C5
x12 VCM VREF_GND VIN VREF EN_VCM[0] EN_VREF_Z[0] Cbtm_0 VDD EN_VSS[0] EN_VIN VSS switch_C5
x13 VCM VIN EN_VCM_DUMMY Cbtm_0_dummy EN_VIN VSS switch_C0_dummy
.ends


* expanding   symbol:  subcells/preamplifier/preamplifier.sym # of pins=9
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/preamplifier/preamplifier.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/preamplifier/preamplifier.sch
.subckt preamplifier IN_N IN_P VDD EN OUT_P OUT_N VSS CAL_P CAL_N
*.ipin VDD
*.ipin VSS
*.ipin IN_P
*.ipin IN_N
*.opin OUT_P
*.opin OUT_N
*.ipin EN
*.ipin CAL_P
*.ipin CAL_N
XM4 net1 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM5 net5 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 OUT_N net5 net9 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM14 OUT_P net5 net10 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM8 net9 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net10 net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net8 EN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 net3 EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net5 EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 EN VSS VSS VDD VDD EN_Z sky130_fd_sc_hd__inv_1
XM20 net6 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM19 VDD OUT_N net6 VSS sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM21 VDD OUT_P net6 VSS sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net12 IN_P net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=24 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM2 net7 IN_N net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=24 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM15 net9 CAL_P net11 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 net10 CAL_N net11 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR6 net2 net3 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM23 net11 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XR3 net8 net2 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[3] rn[0] OUT_N VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[2] rn[1] rn[0] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[1] rn[2] rn[1] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR4[0] common rn[2] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR5 net4 net5 VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM9 OUT_P VSS net7 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT_N VSS net12 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1[3] rp[0] OUT_P VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[2] rp[1] rp[0] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[1] rp[2] rp[1] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR1[0] common rp[2] VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XM11 VDD net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM13 VSS net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM24 net10 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net9 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/latched_comparator/latched_comparator.sym # of pins=7
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/latched_comparator/latched_comparator.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/latched_comparator/latched_comparator.sch
.subckt latched_comparator VDD VIN_P VIN_N EN OUT_P OUT_N VSS
*.ipin VIN_P
*.ipin VIN_N
*.ipin VDD
*.ipin VSS
*.ipin EN
*.opin OUT_N
*.opin OUT_P
x1 EN VSS VSS VDD VDD ENi sky130_fd_sc_hd__buf_4
XM10 net2 ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT_Ni ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 OUT_Ni OUT_Pi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 OUT_Pi OUT_Ni VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT_Ni OUT_Pi net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT_Pi OUT_Ni net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net1 ENi VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM16 net3 VIN_N net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 VIN_P net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 OUT_Pi ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net3 ENi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x4 OUT_Pi VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x5 OUT_Ni VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x6 net5 VSS VSS VDD VDD OUT_N sky130_fd_sc_hd__inv_4
x7 net4 VSS VSS VDD VDD OUT_P sky130_fd_sc_hd__inv_4
XM2 net1 net1 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  subcells/offset_calibration/offset_calibration.sym # of pins=8
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/offset_calibration/offset_calibration.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/offset_calibration/offset_calibration.sch
.subckt offset_calibration VDD CAL_RESULT EN_COMP CAL_P CAL_N EN VSS CAL_CYCLE
*.ipin EN_COMP
*.opin CAL_N
*.opin CAL_P
*.ipin VDD
*.ipin VSS
*.ipin EN
*.ipin CAL_RESULT
*.ipin CAL_CYCLE
XM26 net2 EN_COMPi net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 net1 CAL_RESULTi VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 net2 EN_COMP_Z net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM29 net3 CAL_RESULTi VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 net2 LOAD_CALi CAL_P VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM31 net2 LOAD_CAL_Z CAL_P VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x22 EN net8 net7 VSS VSS VDD VDD LOAD_CAL_Z sky130_fd_sc_hd__nand3_1
x3 LOAD_CAL_Z VSS VSS VDD VDD LOAD_CALi sky130_fd_sc_hd__inv_1
XM32 net5 LOAD_CAL_Z CAL_N VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM33 net5 LOAD_CALi CAL_N VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 net5 EN_COMP_Z net6 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM35 net6 CAL_RESULT_Z VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM36 net5 EN_COMPi net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM37 net4 CAL_RESULT_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM25 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM1 CAL_N EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 CAL_P EN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 CAL_RESULT CAL_CYCLE VSS VSS VDD VDD CAL_RESULT_Z sky130_fd_sc_hd__nand2_1
x4 CAL_RESULT_Z VSS VSS VDD VDD CAL_RESULTi sky130_fd_sc_hd__inv_1
x2 EN_COMP CAL_CYCLE VSS VSS VDD VDD EN_COMP_Z sky130_fd_sc_hd__nand2_1
x5 EN_COMP_Z VSS VSS VDD VDD EN_COMPi sky130_fd_sc_hd__inv_1
x6 EN_COMPi VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_1
x7 CAL_CYCLE VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  subcells/bootstrap/bootstrap.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/bootstrap/bootstrap.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/bootstrap/bootstrap.sch
.subckt bootstrap VDD VSS VIN SW_ON EN VGATE
*.ipin VDD
*.ipin VSS
*.ipin VIN
*.opin VGATE
*.ipin EN
*.opin SW_ON
XM1 VDD VGATE Vtop Vtop sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VGATE EN_Z Vtop Vtop sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 VGATE VDD Vd VSS sky130_fd_pr__nfet_05v0_nvt L=0.9 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vd EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vbottom EN_Z VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vtop Vbottom Vtop Vtop sky130_fd_pr__pfet_01v8 L=15 W=15 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 EN VSS VSS VDD VDD EN_Z sky130_fd_sc_hd__inv_4
XM8 VIN VGATE Vbottom VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 VGATE VDD VGATE_1V8 VSS sky130_fd_pr__nfet_05v0_nvt L=0.9 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 VGATE_1V8 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_2
x3 net1 VSS VSS VDD VDD SW_ON sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  subcells/break_before_make/break_before_make.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/break_before_make/break_before_make.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/break_before_make/break_before_make.sch
.subckt break_before_make EN_VSS_I[10] EN_VSS_I[9] EN_VSS_I[8] EN_VSS_I[7] EN_VSS_I[6] EN_VSS_I[5] EN_VSS_I[4] EN_VSS_I[3]
+ EN_VSS_I[2] EN_VSS_I[1] EN_VSS_I[0] VDD VSS EN_VSS_O[10] EN_VSS_O[9] EN_VSS_O[8] EN_VSS_O[7] EN_VSS_O[6] EN_VSS_O[5] EN_VSS_O[4] EN_VSS_O[3]
+ EN_VSS_O[2] EN_VSS_O[1] EN_VSS_O[0] EN_VREF_Z_O[10] EN_VREF_Z_O[9] EN_VREF_Z_O[8] EN_VREF_Z_O[7] EN_VREF_Z_O[6] EN_VREF_Z_O[5] EN_VREF_Z_O[4]
+ EN_VREF_Z_O[3] EN_VREF_Z_O[2] EN_VREF_Z_O[1] EN_VREF_Z_O[0] EN_VREF_Z_I[10] EN_VREF_Z_I[9] EN_VREF_Z_I[8] EN_VREF_Z_I[7] EN_VREF_Z_I[6]
+ EN_VREF_Z_I[5] EN_VREF_Z_I[4] EN_VREF_Z_I[3] EN_VREF_Z_I[2] EN_VREF_Z_I[1] EN_VREF_Z_I[0]
*.ipin
*+ EN_VSS_I[10],EN_VSS_I[9],EN_VSS_I[8],EN_VSS_I[7],EN_VSS_I[6],EN_VSS_I[5],EN_VSS_I[4],EN_VSS_I[3],EN_VSS_I[2],EN_VSS_I[1],EN_VSS_I[0]
*.ipin
*+ EN_VREF_Z_I[10],EN_VREF_Z_I[9],EN_VREF_Z_I[8],EN_VREF_Z_I[7],EN_VREF_Z_I[6],EN_VREF_Z_I[5],EN_VREF_Z_I[4],EN_VREF_Z_I[3],EN_VREF_Z_I[2],EN_VREF_Z_I[1],EN_VREF_Z_I[0]
*.ipin VDD
*.ipin VSS
*.opin
*+ EN_VSS_O[10],EN_VSS_O[9],EN_VSS_O[8],EN_VSS_O[7],EN_VSS_O[6],EN_VSS_O[5],EN_VSS_O[4],EN_VSS_O[3],EN_VSS_O[2],EN_VSS_O[1],EN_VSS_O[0]
*.opin
*+ EN_VREF_Z_O[10],EN_VREF_Z_O[9],EN_VREF_Z_O[8],EN_VREF_Z_O[7],EN_VREF_Z_O[6],EN_VREF_Z_O[5],EN_VREF_Z_O[4],EN_VREF_Z_O[3],EN_VREF_Z_O[2],EN_VREF_Z_O[1],EN_VREF_Z_O[0]
x1[10] EN_VSS_I[10] EN_VREF_Z_O[10] VSS VSS VDD VDD EN_VSS_O[10] sky130_fd_sc_hd__and2_4
x1[9] EN_VSS_I[9] EN_VREF_Z_O[9] VSS VSS VDD VDD EN_VSS_O[9] sky130_fd_sc_hd__and2_4
x1[8] EN_VSS_I[8] EN_VREF_Z_O[8] VSS VSS VDD VDD EN_VSS_O[8] sky130_fd_sc_hd__and2_4
x1[7] EN_VSS_I[7] EN_VREF_Z_O[7] VSS VSS VDD VDD EN_VSS_O[7] sky130_fd_sc_hd__and2_4
x1[6] EN_VSS_I[6] EN_VREF_Z_O[6] VSS VSS VDD VDD EN_VSS_O[6] sky130_fd_sc_hd__and2_4
x1[5] EN_VSS_I[5] EN_VREF_Z_O[5] VSS VSS VDD VDD EN_VSS_O[5] sky130_fd_sc_hd__and2_4
x1[4] EN_VSS_I[4] EN_VREF_Z_O[4] VSS VSS VDD VDD EN_VSS_O[4] sky130_fd_sc_hd__and2_4
x1[3] EN_VSS_I[3] EN_VREF_Z_O[3] VSS VSS VDD VDD EN_VSS_O[3] sky130_fd_sc_hd__and2_4
x1[2] EN_VSS_I[2] EN_VREF_Z_O[2] VSS VSS VDD VDD EN_VSS_O[2] sky130_fd_sc_hd__and2_4
x1[1] EN_VSS_I[1] EN_VREF_Z_O[1] VSS VSS VDD VDD EN_VSS_O[1] sky130_fd_sc_hd__and2_4
x1[0] EN_VSS_I[0] EN_VREF_Z_O[0] VSS VSS VDD VDD EN_VSS_O[0] sky130_fd_sc_hd__and2_4
x2[10] EN_VSS_O[10] EN_VREF_Z_I[10] VSS VSS VDD VDD EN_VREF_Z_O[10] sky130_fd_sc_hd__or2_4
x2[9] EN_VSS_O[9] EN_VREF_Z_I[9] VSS VSS VDD VDD EN_VREF_Z_O[9] sky130_fd_sc_hd__or2_4
x2[8] EN_VSS_O[8] EN_VREF_Z_I[8] VSS VSS VDD VDD EN_VREF_Z_O[8] sky130_fd_sc_hd__or2_4
x2[7] EN_VSS_O[7] EN_VREF_Z_I[7] VSS VSS VDD VDD EN_VREF_Z_O[7] sky130_fd_sc_hd__or2_4
x2[6] EN_VSS_O[6] EN_VREF_Z_I[6] VSS VSS VDD VDD EN_VREF_Z_O[6] sky130_fd_sc_hd__or2_4
x2[5] EN_VSS_O[5] EN_VREF_Z_I[5] VSS VSS VDD VDD EN_VREF_Z_O[5] sky130_fd_sc_hd__or2_4
x2[4] EN_VSS_O[4] EN_VREF_Z_I[4] VSS VSS VDD VDD EN_VREF_Z_O[4] sky130_fd_sc_hd__or2_4
x2[3] EN_VSS_O[3] EN_VREF_Z_I[3] VSS VSS VDD VDD EN_VREF_Z_O[3] sky130_fd_sc_hd__or2_4
x2[2] EN_VSS_O[2] EN_VREF_Z_I[2] VSS VSS VDD VDD EN_VREF_Z_O[2] sky130_fd_sc_hd__or2_4
x2[1] EN_VSS_O[1] EN_VREF_Z_I[1] VSS VSS VDD VDD EN_VREF_Z_O[1] sky130_fd_sc_hd__or2_4
x2[0] EN_VSS_O[0] EN_VREF_Z_I[0] VSS VSS VDD VDD EN_VREF_Z_O[0] sky130_fd_sc_hd__or2_4
x1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_12
x2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
.ends


* expanding   symbol:  subcells/individual_switches/switch_VCM.sym # of pins=5
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_VCM.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_VCM.sch
.subckt switch_VCM VCM EN_VCM Cbtm VDD VSS
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VSS
*.ipin VDD
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=64 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C10.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C10.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C10.sch
.subckt switch_C10 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=64 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=128 nf=16 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=64 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C9.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C9.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C9.sch
.subckt switch_C9 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=32 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=64 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=32 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C8.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C8.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C8.sch
.subckt switch_C8 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=32 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=16 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C7.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C7.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C7.sch
.subckt switch_C7 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C6.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C6.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C6.sch
.subckt switch_C6 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C5.sym # of pins=11
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C5.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C5.sch
.subckt switch_C5 VCM VREF_GND VIN VREF EN_VCM EN_VREF_Z Cbtm VDD EN_VSS EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VREF_GND
*.ipin VREF
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VDD
*.ipin EN_VSS
*.ipin EN_VREF_Z
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VREF_GND EN_VSS Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Cbtm EN_VREF_Z VREF VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  subcells/individual_switches/switch_C0_dummy.sym # of pins=6
** sym_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C0_dummy.sym
** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/schematic/subcells/individual_switches/switch_C0_dummy.sch
.subckt switch_C0_dummy VCM VIN EN_VCM Cbtm EN_VIN VSS
*.ipin VIN
*.ipin EN_VIN
*.ipin VCM
*.ipin EN_VCM
*.opin Cbtm
*.ipin VSS
XM1 VIN EN_VIN Cbtm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VCM EN_VCM Cbtm VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
