magic
tech sky130A
magscale 1 2
timestamp 1712002891
<< nwell >>
rect 3700 2516 10208 2870
rect 3700 1950 10804 2516
rect 3700 1428 10208 1950
rect 3700 1107 10896 1428
rect 3700 862 10804 1107
rect 3700 364 10208 862
rect 3700 -574 10820 364
rect 3700 -1900 10208 -574
<< pwell >>
rect 10427 2760 10461 2794
rect 10427 2756 10448 2760
rect 10704 2756 10738 2794
rect 10262 2574 10448 2756
rect 10491 2574 10761 2756
rect 10262 1710 10448 1892
rect 10491 1710 10761 1892
rect 10427 1706 10448 1710
rect 10427 1672 10461 1706
rect 10704 1672 10738 1710
rect 10427 1668 10448 1672
rect 10794 1668 10828 1706
rect 10262 1486 10448 1668
rect 10491 1486 10857 1668
rect 10256 622 10442 804
rect 10532 622 10718 804
rect 10256 618 10277 622
rect 10532 618 10553 622
rect 10243 584 10277 618
rect 10519 584 10553 618
rect 10210 -1668 10832 -766
<< nmos >>
rect 10410 -1060 10440 -976
rect 10506 -1060 10536 -976
rect 10602 -1060 10632 -976
rect 10410 -1458 10440 -1374
rect 10506 -1458 10536 -1374
rect 10602 -1458 10632 -1374
<< scnmos >>
rect 10340 2600 10370 2730
rect 10569 2600 10599 2730
rect 10653 2600 10683 2730
rect 10340 1736 10370 1866
rect 10569 1736 10599 1866
rect 10653 1736 10683 1866
rect 10340 1512 10370 1642
rect 10569 1512 10599 1642
rect 10665 1512 10695 1642
rect 10749 1512 10779 1642
rect 10334 648 10364 778
rect 10610 648 10640 778
<< pmos >>
rect 10302 61 10332 145
rect 10398 61 10428 145
rect 10494 61 10524 145
rect 10590 61 10620 145
rect 10302 -355 10332 -271
rect 10398 -355 10428 -271
rect 10494 -355 10524 -271
rect 10590 -355 10620 -271
<< scpmoshvt >>
rect 10340 2280 10370 2480
rect 10569 2280 10599 2480
rect 10653 2280 10683 2480
rect 10340 1986 10370 2186
rect 10569 1986 10599 2186
rect 10653 1986 10683 2186
rect 10340 1192 10370 1392
rect 10569 1192 10599 1392
rect 10665 1192 10695 1392
rect 10749 1192 10779 1392
rect 10334 898 10364 1098
rect 10610 898 10640 1098
<< pmoslvt >>
rect 3896 651 5896 2651
rect 5954 651 7954 2651
rect 8012 651 10012 2651
rect 3896 -1681 5896 319
rect 5954 -1681 7954 319
rect 8012 -1681 10012 319
<< ndiff >>
rect 10288 2714 10340 2730
rect 10288 2680 10296 2714
rect 10330 2680 10340 2714
rect 10288 2646 10340 2680
rect 10288 2612 10296 2646
rect 10330 2612 10340 2646
rect 10288 2600 10340 2612
rect 10370 2714 10422 2730
rect 10370 2680 10380 2714
rect 10414 2680 10422 2714
rect 10370 2646 10422 2680
rect 10370 2612 10380 2646
rect 10414 2612 10422 2646
rect 10370 2600 10422 2612
rect 10517 2718 10569 2730
rect 10517 2684 10525 2718
rect 10559 2684 10569 2718
rect 10517 2650 10569 2684
rect 10517 2616 10525 2650
rect 10559 2616 10569 2650
rect 10517 2600 10569 2616
rect 10599 2600 10653 2730
rect 10683 2718 10735 2730
rect 10683 2684 10693 2718
rect 10727 2684 10735 2718
rect 10683 2650 10735 2684
rect 10683 2616 10693 2650
rect 10727 2616 10735 2650
rect 10683 2600 10735 2616
rect 10288 1854 10340 1866
rect 10288 1820 10296 1854
rect 10330 1820 10340 1854
rect 10288 1786 10340 1820
rect 10288 1752 10296 1786
rect 10330 1752 10340 1786
rect 10288 1736 10340 1752
rect 10370 1854 10422 1866
rect 10370 1820 10380 1854
rect 10414 1820 10422 1854
rect 10370 1786 10422 1820
rect 10370 1752 10380 1786
rect 10414 1752 10422 1786
rect 10370 1736 10422 1752
rect 10517 1850 10569 1866
rect 10517 1816 10525 1850
rect 10559 1816 10569 1850
rect 10517 1782 10569 1816
rect 10517 1748 10525 1782
rect 10559 1748 10569 1782
rect 10517 1736 10569 1748
rect 10599 1736 10653 1866
rect 10683 1850 10735 1866
rect 10683 1816 10693 1850
rect 10727 1816 10735 1850
rect 10683 1782 10735 1816
rect 10683 1748 10693 1782
rect 10727 1748 10735 1782
rect 10683 1736 10735 1748
rect 10288 1626 10340 1642
rect 10288 1592 10296 1626
rect 10330 1592 10340 1626
rect 10288 1558 10340 1592
rect 10288 1524 10296 1558
rect 10330 1524 10340 1558
rect 10288 1512 10340 1524
rect 10370 1626 10422 1642
rect 10370 1592 10380 1626
rect 10414 1592 10422 1626
rect 10370 1558 10422 1592
rect 10370 1524 10380 1558
rect 10414 1524 10422 1558
rect 10370 1512 10422 1524
rect 10517 1630 10569 1642
rect 10517 1596 10525 1630
rect 10559 1596 10569 1630
rect 10517 1562 10569 1596
rect 10517 1528 10525 1562
rect 10559 1528 10569 1562
rect 10517 1512 10569 1528
rect 10599 1512 10665 1642
rect 10695 1512 10749 1642
rect 10779 1624 10831 1642
rect 10779 1590 10789 1624
rect 10823 1590 10831 1624
rect 10779 1512 10831 1590
rect 10282 766 10334 778
rect 10282 732 10290 766
rect 10324 732 10334 766
rect 10282 698 10334 732
rect 10282 664 10290 698
rect 10324 664 10334 698
rect 10282 648 10334 664
rect 10364 766 10416 778
rect 10364 732 10374 766
rect 10408 732 10416 766
rect 10364 698 10416 732
rect 10364 664 10374 698
rect 10408 664 10416 698
rect 10364 648 10416 664
rect 10558 766 10610 778
rect 10558 732 10566 766
rect 10600 732 10610 766
rect 10558 698 10610 732
rect 10558 664 10566 698
rect 10600 664 10610 698
rect 10558 648 10610 664
rect 10640 766 10692 778
rect 10640 732 10650 766
rect 10684 732 10692 766
rect 10640 698 10692 732
rect 10640 664 10650 698
rect 10684 664 10692 698
rect 10640 648 10692 664
rect 10348 -988 10410 -976
rect 10348 -1048 10360 -988
rect 10394 -1048 10410 -988
rect 10348 -1060 10410 -1048
rect 10440 -988 10506 -976
rect 10440 -1048 10456 -988
rect 10490 -1048 10506 -988
rect 10440 -1060 10506 -1048
rect 10536 -988 10602 -976
rect 10536 -1048 10552 -988
rect 10586 -1048 10602 -988
rect 10536 -1060 10602 -1048
rect 10632 -988 10694 -976
rect 10632 -1048 10648 -988
rect 10682 -1048 10694 -988
rect 10632 -1060 10694 -1048
rect 10348 -1386 10410 -1374
rect 10348 -1446 10360 -1386
rect 10394 -1446 10410 -1386
rect 10348 -1458 10410 -1446
rect 10440 -1386 10506 -1374
rect 10440 -1446 10456 -1386
rect 10490 -1446 10506 -1386
rect 10440 -1458 10506 -1446
rect 10536 -1386 10602 -1374
rect 10536 -1446 10552 -1386
rect 10586 -1446 10602 -1386
rect 10536 -1458 10602 -1446
rect 10632 -1386 10694 -1374
rect 10632 -1446 10648 -1386
rect 10682 -1446 10694 -1386
rect 10632 -1458 10694 -1446
<< pdiff >>
rect 3838 2639 3896 2651
rect 3838 663 3850 2639
rect 3884 663 3896 2639
rect 3838 651 3896 663
rect 5896 2639 5954 2651
rect 5896 663 5908 2639
rect 5942 663 5954 2639
rect 5896 651 5954 663
rect 7954 2639 8012 2651
rect 7954 663 7966 2639
rect 8000 663 8012 2639
rect 7954 651 8012 663
rect 10012 2639 10070 2651
rect 10012 663 10024 2639
rect 10058 663 10070 2639
rect 10012 651 10070 663
rect 10288 2462 10340 2480
rect 10288 2428 10296 2462
rect 10330 2428 10340 2462
rect 10288 2394 10340 2428
rect 10288 2360 10296 2394
rect 10330 2360 10340 2394
rect 10288 2326 10340 2360
rect 10288 2292 10296 2326
rect 10330 2292 10340 2326
rect 10288 2280 10340 2292
rect 10370 2462 10422 2480
rect 10370 2428 10380 2462
rect 10414 2428 10422 2462
rect 10370 2394 10422 2428
rect 10370 2360 10380 2394
rect 10414 2360 10422 2394
rect 10370 2326 10422 2360
rect 10370 2292 10380 2326
rect 10414 2292 10422 2326
rect 10370 2280 10422 2292
rect 10517 2462 10569 2480
rect 10517 2428 10525 2462
rect 10559 2428 10569 2462
rect 10517 2394 10569 2428
rect 10517 2360 10525 2394
rect 10559 2360 10569 2394
rect 10517 2326 10569 2360
rect 10517 2292 10525 2326
rect 10559 2292 10569 2326
rect 10517 2280 10569 2292
rect 10599 2462 10653 2480
rect 10599 2428 10609 2462
rect 10643 2428 10653 2462
rect 10599 2394 10653 2428
rect 10599 2360 10609 2394
rect 10643 2360 10653 2394
rect 10599 2326 10653 2360
rect 10599 2292 10609 2326
rect 10643 2292 10653 2326
rect 10599 2280 10653 2292
rect 10683 2462 10735 2480
rect 10683 2428 10693 2462
rect 10727 2428 10735 2462
rect 10683 2394 10735 2428
rect 10683 2360 10693 2394
rect 10727 2360 10735 2394
rect 10683 2326 10735 2360
rect 10683 2292 10693 2326
rect 10727 2292 10735 2326
rect 10683 2280 10735 2292
rect 10288 2174 10340 2186
rect 10288 2140 10296 2174
rect 10330 2140 10340 2174
rect 10288 2106 10340 2140
rect 10288 2072 10296 2106
rect 10330 2072 10340 2106
rect 10288 2038 10340 2072
rect 10288 2004 10296 2038
rect 10330 2004 10340 2038
rect 10288 1986 10340 2004
rect 10370 2174 10422 2186
rect 10370 2140 10380 2174
rect 10414 2140 10422 2174
rect 10370 2106 10422 2140
rect 10370 2072 10380 2106
rect 10414 2072 10422 2106
rect 10370 2038 10422 2072
rect 10370 2004 10380 2038
rect 10414 2004 10422 2038
rect 10370 1986 10422 2004
rect 10517 2174 10569 2186
rect 10517 2140 10525 2174
rect 10559 2140 10569 2174
rect 10517 2106 10569 2140
rect 10517 2072 10525 2106
rect 10559 2072 10569 2106
rect 10517 2038 10569 2072
rect 10517 2004 10525 2038
rect 10559 2004 10569 2038
rect 10517 1986 10569 2004
rect 10599 2174 10653 2186
rect 10599 2140 10609 2174
rect 10643 2140 10653 2174
rect 10599 2106 10653 2140
rect 10599 2072 10609 2106
rect 10643 2072 10653 2106
rect 10599 2038 10653 2072
rect 10599 2004 10609 2038
rect 10643 2004 10653 2038
rect 10599 1986 10653 2004
rect 10683 2174 10735 2186
rect 10683 2140 10693 2174
rect 10727 2140 10735 2174
rect 10683 2106 10735 2140
rect 10683 2072 10693 2106
rect 10727 2072 10735 2106
rect 10683 2038 10735 2072
rect 10683 2004 10693 2038
rect 10727 2004 10735 2038
rect 10683 1986 10735 2004
rect 10288 1374 10340 1392
rect 10288 1340 10296 1374
rect 10330 1340 10340 1374
rect 10288 1306 10340 1340
rect 10288 1272 10296 1306
rect 10330 1272 10340 1306
rect 10288 1238 10340 1272
rect 10288 1204 10296 1238
rect 10330 1204 10340 1238
rect 10288 1192 10340 1204
rect 10370 1374 10422 1392
rect 10370 1340 10380 1374
rect 10414 1340 10422 1374
rect 10370 1306 10422 1340
rect 10370 1272 10380 1306
rect 10414 1272 10422 1306
rect 10370 1238 10422 1272
rect 10370 1204 10380 1238
rect 10414 1204 10422 1238
rect 10370 1192 10422 1204
rect 10517 1374 10569 1392
rect 10517 1340 10525 1374
rect 10559 1340 10569 1374
rect 10517 1306 10569 1340
rect 10517 1272 10525 1306
rect 10559 1272 10569 1306
rect 10517 1238 10569 1272
rect 10517 1204 10525 1238
rect 10559 1204 10569 1238
rect 10517 1192 10569 1204
rect 10599 1306 10665 1392
rect 10599 1272 10621 1306
rect 10655 1272 10665 1306
rect 10599 1238 10665 1272
rect 10599 1204 10621 1238
rect 10655 1204 10665 1238
rect 10599 1192 10665 1204
rect 10695 1374 10749 1392
rect 10695 1340 10705 1374
rect 10739 1340 10749 1374
rect 10695 1306 10749 1340
rect 10695 1272 10705 1306
rect 10739 1272 10749 1306
rect 10695 1238 10749 1272
rect 10695 1204 10705 1238
rect 10739 1204 10749 1238
rect 10695 1192 10749 1204
rect 10779 1374 10831 1392
rect 10779 1340 10789 1374
rect 10823 1340 10831 1374
rect 10779 1306 10831 1340
rect 10779 1272 10789 1306
rect 10823 1272 10831 1306
rect 10779 1238 10831 1272
rect 10779 1204 10789 1238
rect 10823 1204 10831 1238
rect 10779 1192 10831 1204
rect 10282 1086 10334 1098
rect 10282 1052 10290 1086
rect 10324 1052 10334 1086
rect 10282 1018 10334 1052
rect 10282 984 10290 1018
rect 10324 984 10334 1018
rect 10282 950 10334 984
rect 10282 916 10290 950
rect 10324 916 10334 950
rect 10282 898 10334 916
rect 10364 1086 10416 1098
rect 10364 1052 10374 1086
rect 10408 1052 10416 1086
rect 10364 1018 10416 1052
rect 10364 984 10374 1018
rect 10408 984 10416 1018
rect 10364 950 10416 984
rect 10364 916 10374 950
rect 10408 916 10416 950
rect 10364 898 10416 916
rect 10558 1086 10610 1098
rect 10558 1052 10566 1086
rect 10600 1052 10610 1086
rect 10558 1018 10610 1052
rect 10558 984 10566 1018
rect 10600 984 10610 1018
rect 10558 950 10610 984
rect 10558 916 10566 950
rect 10600 916 10610 950
rect 10558 898 10610 916
rect 10640 1086 10692 1098
rect 10640 1052 10650 1086
rect 10684 1052 10692 1086
rect 10640 1018 10692 1052
rect 10640 984 10650 1018
rect 10684 984 10692 1018
rect 10640 950 10692 984
rect 10640 916 10650 950
rect 10684 916 10692 950
rect 10640 898 10692 916
rect 3838 307 3896 319
rect 3838 -1669 3850 307
rect 3884 -1669 3896 307
rect 3838 -1681 3896 -1669
rect 5896 307 5954 319
rect 5896 -1669 5908 307
rect 5942 -1669 5954 307
rect 5896 -1681 5954 -1669
rect 7954 307 8012 319
rect 7954 -1669 7966 307
rect 8000 -1669 8012 307
rect 7954 -1681 8012 -1669
rect 10012 307 10070 319
rect 10012 -1669 10024 307
rect 10058 -1669 10070 307
rect 10012 -1681 10070 -1669
rect 10240 133 10302 145
rect 10240 73 10252 133
rect 10286 73 10302 133
rect 10240 61 10302 73
rect 10332 133 10398 145
rect 10332 73 10348 133
rect 10382 73 10398 133
rect 10332 61 10398 73
rect 10428 133 10494 145
rect 10428 73 10444 133
rect 10478 73 10494 133
rect 10428 61 10494 73
rect 10524 133 10590 145
rect 10524 73 10540 133
rect 10574 73 10590 133
rect 10524 61 10590 73
rect 10620 133 10682 145
rect 10620 73 10636 133
rect 10670 73 10682 133
rect 10620 61 10682 73
rect 10240 -283 10302 -271
rect 10240 -343 10252 -283
rect 10286 -343 10302 -283
rect 10240 -355 10302 -343
rect 10332 -283 10398 -271
rect 10332 -343 10348 -283
rect 10382 -343 10398 -283
rect 10332 -355 10398 -343
rect 10428 -283 10494 -271
rect 10428 -343 10444 -283
rect 10478 -343 10494 -283
rect 10428 -355 10494 -343
rect 10524 -283 10590 -271
rect 10524 -343 10540 -283
rect 10574 -343 10590 -283
rect 10524 -355 10590 -343
rect 10620 -283 10682 -271
rect 10620 -343 10636 -283
rect 10670 -343 10682 -283
rect 10620 -355 10682 -343
<< ndiffc >>
rect 10296 2680 10330 2714
rect 10296 2612 10330 2646
rect 10380 2680 10414 2714
rect 10380 2612 10414 2646
rect 10525 2684 10559 2718
rect 10525 2616 10559 2650
rect 10693 2684 10727 2718
rect 10693 2616 10727 2650
rect 10296 1820 10330 1854
rect 10296 1752 10330 1786
rect 10380 1820 10414 1854
rect 10380 1752 10414 1786
rect 10525 1816 10559 1850
rect 10525 1748 10559 1782
rect 10693 1816 10727 1850
rect 10693 1748 10727 1782
rect 10296 1592 10330 1626
rect 10296 1524 10330 1558
rect 10380 1592 10414 1626
rect 10380 1524 10414 1558
rect 10525 1596 10559 1630
rect 10525 1528 10559 1562
rect 10789 1590 10823 1624
rect 10290 732 10324 766
rect 10290 664 10324 698
rect 10374 732 10408 766
rect 10374 664 10408 698
rect 10566 732 10600 766
rect 10566 664 10600 698
rect 10650 732 10684 766
rect 10650 664 10684 698
rect 10360 -1048 10394 -988
rect 10456 -1048 10490 -988
rect 10552 -1048 10586 -988
rect 10648 -1048 10682 -988
rect 10360 -1446 10394 -1386
rect 10456 -1446 10490 -1386
rect 10552 -1446 10586 -1386
rect 10648 -1446 10682 -1386
<< pdiffc >>
rect 3850 663 3884 2639
rect 5908 663 5942 2639
rect 7966 663 8000 2639
rect 10024 663 10058 2639
rect 10296 2428 10330 2462
rect 10296 2360 10330 2394
rect 10296 2292 10330 2326
rect 10380 2428 10414 2462
rect 10380 2360 10414 2394
rect 10380 2292 10414 2326
rect 10525 2428 10559 2462
rect 10525 2360 10559 2394
rect 10525 2292 10559 2326
rect 10609 2428 10643 2462
rect 10609 2360 10643 2394
rect 10609 2292 10643 2326
rect 10693 2428 10727 2462
rect 10693 2360 10727 2394
rect 10693 2292 10727 2326
rect 10296 2140 10330 2174
rect 10296 2072 10330 2106
rect 10296 2004 10330 2038
rect 10380 2140 10414 2174
rect 10380 2072 10414 2106
rect 10380 2004 10414 2038
rect 10525 2140 10559 2174
rect 10525 2072 10559 2106
rect 10525 2004 10559 2038
rect 10609 2140 10643 2174
rect 10609 2072 10643 2106
rect 10609 2004 10643 2038
rect 10693 2140 10727 2174
rect 10693 2072 10727 2106
rect 10693 2004 10727 2038
rect 10296 1340 10330 1374
rect 10296 1272 10330 1306
rect 10296 1204 10330 1238
rect 10380 1340 10414 1374
rect 10380 1272 10414 1306
rect 10380 1204 10414 1238
rect 10525 1340 10559 1374
rect 10525 1272 10559 1306
rect 10525 1204 10559 1238
rect 10621 1272 10655 1306
rect 10621 1204 10655 1238
rect 10705 1340 10739 1374
rect 10705 1272 10739 1306
rect 10705 1204 10739 1238
rect 10789 1340 10823 1374
rect 10789 1272 10823 1306
rect 10789 1204 10823 1238
rect 10290 1052 10324 1086
rect 10290 984 10324 1018
rect 10290 916 10324 950
rect 10374 1052 10408 1086
rect 10374 984 10408 1018
rect 10374 916 10408 950
rect 10566 1052 10600 1086
rect 10566 984 10600 1018
rect 10566 916 10600 950
rect 10650 1052 10684 1086
rect 10650 984 10684 1018
rect 10650 916 10684 950
rect 3850 -1669 3884 307
rect 5908 -1669 5942 307
rect 7966 -1669 8000 307
rect 10024 -1669 10058 307
rect 10252 73 10286 133
rect 10348 73 10382 133
rect 10444 73 10478 133
rect 10540 73 10574 133
rect 10636 73 10670 133
rect 10252 -343 10286 -283
rect 10348 -343 10382 -283
rect 10444 -343 10478 -283
rect 10540 -343 10574 -283
rect 10636 -343 10670 -283
<< psubdiff >>
rect 10246 -836 10342 -802
rect 10700 -836 10796 -802
rect 10246 -898 10280 -836
rect 10762 -898 10796 -836
rect 10246 -1200 10280 -1138
rect 10762 -1200 10796 -1138
rect 10246 -1234 10342 -1200
rect 10700 -1234 10796 -1200
rect 10246 -1296 10280 -1234
rect 10762 -1296 10796 -1234
rect 10246 -1598 10280 -1536
rect 10762 -1598 10796 -1536
rect 10246 -1632 10342 -1598
rect 10700 -1632 10796 -1598
<< nsubdiff >>
rect 3736 2800 3832 2834
rect 10076 2800 10172 2834
rect 3736 2738 3770 2800
rect 10138 2738 10172 2800
rect 3736 502 3770 564
rect 10138 502 10172 564
rect 3736 468 3832 502
rect 10076 468 10172 502
rect 3736 406 3770 468
rect 10138 406 10172 468
rect 3736 -1830 3770 -1768
rect 10172 294 10234 328
rect 10688 294 10784 328
rect 10750 232 10784 294
rect 10750 -88 10784 -26
rect 10172 -122 10234 -88
rect 10688 -122 10784 -88
rect 10750 -184 10784 -122
rect 10750 -504 10784 -442
rect 10172 -538 10234 -504
rect 10688 -538 10784 -504
rect 10138 -1830 10172 -1768
rect 3736 -1864 3832 -1830
rect 10076 -1864 10172 -1830
<< psubdiffcont >>
rect 10342 -836 10700 -802
rect 10246 -1138 10280 -898
rect 10762 -1138 10796 -898
rect 10342 -1234 10700 -1200
rect 10246 -1536 10280 -1296
rect 10762 -1536 10796 -1296
rect 10342 -1632 10700 -1598
<< nsubdiffcont >>
rect 3832 2800 10076 2834
rect 3736 564 3770 2738
rect 10138 564 10172 2738
rect 3832 468 10076 502
rect 3736 -1768 3770 406
rect 10138 -1768 10172 406
rect 10234 294 10688 328
rect 10750 -26 10784 232
rect 10234 -122 10688 -88
rect 10750 -442 10784 -184
rect 10234 -538 10688 -504
rect 3832 -1864 10076 -1830
<< poly >>
rect 3896 2732 5896 2748
rect 3896 2698 3912 2732
rect 5880 2698 5896 2732
rect 3896 2651 5896 2698
rect 5954 2732 7954 2748
rect 5954 2698 5970 2732
rect 7938 2698 7954 2732
rect 5954 2651 7954 2698
rect 8012 2732 10012 2748
rect 8012 2698 8028 2732
rect 9996 2698 10012 2732
rect 8012 2651 10012 2698
rect 3896 604 5896 651
rect 3896 570 3912 604
rect 5880 570 5896 604
rect 3896 554 5896 570
rect 5954 604 7954 651
rect 5954 570 5970 604
rect 7938 570 7954 604
rect 5954 554 7954 570
rect 8012 604 10012 651
rect 8012 570 8028 604
rect 9996 570 10012 604
rect 8012 554 10012 570
rect 10340 2730 10370 2756
rect 10569 2730 10599 2756
rect 10653 2730 10683 2756
rect 10340 2578 10370 2600
rect 10569 2578 10599 2600
rect 10340 2562 10426 2578
rect 10340 2528 10376 2562
rect 10410 2528 10426 2562
rect 10340 2512 10426 2528
rect 10511 2562 10599 2578
rect 10511 2528 10528 2562
rect 10562 2528 10599 2562
rect 10511 2512 10599 2528
rect 10340 2480 10370 2512
rect 10569 2480 10599 2512
rect 10653 2578 10683 2600
rect 10653 2562 10745 2578
rect 10653 2528 10696 2562
rect 10730 2528 10745 2562
rect 10653 2512 10745 2528
rect 10653 2480 10683 2512
rect 10340 2254 10370 2280
rect 10569 2254 10599 2280
rect 10653 2254 10683 2280
rect 10340 2186 10370 2212
rect 10569 2186 10599 2212
rect 10653 2186 10683 2212
rect 10340 1954 10370 1986
rect 10569 1954 10599 1986
rect 10340 1938 10426 1954
rect 10340 1904 10376 1938
rect 10410 1904 10426 1938
rect 10340 1888 10426 1904
rect 10511 1938 10599 1954
rect 10511 1904 10528 1938
rect 10562 1904 10599 1938
rect 10511 1888 10599 1904
rect 10340 1866 10370 1888
rect 10569 1866 10599 1888
rect 10653 1954 10683 1986
rect 10653 1938 10745 1954
rect 10653 1904 10696 1938
rect 10730 1904 10745 1938
rect 10653 1888 10745 1904
rect 10653 1866 10683 1888
rect 10340 1710 10370 1736
rect 10569 1710 10599 1736
rect 10653 1710 10683 1736
rect 10340 1642 10370 1668
rect 10569 1642 10599 1668
rect 10665 1642 10695 1668
rect 10749 1642 10779 1668
rect 10340 1490 10370 1512
rect 10569 1490 10599 1512
rect 10665 1490 10695 1512
rect 10340 1474 10426 1490
rect 10340 1440 10376 1474
rect 10410 1440 10426 1474
rect 10340 1424 10426 1440
rect 10520 1474 10599 1490
rect 10520 1440 10530 1474
rect 10564 1440 10599 1474
rect 10520 1424 10599 1440
rect 10641 1474 10695 1490
rect 10641 1440 10651 1474
rect 10685 1440 10695 1474
rect 10641 1424 10695 1440
rect 10340 1392 10370 1424
rect 10569 1392 10599 1424
rect 10665 1392 10695 1424
rect 10749 1490 10779 1512
rect 10749 1474 10836 1490
rect 10749 1440 10792 1474
rect 10826 1440 10836 1474
rect 10749 1424 10836 1440
rect 10749 1392 10779 1424
rect 10340 1166 10370 1192
rect 10569 1166 10599 1192
rect 10665 1166 10695 1192
rect 10749 1166 10779 1192
rect 10334 1098 10364 1124
rect 10610 1098 10640 1124
rect 10334 866 10364 898
rect 10610 866 10640 898
rect 10278 850 10364 866
rect 10278 816 10294 850
rect 10328 816 10364 850
rect 10278 800 10364 816
rect 10554 850 10640 866
rect 10554 816 10570 850
rect 10604 816 10640 850
rect 10554 800 10640 816
rect 10334 778 10364 800
rect 10610 778 10640 800
rect 10334 622 10364 648
rect 10610 622 10640 648
rect 3896 400 5896 416
rect 3896 366 3912 400
rect 5880 366 5896 400
rect 3896 319 5896 366
rect 5954 400 7954 416
rect 5954 366 5970 400
rect 7938 366 7954 400
rect 5954 319 7954 366
rect 8012 400 10012 416
rect 8012 366 8028 400
rect 9996 366 10012 400
rect 8012 319 10012 366
rect 3896 -1728 5896 -1681
rect 3896 -1762 3912 -1728
rect 5880 -1762 5896 -1728
rect 3896 -1778 5896 -1762
rect 5954 -1728 7954 -1681
rect 5954 -1762 5970 -1728
rect 7938 -1762 7954 -1728
rect 5954 -1778 7954 -1762
rect 8012 -1728 10012 -1681
rect 8012 -1762 8028 -1728
rect 9996 -1762 10012 -1728
rect 8012 -1778 10012 -1762
rect 10380 226 10446 242
rect 10380 192 10396 226
rect 10430 192 10446 226
rect 10380 176 10446 192
rect 10572 226 10638 242
rect 10572 192 10588 226
rect 10622 192 10638 226
rect 10572 176 10638 192
rect 10302 145 10332 171
rect 10398 145 10428 176
rect 10494 145 10524 171
rect 10590 145 10620 176
rect 10302 30 10332 61
rect 10398 35 10428 61
rect 10494 30 10524 61
rect 10590 35 10620 61
rect 10284 14 10350 30
rect 10284 -20 10300 14
rect 10334 -20 10350 14
rect 10284 -36 10350 -20
rect 10476 14 10542 30
rect 10476 -20 10492 14
rect 10526 -20 10542 14
rect 10476 -36 10542 -20
rect 10284 -190 10350 -174
rect 10284 -224 10300 -190
rect 10334 -224 10350 -190
rect 10284 -240 10350 -224
rect 10476 -190 10542 -174
rect 10476 -224 10492 -190
rect 10526 -224 10542 -190
rect 10476 -240 10542 -224
rect 10302 -271 10332 -240
rect 10398 -271 10428 -245
rect 10494 -271 10524 -240
rect 10590 -271 10620 -245
rect 10302 -381 10332 -355
rect 10398 -386 10428 -355
rect 10494 -381 10524 -355
rect 10590 -386 10620 -355
rect 10380 -402 10446 -386
rect 10380 -436 10396 -402
rect 10430 -436 10446 -402
rect 10380 -452 10446 -436
rect 10572 -402 10638 -386
rect 10572 -436 10588 -402
rect 10622 -436 10638 -402
rect 10572 -452 10638 -436
rect 10392 -904 10458 -888
rect 10392 -938 10408 -904
rect 10442 -938 10458 -904
rect 10392 -954 10458 -938
rect 10584 -904 10650 -888
rect 10584 -938 10600 -904
rect 10634 -938 10650 -904
rect 10410 -976 10440 -954
rect 10506 -976 10536 -950
rect 10584 -954 10650 -938
rect 10602 -976 10632 -954
rect 10410 -1086 10440 -1060
rect 10506 -1082 10536 -1060
rect 10488 -1098 10554 -1082
rect 10602 -1086 10632 -1060
rect 10488 -1132 10504 -1098
rect 10538 -1132 10554 -1098
rect 10488 -1148 10554 -1132
rect 10488 -1302 10554 -1286
rect 10488 -1336 10504 -1302
rect 10538 -1336 10554 -1302
rect 10410 -1374 10440 -1348
rect 10488 -1352 10554 -1336
rect 10506 -1374 10536 -1352
rect 10602 -1374 10632 -1348
rect 10410 -1480 10440 -1458
rect 10392 -1496 10458 -1480
rect 10506 -1484 10536 -1458
rect 10602 -1480 10632 -1458
rect 10392 -1530 10408 -1496
rect 10442 -1530 10458 -1496
rect 10392 -1546 10458 -1530
rect 10584 -1496 10650 -1480
rect 10584 -1530 10600 -1496
rect 10634 -1530 10650 -1496
rect 10584 -1546 10650 -1530
<< polycont >>
rect 3912 2698 5880 2732
rect 5970 2698 7938 2732
rect 8028 2698 9996 2732
rect 3912 570 5880 604
rect 5970 570 7938 604
rect 8028 570 9996 604
rect 10376 2528 10410 2562
rect 10528 2528 10562 2562
rect 10696 2528 10730 2562
rect 10376 1904 10410 1938
rect 10528 1904 10562 1938
rect 10696 1904 10730 1938
rect 10376 1440 10410 1474
rect 10530 1440 10564 1474
rect 10651 1440 10685 1474
rect 10792 1440 10826 1474
rect 10294 816 10328 850
rect 10570 816 10604 850
rect 3912 366 5880 400
rect 5970 366 7938 400
rect 8028 366 9996 400
rect 3912 -1762 5880 -1728
rect 5970 -1762 7938 -1728
rect 8028 -1762 9996 -1728
rect 10396 192 10430 226
rect 10588 192 10622 226
rect 10300 -20 10334 14
rect 10492 -20 10526 14
rect 10300 -224 10334 -190
rect 10492 -224 10526 -190
rect 10396 -436 10430 -402
rect 10588 -436 10622 -402
rect 10408 -938 10442 -904
rect 10600 -938 10634 -904
rect 10504 -1132 10538 -1098
rect 10504 -1336 10538 -1302
rect 10408 -1530 10442 -1496
rect 10600 -1530 10634 -1496
<< locali >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2834 10170 2870
rect 10100 2830 10172 2834
rect 3700 2800 3832 2830
rect 10076 2800 10172 2830
rect 3700 2770 3800 2800
rect 3700 -1770 3710 2770
rect 3780 502 3800 2770
rect 10138 2740 10172 2800
rect 10214 2760 10243 2794
rect 10277 2760 10335 2794
rect 10369 2760 10427 2794
rect 10461 2760 10519 2794
rect 10553 2760 10611 2794
rect 10645 2760 10703 2794
rect 10737 2760 10766 2794
rect 10170 2738 10172 2740
rect 3896 2698 3912 2732
rect 5880 2698 5896 2732
rect 5954 2698 5970 2732
rect 7938 2698 7954 2732
rect 8012 2698 8028 2732
rect 9996 2698 10012 2732
rect 3850 2639 3884 2655
rect 3850 647 3884 663
rect 5908 2639 5942 2655
rect 5908 647 5942 663
rect 7966 2639 8000 2655
rect 7966 647 8000 663
rect 10024 2639 10058 2655
rect 10024 647 10058 663
rect 3896 570 3912 604
rect 5880 570 5896 604
rect 5954 570 5970 604
rect 7938 570 7954 604
rect 8012 570 8028 604
rect 9996 570 10012 604
rect 10280 2714 10346 2726
rect 10280 2680 10296 2714
rect 10330 2680 10346 2714
rect 10280 2646 10346 2680
rect 10280 2612 10296 2646
rect 10330 2612 10346 2646
rect 10280 2600 10346 2612
rect 10380 2714 10426 2760
rect 10414 2680 10426 2714
rect 10380 2646 10426 2680
rect 10414 2612 10426 2646
rect 10280 2480 10326 2600
rect 10380 2596 10426 2612
rect 10507 2718 10646 2726
rect 10507 2684 10525 2718
rect 10559 2684 10646 2718
rect 10507 2650 10646 2684
rect 10507 2616 10525 2650
rect 10559 2616 10646 2650
rect 10507 2600 10646 2616
rect 10687 2718 10749 2760
rect 10687 2684 10693 2718
rect 10727 2684 10749 2718
rect 10687 2650 10749 2684
rect 10687 2616 10693 2650
rect 10727 2616 10749 2650
rect 10687 2600 10749 2616
rect 10577 2512 10578 2562
rect 10612 2480 10646 2600
rect 10280 2470 10346 2480
rect 10330 2410 10346 2470
rect 10280 2394 10346 2410
rect 10280 2360 10296 2394
rect 10330 2360 10346 2394
rect 10280 2326 10346 2360
rect 10280 2292 10296 2326
rect 10330 2292 10346 2326
rect 10280 2284 10346 2292
rect 10380 2462 10422 2478
rect 10414 2428 10422 2462
rect 10380 2394 10422 2428
rect 10414 2360 10422 2394
rect 10380 2326 10422 2360
rect 10414 2292 10422 2326
rect 10380 2250 10422 2292
rect 10507 2462 10559 2478
rect 10507 2428 10525 2462
rect 10507 2394 10559 2428
rect 10507 2360 10525 2394
rect 10507 2326 10559 2360
rect 10507 2292 10525 2326
rect 10507 2250 10559 2292
rect 10593 2462 10659 2480
rect 10593 2428 10609 2462
rect 10643 2428 10659 2462
rect 10593 2410 10659 2428
rect 10593 2350 10600 2410
rect 10650 2350 10659 2410
rect 10593 2326 10659 2350
rect 10593 2292 10609 2326
rect 10643 2292 10659 2326
rect 10593 2284 10659 2292
rect 10693 2462 10749 2478
rect 10727 2428 10749 2462
rect 10693 2394 10749 2428
rect 10727 2360 10749 2394
rect 10693 2326 10749 2360
rect 10727 2292 10749 2326
rect 10693 2250 10749 2292
rect 10214 2216 10243 2250
rect 10277 2216 10335 2250
rect 10369 2216 10427 2250
rect 10461 2216 10519 2250
rect 10553 2216 10611 2250
rect 10645 2216 10703 2250
rect 10737 2216 10766 2250
rect 10280 2174 10346 2182
rect 10280 2140 10296 2174
rect 10330 2140 10346 2174
rect 10280 2127 10346 2140
rect 10280 2072 10296 2077
rect 10330 2072 10346 2127
rect 10280 2038 10346 2072
rect 10280 2004 10296 2038
rect 10330 2004 10346 2038
rect 10280 1986 10346 2004
rect 10380 2174 10422 2216
rect 10414 2140 10422 2174
rect 10380 2106 10422 2140
rect 10414 2072 10422 2106
rect 10380 2038 10422 2072
rect 10414 2004 10422 2038
rect 10380 1988 10422 2004
rect 10507 2174 10559 2216
rect 10507 2140 10525 2174
rect 10507 2106 10559 2140
rect 10507 2072 10525 2106
rect 10507 2038 10559 2072
rect 10507 2004 10525 2038
rect 10507 1988 10559 2004
rect 10593 2174 10659 2182
rect 10593 2140 10609 2174
rect 10643 2140 10659 2174
rect 10593 2106 10659 2140
rect 10593 2072 10609 2106
rect 10643 2072 10659 2106
rect 10593 2038 10659 2072
rect 10593 2004 10609 2038
rect 10643 2004 10659 2038
rect 10593 1986 10659 2004
rect 10693 2174 10749 2216
rect 10727 2140 10749 2174
rect 10693 2106 10749 2140
rect 10727 2072 10749 2106
rect 10693 2038 10749 2072
rect 10727 2004 10749 2038
rect 10693 1988 10749 2004
rect 10280 1866 10326 1986
rect 10360 1904 10362 1952
rect 10423 1904 10426 1952
rect 10280 1854 10346 1866
rect 10280 1820 10296 1854
rect 10330 1820 10346 1854
rect 10280 1786 10346 1820
rect 10280 1752 10296 1786
rect 10330 1752 10346 1786
rect 10280 1740 10346 1752
rect 10380 1854 10426 1870
rect 10612 1866 10646 1986
rect 10414 1820 10426 1854
rect 10380 1786 10426 1820
rect 10414 1752 10426 1786
rect 10380 1706 10426 1752
rect 10507 1850 10646 1866
rect 10507 1838 10525 1850
rect 10559 1838 10646 1850
rect 10507 1789 10519 1838
rect 10580 1789 10646 1838
rect 10507 1782 10646 1789
rect 10507 1748 10525 1782
rect 10559 1748 10646 1782
rect 10507 1740 10646 1748
rect 10687 1850 10749 1866
rect 10687 1816 10693 1850
rect 10727 1816 10749 1850
rect 10687 1782 10749 1816
rect 10687 1748 10693 1782
rect 10727 1748 10749 1782
rect 10687 1706 10749 1748
rect 10214 1672 10243 1706
rect 10277 1672 10335 1706
rect 10369 1672 10427 1706
rect 10461 1672 10519 1706
rect 10553 1672 10611 1706
rect 10645 1672 10703 1706
rect 10737 1672 10795 1706
rect 10829 1672 10858 1706
rect 10280 1626 10346 1638
rect 10280 1592 10296 1626
rect 10330 1592 10346 1626
rect 10280 1580 10346 1592
rect 10340 1520 10346 1580
rect 10280 1512 10346 1520
rect 10380 1626 10426 1672
rect 10414 1592 10426 1626
rect 10380 1558 10426 1592
rect 10414 1524 10426 1558
rect 10509 1630 10755 1638
rect 10509 1596 10525 1630
rect 10559 1604 10755 1630
rect 10559 1596 10629 1604
rect 10509 1570 10629 1596
rect 10663 1570 10755 1604
rect 10789 1624 10840 1672
rect 10823 1590 10840 1624
rect 10789 1574 10840 1590
rect 10509 1562 10575 1570
rect 10509 1528 10525 1562
rect 10559 1528 10575 1562
rect 10509 1524 10575 1528
rect 10280 1392 10326 1512
rect 10380 1508 10426 1524
rect 10610 1490 10685 1536
rect 10610 1430 10620 1490
rect 10680 1474 10685 1490
rect 10680 1430 10685 1440
rect 10610 1424 10685 1430
rect 10280 1374 10346 1392
rect 10719 1390 10755 1570
rect 10792 1500 10836 1540
rect 10792 1474 10800 1500
rect 10792 1430 10800 1440
rect 10792 1424 10836 1430
rect 10280 1340 10296 1374
rect 10330 1340 10346 1374
rect 10280 1306 10346 1340
rect 10280 1272 10296 1306
rect 10330 1272 10346 1306
rect 10280 1238 10346 1272
rect 10280 1204 10296 1238
rect 10330 1204 10346 1238
rect 10280 1196 10346 1204
rect 10380 1374 10422 1390
rect 10414 1340 10422 1374
rect 10380 1306 10422 1340
rect 10414 1272 10422 1306
rect 10380 1238 10422 1272
rect 10414 1204 10422 1238
rect 10380 1162 10422 1204
rect 10509 1374 10755 1390
rect 10509 1340 10525 1374
rect 10559 1356 10705 1374
rect 10559 1340 10575 1356
rect 10509 1306 10575 1340
rect 10689 1340 10705 1356
rect 10739 1340 10755 1374
rect 10509 1272 10525 1306
rect 10559 1272 10575 1306
rect 10509 1238 10575 1272
rect 10509 1204 10525 1238
rect 10559 1204 10575 1238
rect 10509 1196 10575 1204
rect 10609 1306 10655 1322
rect 10609 1272 10621 1306
rect 10609 1238 10655 1272
rect 10609 1204 10621 1238
rect 10609 1162 10655 1204
rect 10689 1306 10755 1340
rect 10689 1272 10705 1306
rect 10739 1272 10755 1306
rect 10689 1238 10755 1272
rect 10689 1204 10705 1238
rect 10739 1204 10755 1238
rect 10689 1196 10755 1204
rect 10789 1374 10840 1390
rect 10823 1340 10840 1374
rect 10789 1306 10840 1340
rect 10823 1272 10840 1306
rect 10789 1238 10840 1272
rect 10823 1204 10840 1238
rect 10789 1162 10840 1204
rect 10214 1128 10243 1162
rect 10277 1128 10335 1162
rect 10369 1128 10427 1162
rect 10461 1128 10519 1162
rect 10553 1128 10611 1162
rect 10645 1128 10703 1162
rect 10737 1128 10795 1162
rect 10829 1128 10858 1162
rect 10282 1086 10324 1128
rect 10282 1052 10290 1086
rect 10282 1018 10324 1052
rect 10282 984 10290 1018
rect 10282 950 10324 984
rect 10282 916 10290 950
rect 10282 900 10324 916
rect 10358 1086 10424 1094
rect 10358 1052 10374 1086
rect 10408 1052 10424 1086
rect 10358 1018 10424 1052
rect 10358 1009 10374 1018
rect 10408 1009 10424 1018
rect 10558 1086 10600 1128
rect 10558 1052 10566 1086
rect 10558 1018 10600 1052
rect 10358 961 10360 1009
rect 10558 984 10566 1018
rect 10358 950 10424 961
rect 10358 916 10374 950
rect 10408 916 10424 950
rect 10358 898 10424 916
rect 10558 950 10600 984
rect 10558 916 10566 950
rect 10558 900 10600 916
rect 10634 1086 10700 1094
rect 10634 1052 10650 1086
rect 10684 1052 10700 1086
rect 10634 1025 10700 1052
rect 10699 977 10700 1025
rect 10634 950 10700 977
rect 10634 916 10650 950
rect 10684 916 10700 950
rect 10634 898 10700 916
rect 10343 816 10344 864
rect 10278 766 10324 782
rect 10378 778 10424 898
rect 10619 816 10620 864
rect 10278 732 10290 766
rect 10278 698 10324 732
rect 10278 664 10290 698
rect 10278 618 10324 664
rect 10358 766 10424 778
rect 10358 732 10374 766
rect 10408 732 10424 766
rect 10358 698 10424 732
rect 10358 664 10374 698
rect 10408 664 10424 698
rect 10358 652 10424 664
rect 10554 766 10600 782
rect 10654 778 10700 898
rect 10554 732 10566 766
rect 10554 698 10600 732
rect 10554 664 10566 698
rect 10554 618 10600 664
rect 10634 766 10700 778
rect 10634 732 10650 766
rect 10684 732 10700 766
rect 10634 698 10700 732
rect 10634 664 10650 698
rect 10684 664 10700 698
rect 10634 652 10700 664
rect 10214 584 10243 618
rect 10277 584 10335 618
rect 10369 584 10427 618
rect 10461 584 10519 618
rect 10553 584 10611 618
rect 10645 584 10703 618
rect 10737 584 10766 618
rect 3780 468 3832 502
rect 10076 468 10130 502
rect 3780 -1770 3800 468
rect 10170 406 10172 564
rect 3896 366 3912 400
rect 5880 366 5896 400
rect 5954 366 5970 400
rect 7938 366 7954 400
rect 8012 366 8028 400
rect 9996 366 10012 400
rect 3850 307 3884 323
rect 3850 -1685 3884 -1669
rect 5908 307 5942 323
rect 5908 -1685 5942 -1669
rect 7966 307 8000 323
rect 7966 -1685 8000 -1669
rect 10024 307 10058 323
rect 10172 294 10234 328
rect 10688 294 10784 328
rect 10750 232 10784 294
rect 10380 192 10396 226
rect 10430 192 10446 226
rect 10572 192 10588 226
rect 10622 192 10638 226
rect 10252 133 10286 149
rect 10252 57 10286 73
rect 10348 133 10382 149
rect 10348 57 10382 73
rect 10444 133 10478 149
rect 10444 57 10478 73
rect 10540 133 10574 149
rect 10540 57 10574 73
rect 10636 133 10670 149
rect 10636 57 10670 73
rect 10284 -20 10300 14
rect 10334 -20 10350 14
rect 10476 -20 10492 14
rect 10526 -20 10542 14
rect 10750 -88 10784 -26
rect 10172 -122 10234 -88
rect 10688 -122 10784 -88
rect 10750 -184 10784 -122
rect 10284 -224 10300 -190
rect 10334 -224 10350 -190
rect 10476 -224 10492 -190
rect 10526 -224 10542 -190
rect 10252 -283 10286 -267
rect 10252 -359 10286 -343
rect 10348 -283 10382 -267
rect 10348 -359 10382 -343
rect 10444 -283 10478 -267
rect 10444 -359 10478 -343
rect 10540 -283 10574 -267
rect 10540 -359 10574 -343
rect 10636 -283 10670 -267
rect 10636 -359 10670 -343
rect 10380 -436 10396 -402
rect 10430 -436 10446 -402
rect 10572 -436 10588 -402
rect 10622 -436 10638 -402
rect 10750 -504 10784 -442
rect 10172 -538 10234 -504
rect 10688 -538 10784 -504
rect 10024 -1685 10058 -1669
rect 3896 -1762 3912 -1728
rect 5880 -1762 5896 -1728
rect 5954 -1762 5970 -1728
rect 7938 -1762 7954 -1728
rect 8012 -1762 8028 -1728
rect 9996 -1762 10012 -1728
rect 3700 -1830 3800 -1770
rect 10246 -830 10250 -802
rect 10310 -802 10340 -770
rect 10310 -830 10342 -802
rect 10246 -836 10342 -830
rect 10700 -836 10796 -802
rect 10246 -898 10280 -836
rect 10762 -898 10796 -836
rect 10392 -938 10408 -904
rect 10442 -938 10458 -904
rect 10584 -938 10600 -904
rect 10634 -938 10650 -904
rect 10360 -988 10394 -972
rect 10360 -1064 10394 -1048
rect 10456 -988 10490 -972
rect 10456 -1064 10490 -1048
rect 10552 -988 10586 -972
rect 10552 -1064 10586 -1048
rect 10648 -988 10682 -972
rect 10648 -1064 10682 -1048
rect 10488 -1132 10504 -1098
rect 10538 -1132 10554 -1098
rect 10246 -1200 10280 -1138
rect 10762 -1200 10796 -1138
rect 10246 -1234 10342 -1200
rect 10700 -1234 10796 -1200
rect 10246 -1296 10280 -1234
rect 10762 -1296 10796 -1234
rect 10488 -1336 10504 -1302
rect 10538 -1336 10554 -1302
rect 10360 -1386 10394 -1370
rect 10360 -1462 10394 -1446
rect 10456 -1386 10490 -1370
rect 10456 -1462 10490 -1446
rect 10552 -1386 10586 -1370
rect 10552 -1462 10586 -1446
rect 10648 -1386 10682 -1370
rect 10648 -1462 10682 -1446
rect 10392 -1530 10408 -1496
rect 10442 -1530 10458 -1496
rect 10584 -1530 10600 -1496
rect 10634 -1530 10650 -1496
rect 10246 -1598 10280 -1536
rect 10762 -1598 10796 -1536
rect 10246 -1632 10342 -1598
rect 10700 -1632 10796 -1598
rect 10138 -1830 10172 -1768
rect 3700 -1840 3832 -1830
rect 10076 -1840 10172 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1864 10172 -1840
rect 10100 -1890 10140 -1864
rect 3700 -1900 10140 -1890
<< viali >>
rect 3830 2834 10100 2870
rect 3830 2830 3832 2834
rect 3832 2830 10076 2834
rect 10076 2830 10100 2834
rect 3710 2738 3780 2770
rect 3710 564 3736 2738
rect 3736 564 3770 2738
rect 3770 564 3780 2738
rect 3710 406 3780 564
rect 10243 2760 10277 2794
rect 10335 2760 10369 2794
rect 10427 2760 10461 2794
rect 10519 2760 10553 2794
rect 10611 2760 10645 2794
rect 10703 2760 10737 2794
rect 10130 2738 10170 2740
rect 3912 2698 5880 2732
rect 5970 2698 7938 2732
rect 8028 2698 9996 2732
rect 3850 663 3884 2639
rect 5908 663 5942 2639
rect 7966 663 8000 2639
rect 10024 663 10058 2639
rect 3912 570 5880 604
rect 5970 570 7938 604
rect 8028 570 9996 604
rect 10130 564 10138 2738
rect 10138 564 10170 2738
rect 10360 2528 10376 2562
rect 10376 2528 10410 2562
rect 10410 2528 10426 2562
rect 10360 2514 10426 2528
rect 10511 2528 10528 2562
rect 10528 2528 10562 2562
rect 10562 2528 10577 2562
rect 10511 2512 10577 2528
rect 10680 2562 10747 2566
rect 10680 2528 10696 2562
rect 10696 2528 10730 2562
rect 10730 2528 10747 2562
rect 10680 2512 10747 2528
rect 10280 2462 10330 2470
rect 10280 2428 10296 2462
rect 10296 2428 10330 2462
rect 10280 2410 10330 2428
rect 10600 2394 10650 2410
rect 10600 2360 10609 2394
rect 10609 2360 10643 2394
rect 10643 2360 10650 2394
rect 10600 2350 10650 2360
rect 10243 2216 10277 2250
rect 10335 2216 10369 2250
rect 10427 2216 10461 2250
rect 10519 2216 10553 2250
rect 10611 2216 10645 2250
rect 10703 2216 10737 2250
rect 10280 2106 10330 2127
rect 10280 2077 10296 2106
rect 10296 2077 10330 2106
rect 10362 1938 10423 1953
rect 10362 1904 10376 1938
rect 10376 1904 10410 1938
rect 10410 1904 10423 1938
rect 10511 1938 10578 1954
rect 10511 1904 10528 1938
rect 10528 1904 10562 1938
rect 10562 1904 10578 1938
rect 10680 1938 10747 1954
rect 10680 1904 10696 1938
rect 10696 1904 10730 1938
rect 10730 1904 10747 1938
rect 10680 1900 10747 1904
rect 10519 1816 10525 1838
rect 10525 1816 10559 1838
rect 10559 1816 10580 1838
rect 10519 1789 10580 1816
rect 10243 1672 10277 1706
rect 10335 1672 10369 1706
rect 10427 1672 10461 1706
rect 10519 1672 10553 1706
rect 10611 1672 10645 1706
rect 10703 1672 10737 1706
rect 10795 1672 10829 1706
rect 10280 1558 10340 1580
rect 10280 1524 10296 1558
rect 10296 1524 10330 1558
rect 10330 1524 10340 1558
rect 10280 1520 10340 1524
rect 10629 1570 10663 1604
rect 10507 1474 10570 1490
rect 10360 1440 10376 1474
rect 10376 1440 10410 1474
rect 10410 1440 10426 1474
rect 10360 1426 10426 1440
rect 10507 1440 10530 1474
rect 10530 1440 10564 1474
rect 10564 1440 10570 1474
rect 10507 1424 10570 1440
rect 10620 1474 10680 1490
rect 10620 1440 10651 1474
rect 10651 1440 10680 1474
rect 10620 1430 10680 1440
rect 10800 1474 10860 1500
rect 10800 1440 10826 1474
rect 10826 1440 10860 1474
rect 10800 1430 10860 1440
rect 10243 1128 10277 1162
rect 10335 1128 10369 1162
rect 10427 1128 10461 1162
rect 10519 1128 10553 1162
rect 10611 1128 10645 1162
rect 10703 1128 10737 1162
rect 10795 1128 10829 1162
rect 10360 984 10374 1009
rect 10374 984 10408 1009
rect 10408 984 10425 1009
rect 10360 961 10425 984
rect 10634 1018 10699 1025
rect 10634 984 10650 1018
rect 10650 984 10684 1018
rect 10684 984 10699 1018
rect 10634 977 10699 984
rect 10278 850 10343 864
rect 10278 816 10294 850
rect 10294 816 10328 850
rect 10328 816 10343 850
rect 10554 850 10619 864
rect 10554 816 10570 850
rect 10570 816 10604 850
rect 10604 816 10619 850
rect 10243 584 10277 618
rect 10335 584 10369 618
rect 10427 584 10461 618
rect 10519 584 10553 618
rect 10611 584 10645 618
rect 10703 584 10737 618
rect 3710 -1768 3736 406
rect 3736 -1768 3770 406
rect 3770 -1768 3780 406
rect 3710 -1770 3780 -1768
rect 10130 406 10170 564
rect 3912 366 5880 400
rect 5970 366 7938 400
rect 8028 366 9996 400
rect 3850 -1669 3884 307
rect 5908 -1669 5942 307
rect 7966 -1669 8000 307
rect 10024 -1669 10058 307
rect 10130 -540 10138 406
rect 10138 -540 10170 406
rect 10396 192 10430 226
rect 10588 192 10622 226
rect 10252 73 10286 133
rect 10348 73 10382 133
rect 10444 73 10478 133
rect 10540 73 10574 133
rect 10636 73 10670 133
rect 10300 -20 10334 14
rect 10492 -20 10526 14
rect 10300 -224 10334 -190
rect 10492 -224 10526 -190
rect 10252 -343 10286 -283
rect 10348 -343 10382 -283
rect 10444 -343 10478 -283
rect 10540 -343 10574 -283
rect 10636 -343 10670 -283
rect 10396 -436 10430 -402
rect 10588 -436 10622 -402
rect 3912 -1762 5880 -1728
rect 5970 -1762 7938 -1728
rect 8028 -1762 9996 -1728
rect 10250 -830 10310 -770
rect 10408 -938 10442 -904
rect 10600 -938 10634 -904
rect 10360 -1048 10394 -988
rect 10456 -1048 10490 -988
rect 10552 -1048 10586 -988
rect 10648 -1048 10682 -988
rect 10504 -1132 10538 -1098
rect 10504 -1336 10538 -1302
rect 10360 -1446 10394 -1386
rect 10456 -1446 10490 -1386
rect 10552 -1446 10586 -1386
rect 10648 -1446 10682 -1386
rect 10408 -1530 10442 -1496
rect 10600 -1530 10634 -1496
rect 3820 -1864 3832 -1840
rect 3832 -1864 10076 -1840
rect 10076 -1864 10100 -1840
rect 3820 -1890 10100 -1864
<< metal1 >>
rect 3700 2870 10170 2900
rect 3700 2830 3830 2870
rect 10100 2830 10170 2870
rect 3700 2810 10170 2830
rect 10210 2810 11700 2900
rect 3700 2770 3800 2810
rect 3700 -1770 3710 2770
rect 3780 1840 3800 2770
rect 10130 2752 10170 2810
rect 10214 2794 10766 2810
rect 10214 2760 10243 2794
rect 10277 2760 10335 2794
rect 10369 2760 10427 2794
rect 10461 2760 10519 2794
rect 10553 2760 10611 2794
rect 10645 2760 10703 2794
rect 10737 2760 10766 2794
rect 6880 2740 6890 2750
rect 3900 2732 6890 2740
rect 6950 2740 6960 2750
rect 10124 2740 10176 2752
rect 6950 2732 10020 2740
rect 3900 2698 3912 2732
rect 5880 2698 5970 2732
rect 7938 2698 8028 2732
rect 9996 2698 10020 2732
rect 3900 2690 6890 2698
rect 6950 2690 10020 2698
rect 3844 2639 3890 2651
rect 3844 1840 3850 2639
rect 3780 1500 3850 1840
rect 3780 -600 3800 1500
rect 3844 663 3850 1500
rect 3884 1840 3890 2639
rect 5902 2639 5948 2651
rect 5902 1840 5908 2639
rect 3884 1500 5908 1840
rect 3884 663 3890 1500
rect 3844 651 3890 663
rect 5902 663 5908 1500
rect 5942 1840 5948 2639
rect 7960 2639 8006 2651
rect 7960 1840 7966 2639
rect 5942 1500 7966 1840
rect 5942 663 5948 1500
rect 5902 651 5948 663
rect 7960 663 7966 1500
rect 8000 1840 8006 2639
rect 10018 2639 10064 2651
rect 10018 1840 10024 2639
rect 8000 1500 10024 1840
rect 8000 663 8006 1500
rect 7960 651 8006 663
rect 10018 663 10024 1500
rect 10058 1840 10064 2639
rect 10124 1840 10130 2740
rect 10058 1500 10130 1840
rect 10058 663 10064 1500
rect 10018 651 10064 663
rect 6880 610 6890 620
rect 3890 604 6890 610
rect 6950 610 6960 620
rect 6950 604 10010 610
rect 3890 570 3912 604
rect 5880 570 5970 604
rect 7938 570 8028 604
rect 9996 570 10010 604
rect 3890 560 6890 570
rect 6950 560 10010 570
rect 6880 410 6890 420
rect 3890 400 6890 410
rect 6950 410 6960 420
rect 6950 400 10010 410
rect 3890 366 3912 400
rect 5880 366 5970 400
rect 7938 366 8028 400
rect 9996 366 10010 400
rect 3890 360 6890 366
rect 6950 360 10010 366
rect 3844 307 3890 319
rect 3844 -600 3850 307
rect 3780 -940 3850 -600
rect 3780 -1770 3800 -940
rect 3844 -1669 3850 -940
rect 3884 -600 3890 307
rect 5902 307 5948 319
rect 5902 -600 5908 307
rect 3884 -940 5908 -600
rect 3884 -1669 3890 -940
rect 3844 -1681 3890 -1669
rect 5902 -1669 5908 -940
rect 5942 -600 5948 307
rect 7960 307 8006 319
rect 7960 -600 7966 307
rect 5942 -940 7966 -600
rect 5942 -1669 5948 -940
rect 5902 -1681 5948 -1669
rect 7960 -1669 7966 -940
rect 8000 -600 8006 307
rect 10018 307 10064 319
rect 9730 70 9740 130
rect 9800 70 9810 130
rect 9750 -460 9790 70
rect 9730 -520 9740 -460
rect 9800 -520 9810 -460
rect 10018 -600 10024 307
rect 8000 -940 10024 -600
rect 8000 -1669 8006 -940
rect 7960 -1681 8006 -1669
rect 10018 -1669 10024 -940
rect 10058 -600 10064 307
rect 10124 -70 10130 1500
rect 10170 2280 10176 2740
rect 10214 2729 10766 2760
rect 10670 2572 10680 2580
rect 10510 2568 10520 2570
rect 10348 2562 10438 2568
rect 10348 2514 10360 2562
rect 10426 2514 10438 2562
rect 10348 2508 10438 2514
rect 10499 2562 10520 2568
rect 10499 2512 10511 2562
rect 10499 2510 10520 2512
rect 10580 2510 10590 2570
rect 10668 2510 10680 2572
rect 10750 2510 10760 2580
rect 11000 2520 11010 2580
rect 11070 2520 11080 2580
rect 10274 2470 10336 2482
rect 10250 2410 10260 2470
rect 10330 2410 10336 2470
rect 10274 2398 10336 2410
rect 10378 2392 10410 2508
rect 10499 2506 10589 2510
rect 10668 2506 10759 2510
rect 10594 2410 10656 2422
rect 10594 2400 10600 2410
rect 10650 2400 10656 2410
rect 10580 2392 10590 2400
rect 10378 2347 10590 2392
rect 10580 2340 10590 2347
rect 10650 2340 10660 2400
rect 10594 2338 10656 2340
rect 10214 2280 10766 2281
rect 10170 2250 10766 2280
rect 10170 2216 10243 2250
rect 10277 2216 10335 2250
rect 10369 2216 10427 2250
rect 10461 2216 10519 2250
rect 10553 2216 10611 2250
rect 10645 2216 10703 2250
rect 10737 2216 10766 2250
rect 10170 2190 10766 2216
rect 10170 1190 10176 2190
rect 10214 2185 10766 2190
rect 10270 2133 10280 2137
rect 10268 2077 10280 2133
rect 10340 2077 10350 2137
rect 10268 2071 10342 2077
rect 11030 1960 11060 2520
rect 11100 2430 11110 2490
rect 11170 2430 11180 2490
rect 10350 1953 10435 1959
rect 10350 1904 10362 1953
rect 10423 1904 10435 1953
rect 10350 1898 10435 1904
rect 10499 1900 10510 1960
rect 10570 1954 10590 1960
rect 10578 1904 10590 1954
rect 10570 1900 10590 1904
rect 10499 1898 10590 1900
rect 10390 1830 10420 1898
rect 10668 1894 10680 1960
rect 10670 1890 10680 1894
rect 10750 1890 10760 1960
rect 11000 1900 11010 1960
rect 11070 1900 11080 1960
rect 10510 1844 10520 1850
rect 10507 1838 10520 1844
rect 10580 1844 10590 1850
rect 10507 1830 10519 1838
rect 10390 1800 10519 1830
rect 10507 1789 10519 1800
rect 10580 1789 10592 1844
rect 10920 1790 10930 1850
rect 10990 1790 11000 1850
rect 10507 1783 10592 1789
rect 10214 1720 10858 1737
rect 10214 1706 10760 1720
rect 10214 1672 10243 1706
rect 10277 1672 10335 1706
rect 10369 1672 10427 1706
rect 10461 1672 10519 1706
rect 10553 1672 10611 1706
rect 10645 1672 10703 1706
rect 10737 1672 10760 1706
rect 10214 1650 10760 1672
rect 10830 1650 10858 1720
rect 10214 1641 10858 1650
rect 10597 1604 10679 1611
rect 10597 1600 10629 1604
rect 10663 1600 10679 1604
rect 10597 1590 10620 1600
rect 10268 1580 10352 1586
rect 10268 1520 10280 1580
rect 10340 1520 10352 1580
rect 10268 1514 10352 1520
rect 10400 1560 10620 1590
rect 10400 1480 10430 1560
rect 10610 1540 10620 1560
rect 10680 1540 10690 1600
rect 10501 1500 10576 1502
rect 10794 1500 10880 1512
rect 10490 1490 10580 1500
rect 10348 1474 10438 1480
rect 10348 1426 10360 1474
rect 10426 1426 10438 1474
rect 10348 1420 10438 1426
rect 10490 1424 10507 1490
rect 10570 1424 10580 1490
rect 10608 1490 10692 1496
rect 10794 1490 10800 1500
rect 10608 1430 10620 1490
rect 10680 1430 10692 1490
rect 10790 1430 10800 1490
rect 10860 1430 10880 1500
rect 10608 1424 10692 1430
rect 10490 1406 10580 1424
rect 10490 1340 10500 1406
rect 10563 1340 10580 1406
rect 10640 1290 10670 1424
rect 10794 1418 10880 1430
rect 10810 1417 10880 1418
rect 10810 1300 10850 1417
rect 10540 1230 10550 1290
rect 10610 1240 10670 1290
rect 10790 1240 10800 1300
rect 10860 1240 10870 1300
rect 10610 1230 10620 1240
rect 10214 1190 10858 1193
rect 10170 1162 10858 1190
rect 10170 1128 10243 1162
rect 10277 1128 10335 1162
rect 10369 1128 10427 1162
rect 10461 1128 10519 1162
rect 10553 1128 10611 1162
rect 10645 1128 10703 1162
rect 10737 1128 10795 1162
rect 10829 1128 10858 1162
rect 10170 1100 10858 1128
rect 10170 150 10176 1100
rect 10214 1097 10858 1100
rect 10622 1030 10711 1031
rect 10350 1015 10360 1020
rect 10348 960 10360 1015
rect 10420 1015 10430 1020
rect 10420 1009 10437 1015
rect 10425 961 10437 1009
rect 10620 970 10630 1030
rect 10700 971 10711 1030
rect 10700 970 10710 971
rect 10420 960 10437 961
rect 10348 955 10437 960
rect 10266 864 10355 870
rect 10266 860 10278 864
rect 10260 816 10278 860
rect 10343 816 10355 864
rect 10260 810 10355 816
rect 10540 810 10550 870
rect 10610 864 10631 870
rect 10619 816 10631 864
rect 10610 810 10631 816
rect 10260 740 10350 810
rect 10260 680 10270 740
rect 10330 690 10350 740
rect 10330 680 10340 690
rect 10214 630 10766 649
rect 10214 618 10690 630
rect 10214 584 10243 618
rect 10277 584 10335 618
rect 10369 584 10427 618
rect 10461 584 10519 618
rect 10553 584 10611 618
rect 10645 584 10690 618
rect 10214 560 10690 584
rect 10760 560 10770 630
rect 10214 553 10766 560
rect 10570 380 10580 440
rect 10640 380 10650 440
rect 10370 180 10380 250
rect 10450 180 10460 250
rect 10590 232 10620 380
rect 10576 226 10634 232
rect 10576 192 10588 226
rect 10622 192 10634 226
rect 10576 186 10634 192
rect 10170 145 10260 150
rect 10170 133 10292 145
rect 10342 142 10388 145
rect 10438 142 10484 145
rect 10170 73 10252 133
rect 10286 73 10292 133
rect 10170 61 10292 73
rect 10328 133 10388 142
rect 10328 132 10348 133
rect 10382 132 10388 133
rect 10328 62 10388 72
rect 10436 133 10496 142
rect 10436 132 10444 133
rect 10478 132 10496 133
rect 10436 62 10496 72
rect 10534 133 10580 145
rect 10534 73 10540 133
rect 10574 73 10580 133
rect 10342 61 10388 62
rect 10438 61 10484 62
rect 10534 61 10580 73
rect 10630 133 10676 145
rect 10630 73 10636 133
rect 10670 110 10676 133
rect 10670 80 10780 110
rect 10670 73 10676 80
rect 10630 61 10676 73
rect 10170 60 10260 61
rect 10170 -70 10176 60
rect 10270 -40 10280 20
rect 10340 -40 10350 20
rect 10480 14 10540 20
rect 10480 -20 10492 14
rect 10526 -20 10540 14
rect 10110 -130 10120 -70
rect 10180 -130 10190 -70
rect 10124 -540 10130 -130
rect 10170 -270 10176 -130
rect 10290 -184 10340 -40
rect 10480 -170 10540 -20
rect 10750 -70 10780 80
rect 10820 70 10830 130
rect 10890 70 10900 130
rect 10730 -130 10740 -70
rect 10800 -130 10810 -70
rect 10288 -190 10346 -184
rect 10288 -224 10300 -190
rect 10334 -224 10346 -190
rect 10288 -230 10346 -224
rect 10470 -230 10480 -170
rect 10540 -230 10550 -170
rect 10170 -271 10260 -270
rect 10170 -283 10292 -271
rect 10170 -343 10252 -283
rect 10286 -343 10292 -283
rect 10170 -355 10292 -343
rect 10328 -280 10388 -270
rect 10328 -343 10348 -340
rect 10382 -343 10388 -340
rect 10328 -350 10388 -343
rect 10436 -280 10496 -270
rect 10436 -343 10444 -340
rect 10478 -343 10496 -340
rect 10436 -350 10496 -343
rect 10534 -283 10580 -271
rect 10534 -343 10540 -283
rect 10574 -343 10580 -283
rect 10342 -355 10388 -350
rect 10438 -355 10484 -350
rect 10534 -355 10580 -343
rect 10630 -283 10676 -271
rect 10630 -343 10636 -283
rect 10670 -300 10676 -283
rect 10750 -300 10780 -130
rect 10670 -330 10780 -300
rect 10670 -343 10676 -330
rect 10630 -355 10676 -343
rect 10170 -360 10260 -355
rect 10170 -440 10176 -360
rect 10170 -540 10180 -440
rect 10370 -460 10380 -390
rect 10450 -460 10460 -390
rect 10576 -402 10634 -396
rect 10576 -436 10588 -402
rect 10622 -436 10634 -402
rect 10576 -442 10634 -436
rect 10124 -600 10180 -540
rect 10590 -580 10620 -442
rect 10058 -940 10180 -600
rect 10560 -640 10570 -580
rect 10630 -640 10640 -580
rect 10240 -670 10330 -660
rect 10240 -730 10260 -670
rect 10320 -730 10330 -670
rect 10730 -730 10740 -670
rect 10800 -730 10810 -670
rect 10240 -764 10330 -730
rect 10238 -770 10330 -764
rect 10238 -830 10250 -770
rect 10310 -830 10330 -770
rect 10580 -830 10590 -770
rect 10650 -830 10660 -770
rect 10238 -836 10330 -830
rect 10240 -840 10330 -836
rect 10390 -930 10400 -870
rect 10460 -930 10470 -870
rect 10600 -898 10630 -830
rect 10588 -904 10646 -898
rect 10396 -938 10408 -930
rect 10442 -938 10454 -930
rect 10058 -1669 10064 -940
rect 10396 -944 10454 -938
rect 10588 -938 10600 -904
rect 10634 -938 10646 -904
rect 10588 -944 10646 -938
rect 10339 -986 10400 -976
rect 10399 -1046 10400 -986
rect 10339 -1048 10360 -1046
rect 10394 -1048 10400 -1046
rect 10339 -1056 10400 -1048
rect 10447 -986 10507 -976
rect 10447 -1048 10456 -1046
rect 10490 -1048 10507 -1046
rect 10447 -1056 10507 -1048
rect 10546 -988 10592 -976
rect 10546 -1048 10552 -988
rect 10586 -1048 10592 -988
rect 10354 -1060 10400 -1056
rect 10450 -1060 10496 -1056
rect 10546 -1060 10592 -1048
rect 10642 -988 10688 -976
rect 10642 -1048 10648 -988
rect 10682 -1000 10688 -988
rect 10740 -1000 10780 -730
rect 10682 -1030 10780 -1000
rect 10682 -1048 10688 -1030
rect 10642 -1060 10688 -1048
rect 10490 -1098 10550 -1090
rect 10490 -1132 10504 -1098
rect 10538 -1132 10550 -1098
rect 10490 -1180 10550 -1132
rect 10480 -1240 10490 -1180
rect 10550 -1240 10560 -1180
rect 10490 -1302 10550 -1240
rect 10490 -1336 10504 -1302
rect 10538 -1336 10550 -1302
rect 10490 -1340 10550 -1336
rect 10492 -1342 10550 -1340
rect 10354 -1376 10400 -1374
rect 10450 -1376 10496 -1374
rect 10339 -1386 10400 -1376
rect 10399 -1446 10400 -1386
rect 10339 -1456 10400 -1446
rect 10447 -1386 10507 -1376
rect 10447 -1456 10507 -1446
rect 10546 -1386 10592 -1374
rect 10546 -1446 10552 -1386
rect 10586 -1446 10592 -1386
rect 10354 -1458 10400 -1456
rect 10450 -1458 10496 -1456
rect 10546 -1458 10592 -1446
rect 10642 -1386 10688 -1374
rect 10642 -1446 10648 -1386
rect 10682 -1400 10688 -1386
rect 10740 -1400 10780 -1030
rect 10840 -990 10870 70
rect 10940 -160 10970 1790
rect 11030 870 11060 1900
rect 11010 810 11020 870
rect 11080 810 11090 870
rect 11020 520 11080 530
rect 11020 450 11080 460
rect 11030 250 11060 450
rect 11010 190 11020 250
rect 11080 190 11090 250
rect 10900 -220 10910 -160
rect 10970 -220 10980 -160
rect 10900 -340 10910 -280
rect 10970 -340 10980 -280
rect 10840 -1050 10850 -990
rect 10910 -1050 10920 -990
rect 10950 -1380 10980 -340
rect 11030 -400 11060 190
rect 11010 -460 11020 -400
rect 11080 -460 11090 -400
rect 11120 -580 11150 2430
rect 11190 2340 11200 2400
rect 11260 2340 11270 2400
rect 11200 430 11230 2340
rect 11270 2087 11280 2147
rect 11340 2087 11350 2147
rect 11290 740 11320 2087
rect 11630 1720 11700 2810
rect 11620 1650 11630 1720
rect 11700 1650 11710 1720
rect 11450 1540 11460 1600
rect 11520 1540 11530 1600
rect 11360 1370 11420 1380
rect 11360 1300 11420 1310
rect 11270 680 11280 740
rect 11340 680 11350 740
rect 11180 370 11190 430
rect 11250 370 11260 430
rect 11080 -640 11090 -580
rect 11150 -640 11160 -580
rect 11010 -910 11020 -850
rect 11080 -910 11090 -850
rect 10682 -1430 10780 -1400
rect 10682 -1446 10688 -1430
rect 10920 -1440 10930 -1380
rect 10990 -1440 11000 -1380
rect 10642 -1458 10688 -1446
rect 11030 -1490 11060 -910
rect 10396 -1496 10454 -1490
rect 10396 -1500 10408 -1496
rect 10442 -1500 10454 -1496
rect 10588 -1496 10646 -1490
rect 10380 -1560 10390 -1500
rect 10450 -1560 10460 -1500
rect 10588 -1530 10600 -1496
rect 10634 -1530 10646 -1496
rect 10588 -1536 10646 -1530
rect 10600 -1630 10630 -1536
rect 11010 -1550 11020 -1490
rect 11080 -1550 11090 -1490
rect 11120 -1630 11150 -640
rect 11200 -760 11230 370
rect 11180 -820 11190 -760
rect 11250 -820 11260 -760
rect 11290 -1190 11320 680
rect 11380 40 11410 1300
rect 11470 520 11500 1540
rect 11540 1490 11600 1500
rect 11540 1420 11600 1430
rect 11440 460 11450 520
rect 11510 460 11520 520
rect 11550 140 11580 1420
rect 11630 630 11700 1650
rect 11620 560 11630 630
rect 11700 560 11710 630
rect 11530 130 11580 140
rect 11500 70 11510 130
rect 11570 70 11580 130
rect 11360 30 11420 40
rect 11360 -40 11420 -30
rect 11550 -860 11580 70
rect 11630 -670 11700 560
rect 11690 -730 11700 -670
rect 11630 -780 11700 -730
rect 11510 -920 11520 -860
rect 11580 -920 11590 -860
rect 11270 -1250 11280 -1190
rect 11340 -1250 11350 -1190
rect 10018 -1681 10064 -1669
rect 10570 -1690 10580 -1630
rect 10640 -1690 10650 -1630
rect 11070 -1690 11080 -1630
rect 11140 -1690 11150 -1630
rect 3700 -1830 3800 -1770
rect 3890 -1728 6890 -1720
rect 6950 -1728 10030 -1720
rect 3890 -1762 3912 -1728
rect 5880 -1762 5970 -1728
rect 7938 -1762 8028 -1728
rect 9996 -1762 10030 -1728
rect 3890 -1780 6890 -1762
rect 6950 -1780 10030 -1762
rect 3700 -1840 10140 -1830
rect 3700 -1890 3820 -1840
rect 10100 -1890 10140 -1840
rect 3700 -1900 10140 -1890
<< via1 >>
rect 6890 2732 6950 2750
rect 6890 2698 6950 2732
rect 6890 2690 6950 2698
rect 6890 604 6950 620
rect 6890 570 6950 604
rect 6890 560 6950 570
rect 6890 400 6950 420
rect 6890 366 6950 400
rect 6890 360 6950 366
rect 9740 70 9800 130
rect 9740 -520 9800 -460
rect 10520 2562 10580 2570
rect 10520 2512 10577 2562
rect 10577 2512 10580 2562
rect 10520 2510 10580 2512
rect 10680 2566 10750 2580
rect 10680 2512 10747 2566
rect 10747 2512 10750 2566
rect 10680 2510 10750 2512
rect 11010 2520 11070 2580
rect 10260 2410 10280 2470
rect 10280 2410 10320 2470
rect 10590 2350 10600 2400
rect 10600 2350 10650 2400
rect 10590 2340 10650 2350
rect 10280 2127 10340 2137
rect 10280 2077 10330 2127
rect 10330 2077 10340 2127
rect 11110 2430 11170 2490
rect 10510 1954 10570 1960
rect 10510 1904 10511 1954
rect 10511 1904 10570 1954
rect 10510 1900 10570 1904
rect 10680 1954 10750 1960
rect 10680 1900 10747 1954
rect 10747 1900 10750 1954
rect 10680 1890 10750 1900
rect 11010 1900 11070 1960
rect 10520 1838 10580 1850
rect 10520 1790 10580 1838
rect 10930 1790 10990 1850
rect 10760 1706 10830 1720
rect 10760 1672 10795 1706
rect 10795 1672 10829 1706
rect 10829 1672 10830 1706
rect 10760 1650 10830 1672
rect 10280 1520 10340 1580
rect 10620 1570 10629 1600
rect 10629 1570 10663 1600
rect 10663 1570 10680 1600
rect 10620 1540 10680 1570
rect 10500 1340 10563 1406
rect 10550 1230 10610 1290
rect 10800 1240 10860 1300
rect 10360 1009 10420 1020
rect 10360 961 10420 1009
rect 10630 1025 10700 1030
rect 10630 977 10634 1025
rect 10634 977 10699 1025
rect 10699 977 10700 1025
rect 10630 970 10700 977
rect 10360 960 10420 961
rect 10550 864 10610 870
rect 10550 816 10554 864
rect 10554 816 10610 864
rect 10550 810 10610 816
rect 10270 680 10330 740
rect 10690 618 10760 630
rect 10690 584 10703 618
rect 10703 584 10737 618
rect 10737 584 10760 618
rect 10690 560 10760 584
rect 10580 380 10640 440
rect 10380 226 10450 250
rect 10380 192 10396 226
rect 10396 192 10430 226
rect 10430 192 10450 226
rect 10380 180 10450 192
rect 10328 73 10348 132
rect 10348 73 10382 132
rect 10382 73 10388 132
rect 10328 72 10388 73
rect 10436 73 10444 132
rect 10444 73 10478 132
rect 10478 73 10496 132
rect 10436 72 10496 73
rect 10280 14 10340 20
rect 10280 -20 10300 14
rect 10300 -20 10334 14
rect 10334 -20 10340 14
rect 10280 -40 10340 -20
rect 10120 -130 10130 -70
rect 10130 -130 10170 -70
rect 10170 -130 10180 -70
rect 10830 70 10890 130
rect 10740 -130 10800 -70
rect 10480 -190 10540 -170
rect 10480 -224 10492 -190
rect 10492 -224 10526 -190
rect 10526 -224 10540 -190
rect 10480 -230 10540 -224
rect 10328 -283 10388 -280
rect 10328 -340 10348 -283
rect 10348 -340 10382 -283
rect 10382 -340 10388 -283
rect 10436 -283 10496 -280
rect 10436 -340 10444 -283
rect 10444 -340 10478 -283
rect 10478 -340 10496 -283
rect 10380 -402 10450 -390
rect 10380 -436 10396 -402
rect 10396 -436 10430 -402
rect 10430 -436 10450 -402
rect 10380 -460 10450 -436
rect 10570 -640 10630 -580
rect 10260 -730 10320 -670
rect 10740 -730 10800 -670
rect 10590 -830 10650 -770
rect 10400 -904 10460 -870
rect 10400 -930 10408 -904
rect 10408 -930 10442 -904
rect 10442 -930 10460 -904
rect 10339 -988 10399 -986
rect 10339 -1046 10360 -988
rect 10360 -1046 10394 -988
rect 10394 -1046 10399 -988
rect 10447 -988 10507 -986
rect 10447 -1046 10456 -988
rect 10456 -1046 10490 -988
rect 10490 -1046 10507 -988
rect 10490 -1240 10550 -1180
rect 10339 -1446 10360 -1386
rect 10360 -1446 10394 -1386
rect 10394 -1446 10399 -1386
rect 10447 -1446 10456 -1386
rect 10456 -1446 10490 -1386
rect 10490 -1446 10507 -1386
rect 11020 810 11080 870
rect 11020 460 11080 520
rect 11020 190 11080 250
rect 10910 -220 10970 -160
rect 10910 -340 10970 -280
rect 10850 -1050 10910 -990
rect 11020 -460 11080 -400
rect 11200 2340 11260 2400
rect 11280 2087 11340 2147
rect 11630 1650 11700 1720
rect 11460 1540 11520 1600
rect 11360 1310 11420 1370
rect 11280 680 11340 740
rect 11190 370 11250 430
rect 11090 -640 11150 -580
rect 11020 -910 11080 -850
rect 10930 -1440 10990 -1380
rect 10390 -1530 10408 -1500
rect 10408 -1530 10442 -1500
rect 10442 -1530 10450 -1500
rect 10390 -1560 10450 -1530
rect 11020 -1550 11080 -1490
rect 11190 -820 11250 -760
rect 11540 1430 11600 1490
rect 11450 460 11510 520
rect 11630 560 11700 630
rect 11510 70 11570 130
rect 11360 -30 11420 30
rect 11630 -730 11690 -670
rect 11520 -920 11580 -860
rect 11280 -1250 11340 -1190
rect 10580 -1690 10640 -1630
rect 11080 -1690 11140 -1630
rect 6890 -1728 6950 -1720
rect 6890 -1762 6950 -1728
rect 6890 -1780 6950 -1762
<< metal2 >>
rect 6890 2750 6950 2760
rect 6890 620 6950 2690
rect 10540 2625 11750 2655
rect 10540 2580 10570 2625
rect 10680 2580 10750 2590
rect 10520 2570 10580 2580
rect 10520 2500 10580 2510
rect 11010 2580 11070 2590
rect 10750 2530 11010 2560
rect 11070 2530 11750 2560
rect 11010 2510 11070 2520
rect 10680 2500 10750 2510
rect 11110 2490 11170 2500
rect 10260 2470 10320 2480
rect 10320 2440 11110 2470
rect 11110 2420 11170 2430
rect 10260 2400 10320 2410
rect 10590 2400 10650 2410
rect 11200 2400 11260 2410
rect 10650 2360 11200 2390
rect 10590 2330 10650 2340
rect 11200 2330 11260 2340
rect 11280 2147 11340 2157
rect 10280 2137 10340 2147
rect 10340 2087 11280 2117
rect 11280 2077 11340 2087
rect 10280 2067 10340 2077
rect 10530 2010 11750 2040
rect 10530 1970 10560 2010
rect 10510 1960 10570 1970
rect 10510 1890 10570 1900
rect 10680 1960 10750 1970
rect 11010 1960 11070 1970
rect 10750 1900 11010 1930
rect 11010 1890 11070 1900
rect 10680 1880 10750 1890
rect 10520 1850 10580 1860
rect 10930 1850 10990 1860
rect 10580 1810 10930 1840
rect 10520 1780 10580 1790
rect 10930 1780 10990 1790
rect 10760 1720 10830 1730
rect 11630 1720 11700 1730
rect 10830 1650 11630 1720
rect 10760 1640 10830 1650
rect 11630 1640 11700 1650
rect 10620 1600 10680 1610
rect 10280 1580 10340 1590
rect 11460 1600 11520 1610
rect 10680 1550 11460 1580
rect 10620 1530 10680 1540
rect 11460 1530 11520 1540
rect 10280 1510 10340 1520
rect 10290 1480 10320 1510
rect 11540 1490 11600 1500
rect 10290 1450 11540 1480
rect 11540 1420 11600 1430
rect 10500 1406 10563 1416
rect 10563 1370 10580 1380
rect 11360 1370 11420 1380
rect 10563 1340 11360 1370
rect 10500 1330 10563 1340
rect 10800 1300 10860 1310
rect 11360 1300 11420 1310
rect 10550 1290 10610 1300
rect 10800 1230 10860 1240
rect 10550 1220 10610 1230
rect 10360 1020 10420 1030
rect 10560 1020 10590 1220
rect 10420 980 10590 1020
rect 10630 1030 10700 1040
rect 10810 1020 10850 1230
rect 10700 980 10850 1020
rect 10630 960 10700 970
rect 10360 950 10420 960
rect 10550 870 10610 880
rect 11020 870 11080 880
rect 10610 820 11020 850
rect 10550 800 10610 810
rect 11020 800 11080 810
rect 10270 740 10330 750
rect 11280 740 11340 750
rect 10330 680 11280 720
rect 10270 670 10330 680
rect 11280 670 11340 680
rect 3610 560 6890 600
rect 10690 630 10760 640
rect 11630 630 11700 640
rect 6950 560 7610 600
rect 6890 550 6950 560
rect 6890 420 6950 430
rect 6890 -290 6950 360
rect 7570 120 7610 560
rect 10760 560 11630 630
rect 10690 550 10760 560
rect 11630 550 11700 560
rect 11020 520 11080 530
rect 11450 520 11510 530
rect 11080 470 11450 500
rect 11020 450 11080 460
rect 11450 450 11510 460
rect 10580 440 10640 450
rect 11190 430 11250 440
rect 10640 390 11190 420
rect 10580 370 10640 380
rect 11190 360 11250 370
rect 10380 250 10450 260
rect 11020 250 11080 260
rect 10450 200 11020 240
rect 11020 180 11080 190
rect 10380 170 10450 180
rect 9740 130 9800 140
rect 7570 80 9740 120
rect 10328 132 10388 142
rect 9800 80 10328 120
rect 9740 60 9800 70
rect 10328 62 10388 72
rect 10436 132 10496 142
rect 10830 130 10890 140
rect 10496 80 10830 120
rect 10436 62 10496 72
rect 10830 60 10890 70
rect 11510 130 11570 140
rect 11510 60 11570 70
rect 11360 30 11420 40
rect 10280 20 10340 30
rect 10340 -20 11360 10
rect 11420 -20 11750 10
rect 11360 -40 11420 -30
rect 10280 -50 10340 -40
rect 10120 -70 10180 -60
rect 10740 -70 10800 -60
rect 10180 -120 10740 -80
rect 10120 -140 10180 -130
rect 10740 -140 10800 -130
rect 10910 -160 10970 -150
rect 10480 -170 10540 -160
rect 10540 -210 10910 -180
rect 10910 -230 10970 -220
rect 10480 -240 10540 -230
rect 10328 -280 10388 -270
rect 3610 -330 10328 -290
rect 6890 -1720 6950 -330
rect 9600 -1400 9640 -330
rect 10328 -350 10388 -340
rect 10436 -280 10496 -270
rect 10910 -280 10970 -270
rect 10496 -330 10910 -300
rect 10436 -350 10496 -340
rect 10910 -350 10970 -340
rect 10380 -390 10450 -380
rect 9740 -460 9800 -450
rect 11020 -400 11080 -390
rect 10450 -450 11020 -410
rect 10380 -470 10450 -460
rect 11020 -470 11080 -460
rect 9740 -530 9800 -520
rect 9750 -1000 9790 -530
rect 10570 -580 10630 -570
rect 11090 -580 11150 -570
rect 10630 -630 11090 -600
rect 10570 -650 10630 -640
rect 11090 -650 11150 -640
rect 10260 -670 10320 -660
rect 10740 -670 10800 -660
rect 10320 -720 10740 -680
rect 10260 -740 10320 -730
rect 11630 -670 11690 -660
rect 10800 -720 11630 -680
rect 10740 -740 10800 -730
rect 11630 -740 11690 -730
rect 11190 -760 11250 -750
rect 10590 -770 10650 -760
rect 10650 -810 11190 -780
rect 11190 -830 11250 -820
rect 10590 -840 10650 -830
rect 11020 -850 11080 -840
rect 10400 -870 10460 -860
rect 10460 -900 11020 -870
rect 11520 -860 11580 -850
rect 11080 -900 11520 -870
rect 11020 -920 11080 -910
rect 11520 -930 11580 -920
rect 10400 -940 10460 -930
rect 10339 -986 10399 -976
rect 9750 -1040 10339 -1000
rect 10339 -1056 10399 -1046
rect 10447 -986 10507 -976
rect 10850 -990 10910 -980
rect 10507 -1030 10850 -1000
rect 10447 -1056 10507 -1046
rect 10850 -1060 10910 -1050
rect 10490 -1180 10550 -1170
rect 11280 -1190 11340 -1180
rect 10550 -1230 11280 -1200
rect 10490 -1250 10550 -1240
rect 11280 -1260 11340 -1250
rect 10339 -1386 10399 -1376
rect 9600 -1440 10339 -1400
rect 10339 -1456 10399 -1446
rect 10447 -1386 10507 -1376
rect 10930 -1380 10990 -1370
rect 10507 -1430 10930 -1390
rect 10447 -1456 10507 -1446
rect 10930 -1450 10990 -1440
rect 11020 -1490 11080 -1480
rect 10390 -1500 10450 -1490
rect 10450 -1550 11020 -1530
rect 10450 -1560 11080 -1550
rect 10390 -1570 10450 -1560
rect 10580 -1630 10640 -1620
rect 11080 -1630 11140 -1620
rect 10640 -1670 11080 -1640
rect 10580 -1700 10640 -1690
rect 11080 -1700 11140 -1690
rect 6890 -1790 6950 -1780
<< labels >>
flabel metal1 11030 305 11060 335 0 FreeSans 80 0 0 0 LOAD_CAL_Z
flabel metal1 10940 300 10970 330 0 FreeSans 80 0 0 0 EN_COMP_Z
flabel metal1 11120 310 11150 340 0 FreeSans 80 0 0 0 CAL_RESULTi
flabel metal1 11200 480 11230 510 0 FreeSans 80 0 0 0 CAL_RESULT_Z
flabel metal1 11290 460 11320 490 0 FreeSans 80 0 0 0 EN_COMPi
rlabel metal2 3610 -330 3650 -290 1 CAL_P
port 3 n
rlabel metal2 3610 560 3650 600 1 CAL_N
port 4 n
rlabel metal1 9980 2820 10140 2880 1 VDD
port 0 n
rlabel metal1 10280 2820 10440 2880 1 VSS
port 6 n
rlabel metal2 11720 2530 11750 2560 1 CAL_CYCLE
port 7 n
rlabel metal2 11720 2625 11750 2655 1 CAL_RESULT
port 1 n
rlabel metal2 11715 2010 11745 2040 1 EN_COMP
port 2 n
rlabel metal2 11715 -20 11745 10 1 EN
port 5 n
<< end >>
