magic
tech sky130A
magscale 1 2
timestamp 1711882560
<< error_p >>
rect -176 5707 -118 5713
rect 20 5707 78 5713
rect -176 5673 -164 5707
rect 20 5673 32 5707
rect -176 5667 -118 5673
rect 20 5667 78 5673
rect -78 4379 -20 4385
rect 118 4379 176 4385
rect -78 4345 -66 4379
rect 118 4345 130 4379
rect -78 4339 -20 4345
rect 118 4339 176 4345
rect -78 4271 -20 4277
rect 118 4271 176 4277
rect -78 4237 -66 4271
rect 118 4237 130 4271
rect -78 4231 -20 4237
rect 118 4231 176 4237
rect -176 2943 -118 2949
rect 20 2943 78 2949
rect -176 2909 -164 2943
rect 20 2909 32 2943
rect -176 2903 -118 2909
rect 20 2903 78 2909
rect -176 2835 -118 2841
rect 20 2835 78 2841
rect -176 2801 -164 2835
rect 20 2801 32 2835
rect -176 2795 -118 2801
rect 20 2795 78 2801
rect -78 1507 -20 1513
rect 118 1507 176 1513
rect -78 1473 -66 1507
rect 118 1473 130 1507
rect -78 1467 -20 1473
rect 118 1467 176 1473
rect -78 1399 -20 1405
rect 118 1399 176 1405
rect -78 1365 -66 1399
rect 118 1365 130 1399
rect -78 1359 -20 1365
rect 118 1359 176 1365
rect -176 71 -118 77
rect 20 71 78 77
rect -176 37 -164 71
rect 20 37 32 71
rect -176 31 -118 37
rect 20 31 78 37
rect -176 -37 -118 -31
rect 20 -37 78 -31
rect -176 -71 -164 -37
rect 20 -71 32 -37
rect -176 -77 -118 -71
rect 20 -77 78 -71
rect -78 -1365 -20 -1359
rect 118 -1365 176 -1359
rect -78 -1399 -66 -1365
rect 118 -1399 130 -1365
rect -78 -1405 -20 -1399
rect 118 -1405 176 -1399
rect -78 -1473 -20 -1467
rect 118 -1473 176 -1467
rect -78 -1507 -66 -1473
rect 118 -1507 130 -1473
rect -78 -1513 -20 -1507
rect 118 -1513 176 -1507
rect -176 -2801 -118 -2795
rect 20 -2801 78 -2795
rect -176 -2835 -164 -2801
rect 20 -2835 32 -2801
rect -176 -2841 -118 -2835
rect 20 -2841 78 -2835
rect -176 -2909 -118 -2903
rect 20 -2909 78 -2903
rect -176 -2943 -164 -2909
rect 20 -2943 32 -2909
rect -176 -2949 -118 -2943
rect 20 -2949 78 -2943
rect -78 -4237 -20 -4231
rect 118 -4237 176 -4231
rect -78 -4271 -66 -4237
rect 118 -4271 130 -4237
rect -78 -4277 -20 -4271
rect 118 -4277 176 -4271
rect -78 -4345 -20 -4339
rect 118 -4345 176 -4339
rect -78 -4379 -66 -4345
rect 118 -4379 130 -4345
rect -78 -4385 -20 -4379
rect 118 -4385 176 -4379
rect -176 -5673 -118 -5667
rect 20 -5673 78 -5667
rect -176 -5707 -164 -5673
rect 20 -5707 32 -5673
rect -176 -5713 -118 -5707
rect 20 -5713 78 -5707
<< nwell >>
rect -363 -5845 363 5845
<< pmos >>
rect -167 4426 -127 5626
rect -69 4426 -29 5626
rect 29 4426 69 5626
rect 127 4426 167 5626
rect -167 2990 -127 4190
rect -69 2990 -29 4190
rect 29 2990 69 4190
rect 127 2990 167 4190
rect -167 1554 -127 2754
rect -69 1554 -29 2754
rect 29 1554 69 2754
rect 127 1554 167 2754
rect -167 118 -127 1318
rect -69 118 -29 1318
rect 29 118 69 1318
rect 127 118 167 1318
rect -167 -1318 -127 -118
rect -69 -1318 -29 -118
rect 29 -1318 69 -118
rect 127 -1318 167 -118
rect -167 -2754 -127 -1554
rect -69 -2754 -29 -1554
rect 29 -2754 69 -1554
rect 127 -2754 167 -1554
rect -167 -4190 -127 -2990
rect -69 -4190 -29 -2990
rect 29 -4190 69 -2990
rect 127 -4190 167 -2990
rect -167 -5626 -127 -4426
rect -69 -5626 -29 -4426
rect 29 -5626 69 -4426
rect 127 -5626 167 -4426
<< pdiff >>
rect -225 5614 -167 5626
rect -225 4438 -213 5614
rect -179 4438 -167 5614
rect -225 4426 -167 4438
rect -127 5614 -69 5626
rect -127 4438 -115 5614
rect -81 4438 -69 5614
rect -127 4426 -69 4438
rect -29 5614 29 5626
rect -29 4438 -17 5614
rect 17 4438 29 5614
rect -29 4426 29 4438
rect 69 5614 127 5626
rect 69 4438 81 5614
rect 115 4438 127 5614
rect 69 4426 127 4438
rect 167 5614 225 5626
rect 167 4438 179 5614
rect 213 4438 225 5614
rect 167 4426 225 4438
rect -225 4178 -167 4190
rect -225 3002 -213 4178
rect -179 3002 -167 4178
rect -225 2990 -167 3002
rect -127 4178 -69 4190
rect -127 3002 -115 4178
rect -81 3002 -69 4178
rect -127 2990 -69 3002
rect -29 4178 29 4190
rect -29 3002 -17 4178
rect 17 3002 29 4178
rect -29 2990 29 3002
rect 69 4178 127 4190
rect 69 3002 81 4178
rect 115 3002 127 4178
rect 69 2990 127 3002
rect 167 4178 225 4190
rect 167 3002 179 4178
rect 213 3002 225 4178
rect 167 2990 225 3002
rect -225 2742 -167 2754
rect -225 1566 -213 2742
rect -179 1566 -167 2742
rect -225 1554 -167 1566
rect -127 2742 -69 2754
rect -127 1566 -115 2742
rect -81 1566 -69 2742
rect -127 1554 -69 1566
rect -29 2742 29 2754
rect -29 1566 -17 2742
rect 17 1566 29 2742
rect -29 1554 29 1566
rect 69 2742 127 2754
rect 69 1566 81 2742
rect 115 1566 127 2742
rect 69 1554 127 1566
rect 167 2742 225 2754
rect 167 1566 179 2742
rect 213 1566 225 2742
rect 167 1554 225 1566
rect -225 1306 -167 1318
rect -225 130 -213 1306
rect -179 130 -167 1306
rect -225 118 -167 130
rect -127 1306 -69 1318
rect -127 130 -115 1306
rect -81 130 -69 1306
rect -127 118 -69 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 69 1306 127 1318
rect 69 130 81 1306
rect 115 130 127 1306
rect 69 118 127 130
rect 167 1306 225 1318
rect 167 130 179 1306
rect 213 130 225 1306
rect 167 118 225 130
rect -225 -130 -167 -118
rect -225 -1306 -213 -130
rect -179 -1306 -167 -130
rect -225 -1318 -167 -1306
rect -127 -130 -69 -118
rect -127 -1306 -115 -130
rect -81 -1306 -69 -130
rect -127 -1318 -69 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 69 -130 127 -118
rect 69 -1306 81 -130
rect 115 -1306 127 -130
rect 69 -1318 127 -1306
rect 167 -130 225 -118
rect 167 -1306 179 -130
rect 213 -1306 225 -130
rect 167 -1318 225 -1306
rect -225 -1566 -167 -1554
rect -225 -2742 -213 -1566
rect -179 -2742 -167 -1566
rect -225 -2754 -167 -2742
rect -127 -1566 -69 -1554
rect -127 -2742 -115 -1566
rect -81 -2742 -69 -1566
rect -127 -2754 -69 -2742
rect -29 -1566 29 -1554
rect -29 -2742 -17 -1566
rect 17 -2742 29 -1566
rect -29 -2754 29 -2742
rect 69 -1566 127 -1554
rect 69 -2742 81 -1566
rect 115 -2742 127 -1566
rect 69 -2754 127 -2742
rect 167 -1566 225 -1554
rect 167 -2742 179 -1566
rect 213 -2742 225 -1566
rect 167 -2754 225 -2742
rect -225 -3002 -167 -2990
rect -225 -4178 -213 -3002
rect -179 -4178 -167 -3002
rect -225 -4190 -167 -4178
rect -127 -3002 -69 -2990
rect -127 -4178 -115 -3002
rect -81 -4178 -69 -3002
rect -127 -4190 -69 -4178
rect -29 -3002 29 -2990
rect -29 -4178 -17 -3002
rect 17 -4178 29 -3002
rect -29 -4190 29 -4178
rect 69 -3002 127 -2990
rect 69 -4178 81 -3002
rect 115 -4178 127 -3002
rect 69 -4190 127 -4178
rect 167 -3002 225 -2990
rect 167 -4178 179 -3002
rect 213 -4178 225 -3002
rect 167 -4190 225 -4178
rect -225 -4438 -167 -4426
rect -225 -5614 -213 -4438
rect -179 -5614 -167 -4438
rect -225 -5626 -167 -5614
rect -127 -4438 -69 -4426
rect -127 -5614 -115 -4438
rect -81 -5614 -69 -4438
rect -127 -5626 -69 -5614
rect -29 -4438 29 -4426
rect -29 -5614 -17 -4438
rect 17 -5614 29 -4438
rect -29 -5626 29 -5614
rect 69 -4438 127 -4426
rect 69 -5614 81 -4438
rect 115 -5614 127 -4438
rect 69 -5626 127 -5614
rect 167 -4438 225 -4426
rect 167 -5614 179 -4438
rect 213 -5614 225 -4438
rect 167 -5626 225 -5614
<< pdiffc >>
rect -213 4438 -179 5614
rect -115 4438 -81 5614
rect -17 4438 17 5614
rect 81 4438 115 5614
rect 179 4438 213 5614
rect -213 3002 -179 4178
rect -115 3002 -81 4178
rect -17 3002 17 4178
rect 81 3002 115 4178
rect 179 3002 213 4178
rect -213 1566 -179 2742
rect -115 1566 -81 2742
rect -17 1566 17 2742
rect 81 1566 115 2742
rect 179 1566 213 2742
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect -213 -2742 -179 -1566
rect -115 -2742 -81 -1566
rect -17 -2742 17 -1566
rect 81 -2742 115 -1566
rect 179 -2742 213 -1566
rect -213 -4178 -179 -3002
rect -115 -4178 -81 -3002
rect -17 -4178 17 -3002
rect 81 -4178 115 -3002
rect 179 -4178 213 -3002
rect -213 -5614 -179 -4438
rect -115 -5614 -81 -4438
rect -17 -5614 17 -4438
rect 81 -5614 115 -4438
rect 179 -5614 213 -4438
<< nsubdiff >>
rect -327 5775 -231 5809
rect 231 5775 327 5809
rect -327 5713 -293 5775
rect 293 5713 327 5775
rect -327 -5775 -293 -5713
rect 293 -5775 327 -5713
rect -327 -5809 -231 -5775
rect 231 -5809 327 -5775
<< nsubdiffcont >>
rect -231 5775 231 5809
rect -327 -5713 -293 5713
rect 293 -5713 327 5713
rect -231 -5809 231 -5775
<< poly >>
rect -180 5707 -114 5723
rect -180 5673 -164 5707
rect -130 5673 -114 5707
rect -180 5657 -114 5673
rect 16 5707 82 5723
rect 16 5673 32 5707
rect 66 5673 82 5707
rect 16 5657 82 5673
rect -167 5626 -127 5657
rect -69 5626 -29 5652
rect 29 5626 69 5657
rect 127 5626 167 5652
rect -167 4400 -127 4426
rect -69 4395 -29 4426
rect 29 4400 69 4426
rect 127 4395 167 4426
rect -82 4379 -16 4395
rect -82 4345 -66 4379
rect -32 4345 -16 4379
rect -82 4329 -16 4345
rect 114 4379 180 4395
rect 114 4345 130 4379
rect 164 4345 180 4379
rect 114 4329 180 4345
rect -82 4271 -16 4287
rect -82 4237 -66 4271
rect -32 4237 -16 4271
rect -82 4221 -16 4237
rect 114 4271 180 4287
rect 114 4237 130 4271
rect 164 4237 180 4271
rect 114 4221 180 4237
rect -167 4190 -127 4216
rect -69 4190 -29 4221
rect 29 4190 69 4216
rect 127 4190 167 4221
rect -167 2959 -127 2990
rect -69 2964 -29 2990
rect 29 2959 69 2990
rect 127 2964 167 2990
rect -180 2943 -114 2959
rect -180 2909 -164 2943
rect -130 2909 -114 2943
rect -180 2893 -114 2909
rect 16 2943 82 2959
rect 16 2909 32 2943
rect 66 2909 82 2943
rect 16 2893 82 2909
rect -180 2835 -114 2851
rect -180 2801 -164 2835
rect -130 2801 -114 2835
rect -180 2785 -114 2801
rect 16 2835 82 2851
rect 16 2801 32 2835
rect 66 2801 82 2835
rect 16 2785 82 2801
rect -167 2754 -127 2785
rect -69 2754 -29 2780
rect 29 2754 69 2785
rect 127 2754 167 2780
rect -167 1528 -127 1554
rect -69 1523 -29 1554
rect 29 1528 69 1554
rect 127 1523 167 1554
rect -82 1507 -16 1523
rect -82 1473 -66 1507
rect -32 1473 -16 1507
rect -82 1457 -16 1473
rect 114 1507 180 1523
rect 114 1473 130 1507
rect 164 1473 180 1507
rect 114 1457 180 1473
rect -82 1399 -16 1415
rect -82 1365 -66 1399
rect -32 1365 -16 1399
rect -82 1349 -16 1365
rect 114 1399 180 1415
rect 114 1365 130 1399
rect 164 1365 180 1399
rect 114 1349 180 1365
rect -167 1318 -127 1344
rect -69 1318 -29 1349
rect 29 1318 69 1344
rect 127 1318 167 1349
rect -167 87 -127 118
rect -69 92 -29 118
rect 29 87 69 118
rect 127 92 167 118
rect -180 71 -114 87
rect -180 37 -164 71
rect -130 37 -114 71
rect -180 21 -114 37
rect 16 71 82 87
rect 16 37 32 71
rect 66 37 82 71
rect 16 21 82 37
rect -180 -37 -114 -21
rect -180 -71 -164 -37
rect -130 -71 -114 -37
rect -180 -87 -114 -71
rect 16 -37 82 -21
rect 16 -71 32 -37
rect 66 -71 82 -37
rect 16 -87 82 -71
rect -167 -118 -127 -87
rect -69 -118 -29 -92
rect 29 -118 69 -87
rect 127 -118 167 -92
rect -167 -1344 -127 -1318
rect -69 -1349 -29 -1318
rect 29 -1344 69 -1318
rect 127 -1349 167 -1318
rect -82 -1365 -16 -1349
rect -82 -1399 -66 -1365
rect -32 -1399 -16 -1365
rect -82 -1415 -16 -1399
rect 114 -1365 180 -1349
rect 114 -1399 130 -1365
rect 164 -1399 180 -1365
rect 114 -1415 180 -1399
rect -82 -1473 -16 -1457
rect -82 -1507 -66 -1473
rect -32 -1507 -16 -1473
rect -82 -1523 -16 -1507
rect 114 -1473 180 -1457
rect 114 -1507 130 -1473
rect 164 -1507 180 -1473
rect 114 -1523 180 -1507
rect -167 -1554 -127 -1528
rect -69 -1554 -29 -1523
rect 29 -1554 69 -1528
rect 127 -1554 167 -1523
rect -167 -2785 -127 -2754
rect -69 -2780 -29 -2754
rect 29 -2785 69 -2754
rect 127 -2780 167 -2754
rect -180 -2801 -114 -2785
rect -180 -2835 -164 -2801
rect -130 -2835 -114 -2801
rect -180 -2851 -114 -2835
rect 16 -2801 82 -2785
rect 16 -2835 32 -2801
rect 66 -2835 82 -2801
rect 16 -2851 82 -2835
rect -180 -2909 -114 -2893
rect -180 -2943 -164 -2909
rect -130 -2943 -114 -2909
rect -180 -2959 -114 -2943
rect 16 -2909 82 -2893
rect 16 -2943 32 -2909
rect 66 -2943 82 -2909
rect 16 -2959 82 -2943
rect -167 -2990 -127 -2959
rect -69 -2990 -29 -2964
rect 29 -2990 69 -2959
rect 127 -2990 167 -2964
rect -167 -4216 -127 -4190
rect -69 -4221 -29 -4190
rect 29 -4216 69 -4190
rect 127 -4221 167 -4190
rect -82 -4237 -16 -4221
rect -82 -4271 -66 -4237
rect -32 -4271 -16 -4237
rect -82 -4287 -16 -4271
rect 114 -4237 180 -4221
rect 114 -4271 130 -4237
rect 164 -4271 180 -4237
rect 114 -4287 180 -4271
rect -82 -4345 -16 -4329
rect -82 -4379 -66 -4345
rect -32 -4379 -16 -4345
rect -82 -4395 -16 -4379
rect 114 -4345 180 -4329
rect 114 -4379 130 -4345
rect 164 -4379 180 -4345
rect 114 -4395 180 -4379
rect -167 -4426 -127 -4400
rect -69 -4426 -29 -4395
rect 29 -4426 69 -4400
rect 127 -4426 167 -4395
rect -167 -5657 -127 -5626
rect -69 -5652 -29 -5626
rect 29 -5657 69 -5626
rect 127 -5652 167 -5626
rect -180 -5673 -114 -5657
rect -180 -5707 -164 -5673
rect -130 -5707 -114 -5673
rect -180 -5723 -114 -5707
rect 16 -5673 82 -5657
rect 16 -5707 32 -5673
rect 66 -5707 82 -5673
rect 16 -5723 82 -5707
<< polycont >>
rect -164 5673 -130 5707
rect 32 5673 66 5707
rect -66 4345 -32 4379
rect 130 4345 164 4379
rect -66 4237 -32 4271
rect 130 4237 164 4271
rect -164 2909 -130 2943
rect 32 2909 66 2943
rect -164 2801 -130 2835
rect 32 2801 66 2835
rect -66 1473 -32 1507
rect 130 1473 164 1507
rect -66 1365 -32 1399
rect 130 1365 164 1399
rect -164 37 -130 71
rect 32 37 66 71
rect -164 -71 -130 -37
rect 32 -71 66 -37
rect -66 -1399 -32 -1365
rect 130 -1399 164 -1365
rect -66 -1507 -32 -1473
rect 130 -1507 164 -1473
rect -164 -2835 -130 -2801
rect 32 -2835 66 -2801
rect -164 -2943 -130 -2909
rect 32 -2943 66 -2909
rect -66 -4271 -32 -4237
rect 130 -4271 164 -4237
rect -66 -4379 -32 -4345
rect 130 -4379 164 -4345
rect -164 -5707 -130 -5673
rect 32 -5707 66 -5673
<< locali >>
rect -327 5775 -231 5809
rect 231 5775 327 5809
rect -327 5713 -293 5775
rect 293 5713 327 5775
rect -180 5673 -164 5707
rect -130 5673 -114 5707
rect 16 5673 32 5707
rect 66 5673 82 5707
rect -213 5614 -179 5630
rect -213 4422 -179 4438
rect -115 5614 -81 5630
rect -115 4422 -81 4438
rect -17 5614 17 5630
rect -17 4422 17 4438
rect 81 5614 115 5630
rect 81 4422 115 4438
rect 179 5614 213 5630
rect 179 4422 213 4438
rect -82 4345 -66 4379
rect -32 4345 -16 4379
rect 114 4345 130 4379
rect 164 4345 180 4379
rect -82 4237 -66 4271
rect -32 4237 -16 4271
rect 114 4237 130 4271
rect 164 4237 180 4271
rect -213 4178 -179 4194
rect -213 2986 -179 3002
rect -115 4178 -81 4194
rect -115 2986 -81 3002
rect -17 4178 17 4194
rect -17 2986 17 3002
rect 81 4178 115 4194
rect 81 2986 115 3002
rect 179 4178 213 4194
rect 179 2986 213 3002
rect -180 2909 -164 2943
rect -130 2909 -114 2943
rect 16 2909 32 2943
rect 66 2909 82 2943
rect -180 2801 -164 2835
rect -130 2801 -114 2835
rect 16 2801 32 2835
rect 66 2801 82 2835
rect -213 2742 -179 2758
rect -213 1550 -179 1566
rect -115 2742 -81 2758
rect -115 1550 -81 1566
rect -17 2742 17 2758
rect -17 1550 17 1566
rect 81 2742 115 2758
rect 81 1550 115 1566
rect 179 2742 213 2758
rect 179 1550 213 1566
rect -82 1473 -66 1507
rect -32 1473 -16 1507
rect 114 1473 130 1507
rect 164 1473 180 1507
rect -82 1365 -66 1399
rect -32 1365 -16 1399
rect 114 1365 130 1399
rect 164 1365 180 1399
rect -213 1306 -179 1322
rect -213 114 -179 130
rect -115 1306 -81 1322
rect -115 114 -81 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 81 1306 115 1322
rect 81 114 115 130
rect 179 1306 213 1322
rect 179 114 213 130
rect -180 37 -164 71
rect -130 37 -114 71
rect 16 37 32 71
rect 66 37 82 71
rect -180 -71 -164 -37
rect -130 -71 -114 -37
rect 16 -71 32 -37
rect 66 -71 82 -37
rect -213 -130 -179 -114
rect -213 -1322 -179 -1306
rect -115 -130 -81 -114
rect -115 -1322 -81 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 81 -130 115 -114
rect 81 -1322 115 -1306
rect 179 -130 213 -114
rect 179 -1322 213 -1306
rect -82 -1399 -66 -1365
rect -32 -1399 -16 -1365
rect 114 -1399 130 -1365
rect 164 -1399 180 -1365
rect -82 -1507 -66 -1473
rect -32 -1507 -16 -1473
rect 114 -1507 130 -1473
rect 164 -1507 180 -1473
rect -213 -1566 -179 -1550
rect -213 -2758 -179 -2742
rect -115 -1566 -81 -1550
rect -115 -2758 -81 -2742
rect -17 -1566 17 -1550
rect -17 -2758 17 -2742
rect 81 -1566 115 -1550
rect 81 -2758 115 -2742
rect 179 -1566 213 -1550
rect 179 -2758 213 -2742
rect -180 -2835 -164 -2801
rect -130 -2835 -114 -2801
rect 16 -2835 32 -2801
rect 66 -2835 82 -2801
rect -180 -2943 -164 -2909
rect -130 -2943 -114 -2909
rect 16 -2943 32 -2909
rect 66 -2943 82 -2909
rect -213 -3002 -179 -2986
rect -213 -4194 -179 -4178
rect -115 -3002 -81 -2986
rect -115 -4194 -81 -4178
rect -17 -3002 17 -2986
rect -17 -4194 17 -4178
rect 81 -3002 115 -2986
rect 81 -4194 115 -4178
rect 179 -3002 213 -2986
rect 179 -4194 213 -4178
rect -82 -4271 -66 -4237
rect -32 -4271 -16 -4237
rect 114 -4271 130 -4237
rect 164 -4271 180 -4237
rect -82 -4379 -66 -4345
rect -32 -4379 -16 -4345
rect 114 -4379 130 -4345
rect 164 -4379 180 -4345
rect -213 -4438 -179 -4422
rect -213 -5630 -179 -5614
rect -115 -4438 -81 -4422
rect -115 -5630 -81 -5614
rect -17 -4438 17 -4422
rect -17 -5630 17 -5614
rect 81 -4438 115 -4422
rect 81 -5630 115 -5614
rect 179 -4438 213 -4422
rect 179 -5630 213 -5614
rect -180 -5707 -164 -5673
rect -130 -5707 -114 -5673
rect 16 -5707 32 -5673
rect 66 -5707 82 -5673
rect -327 -5775 -293 -5713
rect 293 -5775 327 -5713
rect -327 -5809 -231 -5775
rect 231 -5809 327 -5775
<< viali >>
rect -164 5673 -130 5707
rect 32 5673 66 5707
rect -213 4438 -179 5614
rect -115 4438 -81 5614
rect -17 4438 17 5614
rect 81 4438 115 5614
rect 179 4438 213 5614
rect -66 4345 -32 4379
rect 130 4345 164 4379
rect -66 4237 -32 4271
rect 130 4237 164 4271
rect -213 3002 -179 4178
rect -115 3002 -81 4178
rect -17 3002 17 4178
rect 81 3002 115 4178
rect 179 3002 213 4178
rect -164 2909 -130 2943
rect 32 2909 66 2943
rect -164 2801 -130 2835
rect 32 2801 66 2835
rect -213 1566 -179 2742
rect -115 1566 -81 2742
rect -17 1566 17 2742
rect 81 1566 115 2742
rect 179 1566 213 2742
rect -66 1473 -32 1507
rect 130 1473 164 1507
rect -66 1365 -32 1399
rect 130 1365 164 1399
rect -213 130 -179 1306
rect -115 130 -81 1306
rect -17 130 17 1306
rect 81 130 115 1306
rect 179 130 213 1306
rect -164 37 -130 71
rect 32 37 66 71
rect -164 -71 -130 -37
rect 32 -71 66 -37
rect -213 -1306 -179 -130
rect -115 -1306 -81 -130
rect -17 -1306 17 -130
rect 81 -1306 115 -130
rect 179 -1306 213 -130
rect -66 -1399 -32 -1365
rect 130 -1399 164 -1365
rect -66 -1507 -32 -1473
rect 130 -1507 164 -1473
rect -213 -2742 -179 -1566
rect -115 -2742 -81 -1566
rect -17 -2742 17 -1566
rect 81 -2742 115 -1566
rect 179 -2742 213 -1566
rect -164 -2835 -130 -2801
rect 32 -2835 66 -2801
rect -164 -2943 -130 -2909
rect 32 -2943 66 -2909
rect -213 -4178 -179 -3002
rect -115 -4178 -81 -3002
rect -17 -4178 17 -3002
rect 81 -4178 115 -3002
rect 179 -4178 213 -3002
rect -66 -4271 -32 -4237
rect 130 -4271 164 -4237
rect -66 -4379 -32 -4345
rect 130 -4379 164 -4345
rect -213 -5614 -179 -4438
rect -115 -5614 -81 -4438
rect -17 -5614 17 -4438
rect 81 -5614 115 -4438
rect 179 -5614 213 -4438
rect -164 -5707 -130 -5673
rect 32 -5707 66 -5673
<< metal1 >>
rect -176 5707 -118 5713
rect -176 5673 -164 5707
rect -130 5673 -118 5707
rect -176 5667 -118 5673
rect 20 5707 78 5713
rect 20 5673 32 5707
rect 66 5673 78 5707
rect 20 5667 78 5673
rect -219 5614 -173 5626
rect -219 4438 -213 5614
rect -179 4438 -173 5614
rect -219 4426 -173 4438
rect -121 5614 -75 5626
rect -121 4438 -115 5614
rect -81 4438 -75 5614
rect -121 4426 -75 4438
rect -23 5614 23 5626
rect -23 4438 -17 5614
rect 17 4438 23 5614
rect -23 4426 23 4438
rect 75 5614 121 5626
rect 75 4438 81 5614
rect 115 4438 121 5614
rect 75 4426 121 4438
rect 173 5614 219 5626
rect 173 4438 179 5614
rect 213 4438 219 5614
rect 173 4426 219 4438
rect -78 4379 -20 4385
rect -78 4345 -66 4379
rect -32 4345 -20 4379
rect -78 4339 -20 4345
rect 118 4379 176 4385
rect 118 4345 130 4379
rect 164 4345 176 4379
rect 118 4339 176 4345
rect -78 4271 -20 4277
rect -78 4237 -66 4271
rect -32 4237 -20 4271
rect -78 4231 -20 4237
rect 118 4271 176 4277
rect 118 4237 130 4271
rect 164 4237 176 4271
rect 118 4231 176 4237
rect -219 4178 -173 4190
rect -219 3002 -213 4178
rect -179 3002 -173 4178
rect -219 2990 -173 3002
rect -121 4178 -75 4190
rect -121 3002 -115 4178
rect -81 3002 -75 4178
rect -121 2990 -75 3002
rect -23 4178 23 4190
rect -23 3002 -17 4178
rect 17 3002 23 4178
rect -23 2990 23 3002
rect 75 4178 121 4190
rect 75 3002 81 4178
rect 115 3002 121 4178
rect 75 2990 121 3002
rect 173 4178 219 4190
rect 173 3002 179 4178
rect 213 3002 219 4178
rect 173 2990 219 3002
rect -176 2943 -118 2949
rect -176 2909 -164 2943
rect -130 2909 -118 2943
rect -176 2903 -118 2909
rect 20 2943 78 2949
rect 20 2909 32 2943
rect 66 2909 78 2943
rect 20 2903 78 2909
rect -176 2835 -118 2841
rect -176 2801 -164 2835
rect -130 2801 -118 2835
rect -176 2795 -118 2801
rect 20 2835 78 2841
rect 20 2801 32 2835
rect 66 2801 78 2835
rect 20 2795 78 2801
rect -219 2742 -173 2754
rect -219 1566 -213 2742
rect -179 1566 -173 2742
rect -219 1554 -173 1566
rect -121 2742 -75 2754
rect -121 1566 -115 2742
rect -81 1566 -75 2742
rect -121 1554 -75 1566
rect -23 2742 23 2754
rect -23 1566 -17 2742
rect 17 1566 23 2742
rect -23 1554 23 1566
rect 75 2742 121 2754
rect 75 1566 81 2742
rect 115 1566 121 2742
rect 75 1554 121 1566
rect 173 2742 219 2754
rect 173 1566 179 2742
rect 213 1566 219 2742
rect 173 1554 219 1566
rect -78 1507 -20 1513
rect -78 1473 -66 1507
rect -32 1473 -20 1507
rect -78 1467 -20 1473
rect 118 1507 176 1513
rect 118 1473 130 1507
rect 164 1473 176 1507
rect 118 1467 176 1473
rect -78 1399 -20 1405
rect -78 1365 -66 1399
rect -32 1365 -20 1399
rect -78 1359 -20 1365
rect 118 1399 176 1405
rect 118 1365 130 1399
rect 164 1365 176 1399
rect 118 1359 176 1365
rect -219 1306 -173 1318
rect -219 130 -213 1306
rect -179 130 -173 1306
rect -219 118 -173 130
rect -121 1306 -75 1318
rect -121 130 -115 1306
rect -81 130 -75 1306
rect -121 118 -75 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 75 1306 121 1318
rect 75 130 81 1306
rect 115 130 121 1306
rect 75 118 121 130
rect 173 1306 219 1318
rect 173 130 179 1306
rect 213 130 219 1306
rect 173 118 219 130
rect -176 71 -118 77
rect -176 37 -164 71
rect -130 37 -118 71
rect -176 31 -118 37
rect 20 71 78 77
rect 20 37 32 71
rect 66 37 78 71
rect 20 31 78 37
rect -176 -37 -118 -31
rect -176 -71 -164 -37
rect -130 -71 -118 -37
rect -176 -77 -118 -71
rect 20 -37 78 -31
rect 20 -71 32 -37
rect 66 -71 78 -37
rect 20 -77 78 -71
rect -219 -130 -173 -118
rect -219 -1306 -213 -130
rect -179 -1306 -173 -130
rect -219 -1318 -173 -1306
rect -121 -130 -75 -118
rect -121 -1306 -115 -130
rect -81 -1306 -75 -130
rect -121 -1318 -75 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 75 -130 121 -118
rect 75 -1306 81 -130
rect 115 -1306 121 -130
rect 75 -1318 121 -1306
rect 173 -130 219 -118
rect 173 -1306 179 -130
rect 213 -1306 219 -130
rect 173 -1318 219 -1306
rect -78 -1365 -20 -1359
rect -78 -1399 -66 -1365
rect -32 -1399 -20 -1365
rect -78 -1405 -20 -1399
rect 118 -1365 176 -1359
rect 118 -1399 130 -1365
rect 164 -1399 176 -1365
rect 118 -1405 176 -1399
rect -78 -1473 -20 -1467
rect -78 -1507 -66 -1473
rect -32 -1507 -20 -1473
rect -78 -1513 -20 -1507
rect 118 -1473 176 -1467
rect 118 -1507 130 -1473
rect 164 -1507 176 -1473
rect 118 -1513 176 -1507
rect -219 -1566 -173 -1554
rect -219 -2742 -213 -1566
rect -179 -2742 -173 -1566
rect -219 -2754 -173 -2742
rect -121 -1566 -75 -1554
rect -121 -2742 -115 -1566
rect -81 -2742 -75 -1566
rect -121 -2754 -75 -2742
rect -23 -1566 23 -1554
rect -23 -2742 -17 -1566
rect 17 -2742 23 -1566
rect -23 -2754 23 -2742
rect 75 -1566 121 -1554
rect 75 -2742 81 -1566
rect 115 -2742 121 -1566
rect 75 -2754 121 -2742
rect 173 -1566 219 -1554
rect 173 -2742 179 -1566
rect 213 -2742 219 -1566
rect 173 -2754 219 -2742
rect -176 -2801 -118 -2795
rect -176 -2835 -164 -2801
rect -130 -2835 -118 -2801
rect -176 -2841 -118 -2835
rect 20 -2801 78 -2795
rect 20 -2835 32 -2801
rect 66 -2835 78 -2801
rect 20 -2841 78 -2835
rect -176 -2909 -118 -2903
rect -176 -2943 -164 -2909
rect -130 -2943 -118 -2909
rect -176 -2949 -118 -2943
rect 20 -2909 78 -2903
rect 20 -2943 32 -2909
rect 66 -2943 78 -2909
rect 20 -2949 78 -2943
rect -219 -3002 -173 -2990
rect -219 -4178 -213 -3002
rect -179 -4178 -173 -3002
rect -219 -4190 -173 -4178
rect -121 -3002 -75 -2990
rect -121 -4178 -115 -3002
rect -81 -4178 -75 -3002
rect -121 -4190 -75 -4178
rect -23 -3002 23 -2990
rect -23 -4178 -17 -3002
rect 17 -4178 23 -3002
rect -23 -4190 23 -4178
rect 75 -3002 121 -2990
rect 75 -4178 81 -3002
rect 115 -4178 121 -3002
rect 75 -4190 121 -4178
rect 173 -3002 219 -2990
rect 173 -4178 179 -3002
rect 213 -4178 219 -3002
rect 173 -4190 219 -4178
rect -78 -4237 -20 -4231
rect -78 -4271 -66 -4237
rect -32 -4271 -20 -4237
rect -78 -4277 -20 -4271
rect 118 -4237 176 -4231
rect 118 -4271 130 -4237
rect 164 -4271 176 -4237
rect 118 -4277 176 -4271
rect -78 -4345 -20 -4339
rect -78 -4379 -66 -4345
rect -32 -4379 -20 -4345
rect -78 -4385 -20 -4379
rect 118 -4345 176 -4339
rect 118 -4379 130 -4345
rect 164 -4379 176 -4345
rect 118 -4385 176 -4379
rect -219 -4438 -173 -4426
rect -219 -5614 -213 -4438
rect -179 -5614 -173 -4438
rect -219 -5626 -173 -5614
rect -121 -4438 -75 -4426
rect -121 -5614 -115 -4438
rect -81 -5614 -75 -4438
rect -121 -5626 -75 -5614
rect -23 -4438 23 -4426
rect -23 -5614 -17 -4438
rect 17 -5614 23 -4438
rect -23 -5626 23 -5614
rect 75 -4438 121 -4426
rect 75 -5614 81 -4438
rect 115 -5614 121 -4438
rect 75 -5626 121 -5614
rect 173 -4438 219 -4426
rect 173 -5614 179 -4438
rect 213 -5614 219 -4438
rect 173 -5626 219 -5614
rect -176 -5673 -118 -5667
rect -176 -5707 -164 -5673
rect -130 -5707 -118 -5673
rect -176 -5713 -118 -5707
rect 20 -5673 78 -5667
rect 20 -5707 32 -5673
rect 66 -5707 78 -5673
rect 20 -5713 78 -5707
<< properties >>
string FIXED_BBOX -310 -5792 310 5792
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.2 m 8 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
